// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_227 written by SynthGen on 2021/04/05 11:23:26
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_227 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1359, n1419, n1325, n1408, n1365, n1394, n1405, n1399,
 n1380, n1363, n1389, n1313, n1308, n1367, n1348, n1366,
 n1407, n1396, n2022, n2024, n2021, n2029, n2028, n2023,
 n2025, n2026, n2027, n2030, n2019, n2020, n2032, n2031);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1359, n1419, n1325, n1408, n1365, n1394, n1405, n1399,
 n1380, n1363, n1389, n1313, n1308, n1367, n1348, n1366,
 n1407, n1396, n2022, n2024, n2021, n2029, n2028, n2023,
 n2025, n2026, n2027, n2030, n2019, n2020, n2032, n2031;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1309, n1310, n1311, n1312, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1326, n1327, n1328, n1329, n1330, n1331,
 n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
 n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
 n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
 n1357, n1358, n1360, n1361, n1362, n1364, n1368, n1369,
 n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
 n1378, n1379, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1390, n1391, n1392, n1393, n1395, n1397,
 n1398, n1400, n1401, n1402, n1403, n1404, n1406, n1409,
 n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
 n1418, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018;

not  g0 (n57, n8);
buf  g1 (n64, n1);
not  g2 (n42, n2);
buf  g3 (n67, n4);
buf  g4 (n60, n7);
not  g5 (n48, n1);
not  g6 (n46, n1);
buf  g7 (n37, n2);
buf  g8 (n63, n7);
buf  g9 (n33, n5);
not  g10 (n34, n6);
not  g11 (n54, n6);
not  g12 (n50, n8);
not  g13 (n66, n9);
not  g14 (n56, n9);
buf  g15 (n36, n2);
not  g16 (n68, n9);
not  g17 (n58, n4);
not  g18 (n53, n8);
buf  g19 (n52, n7);
not  g20 (n39, n5);
not  g21 (n49, n4);
buf  g22 (n51, n3);
buf  g23 (n43, n3);
buf  g24 (n38, n1);
buf  g25 (n62, n6);
buf  g26 (n65, n7);
buf  g27 (n44, n2);
buf  g28 (n35, n6);
buf  g29 (n61, n5);
not  g30 (n41, n5);
buf  g31 (n47, n9);
not  g32 (n40, n4);
not  g33 (n55, n8);
buf  g34 (n45, n3);
not  g35 (n59, n3);
buf  g36 (n148, n51);
not  g37 (n132, n39);
buf  g38 (n104, n41);
buf  g39 (n163, n36);
not  g40 (n183, n48);
buf  g41 (n128, n61);
not  g42 (n140, n58);
buf  g43 (n113, n52);
buf  g44 (n76, n42);
not  g45 (n151, n48);
not  g46 (n185, n59);
not  g47 (n155, n34);
buf  g48 (n139, n33);
buf  g49 (n170, n63);
not  g50 (n180, n60);
buf  g51 (n95, n61);
not  g52 (n172, n52);
buf  g53 (n111, n51);
buf  g54 (n77, n63);
buf  g55 (n102, n57);
buf  g56 (n190, n54);
buf  g57 (n78, n46);
not  g58 (n165, n51);
not  g59 (n130, n45);
not  g60 (n81, n41);
buf  g61 (n84, n36);
not  g62 (n97, n43);
not  g63 (n193, n54);
not  g64 (n120, n46);
not  g65 (n150, n45);
buf  g66 (n94, n55);
buf  g67 (n116, n49);
buf  g68 (n149, n61);
not  g69 (n74, n55);
not  g70 (n160, n50);
buf  g71 (n112, n35);
buf  g72 (n184, n43);
not  g73 (n106, n40);
buf  g74 (n101, n60);
not  g75 (n147, n42);
not  g76 (n88, n37);
buf  g77 (n131, n49);
buf  g78 (n173, n50);
not  g79 (n91, n42);
buf  g80 (n100, n35);
buf  g81 (n152, n44);
buf  g82 (n98, n59);
not  g83 (n189, n39);
not  g84 (n82, n51);
not  g85 (n187, n62);
not  g86 (n182, n44);
not  g87 (n157, n62);
not  g88 (n127, n59);
not  g89 (n166, n62);
not  g90 (n79, n53);
not  g91 (n123, n53);
not  g92 (n137, n47);
not  g93 (n192, n40);
buf  g94 (n118, n56);
buf  g95 (n121, n46);
buf  g96 (n134, n48);
buf  g97 (n161, n47);
not  g98 (n73, n60);
buf  g99 (n129, n34);
not  g100 (n186, n53);
not  g101 (n144, n42);
buf  g102 (n85, n34);
not  g103 (n110, n58);
not  g104 (n158, n36);
not  g105 (n136, n52);
buf  g106 (n105, n43);
buf  g107 (n75, n38);
not  g108 (n174, n52);
buf  g109 (n176, n44);
not  g110 (n175, n39);
buf  g111 (n159, n45);
buf  g112 (n162, n58);
not  g113 (n154, n59);
not  g114 (n145, n38);
not  g115 (n171, n56);
buf  g116 (n117, n60);
not  g117 (n86, n40);
buf  g118 (n133, n35);
buf  g119 (n167, n57);
buf  g120 (n90, n37);
buf  g121 (n177, n62);
buf  g122 (n181, n35);
not  g123 (n80, n53);
not  g124 (n103, n56);
not  g125 (n146, n56);
buf  g126 (n178, n50);
not  g127 (n87, n37);
not  g128 (n93, n33);
not  g129 (n143, n45);
buf  g130 (n142, n55);
buf  g131 (n71, n54);
buf  g132 (n191, n47);
not  g133 (n107, n40);
not  g134 (n89, n43);
not  g135 (n126, n63);
buf  g136 (n122, n38);
buf  g137 (n72, n33);
buf  g138 (n135, n54);
not  g139 (n115, n58);
buf  g140 (n153, n57);
not  g141 (n108, n38);
buf  g142 (n168, n47);
buf  g143 (n138, n63);
not  g144 (n141, n49);
not  g145 (n114, n41);
not  g146 (n109, n64);
not  g147 (n83, n34);
buf  g148 (n96, n39);
not  g149 (n164, n57);
not  g150 (n119, n46);
not  g151 (n188, n49);
not  g152 (n124, n33);
buf  g153 (n92, n61);
buf  g154 (n169, n44);
buf  g155 (n179, n37);
buf  g156 (n156, n55);
not  g157 (n69, n50);
not  g158 (n70, n41);
buf  g159 (n125, n48);
buf  g160 (n99, n36);
buf  g161 (n200, n90);
not  g162 (n360, n75);
not  g163 (n667, n171);
buf  g164 (n660, n117);
not  g165 (n248, n167);
buf  g166 (n295, n91);
buf  g167 (n212, n180);
buf  g168 (n607, n187);
not  g169 (n328, n167);
not  g170 (n516, n143);
not  g171 (n428, n129);
not  g172 (n491, n171);
buf  g173 (n327, n161);
not  g174 (n333, n125);
not  g175 (n261, n172);
not  g176 (n269, n173);
buf  g177 (n355, n134);
not  g178 (n549, n123);
not  g179 (n488, n160);
not  g180 (n563, n181);
not  g181 (n278, n78);
buf  g182 (n474, n76);
not  g183 (n394, n137);
not  g184 (n230, n169);
not  g185 (n338, n157);
not  g186 (n303, n144);
not  g187 (n460, n149);
buf  g188 (n531, n92);
not  g189 (n341, n92);
not  g190 (n229, n159);
buf  g191 (n283, n116);
buf  g192 (n376, n88);
buf  g193 (n464, n179);
not  g194 (n207, n122);
buf  g195 (n445, n137);
not  g196 (n571, n79);
buf  g197 (n424, n180);
buf  g198 (n511, n112);
not  g199 (n223, n130);
buf  g200 (n203, n103);
buf  g201 (n490, n117);
not  g202 (n357, n91);
not  g203 (n354, n158);
buf  g204 (n621, n69);
buf  g205 (n425, n154);
buf  g206 (n290, n104);
buf  g207 (n204, n169);
not  g208 (n572, n124);
buf  g209 (n492, n185);
buf  g210 (n400, n121);
not  g211 (n663, n147);
buf  g212 (n397, n166);
buf  g213 (n321, n74);
not  g214 (n444, n134);
buf  g215 (n244, n163);
not  g216 (n661, n114);
buf  g217 (n461, n146);
not  g218 (n466, n87);
not  g219 (n544, n118);
not  g220 (n391, n100);
buf  g221 (n503, n91);
buf  g222 (n301, n89);
not  g223 (n656, n156);
buf  g224 (n545, n132);
not  g225 (n489, n167);
buf  g226 (n282, n114);
buf  g227 (n206, n118);
buf  g228 (n243, n79);
buf  g229 (n615, n105);
not  g230 (n408, n140);
not  g231 (n378, n185);
buf  g232 (n548, n172);
not  g233 (n584, n174);
not  g234 (n335, n93);
not  g235 (n476, n166);
buf  g236 (n276, n116);
not  g237 (n440, n80);
buf  g238 (n326, n158);
buf  g239 (n628, n77);
buf  g240 (n277, n166);
buf  g241 (n366, n126);
not  g242 (n219, n106);
not  g243 (n310, n171);
not  g244 (n271, n160);
buf  g245 (n604, n113);
not  g246 (n518, n123);
not  g247 (n555, n113);
buf  g248 (n483, n103);
not  g249 (n287, n174);
not  g250 (n241, n94);
not  g251 (n343, n168);
not  g252 (n612, n95);
not  g253 (n336, n70);
not  g254 (n600, n120);
buf  g255 (n666, n172);
not  g256 (n650, n147);
not  g257 (n358, n86);
not  g258 (n627, n165);
not  g259 (n245, n104);
buf  g260 (n586, n71);
not  g261 (n448, n73);
not  g262 (n349, n133);
not  g263 (n232, n107);
buf  g264 (n469, n180);
not  g265 (n579, n99);
not  g266 (n569, n181);
not  g267 (n194, n106);
buf  g268 (n673, n76);
not  g269 (n345, n141);
buf  g270 (n657, n156);
not  g271 (n455, n184);
not  g272 (n538, n181);
not  g273 (n613, n164);
buf  g274 (n573, n111);
not  g275 (n529, n126);
not  g276 (n433, n186);
not  g277 (n286, n87);
not  g278 (n554, n114);
buf  g279 (n553, n102);
buf  g280 (n668, n184);
buf  g281 (n582, n153);
buf  g282 (n356, n125);
not  g283 (n551, n139);
not  g284 (n405, n128);
buf  g285 (n399, n137);
not  g286 (n209, n149);
buf  g287 (n198, n86);
buf  g288 (n373, n119);
buf  g289 (n382, n72);
not  g290 (n350, n175);
not  g291 (n616, n103);
not  g292 (n514, n182);
not  g293 (n467, n149);
buf  g294 (n452, n145);
buf  g295 (n258, n99);
not  g296 (n380, n147);
not  g297 (n435, n108);
not  g298 (n498, n116);
not  g299 (n669, n109);
buf  g300 (n386, n78);
buf  g301 (n524, n156);
buf  g302 (n462, n182);
not  g303 (n449, n186);
not  g304 (n426, n69);
buf  g305 (n251, n78);
buf  g306 (n504, n135);
not  g307 (n395, n183);
buf  g308 (n371, n176);
buf  g309 (n337, n101);
buf  g310 (n527, n136);
buf  g311 (n329, n158);
buf  g312 (n369, n96);
not  g313 (n353, n97);
buf  g314 (n617, n126);
not  g315 (n671, n110);
buf  g316 (n635, n111);
buf  g317 (n332, n104);
buf  g318 (n305, n127);
not  g319 (n446, n148);
buf  g320 (n252, n100);
buf  g321 (n540, n89);
not  g322 (n228, n94);
not  g323 (n453, n85);
buf  g324 (n606, n136);
buf  g325 (n331, n176);
buf  g326 (n249, n178);
buf  g327 (n471, n79);
buf  g328 (n609, n94);
not  g329 (n562, n132);
buf  g330 (n221, n122);
not  g331 (n642, n170);
not  g332 (n383, n76);
not  g333 (n222, n164);
not  g334 (n557, n82);
buf  g335 (n523, n73);
not  g336 (n525, n83);
not  g337 (n259, n99);
not  g338 (n289, n154);
not  g339 (n316, n108);
not  g340 (n575, n135);
buf  g341 (n659, n157);
buf  g342 (n239, n161);
not  g343 (n567, n168);
buf  g344 (n414, n70);
not  g345 (n296, n82);
not  g346 (n497, n177);
buf  g347 (n533, n181);
buf  g348 (n412, n110);
not  g349 (n318, n185);
buf  g350 (n547, n101);
buf  g351 (n284, n150);
buf  g352 (n515, n134);
buf  g353 (n417, n74);
not  g354 (n441, n77);
not  g355 (n274, n159);
not  g356 (n570, n119);
buf  g357 (n348, n74);
buf  g358 (n447, n87);
buf  g359 (n247, n141);
buf  g360 (n298, n186);
buf  g361 (n513, n76);
not  g362 (n205, n131);
not  g363 (n493, n84);
not  g364 (n478, n138);
buf  g365 (n392, n75);
not  g366 (n377, n98);
not  g367 (n655, n141);
not  g368 (n208, n141);
buf  g369 (n402, n112);
buf  g370 (n591, n113);
buf  g371 (n398, n153);
not  g372 (n450, n124);
not  g373 (n262, n178);
not  g374 (n431, n169);
not  g375 (n599, n164);
not  g376 (n368, n168);
not  g377 (n451, n119);
buf  g378 (n534, n144);
not  g379 (n496, n140);
buf  g380 (n566, n94);
buf  g381 (n434, n99);
not  g382 (n253, n95);
not  g383 (n519, n179);
not  g384 (n201, n120);
buf  g385 (n564, n130);
buf  g386 (n611, n128);
not  g387 (n304, n73);
not  g388 (n587, n160);
buf  g389 (n257, n148);
buf  g390 (n280, n165);
buf  g391 (n231, n154);
not  g392 (n535, n172);
not  g393 (n281, n152);
not  g394 (n324, n145);
buf  g395 (n499, n109);
not  g396 (n211, n95);
not  g397 (n308, n79);
not  g398 (n639, n152);
not  g399 (n517, n128);
not  g400 (n279, n89);
not  g401 (n552, n72);
not  g402 (n605, n175);
not  g403 (n658, n188);
not  g404 (n456, n97);
not  g405 (n590, n102);
buf  g406 (n352, n187);
not  g407 (n665, n165);
buf  g408 (n215, n110);
not  g409 (n195, n157);
not  g410 (n236, n90);
buf  g411 (n644, n127);
buf  g412 (n422, n121);
not  g413 (n472, n170);
buf  g414 (n311, n96);
not  g415 (n463, n186);
buf  g416 (n265, n187);
buf  g417 (n521, n122);
buf  g418 (n436, n140);
not  g419 (n646, n188);
buf  g420 (n539, n182);
not  g421 (n411, n75);
buf  g422 (n583, n142);
buf  g423 (n415, n163);
buf  g424 (n292, n105);
buf  g425 (n420, n83);
buf  g426 (n662, n110);
buf  g427 (n477, n149);
not  g428 (n625, n182);
not  g429 (n294, n82);
buf  g430 (n409, n143);
not  g431 (n473, n139);
buf  g432 (n626, n144);
buf  g433 (n390, n130);
buf  g434 (n220, n70);
not  g435 (n217, n146);
not  g436 (n254, n155);
buf  g437 (n647, n85);
buf  g438 (n481, n97);
buf  g439 (n593, n174);
not  g440 (n653, n140);
buf  g441 (n559, n118);
not  g442 (n260, n169);
buf  g443 (n214, n74);
buf  g444 (n196, n171);
buf  g445 (n300, n73);
not  g446 (n293, n81);
not  g447 (n313, n142);
buf  g448 (n375, n107);
not  g449 (n597, n88);
buf  g450 (n307, n183);
not  g451 (n317, n115);
buf  g452 (n225, n125);
buf  g453 (n309, n134);
not  g454 (n407, n162);
buf  g455 (n631, n111);
buf  g456 (n643, n162);
buf  g457 (n624, n150);
buf  g458 (n528, n109);
buf  g459 (n351, n86);
not  g460 (n306, n84);
not  g461 (n379, n78);
buf  g462 (n648, n167);
buf  g463 (n581, n152);
not  g464 (n346, n83);
buf  g465 (n413, n152);
not  g466 (n427, n80);
not  g467 (n442, n123);
not  g468 (n510, n173);
not  g469 (n410, n183);
not  g470 (n325, n111);
buf  g471 (n598, n162);
not  g472 (n601, n153);
not  g473 (n637, n176);
buf  g474 (n363, n139);
buf  g475 (n302, n75);
buf  g476 (n330, n116);
buf  g477 (n319, n177);
not  g478 (n418, n165);
not  g479 (n640, n154);
not  g480 (n250, n183);
buf  g481 (n482, n170);
not  g482 (n256, n101);
not  g483 (n585, n129);
buf  g484 (n384, n102);
buf  g485 (n588, n95);
not  g486 (n416, n127);
not  g487 (n213, n115);
buf  g488 (n266, n129);
buf  g489 (n475, n131);
buf  g490 (n288, n71);
not  g491 (n505, n187);
not  g492 (n234, n131);
not  g493 (n634, n142);
not  g494 (n226, n151);
not  g495 (n273, n184);
not  g496 (n340, n112);
not  g497 (n596, n174);
not  g498 (n501, n91);
not  g499 (n536, n119);
not  g500 (n361, n161);
not  g501 (n320, n123);
buf  g502 (n419, n166);
not  g503 (n314, n93);
not  g504 (n439, n144);
not  g505 (n502, n179);
not  g506 (n430, n109);
not  g507 (n454, n178);
buf  g508 (n537, n104);
buf  g509 (n576, n98);
buf  g510 (n216, n86);
buf  g511 (n423, n118);
not  g512 (n610, n136);
buf  g513 (n465, n147);
buf  g514 (n556, n122);
buf  g515 (n396, n163);
buf  g516 (n494, n132);
buf  g517 (n237, n173);
not  g518 (n568, n170);
not  g519 (n602, n115);
not  g520 (n458, n146);
not  g521 (n334, n163);
buf  g522 (n509, n162);
not  g523 (n651, n80);
not  g524 (n297, n71);
buf  g525 (n485, n132);
not  g526 (n654, n83);
buf  g527 (n470, n179);
not  g528 (n622, n69);
buf  g529 (n227, n131);
buf  g530 (n370, n84);
not  g531 (n636, n106);
not  g532 (n242, n176);
not  g533 (n233, n145);
not  g534 (n393, n126);
buf  g535 (n255, n112);
buf  g536 (n620, n92);
buf  g537 (n339, n173);
not  g538 (n558, n97);
not  g539 (n438, n150);
not  g540 (n486, n69);
buf  g541 (n578, n160);
buf  g542 (n546, n155);
buf  g543 (n672, n184);
not  g544 (n526, n77);
not  g545 (n291, n77);
not  g546 (n421, n159);
not  g547 (n389, n138);
buf  g548 (n520, n138);
not  g549 (n388, n130);
not  g550 (n268, n177);
buf  g551 (n315, n88);
not  g552 (n618, n71);
buf  g553 (n652, n81);
not  g554 (n638, n178);
not  g555 (n580, n106);
not  g556 (n312, n98);
not  g557 (n614, n72);
buf  g558 (n322, n127);
buf  g559 (n574, n142);
not  g560 (n630, n143);
not  g561 (n344, n96);
not  g562 (n238, n129);
buf  g563 (n565, n151);
not  g564 (n364, n72);
not  g565 (n495, n100);
not  g566 (n619, n107);
not  g567 (n365, n177);
buf  g568 (n542, n180);
not  g569 (n210, n136);
buf  g570 (n272, n84);
buf  g571 (n595, n137);
buf  g572 (n506, n135);
buf  g573 (n632, n175);
buf  g574 (n374, n81);
buf  g575 (n432, n105);
not  g576 (n664, n156);
not  g577 (n670, n90);
buf  g578 (n246, n159);
buf  g579 (n459, n133);
not  g580 (n649, n80);
not  g581 (n385, n185);
not  g582 (n508, n85);
not  g583 (n347, n155);
buf  g584 (n468, n89);
buf  g585 (n641, n146);
not  g586 (n264, n108);
not  g587 (n629, n108);
not  g588 (n530, n103);
buf  g589 (n543, n120);
buf  g590 (n267, n93);
not  g591 (n603, n133);
buf  g592 (n199, n150);
buf  g593 (n359, n124);
not  g594 (n406, n138);
buf  g595 (n577, n135);
buf  g596 (n479, n121);
buf  g597 (n263, n100);
not  g598 (n197, n164);
buf  g599 (n429, n120);
buf  g600 (n323, n139);
not  g601 (n457, n113);
buf  g602 (n608, n82);
not  g603 (n561, n98);
not  g604 (n594, n125);
buf  g605 (n372, n124);
buf  g606 (n522, n90);
not  g607 (n270, n107);
not  g608 (n403, n175);
not  g609 (n592, n128);
buf  g610 (n387, n188);
not  g611 (n240, n81);
not  g612 (n550, n105);
not  g613 (n401, n85);
buf  g614 (n512, n145);
not  g615 (n560, n70);
buf  g616 (n487, n87);
not  g617 (n224, n117);
buf  g618 (n532, n158);
buf  g619 (n541, n121);
not  g620 (n235, n115);
not  g621 (n645, n102);
not  g622 (n342, n148);
buf  g623 (n285, n117);
not  g624 (n437, n157);
buf  g625 (n443, n143);
buf  g626 (n633, n161);
buf  g627 (n507, n101);
not  g628 (n589, n88);
buf  g629 (n202, n92);
buf  g630 (n480, n148);
not  g631 (n218, n151);
buf  g632 (n484, n93);
buf  g633 (n299, n114);
buf  g634 (n623, n188);
not  g635 (n362, n151);
buf  g636 (n500, n155);
buf  g637 (n381, n168);
not  g638 (n275, n96);
not  g639 (n367, n153);
not  g640 (n404, n133);
buf  g641 (n1204, n662);
buf  g642 (n1147, n616);
not  g643 (n1073, n488);
not  g644 (n1201, n662);
not  g645 (n1067, n631);
buf  g646 (n1274, n326);
buf  g647 (n880, n379);
buf  g648 (n1223, n441);
not  g649 (n1183, n510);
not  g650 (n775, n431);
not  g651 (n822, n255);
not  g652 (n1170, n302);
buf  g653 (n1031, n285);
buf  g654 (n942, n269);
buf  g655 (n732, n491);
buf  g656 (n953, n259);
buf  g657 (n800, n489);
not  g658 (n1015, n292);
not  g659 (n864, n248);
buf  g660 (n1236, n583);
buf  g661 (n1174, n370);
buf  g662 (n714, n643);
buf  g663 (n674, n593);
buf  g664 (n1024, n545);
not  g665 (n939, n327);
buf  g666 (n769, n562);
not  g667 (n934, n488);
buf  g668 (n1007, n537);
buf  g669 (n1190, n360);
not  g670 (n1257, n547);
not  g671 (n761, n251);
buf  g672 (n831, n272);
not  g673 (n998, n602);
buf  g674 (n947, n530);
not  g675 (n1180, n385);
not  g676 (n794, n481);
not  g677 (n1193, n353);
buf  g678 (n772, n252);
buf  g679 (n1254, n548);
not  g680 (n1019, n432);
buf  g681 (n784, n432);
not  g682 (n1033, n544);
not  g683 (n1296, n490);
buf  g684 (n1112, n313);
buf  g685 (n811, n526);
not  g686 (n711, n485);
buf  g687 (n762, n449);
buf  g688 (n684, n448);
buf  g689 (n720, n483);
not  g690 (n1069, n591);
not  g691 (n861, n340);
buf  g692 (n1277, n327);
not  g693 (n1253, n585);
not  g694 (n1087, n278);
not  g695 (n1111, n572);
not  g696 (n1049, n568);
not  g697 (n773, n474);
buf  g698 (n923, n461);
not  g699 (n853, n212);
buf  g700 (n1068, n619);
not  g701 (n882, n380);
not  g702 (n1238, n300);
buf  g703 (n1187, n386);
buf  g704 (n1098, n418);
not  g705 (n850, n664);
not  g706 (n1205, n436);
buf  g707 (n852, n422);
not  g708 (n1215, n533);
not  g709 (n890, n457);
buf  g710 (n685, n526);
not  g711 (n1272, n531);
buf  g712 (n952, n261);
buf  g713 (n1291, n527);
buf  g714 (n870, n349);
not  g715 (n983, n366);
buf  g716 (n1262, n550);
buf  g717 (n807, n380);
buf  g718 (n962, n524);
not  g719 (n1000, n344);
buf  g720 (n1138, n503);
not  g721 (n678, n413);
not  g722 (n957, n468);
not  g723 (n989, n483);
buf  g724 (n1171, n594);
buf  g725 (n965, n507);
not  g726 (n716, n308);
not  g727 (n888, n237);
not  g728 (n1284, n373);
not  g729 (n1305, n307);
buf  g730 (n1212, n576);
not  g731 (n1189, n460);
buf  g732 (n781, n357);
not  g733 (n1036, n509);
buf  g734 (n1157, n534);
buf  g735 (n845, n618);
not  g736 (n854, n260);
buf  g737 (n1026, n547);
not  g738 (n1139, n575);
not  g739 (n1005, n548);
buf  g740 (n742, n664);
buf  g741 (n1158, n549);
buf  g742 (n1041, n371);
not  g743 (n760, n583);
buf  g744 (n1125, n260);
buf  g745 (n747, n552);
not  g746 (n1283, n581);
not  g747 (n1259, n456);
not  g748 (n844, n396);
buf  g749 (n799, n385);
buf  g750 (n791, n534);
not  g751 (n1050, n601);
not  g752 (n897, n461);
not  g753 (n839, n633);
not  g754 (n1129, n226);
not  g755 (n721, n241);
not  g756 (n901, n419);
buf  g757 (n1163, n546);
buf  g758 (n833, n651);
buf  g759 (n886, n516);
not  g760 (n1270, n258);
not  g761 (n1121, n498);
not  g762 (n1248, n340);
buf  g763 (n1235, n590);
not  g764 (n697, n194);
not  g765 (n1148, n561);
buf  g766 (n1232, n359);
buf  g767 (n765, n194);
buf  g768 (n759, n417);
buf  g769 (n1243, n567);
not  g770 (n806, n433);
buf  g771 (n948, n379);
buf  g772 (n1058, n630);
not  g773 (n702, n245);
not  g774 (n1197, n350);
buf  g775 (n1079, n355);
not  g776 (n986, n347);
buf  g777 (n1292, n356);
not  g778 (n745, n497);
not  g779 (n1159, n480);
not  g780 (n744, n457);
not  g781 (n804, n603);
buf  g782 (n1186, n569);
not  g783 (n676, n394);
not  g784 (n730, n300);
not  g785 (n900, n576);
not  g786 (n715, n403);
not  g787 (n1255, n211);
buf  g788 (n988, n455);
buf  g789 (n1208, n661);
buf  g790 (n1293, n500);
buf  g791 (n696, n555);
not  g792 (n1221, n342);
not  g793 (n1302, n506);
buf  g794 (n894, n639);
not  g795 (n1074, n580);
buf  g796 (n798, n561);
buf  g797 (n1128, n428);
buf  g798 (n812, n433);
not  g799 (n788, n202);
buf  g800 (n736, n405);
buf  g801 (n1055, n558);
not  g802 (n891, n662);
not  g803 (n789, n209);
not  g804 (n1018, n527);
buf  g805 (n825, n548);
not  g806 (n985, n587);
not  g807 (n677, n303);
not  g808 (n1169, n382);
buf  g809 (n937, n475);
not  g810 (n940, n538);
buf  g811 (n921, n326);
not  g812 (n1116, n558);
not  g813 (n733, n327);
buf  g814 (n911, n605);
buf  g815 (n691, n210);
buf  g816 (n1165, n508);
buf  g817 (n1027, n204);
buf  g818 (n731, n472);
buf  g819 (n1273, n227);
buf  g820 (n680, n287);
buf  g821 (n1130, n638);
buf  g822 (n1135, n201);
buf  g823 (n686, n278);
buf  g824 (n1146, n436);
not  g825 (n1084, n557);
not  g826 (n776, n637);
buf  g827 (n1249, n646);
not  g828 (n902, n606);
not  g829 (n840, n220);
buf  g830 (n1075, n331);
not  g831 (n1188, n393);
buf  g832 (n1127, n320);
not  g833 (n1141, n649);
buf  g834 (n1006, n665);
not  g835 (n827, n500);
buf  g836 (n1251, n264);
not  g837 (n1017, n612);
not  g838 (n1252, n641);
not  g839 (n1172, n450);
not  g840 (n828, n446);
not  g841 (n824, n509);
not  g842 (n1306, n487);
not  g843 (n1271, n614);
not  g844 (n1056, n610);
not  g845 (n838, n357);
not  g846 (n797, n234);
not  g847 (n914, n521);
not  g848 (n846, n412);
not  g849 (n1207, n459);
buf  g850 (n991, n536);
not  g851 (n1156, n218);
buf  g852 (n754, n359);
not  g853 (n1016, n625);
not  g854 (n767, n393);
buf  g855 (n785, n301);
buf  g856 (n1229, n287);
not  g857 (n735, n258);
not  g858 (n1288, n508);
not  g859 (n1009, n383);
not  g860 (n1126, n663);
buf  g861 (n866, n453);
not  g862 (n1286, n508);
not  g863 (n813, n362);
not  g864 (n972, n646);
buf  g865 (n927, n617);
not  g866 (n1168, n659);
not  g867 (n1118, n473);
buf  g868 (n995, n570);
not  g869 (n943, n537);
not  g870 (n1195, n590);
not  g871 (n787, n354);
buf  g872 (n1011, n510);
not  g873 (n1083, n532);
not  g874 (n830, n318);
not  g875 (n795, n554);
buf  g876 (n909, n373);
not  g877 (n1029, n573);
buf  g878 (n722, n549);
not  g879 (n1176, n467);
not  g880 (n1136, n513);
not  g881 (n1153, n434);
buf  g882 (n1088, n631);
buf  g883 (n1239, n429);
buf  g884 (n1061, n606);
not  g885 (n1131, n504);
buf  g886 (n1103, n585);
not  g887 (n763, n376);
not  g888 (n757, n590);
not  g889 (n878, n652);
buf  g890 (n1117, n620);
not  g891 (n933, n655);
buf  g892 (n1295, n350);
not  g893 (n1150, n641);
buf  g894 (n1234, n529);
not  g895 (n837, n198);
not  g896 (n1053, n494);
buf  g897 (n961, n435);
not  g898 (n1022, n299);
not  g899 (n1166, n408);
buf  g900 (n1216, n316);
not  g901 (n862, n537);
not  g902 (n1185, n608);
not  g903 (n1267, n361);
buf  g904 (n768, n536);
not  g905 (n1045, n597);
not  g906 (n774, n619);
not  g907 (n826, n376);
buf  g908 (n1093, n279);
not  g909 (n930, n235);
not  g910 (n740, n271);
buf  g911 (n792, n268);
buf  g912 (n1104, n659);
not  g913 (n692, n552);
not  g914 (n1242, n235);
not  g915 (n750, n581);
not  g916 (n741, n376);
not  g917 (n949, n652);
buf  g918 (n1012, n284);
buf  g919 (n1108, n564);
not  g920 (n1096, n451);
buf  g921 (n938, n411);
not  g922 (n867, n371);
buf  g923 (n778, n493);
not  g924 (n908, n495);
buf  g925 (n1099, n466);
buf  g926 (n1113, n223);
buf  g927 (n782, n666);
not  g928 (n1210, n584);
not  g929 (n1301, n563);
buf  g930 (n1294, n543);
not  g931 (n910, n336);
buf  g932 (n1278, n499);
not  g933 (n1280, n575);
buf  g934 (n941, n311);
not  g935 (n1032, n422);
not  g936 (n1155, n280);
buf  g937 (n1137, n242);
not  g938 (n887, n334);
not  g939 (n699, n665);
not  g940 (n956, n563);
not  g941 (n1152, n505);
not  g942 (n1192, n265);
not  g943 (n1124, n497);
buf  g944 (n932, n646);
not  g945 (n1132, n229);
not  g946 (n918, n221);
buf  g947 (n1106, n567);
or   g948 (n821, n487, n565);
xor  g949 (n996, n427, n613, n642, n640);
xnor g950 (n1091, n529, n495, n580, n334);
and  g951 (n803, n622, n375, n205, n525);
nand g952 (n1085, n615, n565, n457, n362);
xor  g953 (n734, n625, n532, n339, n542);
xnor g954 (n1082, n227, n614, n242, n586);
and  g955 (n1025, n245, n473, n656, n210);
or   g956 (n1122, n421, n424, n535, n338);
and  g957 (n977, n424, n574, n541, n324);
and  g958 (n1162, n476, n597, n647, n617);
or   g959 (n1244, n372, n451, n201, n540);
or   g960 (n1179, n529, n463, n526, n258);
and  g961 (n703, n312, n462, n530, n636);
xor  g962 (n975, n208, n402, n454, n533);
nand g963 (n1037, n319, n635, n648, n580);
nor  g964 (n951, n553, n348, n278, n496);
or   g965 (n842, n356, n539, n357, n566);
nand g966 (n694, n507, n489, n562, n661);
nand g967 (n907, n621, n615, n539, n656);
nand g968 (n978, n232, n455, n238, n513);
xor  g969 (n1047, n654, n294, n265, n414);
xnor g970 (n992, n216, n465, n643, n320);
nor  g971 (n832, n296, n572, n281, n314);
xor  g972 (n1028, n396, n471, n435, n264);
xor  g973 (n1203, n663, n553, n384, n574);
xnor g974 (n1034, n607, n513, n341, n617);
nor  g975 (n857, n288, n595, n637, n262);
nand g976 (n718, n522, n657, n399, n263);
and  g977 (n805, n557, n661, n587, n406);
or   g978 (n1241, n577, n427, n621, n472);
xor  g979 (n979, n593, n219, n560, n259);
and  g980 (n698, n305, n622, n498, n542);
or   g981 (n823, n499, n337, n524, n571);
xor  g982 (n871, n494, n415, n525, n523);
nor  g983 (n1289, n374, n284, n481, n582);
xor  g984 (n879, n667, n407, n316, n578);
or   g985 (n1133, n213, n443, n520, n308);
nand g986 (n884, n405, n502, n601, n249);
nor  g987 (n1281, n197, n212, n564, n341);
or   g988 (n755, n344, n540, n616, n409);
or   g989 (n1003, n416, n592, n391, n559);
and  g990 (n1200, n570, n471, n220, n636);
xor  g991 (n1151, n381, n618, n206, n636);
xor  g992 (n1237, n512, n280, n629, n616);
xnor g993 (n1268, n426, n378, n507, n562);
nor  g994 (n847, n377, n198, n369, n365);
xnor g995 (n924, n276, n640, n516, n253);
or   g996 (n1102, n632, n361, n288, n245);
or   g997 (n1094, n453, n386, n352, n635);
xnor g998 (n1202, n624, n414, n527, n574);
or   g999 (n1046, n332, n597, n415, n544);
xnor g1000 (n958, n626, n239, n506, n627);
nand g1001 (n1266, n390, n476, n450, n647);
or   g1002 (n1043, n390, n283, n249, n506);
xor  g1003 (n920, n464, n528, n293, n484);
nor  g1004 (n1004, n372, n465, n454, n664);
nor  g1005 (n1107, n530, n639, n657, n465);
xnor g1006 (n916, n511, n223, n404, n668);
or   g1007 (n877, n195, n477, n325, n575);
xnor g1008 (n849, n217, n501, n210, n459);
xor  g1009 (n802, n346, n207, n596, n446);
or   g1010 (n1057, n282, n292, n248, n440);
xnor g1011 (n751, n338, n516, n573, n217);
xnor g1012 (n896, n346, n631, n588, n603);
and  g1013 (n1245, n293, n502, n215, n574);
nand g1014 (n1123, n491, n659, n242, n401);
xor  g1015 (n1178, n195, n602, n598, n224);
xor  g1016 (n841, n227, n214, n662, n234);
and  g1017 (n818, n230, n218, n556, n231);
and  g1018 (n967, n420, n269, n318, n215);
nor  g1019 (n708, n428, n304, n467, n642);
and  g1020 (n1071, n462, n272, n664, n283);
xor  g1021 (n1065, n244, n600, n650, n496);
and  g1022 (n860, n241, n543, n458, n304);
xnor g1023 (n1051, n640, n347, n433, n487);
xor  g1024 (n1140, n214, n305, n228, n430);
nand g1025 (n1228, n564, n290, n307, n288);
xnor g1026 (n873, n613, n480, n651, n605);
xor  g1027 (n1224, n617, n497, n246, n535);
nor  g1028 (n1149, n388, n482, n598, n266);
nor  g1029 (n1142, n352, n531, n292, n403);
xor  g1030 (n1198, n250, n626, n651, n211);
xnor g1031 (n710, n524, n271, n360, n269);
xor  g1032 (n1115, n200, n594, n367, n503);
or   g1033 (n926, n594, n622, n641, n539);
and  g1034 (n881, n382, n213, n592, n419);
and  g1035 (n971, n667, n295, n324, n235);
nor  g1036 (n816, n570, n351, n466, n301);
and  g1037 (n1021, n343, n485, n569, n321);
xnor g1038 (n994, n222, n525, n440, n252);
and  g1039 (n1039, n398, n427, n409, n544);
or   g1040 (n981, n391, n632, n563, n634);
or   g1041 (n898, n576, n528, n483, n253);
nand g1042 (n915, n445, n517, n225, n470);
nor  g1043 (n738, n601, n642, n520, n266);
and  g1044 (n1077, n630, n343, n541, n656);
nor  g1045 (n817, n328, n612, n576, n444);
xnor g1046 (n683, n443, n234, n379, n349);
and  g1047 (n700, n416, n440, n265, n231);
nand g1048 (n843, n554, n492, n238, n384);
or   g1049 (n976, n665, n639, n501, n577);
or   g1050 (n709, n322, n481, n639, n398);
nor  g1051 (n1044, n255, n623, n587);
nand g1052 (n969, n332, n203, n489, n545);
xor  g1053 (n728, n374, n513, n626, n416);
xor  g1054 (n1062, n584, n231, n389, n289);
nand g1055 (n945, n502, n545, n546, n666);
xnor g1056 (n743, n279, n628, n203, n579);
nand g1057 (n1089, n287, n423, n552, n318);
and  g1058 (n1191, n609, n549, n222, n610);
xnor g1059 (n1109, n455, n420, n607, n402);
and  g1060 (n793, n658, n660, n566, n530);
nor  g1061 (n689, n275, n511, n356, n239);
xnor g1062 (n913, n322, n631, n573, n329);
xnor g1063 (n869, n392, n325, n538, n536);
nor  g1064 (n770, n329, n589, n644, n246);
or   g1065 (n893, n567, n529, n363, n298);
or   g1066 (n928, n474, n232, n374, n406);
or   g1067 (n1164, n358, n390, n644, n490);
or   g1068 (n987, n509, n510, n531, n309);
xor  g1069 (n829, n330, n603, n550, n657);
nor  g1070 (n1101, n615, n519, n448, n508);
xor  g1071 (n705, n236, n444, n492, n611);
nor  g1072 (n1260, n368, n568, n205, n605);
or   g1073 (n1080, n666, n479, n599, n504);
or   g1074 (n865, n303, n488, n425, n498);
nand g1075 (n1048, n279, n521, n533, n397);
nor  g1076 (n858, n503, n504, n600, n247);
nor  g1077 (n1086, n290, n438, n600, n451);
nor  g1078 (n964, n226, n647, n404, n634);
nor  g1079 (n695, n586, n604, n616, n353);
xor  g1080 (n1052, n475, n493, n435, n309);
xor  g1081 (n1010, n239, n645, n442, n262);
xor  g1082 (n1290, n456, n445, n407, n270);
xnor g1083 (n1144, n406, n439, n313, n216);
xnor g1084 (n1298, n518, n593, n423, n408);
or   g1085 (n723, n371, n609, n360, n370);
and  g1086 (n999, n246, n241, n546, n355);
nand g1087 (n1184, n591, n472, n522, n314);
xor  g1088 (n856, n335, n559, n629, n200);
or   g1089 (n906, n620, n468, n375, n667);
nor  g1090 (n1275, n467, n436, n524, n586);
xnor g1091 (n1240, n389, n577, n237, n589);
and  g1092 (n727, n658, n302, n291, n648);
nor  g1093 (n790, n654, n375, n306, n476);
nand g1094 (n968, n233, n640, n614, n295);
or   g1095 (n1120, n250, n447, n251, n648);
xnor g1096 (n779, n553, n518, n495, n470);
xor  g1097 (n859, n470, n458, n229, n273);
and  g1098 (n820, n583, n607, n599, n262);
nor  g1099 (n1160, n211, n257, n196, n395);
xnor g1100 (n931, n315, n633, n500, n654);
xor  g1101 (n681, n502, n625, n547, n453);
nor  g1102 (n1269, n571, n326, n342, n652);
or   g1103 (n1219, n335, n447, n229, n532);
nor  g1104 (n835, n209, n209, n256, n604);
nor  g1105 (n726, n517, n348, n388, n395);
and  g1106 (n980, n535, n303, n491, n512);
or   g1107 (n868, n382, n422, n385, n541);
xnor g1108 (n693, n215, n638, n421, n297);
nor  g1109 (n737, n222, n543, n459, n412);
nand g1110 (n758, n207, n660, n523, n315);
xnor g1111 (n1217, n514, n638, n458, n238);
nor  g1112 (n1173, n598, n236, n311, n558);
or   g1113 (n724, n243, n346, n333, n214);
or   g1114 (n1285, n487, n264, n256, n551);
nor  g1115 (n1070, n466, n635, n663, n282);
xor  g1116 (n706, n352, n620, n545, n413);
nor  g1117 (n1035, n339, n399, n198, n197);
nand g1118 (n766, n381, n469, n417, n637);
and  g1119 (n1211, n368, n590, n283, n627);
xnor g1120 (n936, n329, n270, n551, n354);
xnor g1121 (n1276, n469, n650, n626, n212);
and  g1122 (n1233, n366, n527, n522, n606);
or   g1123 (n717, n392, n557, n645, n471);
nand g1124 (n1076, n525, n349, n655, n537);
and  g1125 (n780, n341, n253, n217, n409);
and  g1126 (n1090, n539, n478, n595, n582);
xnor g1127 (n912, n598, n339, n514, n237);
nand g1128 (n810, n332, n263, n257, n522);
and  g1129 (n771, n503, n653, n331, n420);
xnor g1130 (n1078, n547, n397, n314, n496);
and  g1131 (n1063, n500, n532, n490, n542);
or   g1132 (n917, n649, n606, n568, n267);
nand g1133 (n929, n304, n634, n504, n610);
xnor g1134 (n752, n270, n347, n251, n591);
nand g1135 (n1002, n443, n306, n589, n659);
xnor g1136 (n1227, n200, n228, n225, n540);
nor  g1137 (n713, n660, n280, n232, n515);
nor  g1138 (n834, n653, n423, n493, n482);
or   g1139 (n707, n611, n308, n244, n560);
xor  g1140 (n1054, n515, n650, n431, n534);
nor  g1141 (n960, n597, n483, n560, n413);
or   g1142 (n1110, n315, n351, n604, n286);
and  g1143 (n1299, n400, n337, n646, n355);
nor  g1144 (n1161, n464, n494, n381, n387);
xor  g1145 (n1175, n260, n498, n521, n195);
xor  g1146 (n756, n310, n515, n311, n600);
and  g1147 (n1100, n577, n221, n199, n444);
or   g1148 (n970, n437, n328, n221, n225);
and  g1149 (n872, n439, n594, n383, n549);
nor  g1150 (n1226, n307, n401, n516, n561);
nand g1151 (n863, n384, n634, n243, n538);
and  g1152 (n899, n573, n492, n336, n319);
xor  g1153 (n712, n223, n592, n257, n452);
xnor g1154 (n749, n410, n219, n555, n660);
or   g1155 (n984, n644, n507, n296, n541);
or   g1156 (n959, n557, n570, n480, n236);
or   g1157 (n1038, n430, n358, n528, n563);
xnor g1158 (n1182, n250, n395, n201, n578);
and  g1159 (n1279, n625, n254, n521, n648);
and  g1160 (n704, n627, n194, n448, n266);
xnor g1161 (n719, n407, n367, n589, n274);
and  g1162 (n801, n559, n197, n437, n377);
xor  g1163 (n876, n658, n593, n560, n431);
xnor g1164 (n1300, n285, n544, n401, n585);
xor  g1165 (n883, n608, n555, n484, n567);
and  g1166 (n1119, n556, n474, n566, n249);
nor  g1167 (n950, n581, n542, n636, n267);
or   g1168 (n1167, n477, n628, n603, n526);
nor  g1169 (n1040, n400, n312, n515, n389);
nand g1170 (n1023, n338, n643, n322, n632);
nor  g1171 (n796, n571, n365, n437, n647);
and  g1172 (n1097, n538, n601, n226, n482);
xor  g1173 (n725, n452, n429, n216, n599);
xnor g1174 (n1134, n334, n224, n272, n312);
xnor g1175 (n1247, n536, n452, n313, n403);
xor  g1176 (n1209, n386, n321, n377, n621);
nand g1177 (n851, n387, n240, n464, n319);
xnor g1178 (n903, n276, n333, n495, n584);
xor  g1179 (n1145, n438, n316, n587, n410);
xnor g1180 (n889, n275, n337, n551, n494);
or   g1181 (n1114, n579, n578, n552, n460);
nor  g1182 (n954, n364, n613, n259, n233);
and  g1183 (n836, n298, n614, n441, n657);
nor  g1184 (n922, n628, n432, n310, n429);
and  g1185 (n748, n393, n363, n203, n523);
or   g1186 (n777, n290, n608, n419, n641);
or   g1187 (n815, n535, n665, n588, n348);
and  g1188 (n1042, n445, n363, n405, n196);
xor  g1189 (n679, n629, n533, n492, n294);
or   g1190 (n855, n276, n298, n596, n421);
nor  g1191 (n1066, n378, n565, n543);
xor  g1192 (n1081, n621, n268, n309, n302);
xor  g1193 (n1287, n633, n612, n463, n486);
xor  g1194 (n966, n497, n398, n450, n619);
nand g1195 (n687, n428, n323, n592, n568);
or   g1196 (n753, n218, n638, n449, n252);
or   g1197 (n1264, n628, n208, n425, n330);
or   g1198 (n1013, n528, n281, n369, n284);
nand g1199 (n809, n499, n637, n324, n299);
nor  g1200 (n997, n642, n645, n305, n478);
and  g1201 (n990, n282, n268, n359, n501);
and  g1202 (n955, n248, n206, n604, n486);
xor  g1203 (n1014, n566, n512, n317, n571);
xor  g1204 (n1256, n442, n596, n572, n294);
xnor g1205 (n1220, n556, n418, n651, n479);
and  g1206 (n1230, n297, n514, n486, n582);
xor  g1207 (n1231, n523, n364, n372, n417);
xnor g1208 (n786, n618, n373, n654, n519);
nor  g1209 (n1154, n475, n383, n402, n623);
xnor g1210 (n1143, n430, n345, n354, n666);
xnor g1211 (n1095, n286, n342, n425, n202);
nand g1212 (n1263, n622, n220, n564, n244);
xor  g1213 (n885, n653, n396, n485, n608);
xor  g1214 (n701, n439, n602, n496);
nand g1215 (n1265, n519, n387, n649, n572);
or   g1216 (n1282, n579, n473, n620, n551);
nor  g1217 (n1303, n478, n520, n291, n412);
xor  g1218 (n904, n584, n619, n205, n643);
xor  g1219 (n848, n331, n358, n414, n596);
or   g1220 (n1258, n335, n548, n463, n493);
xnor g1221 (n1206, n350, n267, n394, n295);
and  g1222 (n1199, n306, n505, n661, n461);
xor  g1223 (n1225, n399, n449, n207, n580);
nand g1224 (n1072, n477, n658, n274, n514);
xor  g1225 (n892, n196, n274, n208, n578);
nor  g1226 (n1177, n456, n519, n273, n479);
nor  g1227 (n935, n366, n599, n289, n362);
nand g1228 (n1196, n273, n635, n650, n663);
or   g1229 (n982, n554, n394, n489, n441);
nor  g1230 (n819, n369, n345, n275, n228);
xor  g1231 (n1020, n240, n581, n410, n645);
xor  g1232 (n963, n501, n325, n404, n277);
xor  g1233 (n974, n591, n505, n585, n468);
nor  g1234 (n690, n368, n286, n615, n323);
and  g1235 (n814, n630, n534, n199, n484);
xor  g1236 (n973, n277, n595, n353, n378);
nand g1237 (n1304, n301, n240, n609, n575);
and  g1238 (n946, n562, n462, n219, n388);
nor  g1239 (n783, n520, n469, n300, n655);
xor  g1240 (n1214, n488, n293, n365, n484);
or   g1241 (n925, n649, n559, n460, n490);
nand g1242 (n1008, n263, n632, n391, n446);
xnor g1243 (n874, n408, n442, n434, n328);
xor  g1244 (n688, n340, n509, n624, n482);
nor  g1245 (n1064, n296, n254, n285, n202);
nor  g1246 (n1105, n411, n361, n629, n281);
or   g1247 (n1297, n555, n644, n392, n518);
and  g1248 (n1261, n511, n204, n553, n582);
xor  g1249 (n895, n230, n561, n618, n554);
xor  g1250 (n1030, n299, n485, n247, n310);
and  g1251 (n808, n655, n486, n605, n344);
xor  g1252 (n1092, n277, n297, n517, n511);
nor  g1253 (n944, n424, n595, n336, n438);
and  g1254 (n875, n512, n579, n330, n633);
nor  g1255 (n1218, n204, n623, n627, n426);
and  g1256 (n764, n556, n323, n317, n247);
nand g1257 (n1246, n367, n351, n611, n447);
xnor g1258 (n1060, n558, n426, n540, n454);
nand g1259 (n1001, n434, n652, n624, n233);
and  g1260 (n729, n499, n255, n291, n317);
and  g1261 (n1222, n611, n320, n415, n199);
nand g1262 (n682, n370, n491, n612, n380);
nand g1263 (n905, n256, n550, n243, n506);
xor  g1264 (n675, n343, n230, n289, n411);
xnor g1265 (n1181, n588, n546, n364, n518);
nor  g1266 (n1059, n656, n624, n224, n418);
and  g1267 (n746, n345, n254, n531, n653);
nand g1268 (n1194, n588, n321, n510, n569);
and  g1269 (n1213, n667, n397, n505, n213);
nand g1270 (n993, n569, n550, n517, n271);
nand g1271 (n919, n609, n610, n400, n630);
xnor g1272 (n1250, n261, n607, n613, n206);
or   g1273 (n739, n333, n583, n261, n586);
nand g1274 (n1387, n1035, n1008, n889, n851);
and  g1275 (n1321, n908, n676, n1144, n1190);
or   g1276 (n1360, n795, n785, n801, n1033);
nand g1277 (n1423, n1101, n996, n997, n1169);
and  g1278 (n1372, n727, n780, n1106, n781);
xor  g1279 (n1431, n755, n1052, n933, n1181);
xor  g1280 (n1370, n721, n811, n765, n715);
nor  g1281 (n1369, n698, n834, n748, n965);
nor  g1282 (n1402, n1125, n799, n1166, n1150);
nor  g1283 (n1361, n978, n1107, n722, n754);
or   g1284 (n1343, n1063, n905, n1177, n869);
nand g1285 (n1324, n890, n1149, n880, n803);
nand g1286 (n1359, n1090, n903, n1045, n995);
xor  g1287 (n1331, n981, n777, n720, n1104);
and  g1288 (n1334, n974, n1119, n952, n861);
xor  g1289 (n1325, n929, n1178, n1188, n967);
nand g1290 (n1404, n953, n912, n973, n787);
or   g1291 (n1437, n977, n1088, n691, n984);
or   g1292 (n1337, n1124, n959, n1185, n1162);
or   g1293 (n1385, n769, n1015, n1157, n809);
xnor g1294 (n1340, n700, n876, n778, n786);
xor  g1295 (n1384, n1198, n773, n1002, n800);
or   g1296 (n1418, n897, n838, n1103, n1203);
xnor g1297 (n1414, n979, n687, n1174, n716);
or   g1298 (n1347, n1086, n839, n1018, n1006);
nor  g1299 (n1427, n775, n848, n1175, n833);
and  g1300 (n1394, n919, n1095, n988, n759);
and  g1301 (n1438, n1154, n925, n793, n751);
and  g1302 (n1326, n1102, n852, n1099, n990);
or   g1303 (n1401, n961, n744, n1130, n1011);
and  g1304 (n1426, n900, n766, n746, n872);
or   g1305 (n1390, n709, n918, n1205, n937);
nand g1306 (n1311, n854, n936, n960, n914);
nor  g1307 (n1417, n1009, n1065, n899, n845);
xnor g1308 (n1318, n949, n1056, n913, n926);
xnor g1309 (n1429, n1025, n1084, n734, n843);
nor  g1310 (n1351, n1014, n794, n837, n817);
or   g1311 (n1395, n946, n901, n878, n1127);
xor  g1312 (n1408, n1078, n868, n860, n823);
and  g1313 (n1368, n761, n699, n1165, n1044);
nor  g1314 (n1333, n1028, n694, n808, n742);
xnor g1315 (n1435, n948, n877, n713, n920);
and  g1316 (n1422, n1022, n941, n1168, n1030);
xor  g1317 (n1355, n940, n688, n681, n1024);
nand g1318 (n1350, n1046, n782, n832, n856);
and  g1319 (n1400, n1121, n1069, n682, n1191);
nand g1320 (n1354, n1094, n745, n1032, n791);
xnor g1321 (n1389, n1019, n911, n675, n693);
and  g1322 (n1412, n760, n772, n1079, n1055);
xnor g1323 (n1439, n1036, n708, n707, n870);
and  g1324 (n1348, n1195, n1058, n1005, n942);
and  g1325 (n1339, n1096, n1135, n1012, n1139);
xor  g1326 (n1344, n1070, n739, n1117, n726);
nand g1327 (n1425, n762, n714, n1161, n1097);
nand g1328 (n1378, n1176, n1129, n1179, n767);
xor  g1329 (n1397, n1192, n758, n821, n686);
nor  g1330 (n1317, n874, n1141, n1077, n902);
xnor g1331 (n1399, n898, n969, n1193, n805);
nor  g1332 (n1428, n887, n1093, n1082, n704);
xnor g1333 (n1380, n1145, n958, n830, n1120);
nand g1334 (n1433, n740, n999, n696, n951);
or   g1335 (n1379, n944, n964, n807, n1039);
and  g1336 (n1349, n1142, n1118, n883, n757);
xnor g1337 (n1329, n1110, n895, n1187, n894);
and  g1338 (n1430, n994, n1051, n678, n1076);
nand g1339 (n1403, n982, n975, n692, n892);
nor  g1340 (n1320, n886, n683, n989, n1038);
nor  g1341 (n1367, n1074, n737, n863, n966);
nand g1342 (n1406, n1001, n1000, n1137, n827);
and  g1343 (n1352, n888, n1010, n702, n935);
nor  g1344 (n1328, n1172, n1072, n1043, n1153);
nand g1345 (n1420, n938, n836, n1048, n743);
nor  g1346 (n1377, n738, n904, n906, n1171);
xnor g1347 (n1407, n1136, n840, n701, n1059);
and  g1348 (n1312, n985, n1004, n1021, n814);
or   g1349 (n1313, n689, n828, n1003, n818);
nand g1350 (n1410, n865, n790, n789, n1123);
nand g1351 (n1436, n1204, n1112, n719, n1116);
xnor g1352 (n1373, n695, n1156, n764, n1049);
or   g1353 (n1366, n857, n813, n1054, n932);
nand g1354 (n1323, n1023, n939, n806, n690);
nand g1355 (n1388, n1183, n879, n776, n1068);
and  g1356 (n1382, n835, n788, n991, n1133);
xnor g1357 (n1332, n752, n712, n1199, n923);
xnor g1358 (n1358, n674, n1131, n916, n1189);
and  g1359 (n1346, n822, n1031, n1053, n749);
nor  g1360 (n1357, n987, n921, n1075, n680);
xnor g1361 (n1413, n1115, n797, n1186, n972);
xnor g1362 (n1322, n1138, n980, n1151, n1085);
nor  g1363 (n1335, n779, n710, n774, n1066);
or   g1364 (n1396, n1146, n1060, n677, n829);
nand g1365 (n1307, n1184, n1197, n810, n1122);
or   g1366 (n1381, n1167, n1170, n842, n763);
and  g1367 (n1386, n1100, n697, n873, n1108);
nor  g1368 (n1336, n922, n907, n893, n846);
nor  g1369 (n1375, n957, n1113, n867, n986);
xor  g1370 (n1392, n1109, n825, n705, n849);
xnor g1371 (n1393, n1182, n1062, n956, n1041);
or   g1372 (n1341, n1147, n1134, n924, n768);
and  g1373 (n1308, n750, n819, n1201, n882);
nor  g1374 (n1416, n753, n1020, n816, n862);
nand g1375 (n1314, n1126, n1037, n812, n934);
or   g1376 (n1310, n1029, n1026, n1180, n864);
or   g1377 (n1316, n844, n1089, n1061, n1111);
or   g1378 (n1365, n747, n885, n976, n815);
or   g1379 (n1345, n729, n1105, n733, n1158);
nor  g1380 (n1371, n1091, n928, n1027, n1071);
nand g1381 (n1424, n1160, n855, n728, n1114);
xnor g1382 (n1309, n820, n871, n968, n1163);
xor  g1383 (n1376, n884, n947, n826, n943);
nor  g1384 (n1364, n998, n684, n1057, n756);
or   g1385 (n1432, n804, n917, n910, n1098);
and  g1386 (n1391, n770, n1047, n1007, n792);
nor  g1387 (n1315, n927, n1132, n1155, n1140);
nand g1388 (n1419, n703, n711, n881, n824);
and  g1389 (n1353, n741, n679, n1128, n718);
nor  g1390 (n1330, n1196, n1092, n1200, n963);
xnor g1391 (n1374, n970, n850, n1159, n1202);
nand g1392 (n1434, n1016, n1017, n930, n1081);
xor  g1393 (n1319, n841, n796, n993, n802);
nor  g1394 (n1383, n866, n847, n706, n1067);
xor  g1395 (n1421, n771, n945, n1173, n1073);
and  g1396 (n1363, n1064, n950, n915, n831);
or   g1397 (n1398, n955, n723, n731, n1083);
or   g1398 (n1405, n962, n1042, n730, n732);
xor  g1399 (n1362, n859, n1087, n725, n1148);
xnor g1400 (n1411, n853, n1040, n1164, n1080);
nor  g1401 (n1415, n784, n798, n1013, n1034);
and  g1402 (n1356, n992, n875, n1152, n896);
or   g1403 (n1342, n736, n954, n983, n891);
nor  g1404 (n1327, n783, n717, n858, n1050);
nand g1405 (n1409, n1194, n931, n685, n1143);
xnor g1406 (n1338, n735, n724, n909, n971);
not  g1407 (n1445, n1316);
not  g1408 (n1450, n1313);
buf  g1409 (n1448, n1318);
buf  g1410 (n1453, n1315);
buf  g1411 (n1447, n1321);
buf  g1412 (n1454, n1314);
not  g1413 (n1441, n1319);
buf  g1414 (n1452, n1312);
buf  g1415 (n1451, n1320);
buf  g1416 (n1449, n1317);
buf  g1417 (n1440, n1309);
buf  g1418 (n1442, n1323);
not  g1419 (n1443, n1310);
not  g1420 (n1455, n1311);
buf  g1421 (n1446, n1322);
buf  g1422 (n1444, n1324);
nand g1423 (n1457, n1446, n1252, n1275, n1229);
nand g1424 (n1472, n1227, n1254, n1286, n1277);
or   g1425 (n1465, n1239, n1238, n1220, n1206);
nor  g1426 (n1470, n1283, n1442, n1251, n1273);
and  g1427 (n1474, n1233, n1221, n1266, n1215);
or   g1428 (n1466, n1207, n1228, n1237, n1281);
or   g1429 (n1456, n1257, n1282, n1443, n1211);
xor  g1430 (n1461, n1270, n1224, n1263, n1267);
xor  g1431 (n1478, n1440, n1249, n1250, n1242);
xnor g1432 (n1476, n1441, n1280, n1446, n1271);
xnor g1433 (n1460, n1272, n1231, n1285, n1265);
or   g1434 (n1480, n1258, n1261, n1244, n1445);
or   g1435 (n1481, n1274, n1218, n1222, n1278);
nand g1436 (n1458, n1216, n1245, n1225, n1284);
nor  g1437 (n1469, n1443, n1441, n1241, n1243);
nor  g1438 (n1464, n1445, n1441, n1255, n1259);
nand g1439 (n1479, n1269, n1445, n1276, n1444);
nand g1440 (n1473, n1219, n1440, n1208, n1246);
nand g1441 (n1462, n1446, n1232, n1440, n1230);
and  g1442 (n1463, n1444, n1442, n1235, n1264);
and  g1443 (n1477, n1226, n1268, n1240, n1223);
or   g1444 (n1468, n1279, n1442, n1213, n1253);
xor  g1445 (n1471, n1210, n1444, n1445, n1256);
and  g1446 (n1475, n1443, n1442, n1236, n1247);
xnor g1447 (n1459, n1443, n1262, n1212, n1217);
nand g1448 (n1482, n1214, n1444, n1440, n1209);
xor  g1449 (n1467, n1260, n1248, n1234, n1441);
and  g1450 (n1485, n1381, n1458, n1379, n1386);
xnor g1451 (n1510, n1392, n1341, n1367, n1345);
nand g1452 (n1488, n1359, n1460, n1344, n1374);
xor  g1453 (n1509, n1457, n1399, n1372, n1401);
xor  g1454 (n1508, n1460, n1395, n1360, n1380);
or   g1455 (n1489, n1403, n1327, n1349, n1456);
xnor g1456 (n1506, n1394, n1456, n1350, n1337);
nor  g1457 (n1492, n1370, n1414, n1354, n1463);
or   g1458 (n1486, n1365, n1389, n1364, n1405);
xnor g1459 (n1496, n1413, n1407, n1368, n1366);
nand g1460 (n1505, n1390, n1397, n1460, n1457);
nor  g1461 (n1512, n1362, n1339, n1459, n1461);
and  g1462 (n1497, n1373, n1347, n1356, n1334);
nand g1463 (n1495, n1343, n1363, n1329, n1353);
nand g1464 (n1483, n1402, n1382, n1383, n1378);
or   g1465 (n1498, n1459, n1338, n1351, n1461);
xnor g1466 (n1511, n1461, n1336, n1400, n1462);
nor  g1467 (n1491, n1328, n1342, n1325, n1398);
xnor g1468 (n1494, n1369, n1457, n1375, n1396);
or   g1469 (n1504, n1459, n1332, n1411, n1333);
and  g1470 (n1502, n1461, n1387, n1404, n1410);
and  g1471 (n1493, n1409, n1412, n1456, n1331);
and  g1472 (n1500, n1458, n1330, n1335, n1462);
and  g1473 (n1503, n1459, n1376, n1361, n1348);
xnor g1474 (n1501, n1457, n1458, n1391, n1326);
xor  g1475 (n1490, n1355, n1460, n1358, n1340);
nor  g1476 (n1507, n1352, n1357, n1377, n1384);
and  g1477 (n1487, n1462, n1458, n1463, n1456);
xor  g1478 (n1484, n1385, n1393, n1346, n1371);
xor  g1479 (n1499, n1408, n1388, n1462, n1406);
not  g1480 (n1552, n192);
not  g1481 (n1527, n11);
not  g1482 (n1526, n190);
buf  g1483 (n1531, n1464);
nor  g1484 (n1548, n1486, n1455);
and  g1485 (n1513, n1506, n1451, n1511, n193);
xnor g1486 (n1514, n1295, n1448, n1511, n1505);
and  g1487 (n1539, n668, n1449, n193, n1464);
and  g1488 (n1550, n1501, n1466, n1465, n1447);
or   g1489 (n1537, n1484, n1508, n1453, n1507);
nor  g1490 (n1542, n1450, n1503, n1485, n1449);
or   g1491 (n1524, n1512, n1292, n1450, n1509);
xnor g1492 (n1547, n191, n1448, n1453, n1492);
nor  g1493 (n1519, n1491, n1504, n1502, n1510);
nor  g1494 (n1518, n64, n11, n1490, n1448);
nor  g1495 (n1515, n1466, n668, n10, n1287);
xor  g1496 (n1535, n1487, n668, n10, n1504);
xor  g1497 (n1525, n1464, n669, n1512, n1415);
nand g1498 (n1534, n190, n1483, n1464, n1451);
and  g1499 (n1520, n192, n190, n669, n189);
xnor g1500 (n1540, n11, n65, n1465, n189);
xnor g1501 (n1541, n64, n191, n1453, n1455);
nand g1502 (n1532, n191, n1454, n1499, n1505);
xnor g1503 (n1538, n1450, n1495, n1289, n1452);
or   g1504 (n1529, n1455, n192, n11, n1497);
nor  g1505 (n1536, n10, n1452, n1489, n1291);
or   g1506 (n1528, n1510, n1509, n1508, n1452);
and  g1507 (n1543, n1447, n1500, n1506, n1296);
nand g1508 (n1517, n1496, n1290, n12, n1455);
and  g1509 (n1533, n65, n189, n1449, n1507);
nand g1510 (n1549, n1493, n1299, n1463, n1450);
nor  g1511 (n1551, n1297, n1298, n1453, n1498);
xor  g1512 (n1523, n669, n1463, n1451, n1300);
or   g1513 (n1516, n1301, n1454, n1446, n1447);
xnor g1514 (n1546, n1452, n1503, n10, n1449);
or   g1515 (n1545, n64, n1293, n1288, n1465);
or   g1516 (n1522, n189, n1451, n1302, n191);
or   g1517 (n1521, n1465, n1454, n1294, n65);
xor  g1518 (n1544, n192, n1494, n190, n1488);
nand g1519 (n1530, n65, n1447, n1454, n1448);
buf  g1520 (n1575, n1547);
buf  g1521 (n1665, n1537);
not  g1522 (n1708, n1548);
buf  g1523 (n1693, n1527);
buf  g1524 (n1650, n30);
not  g1525 (n1689, n1540);
buf  g1526 (n1660, n17);
buf  g1527 (n1561, n1551);
buf  g1528 (n1656, n1469);
buf  g1529 (n1620, n1536);
not  g1530 (n1574, n1470);
not  g1531 (n1572, n29);
buf  g1532 (n1566, n21);
not  g1533 (n1648, n1524);
buf  g1534 (n1638, n22);
buf  g1535 (n1647, n1478);
buf  g1536 (n1663, n1478);
not  g1537 (n1707, n1532);
not  g1538 (n1587, n1479);
not  g1539 (n1674, n1516);
buf  g1540 (n1629, n31);
not  g1541 (n1664, n19);
not  g1542 (n1591, n1541);
buf  g1543 (n1560, n28);
buf  g1544 (n1642, n32);
buf  g1545 (n1576, n24);
not  g1546 (n1617, n1514);
buf  g1547 (n1643, n1524);
not  g1548 (n1634, n1467);
buf  g1549 (n1652, n1542);
buf  g1550 (n1627, n1547);
buf  g1551 (n1631, n1523);
not  g1552 (n1635, n1470);
buf  g1553 (n1659, n1531);
buf  g1554 (n1622, n25);
buf  g1555 (n1555, n1538);
not  g1556 (n1646, n1475);
buf  g1557 (n1700, n16);
buf  g1558 (n1640, n21);
buf  g1559 (n1625, n1517);
buf  g1560 (n1563, n31);
buf  g1561 (n1711, n14);
not  g1562 (n1583, n1518);
buf  g1563 (n1600, n1548);
not  g1564 (n1585, n1544);
buf  g1565 (n1614, n22);
not  g1566 (n1559, n1518);
buf  g1567 (n1691, n16);
buf  g1568 (n1655, n19);
buf  g1569 (n1662, n1543);
buf  g1570 (n1606, n28);
not  g1571 (n1694, n1477);
buf  g1572 (n1666, n20);
buf  g1573 (n1658, n1546);
not  g1574 (n1599, n1530);
buf  g1575 (n1564, n29);
buf  g1576 (n1688, n1526);
buf  g1577 (n1567, n17);
buf  g1578 (n1613, n30);
buf  g1579 (n1710, n1517);
not  g1580 (n1675, n1477);
buf  g1581 (n1582, n1530);
buf  g1582 (n1651, n1473);
buf  g1583 (n1624, n1480);
buf  g1584 (n1702, n24);
buf  g1585 (n1667, n1474);
buf  g1586 (n1712, n1546);
not  g1587 (n1696, n26);
buf  g1588 (n1657, n1468);
buf  g1589 (n1578, n1538);
not  g1590 (n1581, n1548);
buf  g1591 (n1679, n66);
buf  g1592 (n1593, n1532);
not  g1593 (n1568, n1471);
buf  g1594 (n1597, n1533);
buf  g1595 (n1706, n32);
buf  g1596 (n1616, n22);
buf  g1597 (n1698, n26);
buf  g1598 (n1697, n1479);
buf  g1599 (n1601, n15);
not  g1600 (n1681, n1541);
buf  g1601 (n1586, n18);
not  g1602 (n1579, n1547);
buf  g1603 (n1569, n1515);
buf  g1604 (n1670, n1552);
not  g1605 (n1612, n1521);
buf  g1606 (n1703, n1519);
not  g1607 (n1577, n15);
not  g1608 (n1595, n12);
buf  g1609 (n1628, n1536);
not  g1610 (n1654, n1530);
not  g1611 (n1603, n1531);
not  g1612 (n1641, n29);
buf  g1613 (n1686, n1516);
not  g1614 (n1678, n19);
not  g1615 (n1623, n1531);
buf  g1616 (n1604, n1468);
buf  g1617 (n1699, n27);
not  g1618 (n1690, n1533);
not  g1619 (n1671, n1544);
buf  g1620 (n1571, n1537);
buf  g1621 (n1639, n13);
not  g1622 (n1632, n1551);
not  g1623 (n1589, n14);
not  g1624 (n1645, n1525);
buf  g1625 (n1615, n66);
not  g1626 (n1621, n1466);
buf  g1627 (n1683, n1480);
nand g1628 (n1704, n1552, n1546, n1472, n1521);
xnor g1629 (n1562, n1552, n1544, n1533, n1479);
or   g1630 (n1669, n1532, n1476, n1536, n67);
and  g1631 (n1598, n1545, n1531, n1539, n1520);
nand g1632 (n1556, n26, n1532, n1467, n1471);
xor  g1633 (n1580, n30, n20, n32, n67);
xor  g1634 (n1676, n1528, n23, n1539, n1517);
xor  g1635 (n1611, n1515, n1518, n1539, n1523);
xnor g1636 (n1653, n1551, n18, n1524, n1545);
nand g1637 (n1588, n1545, n31, n1549, n1473);
xor  g1638 (n1677, n1470, n1480, n1529);
nor  g1639 (n1705, n1520, n1475, n1473, n1469);
xnor g1640 (n1610, n1545, n21, n14, n25);
nor  g1641 (n1633, n1481, n1514, n1542, n1534);
and  g1642 (n1672, n17, n15, n1550, n1538);
or   g1643 (n1685, n1477, n1526, n1533, n13);
nand g1644 (n1609, n24, n1514, n1544, n18);
or   g1645 (n1668, n23, n1528, n1540, n1542);
xnor g1646 (n1626, n1551, n18, n1539, n29);
and  g1647 (n1590, n1467, n1522, n1473, n24);
xnor g1648 (n1558, n1472, n15, n1524, n1482);
or   g1649 (n1673, n1518, n19, n1482, n1535);
or   g1650 (n1630, n1527, n1534, n23, n1535);
and  g1651 (n1554, n1550, n1543, n1481, n16);
xor  g1652 (n1602, n66, n1474, n1513, n1476);
nor  g1653 (n1584, n1550, n1528, n1516, n25);
xor  g1654 (n1637, n1535, n66, n1475, n1478);
xor  g1655 (n1573, n1467, n1536, n1519, n1475);
nand g1656 (n1644, n1519, n1530, n25, n1549);
xor  g1657 (n1687, n1468, n28, n1534, n1472);
and  g1658 (n1594, n17, n1529, n1522, n1474);
or   g1659 (n1684, n1525, n1478, n1481, n1482);
xnor g1660 (n1619, n1547, n1543, n1529, n1542);
nor  g1661 (n1709, n1525, n1527, n1481, n1482);
nand g1662 (n1701, n1538, n1521, n1517, n1468);
nor  g1663 (n1636, n1522, n1540, n1476, n1477);
xor  g1664 (n1553, n1516, n1541, n1469, n1550);
xnor g1665 (n1557, n30, n1525, n1527, n1546);
and  g1666 (n1592, n1523, n21, n20, n1549);
xor  g1667 (n1695, n20, n1526, n1537, n1471);
nand g1668 (n1692, n22, n1552, n26, n1540);
and  g1669 (n1570, n32, n27, n1522, n1479);
nor  g1670 (n1596, n1466, n1470, n1515, n14);
or   g1671 (n1565, n31, n1513, n12, n1514);
nand g1672 (n1607, n1521, n1474, n1513, n28);
nor  g1673 (n1682, n1534, n1471, n1537, n27);
and  g1674 (n1680, n16, n13, n1513, n1476);
nor  g1675 (n1605, n1549, n13, n1520);
nor  g1676 (n1608, n1469, n23, n1526, n1528);
or   g1677 (n1661, n12, n1523, n1472, n1543);
and  g1678 (n1649, n27, n1548, n67, n1519);
xor  g1679 (n1618, n1529, n1541, n1535, n1515);
xor  g1680 (n1771, n1622, n1575, n1557, n1612);
and  g1681 (n1756, n1579, n1670, n1583, n1573);
xor  g1682 (n1774, n1644, n1665, n1566, n1652);
nor  g1683 (n1777, n1554, n1631, n1582, n1651);
or   g1684 (n1744, n1627, n1576, n1560, n1618);
xor  g1685 (n1793, n1602, n1632, n1585, n1665);
xor  g1686 (n1788, n1599, n1646, n1615, n1604);
nor  g1687 (n1729, n1573, n1632, n1584, n1628);
nand g1688 (n1751, n1559, n1658, n1617, n1645);
nand g1689 (n1769, n1603, n1625, n1650, n1651);
nand g1690 (n1736, n1568, n1568, n1604, n1605);
and  g1691 (n1734, n1635, n1647, n1667, n1596);
xnor g1692 (n1783, n1662, n1584, n1620, n1646);
and  g1693 (n1801, n1628, n1594, n1635, n1571);
and  g1694 (n1779, n1588, n1648, n1611, n1612);
xor  g1695 (n1721, n1610, n1661, n1567, n1657);
nor  g1696 (n1764, n1609, n1577, n1660, n1644);
xnor g1697 (n1730, n1594, n1663, n1646, n1658);
xor  g1698 (n1775, n1616, n1663, n1654, n1664);
nand g1699 (n1767, n1672, n1648, n1624, n1615);
and  g1700 (n1718, n1594, n1607, n1591, n1569);
xnor g1701 (n1761, n1636, n1624, n1625, n1607);
nor  g1702 (n1713, n1655, n1558, n1587, n1610);
xor  g1703 (n1726, n1622, n1640, n1645, n1653);
nor  g1704 (n1762, n1555, n1634, n1581, n1606);
and  g1705 (n1765, n1622, n1603, n1633, n1627);
xor  g1706 (n1768, n1644, n1611, n1629, n1660);
xnor g1707 (n1731, n1586, n1617, n1565, n1663);
xor  g1708 (n1716, n1565, n1563, n1557, n1609);
nand g1709 (n1732, n1561, n1655, n1595, n1562);
nand g1710 (n1720, n1592, n1595, n1580);
xor  g1711 (n1778, n1566, n1574, n1596, n1632);
xnor g1712 (n1727, n1563, n1619, n1581, n1659);
nor  g1713 (n1766, n1613, n1553, n1592, n1669);
and  g1714 (n1750, n1607, n1558, n1591, n1608);
nand g1715 (n1745, n1601, n1627, n1617, n1609);
nand g1716 (n1757, n1567, n1588, n1579, n1666);
xor  g1717 (n1780, n1561, n1642, n1569, n1611);
xor  g1718 (n1752, n1571, n1637, n1642, n1640);
nor  g1719 (n1743, n1643, n1621, n1638, n1624);
nor  g1720 (n1795, n1638, n1621, n1595, n1648);
nor  g1721 (n1776, n1600, n1568, n1564, n1639);
nor  g1722 (n1738, n1571, n1623, n1638, n1588);
xor  g1723 (n1749, n1572, n1625, n1652, n1618);
and  g1724 (n1737, n1605, n1585, n1637, n1657);
xor  g1725 (n1794, n1560, n1664, n1599, n1575);
xor  g1726 (n1799, n1559, n1596, n1634, n1572);
or   g1727 (n1770, n1629, n1641, n1586, n1667);
and  g1728 (n1787, n1654, n1650, n1626, n1583);
and  g1729 (n1785, n1601, n1649, n1598, n1615);
nand g1730 (n1758, n1660, n1554, n1636, n1572);
xor  g1731 (n1733, n1656, n1556, n1619, n1672);
xnor g1732 (n1724, n1619, n1658, n1579, n1636);
nor  g1733 (n1763, n1661, n1593, n1567, n1604);
and  g1734 (n1796, n1612, n1671, n1647, n1645);
and  g1735 (n1791, n1601, n1643, n1562, n1578);
nand g1736 (n1797, n1587, n1582, n1635, n1637);
xor  g1737 (n1754, n1664, n1651, n1653, n1643);
nand g1738 (n1717, n1600, n1672, n1606, n1613);
nand g1739 (n1782, n1583, n1661, n1671, n1564);
nor  g1740 (n1781, n1620, n1593, n1614, n1566);
xor  g1741 (n1798, n1621, n1563, n1591, n1598);
xnor g1742 (n1740, n1662, n1629, n1597, n1577);
nand g1743 (n1728, n1650, n1616, n1633, n1555);
nand g1744 (n1725, n1593, n1578, n1597, n1576);
or   g1745 (n1715, n1630, n1641, n1589, n1631);
or   g1746 (n1735, n1580, n1590, n1608, n1570);
xnor g1747 (n1748, n1589, n1565, n1630, n1639);
nand g1748 (n1747, n1559, n1561, n1556, n1655);
xnor g1749 (n1786, n1669, n1574, n1626, n1647);
xnor g1750 (n1784, n1603, n1659, n1640, n1558);
xor  g1751 (n1742, n1641, n1631, n1628, n1575);
or   g1752 (n1746, n1560, n1584, n1614, n1618);
nor  g1753 (n1790, n1573, n1670, n1639, n1582);
xnor g1754 (n1739, n1620, n1668, n1666, n1587);
nor  g1755 (n1741, n1614, n1562, n1574, n1606);
and  g1756 (n1792, n1585, n1557, n1608, n1570);
or   g1757 (n1772, n1553, n1667, n1605, n1626);
xor  g1758 (n1800, n1576, n1581, n1592, n1671);
and  g1759 (n1753, n1666, n1654, n1564, n1590);
or   g1760 (n1789, n1669, n1623, n1613, n1662);
nor  g1761 (n1723, n1586, n1656, n1602, n1642);
nand g1762 (n1714, n1649, n1599, n1590, n1623);
nand g1763 (n1719, n1656, n1630, n1602, n1600);
nor  g1764 (n1755, n1668, n1653, n1649, n1652);
xor  g1765 (n1722, n1589, n1665, n1657, n1578);
xor  g1766 (n1759, n1616, n1633, n1577, n1570);
nor  g1767 (n1773, n1668, n1569, n1670, n1634);
nor  g1768 (n1760, n1597, n1610, n1598, n1659);
buf  g1769 (n1803, n1722);
buf  g1770 (n1804, n1720);
not  g1771 (n1807, n1724);
buf  g1772 (n1806, n1713);
and  g1773 (n1802, n1717, n1723, n1714, n1721);
and  g1774 (n1805, n1715, n1718, n1719, n1716);
not  g1775 (n1819, n1804);
buf  g1776 (n1810, n1804);
buf  g1777 (n1812, n1805);
not  g1778 (n1809, n1802);
buf  g1779 (n1818, n1803);
not  g1780 (n1808, n1804);
not  g1781 (n1814, n1806);
not  g1782 (n1811, n1805);
buf  g1783 (n1813, n1803);
not  g1784 (n1815, n1803);
not  g1785 (n1817, n1805);
not  g1786 (n1816, n1802);
not  g1787 (n1821, n1808);
not  g1788 (n1822, n1809);
not  g1789 (n1823, n1303);
not  g1790 (n1825, n1808);
buf  g1791 (n1820, n1809);
not  g1792 (n1826, n1808);
xnor g1793 (n1824, n1809, n1808);
buf  g1794 (n1831, n1822);
buf  g1795 (n1835, n1823);
buf  g1796 (n1841, n1821);
buf  g1797 (n1827, n1826);
buf  g1798 (n1844, n1824);
not  g1799 (n1850, n1825);
buf  g1800 (n1853, n1821);
buf  g1801 (n1854, n1821);
buf  g1802 (n1834, n1823);
buf  g1803 (n1840, n1825);
not  g1804 (n1838, n1826);
not  g1805 (n1832, n1820);
not  g1806 (n1836, n1825);
not  g1807 (n1846, n1820);
buf  g1808 (n1848, n1824);
not  g1809 (n1845, n1825);
not  g1810 (n1852, n1824);
buf  g1811 (n1830, n1822);
not  g1812 (n1839, n1822);
not  g1813 (n1833, n1820);
buf  g1814 (n1829, n1826);
buf  g1815 (n1837, n1823);
buf  g1816 (n1842, n1822);
buf  g1817 (n1849, n1823);
buf  g1818 (n1847, n1821);
buf  g1819 (n1828, n1826);
buf  g1820 (n1851, n1820);
buf  g1821 (n1843, n1824);
not  g1822 (n1869, n1833);
xnor g1823 (n1855, n1846, n1828, n1833);
and  g1824 (n1882, n1813, n1844, n1838, n1819);
and  g1825 (n1871, n1819, n1846, n1831, n1827);
or   g1826 (n1865, n1833, n1840, n1416);
and  g1827 (n1868, n1829, n1814, n1815, n1843);
and  g1828 (n1877, n1827, n1839, n1818, n1842);
nor  g1829 (n1883, n1839, n1845, n1848, n1838);
or   g1830 (n1890, n1832, n1819, n1818, n1834);
and  g1831 (n1864, n1811, n1851, n1849, n1847);
and  g1832 (n1875, n1815, n1838, n1850, n1837);
xnor g1833 (n1862, n1835, n1842, n1844, n1839);
nor  g1834 (n1873, n1846, n1840, n1816, n1837);
nand g1835 (n1879, n1813, n1811, n1827, n1836);
xnor g1836 (n1874, n1847, n1849, n1836);
nand g1837 (n1866, n1811, n1850, n1831, n1817);
xor  g1838 (n1861, n1835, n1841, n1814, n1817);
xnor g1839 (n1867, n1814, n1818, n1417, n1816);
nand g1840 (n1888, n1830, n1816, n1829);
and  g1841 (n1857, n1848, n1813, n1837, n1845);
xnor g1842 (n1859, n1841, n1843, n1847, n1832);
xnor g1843 (n1884, n1831, n1810, n1818, n1834);
and  g1844 (n1886, n1848, n1830, n1833, n1840);
xnor g1845 (n1872, n1842, n1814, n1810, n1831);
xnor g1846 (n1860, n1809, n1827, n1836, n1835);
or   g1847 (n1870, n1845, n1830, n1841, n1811);
nor  g1848 (n1881, n1850, n1842, n1832, n1836);
nand g1849 (n1887, n1830, n1816, n1817);
xnor g1850 (n1863, n1844, n1848, n1812, n1834);
or   g1851 (n1889, n1829, n1847, n1843, n1810);
or   g1852 (n1876, n1828, n1835, n1844, n1841);
and  g1853 (n1858, n1834, n1812, n1837);
or   g1854 (n1878, n1810, n1812, n1849, n1828);
or   g1855 (n1856, n1828, n1815, n1819, n1845);
xnor g1856 (n1885, n1846, n1839, n1843, n1850);
nand g1857 (n1880, n1832, n1813, n1838, n1815);
not  g1858 (n1894, n1856);
buf  g1859 (n1892, n1858);
buf  g1860 (n1893, n1855);
not  g1861 (n1891, n1857);
and  g1862 (n1902, n671, n1853, n1428, n670);
xor  g1863 (n1898, n672, n1894, n1893, n1432);
and  g1864 (n1905, n1851, n1854, n1427, n1433);
xnor g1865 (n1904, n1854, n1892, n1851, n1421);
nand g1866 (n1907, n1853, n1893, n1422);
xnor g1867 (n1895, n673, n1425, n1853, n670);
and  g1868 (n1909, n672, n1424, n1891, n1852);
xnor g1869 (n1901, n1420, n670, n1431, n1852);
or   g1870 (n1903, n1304, n1853, n1419, n1418);
nor  g1871 (n1908, n1893, n1891, n1434);
xor  g1872 (n1910, n669, n1852, n672, n1429);
xnor g1873 (n1896, n671, n1852, n1854, n672);
xor  g1874 (n1897, n1894, n673, n1891, n1423);
xor  g1875 (n1900, n1894, n1426, n671, n1854);
or   g1876 (n1899, n670, n1892, n1894);
nand g1877 (n1906, n1851, n671, n1892, n1430);
nor  g1878 (n1919, n68, n1910, n1906);
xnor g1879 (n1918, n1437, n1861, n1869);
nor  g1880 (n1923, n1435, n1863, n1884);
and  g1881 (n1922, n1905, n1910, n1867);
and  g1882 (n1913, n1874, n1877, n1909);
nor  g1883 (n1926, n1864, n1900, n1885);
nor  g1884 (n1927, n1876, n1865, n1887);
nor  g1885 (n1921, n1872, n1878, n1883);
xnor g1886 (n1912, n1860, n1908, n68);
nand g1887 (n1924, n1890, n193, n68);
xor  g1888 (n1925, n1898, n1880, n1895);
or   g1889 (n1929, n1907, n1899, n1889);
and  g1890 (n1914, n1902, n1908, n1868);
xnor g1891 (n1915, n1866, n1879, n1862);
and  g1892 (n1917, n1901, n1909, n1439);
xnor g1893 (n1911, n1896, n1897, n1859);
nor  g1894 (n1928, n1873, n1903, n1875, n1882);
xnor g1895 (n1916, n1871, n1886, n1870, n67);
xor  g1896 (n1920, n193, n68, n1888, n1438);
nor  g1897 (n1930, n1881, n1907, n1904, n1436);
or   g1898 (n1967, n1694, n1700, n1921, n1928);
nor  g1899 (n1944, n1682, n1693, n1705, n1695);
and  g1900 (n1960, n1683, n1912, n1694, n1681);
xor  g1901 (n1933, n1711, n1673, n1929, n1690);
xor  g1902 (n1958, n1688, n1701, n1920, n1673);
or   g1903 (n1968, n1676, n1916, n1696, n1701);
nor  g1904 (n1964, n1923, n1675, n1928, n1698);
nand g1905 (n1950, n1687, n1926, n1674, n1673);
xnor g1906 (n1954, n1923, n1680, n1699, n1708);
nor  g1907 (n1965, n1679, n1710, n1915);
nand g1908 (n1936, n1916, n1924, n1680, n1697);
xor  g1909 (n1959, n1688, n1930, n1681, n1693);
or   g1910 (n1962, n1696, n1682, n1674, n1683);
nor  g1911 (n1955, n1929, n1700, n1702, n1926);
nand g1912 (n1956, n1922, n1911, n1913);
nand g1913 (n1945, n1921, n1685, n1696, n1707);
xnor g1914 (n1951, n1925, n1703, n1677, n1919);
xor  g1915 (n1952, n1686, n1708, n1914, n1694);
and  g1916 (n1961, n1684, n1706, n1693, n1678);
or   g1917 (n1963, n1709, n1699, n1686, n1691);
xor  g1918 (n1946, n1917, n1689, n1703, n1709);
or   g1919 (n1932, n1680, n1929, n1706, n1927);
nor  g1920 (n1937, n1684, n1695, n1918, n1682);
nor  g1921 (n1935, n1681, n1706, n1703, n1690);
nand g1922 (n1942, n1684, n1702, n1697, n1920);
xnor g1923 (n1966, n1704, n1924, n1918, n1697);
nor  g1924 (n1949, n1686, n1927, n1683, n1679);
xnor g1925 (n1934, n1712, n1914, n1704, n1701);
or   g1926 (n1943, n1687, n1687, n1700, n1702);
and  g1927 (n1939, n1692, n1689, n1691, n1925);
xnor g1928 (n1948, n1699, n1691, n1705, n1710);
nor  g1929 (n1947, n1709, n1930, n1698, n1688);
or   g1930 (n1941, n1679, n1919, n1917, n1707);
xnor g1931 (n1957, n1922, n1711, n1698, n1677);
and  g1932 (n1970, n1675, n1915, n1707, n1678);
or   g1933 (n1969, n1695, n1676, n1930, n1708);
or   g1934 (n1938, n1689, n1678, n1705, n1676);
xor  g1935 (n1931, n1704, n1677, n1692, n1712);
nand g1936 (n1953, n1690, n1674, n1711, n1675);
xor  g1937 (n1940, n1685, n1685, n1712, n1692);
and  g1938 (n1985, n1730, n1959, n1946, n1962);
or   g1939 (n2005, n1777, n1965, n1800);
nor  g1940 (n1977, n1933, n1725, n1757, n1944);
xor  g1941 (n2009, n1955, n1958, n1942, n1774);
nor  g1942 (n1986, n673, n1745, n1969, n1779);
nand g1943 (n2000, n1732, n1769, n1948, n1947);
or   g1944 (n1998, n1945, n1750, n1969);
or   g1945 (n1993, n1932, n1739, n1953, n1934);
xnor g1946 (n1976, n1776, n1944, n1966, n1941);
xor  g1947 (n1987, n1738, n1962, n1788, n1787);
xor  g1948 (n1979, n1963, n1952, n1939, n1957);
xor  g1949 (n2010, n1764, n1970, n1763, n1933);
nor  g1950 (n2002, n1784, n1749, n1940, n1798);
xor  g1951 (n2018, n1786, n1947, n1746, n1968);
xnor g1952 (n2007, n1939, n1729, n1942, n1781);
nor  g1953 (n1997, n1940, n1968, n1736, n1943);
xor  g1954 (n2004, n1943, n1743, n1951, n1963);
nor  g1955 (n1984, n1956, n1950, n1958, n1935);
nand g1956 (n2006, n1759, n1946, n1937, n1748);
or   g1957 (n1980, n1961, n1948, n1744);
xnor g1958 (n2003, n1791, n1964, n1959, n1954);
and  g1959 (n1972, n1931, n1954, n1951, n1956);
nor  g1960 (n1988, n1735, n1967, n1726, n1953);
or   g1961 (n1992, n1967, n1932, n1961, n1797);
xor  g1962 (n1982, n1773, n1944, n1772, n1767);
xor  g1963 (n1990, n1782, n1742, n1949);
xor  g1964 (n1991, n1790, n1943, n1799, n1728);
xor  g1965 (n2013, n1970, n1747, n1952, n1958);
xor  g1966 (n2017, n1938, n1795, n1771, n1964);
xnor g1967 (n2011, n1952, n1931, n1960, n1789);
or   g1968 (n1978, n1794, n1966, n1945, n1960);
and  g1969 (n1973, n1796, n1951, n1938, n1970);
or   g1970 (n2016, n1942, n1783, n1954, n1792);
nor  g1971 (n2001, n1936, n1727, n1955, n1934);
nand g1972 (n1975, n1737, n1955, n1785, n1741);
nand g1973 (n1995, n1961, n1939, n1766, n1966);
nand g1974 (n1996, n1964, n1960, n1770, n1936);
nand g1975 (n1974, n1778, n1793, n1967, n1947);
xor  g1976 (n2008, n1753, n1957, n1761, n1963);
or   g1977 (n2012, n1941, n1953, n1956, n1775);
nand g1978 (n1989, n1765, n1937, n1755, n1962);
nand g1979 (n2015, n1938, n1945, n1965, n1959);
nor  g1980 (n1999, n1968, n1937, n1950, n1801);
or   g1981 (n1983, n1751, n1768, n1758, n1957);
and  g1982 (n1981, n1780, n1754, n1733, n1946);
nand g1983 (n1971, n1949, n1760, n1950, n1941);
nand g1984 (n2014, n1740, n1762, n1734, n1756);
or   g1985 (n1994, n1940, n1935, n1731, n1752);
and  g1986 (n2020, n1993, n1807, n2000, n1991);
xor  g1987 (n2024, n2004, n673, n2006, n1806);
xnor g1988 (n2025, n1992, n1997, n1990, n2011);
or   g1989 (n2023, n2010, n1994, n1999, n2007);
xor  g1990 (n2027, n1806, n2003, n2008, n1979);
xnor g1991 (n2029, n2017, n1974, n2002, n1995);
xor  g1992 (n2031, n1980, n1305, n2016, n2012);
nor  g1993 (n2021, n1998, n1996, n1984, n1972);
and  g1994 (n2032, n1807, n1985, n1982, n1987);
or   g1995 (n2022, n1306, n1978, n2009, n1973);
and  g1996 (n2026, n1989, n1976, n1986, n1977);
and  g1997 (n2030, n2001, n1981, n1988, n2015);
nor  g1998 (n2028, n1971, n1983, n2014, n2013);
and  g1999 (n2019, n2005, n2018, n1807, n1975);
endmodule
