

module Stat_100_41
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n131,
  n117,
  n108,
  n125,
  n121,
  n130,
  n118,
  n102,
  n116,
  n110,
  n124,
  n128,
  n122,
  n114,
  n104,
  n109,
  n113,
  n123,
  n101,
  n127,
  n105,
  n119,
  n103,
  n120,
  n106,
  n132,
  n129,
  n107,
  n126,
  n111,
  n115,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n112;output n131;output n117;output n108;output n125;output n121;output n130;output n118;output n102;output n116;output n110;output n124;output n128;output n122;output n114;output n104;output n109;output n113;output n123;output n101;output n127;output n105;output n119;output n103;output n120;output n106;output n132;output n129;output n107;output n126;output n111;output n115;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n40,
    n4
  );


  not
  g1
  (
    KeyWire_0_29,
    n2
  );


  not
  g2
  (
    KeyWire_0_11,
    n3
  );


  buf
  g3
  (
    KeyWire_0_25,
    n3
  );


  buf
  g4
  (
    n35,
    n2
  );


  not
  g5
  (
    n41,
    n1
  );


  buf
  g6
  (
    KeyWire_0_7,
    n3
  );


  not
  g7
  (
    n38,
    n4
  );


  buf
  g8
  (
    n36,
    n1
  );


  not
  g9
  (
    n43,
    n1
  );


  buf
  g10
  (
    n33,
    n2
  );


  not
  g11
  (
    KeyWire_0_16,
    n4
  );


  not
  g12
  (
    KeyWire_0_0,
    n13
  );


  buf
  g13
  (
    n66,
    n15
  );


  buf
  g14
  (
    KeyWire_0_14,
    n27
  );


  not
  g15
  (
    KeyWire_0_10,
    n8
  );


  not
  g16
  (
    n51,
    n31
  );


  not
  g17
  (
    n73,
    n33
  );


  buf
  g18
  (
    n71,
    n31
  );


  not
  g19
  (
    KeyWire_0_30,
    n19
  );


  or
  g20
  (
    n61,
    n11,
    n21,
    n18,
    n42
  );


  nor
  g21
  (
    KeyWire_0_12,
    n22,
    n41,
    n36,
    n18
  );


  nand
  g22
  (
    KeyWire_0_8,
    n35,
    n17,
    n25,
    n20
  );


  nand
  g23
  (
    n45,
    n37,
    n39,
    n42,
    n43
  );


  nor
  g24
  (
    KeyWire_0_6,
    n22,
    n19,
    n35,
    n44
  );


  or
  g25
  (
    KeyWire_0_9,
    n18,
    n13,
    n7,
    n28
  );


  xor
  g26
  (
    n60,
    n43,
    n30,
    n39,
    n38
  );


  xor
  g27
  (
    n49,
    n29,
    n24,
    n6,
    n26
  );


  nor
  g28
  (
    n65,
    n40,
    n14,
    n9,
    n11
  );


  and
  g29
  (
    KeyWire_0_18,
    n7,
    n16,
    n10,
    n19
  );


  or
  g30
  (
    KeyWire_0_4,
    n9,
    n35,
    n16,
    n42
  );


  and
  g31
  (
    n69,
    n29,
    n41,
    n37,
    n20
  );


  and
  g32
  (
    KeyWire_0_23,
    n37,
    n44,
    n23,
    n27
  );


  nand
  g33
  (
    KeyWire_0_26,
    n32,
    n25,
    n34,
    n5
  );


  and
  g34
  (
    n52,
    n14,
    n38,
    n44,
    n8
  );


  xor
  g35
  (
    n55,
    n9,
    n23,
    n22,
    n15
  );


  and
  g36
  (
    KeyWire_0_3,
    n17,
    n6,
    n33,
    n43
  );


  nand
  g37
  (
    n47,
    n12,
    n24,
    n5,
    n26
  );


  or
  g38
  (
    KeyWire_0_1,
    n24,
    n16,
    n32,
    n13
  );


  and
  g39
  (
    n48,
    n29,
    n11,
    n7,
    n26
  );


  nand
  g40
  (
    n46,
    n30,
    n36,
    n40,
    n6
  );


  nor
  g41
  (
    n56,
    n30,
    n39,
    n21,
    n10
  );


  nand
  g42
  (
    n54,
    n25,
    n10,
    n41,
    n31
  );


  nand
  g43
  (
    n67,
    n14,
    n15,
    n5,
    n8
  );


  nor
  g44
  (
    n57,
    n38,
    n27,
    n36,
    n32
  );


  and
  g45
  (
    KeyWire_0_5,
    n17,
    n34,
    n33,
    n20
  );


  xor
  g46
  (
    n77,
    n28,
    n23,
    n12,
    n40
  );


  xor
  g47
  (
    KeyWire_0_27,
    n34,
    n21,
    n12,
    n28
  );


  buf
  g48
  (
    KeyWire_0_13,
    n45
  );


  not
  g49
  (
    n84,
    n49
  );


  buf
  g50
  (
    n81,
    n48
  );


  buf
  g51
  (
    n92,
    n45
  );


  buf
  g52
  (
    n83,
    n46
  );


  buf
  g53
  (
    n91,
    n48
  );


  buf
  g54
  (
    n85,
    n46
  );


  not
  g55
  (
    n90,
    n50
  );


  buf
  g56
  (
    KeyWire_0_2,
    n50
  );


  buf
  g57
  (
    n89,
    n49
  );


  buf
  g58
  (
    KeyWire_0_22,
    n51
  );


  not
  g59
  (
    n88,
    n51
  );


  buf
  g60
  (
    n86,
    n48
  );


  buf
  g61
  (
    KeyWire_0_15,
    n50
  );


  not
  g62
  (
    n98,
    n46
  );


  buf
  g63
  (
    n93,
    n45
  );


  buf
  g64
  (
    n87,
    n47
  );


  not
  g65
  (
    n97,
    n47
  );


  not
  g66
  (
    KeyWire_0_31,
    n47
  );


  not
  g67
  (
    n95,
    n49
  );


  or
  g68
  (
    KeyWire_0_17,
    n97,
    n64,
    n98,
    n70
  );


  xnor
  g69
  (
    n102,
    n60,
    n80,
    n95
  );


  or
  g70
  (
    n125,
    n78,
    n74,
    n71,
    n77
  );


  or
  g71
  (
    n130,
    n57,
    n63,
    n69,
    n99
  );


  xnor
  g72
  (
    n121,
    n88,
    n56,
    n72,
    n58
  );


  or
  g73
  (
    n128,
    n70,
    n91,
    n94,
    n60
  );


  or
  g74
  (
    n113,
    n71,
    n54,
    n51,
    n59
  );


  nand
  g75
  (
    KeyWire_0_21,
    n86,
    n94,
    n62
  );


  nand
  g76
  (
    n129,
    n82,
    n75,
    n52,
    n61
  );


  and
  g77
  (
    n112,
    n62,
    n85,
    n54,
    n75
  );


  xor
  g78
  (
    n108,
    n59,
    n79,
    n68,
    n91
  );


  xor
  g79
  (
    n114,
    n69,
    n92,
    n53,
    n65
  );


  xor
  g80
  (
    n119,
    n83,
    n91,
    n60,
    n68
  );


  nand
  g81
  (
    KeyWire_0_20,
    n74,
    n72,
    n89,
    n65
  );


  xor
  g82
  (
    n105,
    n68,
    n64,
    n81,
    n92
  );


  xnor
  g83
  (
    n110,
    n53,
    n92,
    n99,
    n98
  );


  or
  g84
  (
    KeyWire_0_24,
    n56,
    n56,
    n61,
    n66
  );


  nand
  g85
  (
    n106,
    n65,
    n99,
    n93,
    n74
  );


  nand
  g86
  (
    n118,
    n73,
    n55,
    n78,
    n76
  );


  xnor
  g87
  (
    n123,
    n95,
    n87,
    n71,
    n55
  );


  nor
  g88
  (
    n107,
    n97,
    n70,
    n84,
    n79
  );


  nor
  g89
  (
    n103,
    n58,
    n77,
    n66,
    n52
  );


  nand
  g90
  (
    n122,
    n63,
    n80,
    n59,
    n93
  );


  nand
  g91
  (
    n109,
    n64,
    n72,
    n100,
    n57
  );


  nor
  g92
  (
    KeyWire_0_19,
    n58,
    n67,
    n73,
    n66
  );


  xor
  g93
  (
    n117,
    n100,
    n73,
    n80,
    n96
  );


  and
  g94
  (
    n124,
    n54,
    n67,
    n90,
    n61
  );


  xnor
  g95
  (
    KeyWire_0_28,
    n76,
    n75,
    n52,
    n53
  );


  or
  g96
  (
    n132,
    n67,
    n93,
    n96,
    n78
  );


  or
  g97
  (
    n131,
    n98,
    n96,
    n94,
    n79
  );


  nor
  g98
  (
    n116,
    n69,
    n97,
    n57,
    n100
  );


  or
  g99
  (
    n127,
    n55,
    n76,
    n63,
    n77
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n59,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n79,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n82,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n70,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n58,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n68,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n80,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n37,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n78,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n74,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n72,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n34,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n64,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n96,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n76,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n100,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n44,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n120,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n50,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n126,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n104,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n115,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n94,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n53,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n101,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n42,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n63,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n62,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n111,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n39,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n75,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n99,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

