

module Stat_2068_22_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n1300,
  n1261,
  n1285,
  n1276,
  n1264,
  n1287,
  n1269,
  n1299,
  n1272,
  n1289,
  n1278,
  n1294,
  n1275,
  n1265,
  n1283,
  n1280,
  n1262,
  n1286,
  n1267,
  n1293,
  n1297,
  n1296,
  n1281,
  n1277,
  n1303,
  n1273,
  n1365,
  n1382,
  n1383,
  n1372,
  n1381,
  n1374,
  n1384,
  n1377,
  n1369,
  n2095,
  n2088,
  n2098,
  n2087,
  n2089,
  n2090,
  n2091,
  n2092,
  n2093,
  n2097,
  n2094,
  n2096,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1300;output n1261;output n1285;output n1276;output n1264;output n1287;output n1269;output n1299;output n1272;output n1289;output n1278;output n1294;output n1275;output n1265;output n1283;output n1280;output n1262;output n1286;output n1267;output n1293;output n1297;output n1296;output n1281;output n1277;output n1303;output n1273;output n1365;output n1382;output n1383;output n1372;output n1381;output n1374;output n1384;output n1377;output n1369;output n2095;output n2088;output n2098;output n2087;output n2089;output n2090;output n2091;output n2092;output n2093;output n2097;output n2094;output n2096;
  wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1263;wire n1266;wire n1268;wire n1270;wire n1271;wire n1274;wire n1279;wire n1282;wire n1284;wire n1288;wire n1290;wire n1291;wire n1292;wire n1295;wire n1298;wire n1301;wire n1302;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1366;wire n1367;wire n1368;wire n1370;wire n1371;wire n1373;wire n1375;wire n1376;wire n1378;wire n1379;wire n1380;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n67,
    n20
  );


  buf
  g1
  (
    n32,
    n3
  );


  not
  g2
  (
    n133,
    n30
  );


  not
  g3
  (
    n135,
    n21
  );


  not
  g4
  (
    n65,
    n10
  );


  buf
  g5
  (
    n42,
    n13
  );


  not
  g6
  (
    n64,
    n17
  );


  not
  g7
  (
    n103,
    n16
  );


  not
  g8
  (
    n89,
    n11
  );


  buf
  g9
  (
    n117,
    n7
  );


  not
  g10
  (
    n84,
    n1
  );


  buf
  g11
  (
    n54,
    n23
  );


  buf
  g12
  (
    n137,
    n2
  );


  not
  g13
  (
    n141,
    n4
  );


  buf
  g14
  (
    n98,
    n1
  );


  not
  g15
  (
    n114,
    n26
  );


  not
  g16
  (
    n73,
    n14
  );


  not
  g17
  (
    n33,
    n11
  );


  not
  g18
  (
    n68,
    n6
  );


  buf
  g19
  (
    n92,
    n23
  );


  not
  g20
  (
    n34,
    n19
  );


  buf
  g21
  (
    n118,
    n17
  );


  buf
  g22
  (
    n150,
    n15
  );


  buf
  g23
  (
    n124,
    n8
  );


  buf
  g24
  (
    KeyWire_0_22,
    n22
  );


  not
  g25
  (
    n112,
    n17
  );


  not
  g26
  (
    n76,
    n7
  );


  buf
  g27
  (
    n121,
    n27
  );


  not
  g28
  (
    n142,
    n5
  );


  buf
  g29
  (
    n72,
    n22
  );


  buf
  g30
  (
    n96,
    n30
  );


  not
  g31
  (
    KeyWire_0_21,
    n24
  );


  buf
  g32
  (
    n46,
    n18
  );


  buf
  g33
  (
    n138,
    n22
  );


  buf
  g34
  (
    n36,
    n6
  );


  not
  g35
  (
    n31,
    n2
  );


  buf
  g36
  (
    n108,
    n29
  );


  buf
  g37
  (
    n49,
    n10
  );


  not
  g38
  (
    n58,
    n10
  );


  buf
  g39
  (
    n93,
    n20
  );


  not
  g40
  (
    n44,
    n3
  );


  buf
  g41
  (
    n47,
    n21
  );


  not
  g42
  (
    n60,
    n25
  );


  not
  g43
  (
    n125,
    n26
  );


  not
  g44
  (
    n102,
    n20
  );


  buf
  g45
  (
    n110,
    n5
  );


  buf
  g46
  (
    n51,
    n12
  );


  not
  g47
  (
    KeyWire_0_15,
    n28
  );


  buf
  g48
  (
    n74,
    n15
  );


  buf
  g49
  (
    n80,
    n27
  );


  not
  g50
  (
    n55,
    n19
  );


  not
  g51
  (
    n97,
    n16
  );


  buf
  g52
  (
    n50,
    n18
  );


  not
  g53
  (
    n120,
    n28
  );


  buf
  g54
  (
    n56,
    n9
  );


  buf
  g55
  (
    n109,
    n4
  );


  buf
  g56
  (
    n61,
    n20
  );


  not
  g57
  (
    n94,
    n27
  );


  buf
  g58
  (
    n106,
    n25
  );


  not
  g59
  (
    n107,
    n18
  );


  not
  g60
  (
    n126,
    n16
  );


  not
  g61
  (
    n59,
    n29
  );


  buf
  g62
  (
    n88,
    n15
  );


  buf
  g63
  (
    n45,
    n8
  );


  not
  g64
  (
    n91,
    n24
  );


  buf
  g65
  (
    n143,
    n10
  );


  not
  g66
  (
    n41,
    n6
  );


  buf
  g67
  (
    n129,
    n1
  );


  buf
  g68
  (
    n148,
    n25
  );


  not
  g69
  (
    n39,
    n4
  );


  not
  g70
  (
    n35,
    n5
  );


  buf
  g71
  (
    n85,
    n9
  );


  not
  g72
  (
    n53,
    n15
  );


  not
  g73
  (
    n63,
    n19
  );


  buf
  g74
  (
    n115,
    n9
  );


  buf
  g75
  (
    n71,
    n1
  );


  buf
  g76
  (
    n69,
    n8
  );


  buf
  g77
  (
    n147,
    n23
  );


  buf
  g78
  (
    n38,
    n23
  );


  not
  g79
  (
    n101,
    n2
  );


  buf
  g80
  (
    n90,
    n14
  );


  buf
  g81
  (
    n62,
    n11
  );


  not
  g82
  (
    n131,
    n7
  );


  buf
  g83
  (
    n136,
    n25
  );


  not
  g84
  (
    n100,
    n28
  );


  not
  g85
  (
    n87,
    n19
  );


  not
  g86
  (
    n128,
    n24
  );


  buf
  g87
  (
    n104,
    n30
  );


  buf
  g88
  (
    n140,
    n13
  );


  buf
  g89
  (
    n132,
    n24
  );


  not
  g90
  (
    n52,
    n3
  );


  not
  g91
  (
    n134,
    n12
  );


  not
  g92
  (
    n123,
    n11
  );


  buf
  g93
  (
    n139,
    n12
  );


  not
  g94
  (
    n78,
    n17
  );


  buf
  g95
  (
    n77,
    n14
  );


  not
  g96
  (
    n122,
    n14
  );


  buf
  g97
  (
    n37,
    n4
  );


  buf
  g98
  (
    n95,
    n6
  );


  buf
  g99
  (
    n145,
    n13
  );


  buf
  g100
  (
    n57,
    n12
  );


  buf
  g101
  (
    n144,
    n2
  );


  buf
  g102
  (
    n113,
    n9
  );


  buf
  g103
  (
    n130,
    n28
  );


  buf
  g104
  (
    n149,
    n5
  );


  not
  g105
  (
    n70,
    n7
  );


  not
  g106
  (
    n75,
    n29
  );


  buf
  g107
  (
    n99,
    n29
  );


  not
  g108
  (
    n146,
    n26
  );


  buf
  g109
  (
    n111,
    n22
  );


  not
  g110
  (
    n81,
    n13
  );


  not
  g111
  (
    n83,
    n18
  );


  not
  g112
  (
    n116,
    n21
  );


  not
  g113
  (
    n119,
    n26
  );


  buf
  g114
  (
    n127,
    n21
  );


  buf
  g115
  (
    n43,
    n3
  );


  buf
  g116
  (
    n79,
    n30
  );


  not
  g117
  (
    n66,
    n27
  );


  not
  g118
  (
    KeyWire_0_2,
    n16
  );


  buf
  g119
  (
    n86,
    n8
  );


  not
  g120
  (
    n227,
    n85
  );


  not
  g121
  (
    n244,
    n75
  );


  not
  g122
  (
    n463,
    n83
  );


  not
  g123
  (
    n513,
    n36
  );


  not
  g124
  (
    n165,
    n121
  );


  buf
  g125
  (
    n467,
    n108
  );


  buf
  g126
  (
    n461,
    n85
  );


  not
  g127
  (
    n402,
    n108
  );


  buf
  g128
  (
    n597,
    n58
  );


  buf
  g129
  (
    n283,
    n92
  );


  buf
  g130
  (
    n559,
    n141
  );


  not
  g131
  (
    n213,
    n71
  );


  not
  g132
  (
    n560,
    n144
  );


  not
  g133
  (
    n242,
    n37
  );


  buf
  g134
  (
    n486,
    n79
  );


  not
  g135
  (
    n366,
    n107
  );


  buf
  g136
  (
    n552,
    n69
  );


  not
  g137
  (
    n209,
    n32
  );


  not
  g138
  (
    n306,
    n139
  );


  buf
  g139
  (
    n528,
    n45
  );


  buf
  g140
  (
    n501,
    n116
  );


  buf
  g141
  (
    n553,
    n136
  );


  not
  g142
  (
    n293,
    n103
  );


  buf
  g143
  (
    n404,
    n102
  );


  buf
  g144
  (
    n427,
    n64
  );


  buf
  g145
  (
    n511,
    n50
  );


  buf
  g146
  (
    n519,
    n105
  );


  buf
  g147
  (
    n415,
    n46
  );


  not
  g148
  (
    n436,
    n143
  );


  buf
  g149
  (
    n545,
    n66
  );


  buf
  g150
  (
    n155,
    n88
  );


  not
  g151
  (
    n591,
    n86
  );


  not
  g152
  (
    n162,
    n106
  );


  buf
  g153
  (
    n389,
    n84
  );


  not
  g154
  (
    n580,
    n101
  );


  not
  g155
  (
    n367,
    n67
  );


  buf
  g156
  (
    n369,
    n35
  );


  buf
  g157
  (
    n157,
    n31
  );


  not
  g158
  (
    n601,
    n89
  );


  buf
  g159
  (
    n495,
    n100
  );


  buf
  g160
  (
    n193,
    n98
  );


  buf
  g161
  (
    n605,
    n60
  );


  buf
  g162
  (
    n466,
    n82
  );


  not
  g163
  (
    n252,
    n66
  );


  buf
  g164
  (
    n421,
    n139
  );


  not
  g165
  (
    n212,
    n93
  );


  not
  g166
  (
    n592,
    n53
  );


  not
  g167
  (
    n181,
    n123
  );


  buf
  g168
  (
    n422,
    n52
  );


  buf
  g169
  (
    n454,
    n35
  );


  not
  g170
  (
    n185,
    n119
  );


  buf
  g171
  (
    n465,
    n114
  );


  buf
  g172
  (
    n507,
    n125
  );


  not
  g173
  (
    n310,
    n74
  );


  not
  g174
  (
    n362,
    n99
  );


  not
  g175
  (
    n243,
    n45
  );


  not
  g176
  (
    n566,
    n114
  );


  not
  g177
  (
    n499,
    n42
  );


  buf
  g178
  (
    n236,
    n142
  );


  not
  g179
  (
    n285,
    n33
  );


  buf
  g180
  (
    n479,
    n65
  );


  buf
  g181
  (
    n319,
    n91
  );


  buf
  g182
  (
    n260,
    n53
  );


  buf
  g183
  (
    n448,
    n126
  );


  buf
  g184
  (
    n224,
    n80
  );


  not
  g185
  (
    KeyWire_0_19,
    n128
  );


  buf
  g186
  (
    n583,
    n73
  );


  not
  g187
  (
    n251,
    n138
  );


  buf
  g188
  (
    n468,
    n43
  );


  not
  g189
  (
    n456,
    n140
  );


  not
  g190
  (
    n284,
    n104
  );


  buf
  g191
  (
    n523,
    n72
  );


  not
  g192
  (
    n378,
    n130
  );


  not
  g193
  (
    n270,
    n112
  );


  buf
  g194
  (
    n175,
    n42
  );


  buf
  g195
  (
    n584,
    n41
  );


  buf
  g196
  (
    n573,
    n126
  );


  not
  g197
  (
    n277,
    n34
  );


  buf
  g198
  (
    n163,
    n72
  );


  buf
  g199
  (
    KeyWire_0_4,
    n78
  );


  not
  g200
  (
    n509,
    n133
  );


  buf
  g201
  (
    n439,
    n126
  );


  not
  g202
  (
    n401,
    n78
  );


  not
  g203
  (
    n409,
    n39
  );


  not
  g204
  (
    n491,
    n46
  );


  not
  g205
  (
    n506,
    n112
  );


  buf
  g206
  (
    n395,
    n54
  );


  buf
  g207
  (
    n254,
    n104
  );


  not
  g208
  (
    n291,
    n136
  );


  buf
  g209
  (
    n354,
    n47
  );


  not
  g210
  (
    n267,
    n57
  );


  buf
  g211
  (
    n297,
    n61
  );


  not
  g212
  (
    n426,
    n131
  );


  buf
  g213
  (
    n218,
    n115
  );


  buf
  g214
  (
    n535,
    n135
  );


  not
  g215
  (
    n237,
    n49
  );


  not
  g216
  (
    n200,
    n105
  );


  buf
  g217
  (
    n440,
    n137
  );


  buf
  g218
  (
    n177,
    n143
  );


  buf
  g219
  (
    n159,
    n101
  );


  not
  g220
  (
    n292,
    n131
  );


  buf
  g221
  (
    n544,
    n107
  );


  buf
  g222
  (
    n525,
    n34
  );


  not
  g223
  (
    n205,
    n116
  );


  not
  g224
  (
    n450,
    n55
  );


  not
  g225
  (
    n432,
    n98
  );


  buf
  g226
  (
    n392,
    n68
  );


  buf
  g227
  (
    n517,
    n126
  );


  buf
  g228
  (
    n555,
    n119
  );


  not
  g229
  (
    n576,
    n110
  );


  buf
  g230
  (
    n223,
    n85
  );


  not
  g231
  (
    n249,
    n143
  );


  not
  g232
  (
    n203,
    n44
  );


  buf
  g233
  (
    n444,
    n132
  );


  buf
  g234
  (
    n430,
    n101
  );


  buf
  g235
  (
    n483,
    n103
  );


  buf
  g236
  (
    n539,
    n62
  );


  buf
  g237
  (
    n323,
    n113
  );


  buf
  g238
  (
    n348,
    n86
  );


  buf
  g239
  (
    n569,
    n107
  );


  not
  g240
  (
    n289,
    n132
  );


  buf
  g241
  (
    n315,
    n40
  );


  not
  g242
  (
    n320,
    n122
  );


  not
  g243
  (
    n529,
    n139
  );


  buf
  g244
  (
    n424,
    n129
  );


  not
  g245
  (
    n441,
    n77
  );


  not
  g246
  (
    n337,
    n43
  );


  buf
  g247
  (
    n373,
    n57
  );


  not
  g248
  (
    n184,
    n90
  );


  buf
  g249
  (
    n418,
    n114
  );


  buf
  g250
  (
    n356,
    n68
  );


  not
  g251
  (
    n384,
    n123
  );


  buf
  g252
  (
    n229,
    n62
  );


  buf
  g253
  (
    n462,
    n133
  );


  buf
  g254
  (
    n302,
    n47
  );


  not
  g255
  (
    n253,
    n106
  );


  not
  g256
  (
    n408,
    n109
  );


  buf
  g257
  (
    n547,
    n31
  );


  buf
  g258
  (
    n590,
    n57
  );


  buf
  g259
  (
    n433,
    n58
  );


  not
  g260
  (
    n282,
    n64
  );


  buf
  g261
  (
    n264,
    n77
  );


  not
  g262
  (
    n370,
    n75
  );


  buf
  g263
  (
    n385,
    n37
  );


  not
  g264
  (
    n346,
    n78
  );


  buf
  g265
  (
    n480,
    n74
  );


  not
  g266
  (
    n188,
    n137
  );


  not
  g267
  (
    n574,
    n118
  );


  not
  g268
  (
    n311,
    n47
  );


  not
  g269
  (
    n464,
    n52
  );


  buf
  g270
  (
    n414,
    n109
  );


  buf
  g271
  (
    n363,
    n33
  );


  not
  g272
  (
    n508,
    n76
  );


  buf
  g273
  (
    n296,
    n34
  );


  buf
  g274
  (
    n295,
    n97
  );


  buf
  g275
  (
    n156,
    n139
  );


  buf
  g276
  (
    n561,
    n94
  );


  not
  g277
  (
    n562,
    n133
  );


  not
  g278
  (
    n210,
    n39
  );


  buf
  g279
  (
    n220,
    n94
  );


  buf
  g280
  (
    n231,
    n117
  );


  buf
  g281
  (
    n393,
    n56
  );


  buf
  g282
  (
    n215,
    n38
  );


  not
  g283
  (
    n411,
    n69
  );


  not
  g284
  (
    n504,
    n64
  );


  not
  g285
  (
    n279,
    n130
  );


  not
  g286
  (
    n376,
    n32
  );


  not
  g287
  (
    n221,
    n74
  );


  buf
  g288
  (
    n326,
    n90
  );


  buf
  g289
  (
    n299,
    n108
  );


  buf
  g290
  (
    n204,
    n88
  );


  not
  g291
  (
    n412,
    n117
  );


  not
  g292
  (
    n485,
    n36
  );


  not
  g293
  (
    n546,
    n76
  );


  not
  g294
  (
    n298,
    n107
  );


  buf
  g295
  (
    n338,
    n87
  );


  not
  g296
  (
    n405,
    n109
  );


  buf
  g297
  (
    n154,
    n56
  );


  not
  g298
  (
    n452,
    n127
  );


  buf
  g299
  (
    n558,
    n62
  );


  buf
  g300
  (
    n312,
    n59
  );


  buf
  g301
  (
    n374,
    n43
  );


  buf
  g302
  (
    n358,
    n118
  );


  buf
  g303
  (
    n304,
    n140
  );


  buf
  g304
  (
    n365,
    n142
  );


  not
  g305
  (
    n275,
    n124
  );


  not
  g306
  (
    n322,
    n77
  );


  not
  g307
  (
    n241,
    n51
  );


  not
  g308
  (
    n457,
    n88
  );


  not
  g309
  (
    n271,
    n33
  );


  not
  g310
  (
    n478,
    n110
  );


  not
  g311
  (
    n214,
    n36
  );


  not
  g312
  (
    n589,
    n84
  );


  not
  g313
  (
    n470,
    n120
  );


  buf
  g314
  (
    n161,
    n137
  );


  not
  g315
  (
    n153,
    n73
  );


  not
  g316
  (
    n600,
    n109
  );


  not
  g317
  (
    n488,
    n72
  );


  buf
  g318
  (
    n342,
    n89
  );


  buf
  g319
  (
    n531,
    n37
  );


  not
  g320
  (
    n476,
    n105
  );


  buf
  g321
  (
    n554,
    n96
  );


  buf
  g322
  (
    n194,
    n120
  );


  buf
  g323
  (
    n208,
    n117
  );


  buf
  g324
  (
    n572,
    n35
  );


  buf
  g325
  (
    n331,
    n106
  );


  buf
  g326
  (
    n364,
    n40
  );


  buf
  g327
  (
    n190,
    n73
  );


  not
  g328
  (
    n187,
    n62
  );


  not
  g329
  (
    n556,
    n71
  );


  not
  g330
  (
    n514,
    n67
  );


  not
  g331
  (
    n413,
    n83
  );


  buf
  g332
  (
    n276,
    n82
  );


  not
  g333
  (
    n330,
    n93
  );


  buf
  g334
  (
    n602,
    n92
  );


  buf
  g335
  (
    n341,
    n95
  );


  not
  g336
  (
    n334,
    n61
  );


  buf
  g337
  (
    n472,
    n134
  );


  not
  g338
  (
    n381,
    n132
  );


  buf
  g339
  (
    n186,
    n35
  );


  not
  g340
  (
    n327,
    n89
  );


  not
  g341
  (
    n325,
    n41
  );


  buf
  g342
  (
    n172,
    n134
  );


  not
  g343
  (
    n459,
    n52
  );


  buf
  g344
  (
    KeyWire_0_30,
    n56
  );


  not
  g345
  (
    n564,
    n50
  );


  buf
  g346
  (
    n570,
    n79
  );


  buf
  g347
  (
    n451,
    n110
  );


  buf
  g348
  (
    n429,
    n122
  );


  not
  g349
  (
    n280,
    n119
  );


  buf
  g350
  (
    n522,
    n48
  );


  buf
  g351
  (
    n567,
    n55
  );


  not
  g352
  (
    n178,
    n140
  );


  buf
  g353
  (
    n386,
    n55
  );


  not
  g354
  (
    n192,
    n67
  );


  not
  g355
  (
    n353,
    n95
  );


  buf
  g356
  (
    n526,
    n93
  );


  not
  g357
  (
    n189,
    n53
  );


  not
  g358
  (
    n520,
    n39
  );


  not
  g359
  (
    n173,
    n140
  );


  not
  g360
  (
    n332,
    n32
  );


  buf
  g361
  (
    n582,
    n51
  );


  buf
  g362
  (
    n216,
    n115
  );


  buf
  g363
  (
    n489,
    n113
  );


  not
  g364
  (
    n383,
    n42
  );


  buf
  g365
  (
    n375,
    n102
  );


  not
  g366
  (
    KeyWire_0_8,
    n60
  );


  not
  g367
  (
    n434,
    n118
  );


  buf
  g368
  (
    n417,
    n111
  );


  not
  g369
  (
    n536,
    n102
  );


  buf
  g370
  (
    n349,
    n98
  );


  not
  g371
  (
    n391,
    n44
  );


  not
  g372
  (
    n586,
    n59
  );


  buf
  g373
  (
    n226,
    n55
  );


  not
  g374
  (
    n577,
    n128
  );


  buf
  g375
  (
    n183,
    n56
  );


  not
  g376
  (
    n598,
    n130
  );


  buf
  g377
  (
    n256,
    n128
  );


  not
  g378
  (
    n222,
    n41
  );


  buf
  g379
  (
    n477,
    n63
  );


  not
  g380
  (
    n446,
    n141
  );


  buf
  g381
  (
    n578,
    n127
  );


  buf
  g382
  (
    n387,
    n61
  );


  not
  g383
  (
    n281,
    n65
  );


  not
  g384
  (
    n388,
    n118
  );


  buf
  g385
  (
    n169,
    n84
  );


  buf
  g386
  (
    n596,
    n111
  );


  not
  g387
  (
    n211,
    n87
  );


  buf
  g388
  (
    n359,
    n116
  );


  buf
  g389
  (
    n435,
    n134
  );


  buf
  g390
  (
    n581,
    n84
  );


  not
  g391
  (
    n599,
    n135
  );


  buf
  g392
  (
    n443,
    n33
  );


  buf
  g393
  (
    n355,
    n89
  );


  buf
  g394
  (
    n329,
    n86
  );


  buf
  g395
  (
    n288,
    n58
  );


  buf
  g396
  (
    n345,
    n68
  );


  buf
  g397
  (
    KeyWire_0_26,
    n95
  );


  buf
  g398
  (
    n447,
    n91
  );


  not
  g399
  (
    n371,
    n71
  );


  buf
  g400
  (
    n431,
    n80
  );


  buf
  g401
  (
    n420,
    n113
  );


  not
  g402
  (
    n471,
    n96
  );


  not
  g403
  (
    n449,
    n70
  );


  not
  g404
  (
    n350,
    n135
  );


  buf
  g405
  (
    n557,
    n97
  );


  buf
  g406
  (
    n542,
    n138
  );


  buf
  g407
  (
    n232,
    n130
  );


  buf
  g408
  (
    n294,
    n96
  );


  buf
  g409
  (
    n168,
    n43
  );


  not
  g410
  (
    n152,
    n113
  );


  not
  g411
  (
    n518,
    n90
  );


  buf
  g412
  (
    n151,
    n91
  );


  not
  g413
  (
    n246,
    n110
  );


  buf
  g414
  (
    n274,
    n34
  );


  buf
  g415
  (
    n245,
    n82
  );


  buf
  g416
  (
    n594,
    n49
  );


  buf
  g417
  (
    n423,
    n123
  );


  not
  g418
  (
    n160,
    n73
  );


  not
  g419
  (
    n534,
    n92
  );


  buf
  g420
  (
    n368,
    n93
  );


  not
  g421
  (
    n540,
    n87
  );


  buf
  g422
  (
    n217,
    n60
  );


  not
  g423
  (
    n352,
    n100
  );


  buf
  g424
  (
    n503,
    n111
  );


  not
  g425
  (
    n484,
    n104
  );


  not
  g426
  (
    n196,
    n75
  );


  not
  g427
  (
    n230,
    n31
  );


  buf
  g428
  (
    n530,
    n86
  );


  buf
  g429
  (
    n551,
    n67
  );


  buf
  g430
  (
    n266,
    n51
  );


  not
  g431
  (
    n233,
    n75
  );


  buf
  g432
  (
    n228,
    n63
  );


  buf
  g433
  (
    n307,
    n54
  );


  buf
  g434
  (
    n317,
    n115
  );


  buf
  g435
  (
    n541,
    n57
  );


  not
  g436
  (
    n176,
    n98
  );


  not
  g437
  (
    n516,
    n92
  );


  buf
  g438
  (
    n335,
    n66
  );


  buf
  g439
  (
    n593,
    n64
  );


  buf
  g440
  (
    n397,
    n44
  );


  not
  g441
  (
    n170,
    n81
  );


  buf
  g442
  (
    n278,
    n100
  );


  not
  g443
  (
    n498,
    n53
  );


  not
  g444
  (
    n500,
    n74
  );


  buf
  g445
  (
    n261,
    n144
  );


  not
  g446
  (
    n328,
    n111
  );


  not
  g447
  (
    n238,
    n121
  );


  buf
  g448
  (
    n336,
    n112
  );


  not
  g449
  (
    n313,
    n79
  );


  not
  g450
  (
    n604,
    n87
  );


  not
  g451
  (
    n533,
    n51
  );


  not
  g452
  (
    n512,
    n138
  );


  buf
  g453
  (
    n287,
    n129
  );


  not
  g454
  (
    n406,
    n38
  );


  not
  g455
  (
    n180,
    n95
  );


  buf
  g456
  (
    n399,
    n81
  );


  buf
  g457
  (
    n390,
    n46
  );


  buf
  g458
  (
    n191,
    n63
  );


  buf
  g459
  (
    n248,
    n61
  );


  not
  g460
  (
    n497,
    n54
  );


  not
  g461
  (
    n262,
    n121
  );


  buf
  g462
  (
    n309,
    n58
  );


  not
  g463
  (
    n321,
    n40
  );


  not
  g464
  (
    n532,
    n132
  );


  buf
  g465
  (
    n372,
    n141
  );


  not
  g466
  (
    n537,
    n71
  );


  not
  g467
  (
    n460,
    n138
  );


  not
  g468
  (
    n344,
    n39
  );


  buf
  g469
  (
    n197,
    n81
  );


  buf
  g470
  (
    n206,
    n91
  );


  buf
  g471
  (
    n357,
    n83
  );


  buf
  g472
  (
    n481,
    n68
  );


  not
  g473
  (
    n239,
    n121
  );


  not
  g474
  (
    n174,
    n134
  );


  buf
  g475
  (
    n407,
    n137
  );


  buf
  g476
  (
    n360,
    n48
  );


  buf
  g477
  (
    n377,
    n106
  );


  not
  g478
  (
    n259,
    n122
  );


  buf
  g479
  (
    n225,
    n117
  );


  not
  g480
  (
    n585,
    n94
  );


  buf
  g481
  (
    n171,
    n103
  );


  buf
  g482
  (
    n548,
    n77
  );


  buf
  g483
  (
    n527,
    n45
  );


  not
  g484
  (
    n575,
    n128
  );


  buf
  g485
  (
    n453,
    n127
  );


  not
  g486
  (
    n588,
    n32
  );


  not
  g487
  (
    n250,
    n120
  );


  not
  g488
  (
    n164,
    n103
  );


  not
  g489
  (
    n201,
    n141
  );


  buf
  g490
  (
    n515,
    n70
  );


  not
  g491
  (
    n219,
    n46
  );


  buf
  g492
  (
    n455,
    n124
  );


  buf
  g493
  (
    n361,
    n38
  );


  buf
  g494
  (
    n469,
    n41
  );


  not
  g495
  (
    n425,
    n45
  );


  not
  g496
  (
    n487,
    n76
  );


  buf
  g497
  (
    n286,
    n99
  );


  not
  g498
  (
    n303,
    n142
  );


  buf
  g499
  (
    n268,
    n99
  );


  buf
  g500
  (
    KeyWire_0_9,
    n59
  );


  buf
  g501
  (
    n543,
    n135
  );


  not
  g502
  (
    n549,
    n114
  );


  not
  g503
  (
    n300,
    n78
  );


  not
  g504
  (
    n394,
    n142
  );


  not
  g505
  (
    n438,
    n112
  );


  buf
  g506
  (
    n492,
    n49
  );


  buf
  g507
  (
    n301,
    n38
  );


  not
  g508
  (
    n396,
    n70
  );


  not
  g509
  (
    n550,
    n97
  );


  not
  g510
  (
    n240,
    n40
  );


  buf
  g511
  (
    n343,
    n99
  );


  not
  g512
  (
    n255,
    n131
  );


  buf
  g513
  (
    n490,
    n80
  );


  buf
  g514
  (
    n473,
    n37
  );


  not
  g515
  (
    n382,
    n124
  );


  buf
  g516
  (
    n563,
    n90
  );


  not
  g517
  (
    n403,
    n123
  );


  not
  g518
  (
    n445,
    n48
  );


  buf
  g519
  (
    n263,
    n63
  );


  buf
  g520
  (
    n505,
    n50
  );


  buf
  g521
  (
    n167,
    n102
  );


  buf
  g522
  (
    n571,
    n129
  );


  buf
  g523
  (
    n380,
    n69
  );


  buf
  g524
  (
    n524,
    n48
  );


  not
  g525
  (
    n202,
    n65
  );


  buf
  g526
  (
    n416,
    n31
  );


  buf
  g527
  (
    n442,
    n49
  );


  buf
  g528
  (
    n305,
    n54
  );


  not
  g529
  (
    n308,
    n122
  );


  not
  g530
  (
    n595,
    n108
  );


  buf
  g531
  (
    n158,
    n85
  );


  not
  g532
  (
    n333,
    n44
  );


  not
  g533
  (
    n400,
    n52
  );


  not
  g534
  (
    n579,
    n120
  );


  buf
  g535
  (
    n166,
    n72
  );


  buf
  g536
  (
    n195,
    n47
  );


  not
  g537
  (
    n493,
    n115
  );


  not
  g538
  (
    n474,
    n97
  );


  buf
  g539
  (
    n437,
    n50
  );


  not
  g540
  (
    n340,
    n81
  );


  not
  g541
  (
    n419,
    n42
  );


  not
  g542
  (
    n482,
    n96
  );


  not
  g543
  (
    n324,
    n143
  );


  not
  g544
  (
    n258,
    n69
  );


  buf
  g545
  (
    n458,
    n101
  );


  buf
  g546
  (
    n398,
    n136
  );


  buf
  g547
  (
    n199,
    n104
  );


  not
  g548
  (
    n290,
    n36
  );


  buf
  g549
  (
    n494,
    n79
  );


  not
  g550
  (
    n234,
    n136
  );


  not
  g551
  (
    n587,
    n124
  );


  not
  g552
  (
    n257,
    n125
  );


  buf
  g553
  (
    n273,
    n76
  );


  not
  g554
  (
    n207,
    n129
  );


  not
  g555
  (
    n521,
    n100
  );


  buf
  g556
  (
    n475,
    n60
  );


  not
  g557
  (
    n538,
    n105
  );


  buf
  g558
  (
    n568,
    n70
  );


  buf
  g559
  (
    n272,
    n125
  );


  not
  g560
  (
    n198,
    n83
  );


  buf
  g561
  (
    n565,
    n65
  );


  not
  g562
  (
    n314,
    n127
  );


  buf
  g563
  (
    n247,
    n131
  );


  not
  g564
  (
    n510,
    n133
  );


  not
  g565
  (
    n496,
    n94
  );


  not
  g566
  (
    n428,
    n82
  );


  not
  g567
  (
    n316,
    n125
  );


  buf
  g568
  (
    n603,
    n59
  );


  buf
  g569
  (
    n179,
    n116
  );


  not
  g570
  (
    n265,
    n80
  );


  buf
  g571
  (
    n318,
    n88
  );


  not
  g572
  (
    n379,
    n66
  );


  buf
  g573
  (
    n502,
    n144
  );


  buf
  g574
  (
    n182,
    n119
  );


  not
  g575
  (
    n890,
    n352
  );


  not
  g576
  (
    n806,
    n340
  );


  buf
  g577
  (
    n726,
    n520
  );


  buf
  g578
  (
    n939,
    n542
  );


  not
  g579
  (
    n1209,
    n581
  );


  not
  g580
  (
    n1128,
    n396
  );


  not
  g581
  (
    n955,
    n283
  );


  not
  g582
  (
    n752,
    n399
  );


  not
  g583
  (
    n815,
    n543
  );


  not
  g584
  (
    n796,
    n316
  );


  buf
  g585
  (
    n944,
    n541
  );


  not
  g586
  (
    n694,
    n183
  );


  not
  g587
  (
    n965,
    n532
  );


  buf
  g588
  (
    n630,
    n240
  );


  not
  g589
  (
    n672,
    n157
  );


  buf
  g590
  (
    n804,
    n422
  );


  not
  g591
  (
    n715,
    n544
  );


  buf
  g592
  (
    n949,
    n412
  );


  buf
  g593
  (
    n807,
    n529
  );


  not
  g594
  (
    n1057,
    n176
  );


  buf
  g595
  (
    n654,
    n314
  );


  buf
  g596
  (
    n972,
    n342
  );


  buf
  g597
  (
    n812,
    n331
  );


  buf
  g598
  (
    n1175,
    n239
  );


  not
  g599
  (
    n960,
    n571
  );


  not
  g600
  (
    n779,
    n567
  );


  not
  g601
  (
    n612,
    n476
  );


  buf
  g602
  (
    n1031,
    n300
  );


  not
  g603
  (
    n943,
    n432
  );


  not
  g604
  (
    n725,
    n405
  );


  buf
  g605
  (
    n938,
    n161
  );


  buf
  g606
  (
    n1143,
    n370
  );


  not
  g607
  (
    n1086,
    n397
  );


  buf
  g608
  (
    n1145,
    n426
  );


  buf
  g609
  (
    n1046,
    n393
  );


  buf
  g610
  (
    n936,
    n155
  );


  buf
  g611
  (
    n1197,
    n227
  );


  not
  g612
  (
    n822,
    n210
  );


  buf
  g613
  (
    n825,
    n263
  );


  not
  g614
  (
    n1189,
    n344
  );


  not
  g615
  (
    n1111,
    n528
  );


  not
  g616
  (
    n625,
    n542
  );


  not
  g617
  (
    n728,
    n216
  );


  buf
  g618
  (
    n1093,
    n434
  );


  not
  g619
  (
    KeyWire_0_1,
    n315
  );


  buf
  g620
  (
    n1157,
    n482
  );


  buf
  g621
  (
    n1094,
    n369
  );


  buf
  g622
  (
    n865,
    n518
  );


  not
  g623
  (
    n977,
    n176
  );


  not
  g624
  (
    n813,
    n295
  );


  not
  g625
  (
    n787,
    n181
  );


  buf
  g626
  (
    n1014,
    n451
  );


  not
  g627
  (
    n792,
    n473
  );


  not
  g628
  (
    n1098,
    n301
  );


  not
  g629
  (
    n1121,
    n296
  );


  not
  g630
  (
    n862,
    n269
  );


  not
  g631
  (
    KeyWire_0_13,
    n358
  );


  buf
  g632
  (
    n1119,
    n199
  );


  not
  g633
  (
    n799,
    n232
  );


  buf
  g634
  (
    n986,
    n170
  );


  buf
  g635
  (
    n1202,
    n376
  );


  buf
  g636
  (
    n864,
    n522
  );


  not
  g637
  (
    n629,
    n580
  );


  buf
  g638
  (
    n1092,
    n206
  );


  not
  g639
  (
    n662,
    n389
  );


  buf
  g640
  (
    n1015,
    n568
  );


  buf
  g641
  (
    n942,
    n307
  );


  not
  g642
  (
    n719,
    n248
  );


  buf
  g643
  (
    n782,
    n512
  );


  not
  g644
  (
    n789,
    n307
  );


  buf
  g645
  (
    n1068,
    n430
  );


  not
  g646
  (
    n1196,
    n521
  );


  not
  g647
  (
    n895,
    n506
  );


  not
  g648
  (
    n985,
    n414
  );


  buf
  g649
  (
    n772,
    n238
  );


  not
  g650
  (
    n994,
    n359
  );


  buf
  g651
  (
    n683,
    n509
  );


  not
  g652
  (
    n912,
    n510
  );


  buf
  g653
  (
    n1027,
    n198
  );


  not
  g654
  (
    n1091,
    n303
  );


  not
  g655
  (
    n622,
    n548
  );


  not
  g656
  (
    n899,
    n229
  );


  buf
  g657
  (
    n1076,
    n437
  );


  buf
  g658
  (
    n1186,
    n465
  );


  buf
  g659
  (
    n1019,
    n257
  );


  not
  g660
  (
    n717,
    n500
  );


  not
  g661
  (
    n671,
    n454
  );


  not
  g662
  (
    n785,
    n282
  );


  not
  g663
  (
    n661,
    n447
  );


  buf
  g664
  (
    n722,
    n278
  );


  buf
  g665
  (
    n742,
    n393
  );


  buf
  g666
  (
    n1142,
    n197
  );


  not
  g667
  (
    n729,
    n542
  );


  not
  g668
  (
    n983,
    n338
  );


  buf
  g669
  (
    n664,
    n218
  );


  not
  g670
  (
    n1132,
    n434
  );


  not
  g671
  (
    n699,
    n318
  );


  not
  g672
  (
    n823,
    n582
  );


  not
  g673
  (
    n831,
    n341
  );


  not
  g674
  (
    n993,
    n404
  );


  not
  g675
  (
    n829,
    n447
  );


  not
  g676
  (
    n790,
    n353
  );


  not
  g677
  (
    n1165,
    n177
  );


  not
  g678
  (
    n1110,
    n240
  );


  buf
  g679
  (
    n933,
    n293
  );


  not
  g680
  (
    n866,
    n567
  );


  not
  g681
  (
    n875,
    n446
  );


  not
  g682
  (
    n1122,
    n445
  );


  not
  g683
  (
    n709,
    n335
  );


  buf
  g684
  (
    n1047,
    n280
  );


  not
  g685
  (
    n1208,
    n503
  );


  not
  g686
  (
    n843,
    n169
  );


  buf
  g687
  (
    n1069,
    n427
  );


  not
  g688
  (
    n735,
    n412
  );


  buf
  g689
  (
    n665,
    n460
  );


  not
  g690
  (
    n844,
    n347
  );


  not
  g691
  (
    n1127,
    n151
  );


  not
  g692
  (
    n973,
    n305
  );


  buf
  g693
  (
    n1151,
    n492
  );


  not
  g694
  (
    KeyWire_0_5,
    n487
  );


  buf
  g695
  (
    n1077,
    n276
  );


  not
  g696
  (
    n1003,
    n259
  );


  buf
  g697
  (
    n774,
    n214
  );


  buf
  g698
  (
    n1037,
    n227
  );


  buf
  g699
  (
    n915,
    n180
  );


  not
  g700
  (
    n921,
    n298
  );


  buf
  g701
  (
    n1039,
    n478
  );


  buf
  g702
  (
    n712,
    n549
  );


  not
  g703
  (
    n763,
    n476
  );


  buf
  g704
  (
    n889,
    n202
  );


  buf
  g705
  (
    n833,
    n529
  );


  buf
  g706
  (
    n777,
    n550
  );


  not
  g707
  (
    n1169,
    n567
  );


  buf
  g708
  (
    n966,
    n271
  );


  not
  g709
  (
    n1007,
    n484
  );


  not
  g710
  (
    n940,
    n288
  );


  not
  g711
  (
    n1080,
    n442
  );


  buf
  g712
  (
    n801,
    n252
  );


  buf
  g713
  (
    n1156,
    n300
  );


  buf
  g714
  (
    n1041,
    n569
  );


  not
  g715
  (
    n981,
    n501
  );


  buf
  g716
  (
    n1192,
    n534
  );


  buf
  g717
  (
    n743,
    n523
  );


  not
  g718
  (
    n1009,
    n500
  );


  not
  g719
  (
    n882,
    n208
  );


  not
  g720
  (
    n1067,
    n252
  );


  buf
  g721
  (
    n759,
    n455
  );


  buf
  g722
  (
    n702,
    n408
  );


  buf
  g723
  (
    n1082,
    n260
  );


  not
  g724
  (
    n828,
    n266
  );


  buf
  g725
  (
    n1190,
    n264
  );


  not
  g726
  (
    n618,
    n430
  );


  not
  g727
  (
    n818,
    n492
  );


  not
  g728
  (
    n928,
    n251
  );


  not
  g729
  (
    n1164,
    n514
  );


  buf
  g730
  (
    n1021,
    n179
  );


  buf
  g731
  (
    n927,
    n375
  );


  buf
  g732
  (
    n892,
    n207
  );


  buf
  g733
  (
    n1062,
    n251
  );


  not
  g734
  (
    n860,
    n573
  );


  buf
  g735
  (
    n810,
    n336
  );


  buf
  g736
  (
    n1066,
    n243
  );


  buf
  g737
  (
    n614,
    n283
  );


  buf
  g738
  (
    n1084,
    n205
  );


  not
  g739
  (
    n1171,
    n280
  );


  buf
  g740
  (
    n1089,
    n343
  );


  not
  g741
  (
    n1065,
    n236
  );


  buf
  g742
  (
    n998,
    n405
  );


  buf
  g743
  (
    n1042,
    n333
  );


  not
  g744
  (
    n677,
    n326
  );


  buf
  g745
  (
    n929,
    n583
  );


  buf
  g746
  (
    n1123,
    n506
  );


  buf
  g747
  (
    n765,
    n565
  );


  not
  g748
  (
    n624,
    n357
  );


  not
  g749
  (
    n623,
    n270
  );


  buf
  g750
  (
    n1207,
    n444
  );


  not
  g751
  (
    n633,
    n233
  );


  not
  g752
  (
    n658,
    n533
  );


  not
  g753
  (
    n1136,
    n319
  );


  buf
  g754
  (
    n1180,
    n462
  );


  not
  g755
  (
    n857,
    n229
  );


  not
  g756
  (
    n989,
    n282
  );


  buf
  g757
  (
    n1187,
    n569
  );


  not
  g758
  (
    n746,
    n443
  );


  not
  g759
  (
    n1061,
    n416
  );


  buf
  g760
  (
    n838,
    n240
  );


  not
  g761
  (
    n1166,
    n231
  );


  not
  g762
  (
    n754,
    n382
  );


  buf
  g763
  (
    n649,
    n479
  );


  not
  g764
  (
    n737,
    n507
  );


  buf
  g765
  (
    n903,
    n194
  );


  buf
  g766
  (
    n657,
    n199
  );


  not
  g767
  (
    n1144,
    n152
  );


  buf
  g768
  (
    n1102,
    n292
  );


  buf
  g769
  (
    n1135,
    n486
  );


  not
  g770
  (
    n1001,
    n577
  );


  buf
  g771
  (
    n888,
    n438
  );


  not
  g772
  (
    n755,
    n356
  );


  not
  g773
  (
    n736,
    n203
  );


  not
  g774
  (
    n617,
    n272
  );


  not
  g775
  (
    n1035,
    n552
  );


  not
  g776
  (
    n837,
    n446
  );


  buf
  g777
  (
    n1058,
    n285
  );


  buf
  g778
  (
    n1017,
    n540
  );


  buf
  g779
  (
    n934,
    n225
  );


  not
  g780
  (
    n637,
    n537
  );


  buf
  g781
  (
    n747,
    n281
  );


  buf
  g782
  (
    n1056,
    n260
  );


  not
  g783
  (
    n780,
    n560
  );


  not
  g784
  (
    n1181,
    n489
  );


  not
  g785
  (
    n879,
    n414
  );


  buf
  g786
  (
    n668,
    n489
  );


  buf
  g787
  (
    n1200,
    n477
  );


  buf
  g788
  (
    n853,
    n236
  );


  buf
  g789
  (
    n731,
    n559
  );


  buf
  g790
  (
    n920,
    n297
  );


  buf
  g791
  (
    n647,
    n365
  );


  not
  g792
  (
    n845,
    n251
  );


  nor
  g793
  (
    n886,
    n399,
    n206
  );


  and
  g794
  (
    n734,
    n510,
    n164,
    n524,
    n185
  );


  or
  g795
  (
    n867,
    n431,
    n192,
    n540,
    n188
  );


  nand
  g796
  (
    n773,
    n288,
    n381,
    n585,
    n531
  );


  nand
  g797
  (
    n1115,
    n294,
    n196,
    n343,
    n501
  );


  or
  g798
  (
    n877,
    n198,
    n281,
    n394,
    n494
  );


  and
  g799
  (
    n1126,
    n480,
    n329,
    n210,
    n452
  );


  xnor
  g800
  (
    n659,
    n453,
    n524,
    n420,
    n476
  );


  and
  g801
  (
    n643,
    n262,
    n321,
    n375,
    n473
  );


  nor
  g802
  (
    n800,
    n581,
    n228,
    n432,
    n213
  );


  xor
  g803
  (
    n996,
    n219,
    n210,
    n545,
    n580
  );


  nand
  g804
  (
    n766,
    n340,
    n362,
    n287,
    n415
  );


  xor
  g805
  (
    n863,
    n244,
    n502,
    n354,
    n451
  );


  nor
  g806
  (
    n655,
    n461,
    n221,
    n353,
    n556
  );


  xnor
  g807
  (
    n1063,
    n179,
    n522,
    n363,
    n266
  );


  nor
  g808
  (
    n1000,
    n369,
    n457,
    n490,
    n422
  );


  nand
  g809
  (
    n846,
    n354,
    n396,
    n189,
    n565
  );


  and
  g810
  (
    n1182,
    n494,
    n515,
    n191,
    n470
  );


  nand
  g811
  (
    n1124,
    n380,
    n189,
    n361,
    n509
  );


  nor
  g812
  (
    n1020,
    n300,
    n234,
    n173,
    n155
  );


  or
  g813
  (
    n1118,
    n293,
    n298,
    n580,
    n505
  );


  and
  g814
  (
    n914,
    n474,
    n223,
    n242,
    n567
  );


  nand
  g815
  (
    n1194,
    n531,
    n161,
    n416,
    n202
  );


  xnor
  g816
  (
    n1051,
    n563,
    n273,
    n546,
    n484
  );


  nand
  g817
  (
    n1204,
    n505,
    n422,
    n371,
    n513
  );


  nor
  g818
  (
    n1198,
    n417,
    n286,
    n231,
    n281
  );


  xnor
  g819
  (
    n945,
    n401,
    n452,
    n442,
    n469
  );


  xor
  g820
  (
    n1044,
    n344,
    n549,
    n299,
    n311
  );


  and
  g821
  (
    n1054,
    n463,
    n413,
    n338,
    n398
  );


  and
  g822
  (
    n703,
    n284,
    n517,
    n370,
    n453
  );


  and
  g823
  (
    n835,
    n452,
    n508,
    n375,
    n298
  );


  xor
  g824
  (
    n648,
    n312,
    n203,
    n409,
    n263
  );


  xor
  g825
  (
    n701,
    n458,
    n499,
    n204,
    n554
  );


  xnor
  g826
  (
    n1173,
    n277,
    n584,
    n376,
    n338
  );


  xor
  g827
  (
    n695,
    n318,
    n533,
    n483,
    n249
  );


  and
  g828
  (
    n707,
    n434,
    n450,
    n332,
    n419
  );


  and
  g829
  (
    n721,
    n281,
    n518,
    n522,
    n165
  );


  or
  g830
  (
    n1026,
    n520,
    n345,
    n435,
    n402
  );


  and
  g831
  (
    n1140,
    n171,
    n349,
    n385,
    n231
  );


  nor
  g832
  (
    n871,
    n274,
    n557,
    n168,
    n214
  );


  xnor
  g833
  (
    n689,
    n291,
    n421,
    n249,
    n223
  );


  nor
  g834
  (
    n840,
    n519,
    n216,
    n475,
    n514
  );


  nor
  g835
  (
    n1012,
    n259,
    n272,
    n196,
    n587
  );


  nor
  g836
  (
    n1087,
    n577,
    n484,
    n256,
    n497
  );


  xnor
  g837
  (
    n1013,
    n382,
    n278,
    n202,
    n189
  );


  and
  g838
  (
    n770,
    n200,
    n584,
    n499,
    n481
  );


  xnor
  g839
  (
    n1147,
    n423,
    n357,
    n400,
    n297
  );


  and
  g840
  (
    n724,
    n209,
    n246,
    n416,
    n251
  );


  xor
  g841
  (
    n900,
    n195,
    n553,
    n172,
    n520
  );


  nand
  g842
  (
    n1141,
    n433,
    n398,
    n573,
    n204
  );


  or
  g843
  (
    n786,
    n157,
    n536,
    n527,
    n288
  );


  nand
  g844
  (
    n1095,
    n191,
    n498,
    n196,
    n379
  );


  xnor
  g845
  (
    n1150,
    n469,
    n410,
    n153,
    n400
  );


  and
  g846
  (
    n852,
    n513,
    n468,
    n416,
    n174
  );


  or
  g847
  (
    n1158,
    n272,
    n247,
    n299,
    n384
  );


  xnor
  g848
  (
    n941,
    n589,
    n271,
    n550,
    n202
  );


  nand
  g849
  (
    KeyWire_0_20,
    n472,
    n566,
    n491,
    n164
  );


  nand
  g850
  (
    n788,
    n304,
    n467,
    n200,
    n343
  );


  nor
  g851
  (
    n656,
    n530,
    n498,
    n529,
    n156
  );


  xor
  g852
  (
    n854,
    n375,
    n155,
    n323,
    n366
  );


  nor
  g853
  (
    n741,
    n571,
    n205,
    n426,
    n369
  );


  xnor
  g854
  (
    n758,
    n468,
    n297,
    n233,
    n160
  );


  xor
  g855
  (
    n1163,
    n462,
    n212,
    n377,
    n511
  );


  nor
  g856
  (
    n1139,
    n439,
    n194,
    n319,
    n470
  );


  xor
  g857
  (
    n1078,
    n439,
    n433,
    n229,
    n444
  );


  xnor
  g858
  (
    n760,
    n192,
    n483,
    n534,
    n259
  );


  and
  g859
  (
    n883,
    n483,
    n448,
    n586,
    n522
  );


  xor
  g860
  (
    n1018,
    n579,
    n187,
    n256,
    n539
  );


  and
  g861
  (
    n1199,
    n427,
    n527,
    n431,
    n274
  );


  nand
  g862
  (
    n1206,
    n431,
    n351,
    n253,
    n188
  );


  or
  g863
  (
    n1130,
    n215,
    n191,
    n491,
    n562
  );


  and
  g864
  (
    n628,
    n405,
    n429,
    n512,
    n265
  );


  xnor
  g865
  (
    n1100,
    n547,
    n322,
    n504,
    n175
  );


  nor
  g866
  (
    n733,
    n371,
    n334,
    n220,
    n542
  );


  and
  g867
  (
    n1195,
    n560,
    n572,
    n564,
    n383
  );


  and
  g868
  (
    n1079,
    n334,
    n327,
    n529,
    n520
  );


  nand
  g869
  (
    n874,
    n473,
    n318,
    n256,
    n224
  );


  xor
  g870
  (
    n1081,
    n538,
    n488,
    n325,
    n589
  );


  or
  g871
  (
    n615,
    n219,
    n286,
    n287
  );


  or
  g872
  (
    n693,
    n493,
    n238,
    n402,
    n359
  );


  xnor
  g873
  (
    n902,
    n470,
    n185,
    n315,
    n590
  );


  nand
  g874
  (
    n894,
    n386,
    n311,
    n252,
    n339
  );


  nor
  g875
  (
    n1153,
    n500,
    n584,
    n156,
    n352
  );


  xor
  g876
  (
    n607,
    n425,
    n335,
    n365,
    n377
  );


  nor
  g877
  (
    n1016,
    n405,
    n397,
    n222,
    n536
  );


  nand
  g878
  (
    n764,
    n242,
    n582,
    n197,
    n404
  );


  nor
  g879
  (
    n716,
    n539,
    n349,
    n581,
    n569
  );


  or
  g880
  (
    n1179,
    n548,
    n583,
    n559,
    n272
  );


  xnor
  g881
  (
    n911,
    n154,
    n207,
    n555,
    n220
  );


  xnor
  g882
  (
    n1154,
    n336,
    n564,
    n316,
    n364
  );


  xnor
  g883
  (
    n963,
    n492,
    n230,
    n214,
    n295
  );


  nor
  g884
  (
    n969,
    n238,
    n574,
    n373,
    n227
  );


  and
  g885
  (
    n1129,
    n383,
    n217,
    n245,
    n151
  );


  nand
  g886
  (
    n982,
    n239,
    n249,
    n330,
    n541
  );


  nor
  g887
  (
    n904,
    n556,
    n362,
    n544,
    n366
  );


  xnor
  g888
  (
    n1148,
    n194,
    n561,
    n466,
    n311
  );


  xnor
  g889
  (
    n1075,
    n178,
    n203,
    n160,
    n523
  );


  nand
  g890
  (
    n901,
    n226,
    n451,
    n523,
    n279
  );


  xor
  g891
  (
    n1170,
    n367,
    n248,
    n555,
    n415
  );


  nand
  g892
  (
    n1193,
    n515,
    n496,
    n557,
    n406
  );


  and
  g893
  (
    n1045,
    n410,
    n208,
    n252,
    n508
  );


  xor
  g894
  (
    n1088,
    n583,
    n437,
    n380,
    n531
  );


  nor
  g895
  (
    n1025,
    n544,
    n366,
    n159,
    n515
  );


  or
  g896
  (
    n1083,
    n437,
    n524,
    n487,
    n302
  );


  xor
  g897
  (
    n896,
    n413,
    n512,
    n515,
    n417
  );


  nand
  g898
  (
    n700,
    n385,
    n578,
    n574,
    n439
  );


  nor
  g899
  (
    n1073,
    n224,
    n517,
    n232,
    n331
  );


  xnor
  g900
  (
    n682,
    n582,
    n392,
    n355,
    n363
  );


  xnor
  g901
  (
    n727,
    n241,
    n373,
    n590,
    n419
  );


  xor
  g902
  (
    n1024,
    n455,
    n166,
    n519,
    n450
  );


  xor
  g903
  (
    n1131,
    n153,
    n424,
    n503,
    n390
  );


  nand
  g904
  (
    n820,
    n575,
    n367,
    n278,
    n236
  );


  and
  g905
  (
    n832,
    n430,
    n395,
    n558,
    n468
  );


  and
  g906
  (
    n819,
    n434,
    n408,
    n374,
    n320
  );


  xor
  g907
  (
    n930,
    n161,
    n336,
    n339,
    n332
  );


  nor
  g908
  (
    n891,
    n376,
    n365,
    n438,
    n441
  );


  and
  g909
  (
    n626,
    n291,
    n495,
    n237,
    n498
  );


  xor
  g910
  (
    n681,
    n328,
    n406,
    n486,
    n351
  );


  xor
  g911
  (
    n881,
    n299,
    n383,
    n449,
    n408
  );


  nand
  g912
  (
    n980,
    n330,
    n289,
    n561,
    n356
  );


  nand
  g913
  (
    n954,
    n244,
    n233,
    n570,
    n586
  );


  nor
  g914
  (
    n1176,
    n423,
    n407,
    n526,
    n555
  );


  and
  g915
  (
    n893,
    n279,
    n578,
    n463,
    n406
  );


  and
  g916
  (
    n872,
    n175,
    n178,
    n543,
    n271
  );


  xnor
  g917
  (
    n984,
    n290,
    n508,
    n160,
    n425
  );


  xnor
  g918
  (
    n1072,
    n577,
    n355,
    n563,
    n293
  );


  xor
  g919
  (
    n1104,
    n225,
    n505,
    n244,
    n482
  );


  xor
  g920
  (
    n1034,
    n307,
    n554,
    n190,
    n558
  );


  and
  g921
  (
    n687,
    n216,
    n290,
    n459,
    n324
  );


  nand
  g922
  (
    n811,
    n228,
    n358,
    n156,
    n456
  );


  xnor
  g923
  (
    n710,
    n329,
    n525,
    n456,
    n507
  );


  xor
  g924
  (
    n690,
    n328,
    n310,
    n196,
    n319
  );


  xnor
  g925
  (
    n691,
    n180,
    n461,
    n551,
    n267
  );


  nand
  g926
  (
    n723,
    n509,
    n207,
    n296,
    n471
  );


  xnor
  g927
  (
    n791,
    n360,
    n237,
    n164,
    n350
  );


  xor
  g928
  (
    n1152,
    n293,
    n474,
    n564,
    n580
  );


  or
  g929
  (
    n611,
    n491,
    n277,
    n377,
    n288
  );


  xnor
  g930
  (
    n919,
    n548,
    n453,
    n286,
    n415
  );


  or
  g931
  (
    n1090,
    n438,
    n257,
    n187,
    n201
  );


  xor
  g932
  (
    n776,
    n513,
    n332,
    n168,
    n258
  );


  and
  g933
  (
    n923,
    n395,
    n365,
    n224,
    n575
  );


  nor
  g934
  (
    n609,
    n541,
    n313,
    n429,
    n532
  );


  xor
  g935
  (
    n610,
    n376,
    n205,
    n280,
    n181
  );


  nand
  g936
  (
    n842,
    n389,
    n527,
    n220,
    n587
  );


  nor
  g937
  (
    n909,
    n406,
    n423,
    n217,
    n464
  );


  and
  g938
  (
    n1030,
    n560,
    n464,
    n559,
    n270
  );


  nor
  g939
  (
    n848,
    n485,
    n323,
    n569,
    n183
  );


  or
  g940
  (
    n834,
    n158,
    n255,
    n558,
    n519
  );


  nand
  g941
  (
    n638,
    n353,
    n294,
    n305,
    n276
  );


  xnor
  g942
  (
    n935,
    n374,
    n358,
    n537,
    n175
  );


  nor
  g943
  (
    n1114,
    n474,
    n304,
    n470,
    n467
  );


  and
  g944
  (
    n1097,
    n324,
    n152,
    n459,
    n518
  );


  xnor
  g945
  (
    n667,
    n463,
    n361,
    n379,
    n250
  );


  xnor
  g946
  (
    n713,
    n492,
    n387,
    n465,
    n477
  );


  nand
  g947
  (
    KeyWire_0_10,
    n423,
    n426,
    n261,
    n290
  );


  xnor
  g948
  (
    n1146,
    n305,
    n414,
    n494,
    n478
  );


  nand
  g949
  (
    n1162,
    n263,
    n426,
    n186,
    n322
  );


  nand
  g950
  (
    n898,
    n479,
    n430,
    n349,
    n433
  );


  xor
  g951
  (
    n1008,
    n306,
    n381,
    n195,
    n404
  );


  nand
  g952
  (
    n917,
    n472,
    n495,
    n524,
    n286
  );


  xnor
  g953
  (
    n952,
    n184,
    n248,
    n395,
    n566
  );


  xnor
  g954
  (
    n913,
    n538,
    n561,
    n462,
    n579
  );


  and
  g955
  (
    n830,
    n282,
    n491,
    n409,
    n471
  );


  and
  g956
  (
    KeyWire_0_14,
    n250,
    n418,
    n234,
    n242
  );


  xnor
  g957
  (
    n1106,
    n466,
    n581,
    n314,
    n323
  );


  nand
  g958
  (
    n711,
    n528,
    n389,
    n213,
    n367
  );


  or
  g959
  (
    n793,
    n245,
    n319,
    n277,
    n306
  );


  or
  g960
  (
    n718,
    n417,
    n450,
    n468,
    n228
  );


  nand
  g961
  (
    n696,
    n315,
    n158,
    n485,
    n582
  );


  or
  g962
  (
    n680,
    n458,
    n309,
    n549,
    n246
  );


  and
  g963
  (
    n880,
    n521,
    n254,
    n475,
    n186
  );


  xor
  g964
  (
    n856,
    n151,
    n164,
    n526,
    n516
  );


  xor
  g965
  (
    n1002,
    n528,
    n400,
    n457,
    n176
  );


  and
  g966
  (
    n1085,
    n363,
    n284,
    n521,
    n461
  );


  xnor
  g967
  (
    n1107,
    n479,
    n189,
    n506,
    n182
  );


  xor
  g968
  (
    n1191,
    n200,
    n453,
    n208,
    n314
  );


  nand
  g969
  (
    n836,
    n199,
    n374,
    n588,
    n479
  );


  xnor
  g970
  (
    n1161,
    n271,
    n497,
    n345,
    n249
  );


  and
  g971
  (
    n962,
    n465,
    n253,
    n225,
    n193
  );


  nand
  g972
  (
    n606,
    n234,
    n409,
    n176,
    n428
  );


  xor
  g973
  (
    n1043,
    n402,
    n346,
    n589,
    n354
  );


  or
  g974
  (
    n878,
    n481,
    n412,
    n151,
    n358
  );


  xor
  g975
  (
    n1050,
    n195,
    n181,
    n243,
    n586
  );


  nor
  g976
  (
    n805,
    n463,
    n279,
    n420,
    n337
  );


  xor
  g977
  (
    n794,
    n504,
    n184,
    n574,
    n584
  );


  or
  g978
  (
    n931,
    n480,
    n562,
    n362,
    n568
  );


  or
  g979
  (
    n714,
    n239,
    n273,
    n292,
    n552
  );


  or
  g980
  (
    n1134,
    n485,
    n565,
    n231,
    n209
  );


  xor
  g981
  (
    n744,
    n410,
    n435,
    n247,
    n359
  );


  xnor
  g982
  (
    n1120,
    n481,
    n454,
    n540,
    n294
  );


  xnor
  g983
  (
    n868,
    n562,
    n344,
    n422,
    n357
  );


  xor
  g984
  (
    n650,
    n425,
    n586,
    n399,
    n246
  );


  xor
  g985
  (
    n958,
    n194,
    n533,
    n471,
    n264
  );


  xnor
  g986
  (
    n1074,
    n381,
    n226,
    n357,
    n532
  );


  xor
  g987
  (
    n1112,
    n210,
    n356,
    n448,
    n544
  );


  nand
  g988
  (
    n951,
    n283,
    n483,
    n509,
    n217
  );


  and
  g989
  (
    n1070,
    n333,
    n559,
    n335,
    n162
  );


  nand
  g990
  (
    n639,
    n333,
    n180,
    n340,
    n488
  );


  or
  g991
  (
    n808,
    n380,
    n525,
    n364,
    n446
  );


  xor
  g992
  (
    n1125,
    n431,
    n502,
    n420,
    n153
  );


  and
  g993
  (
    n1029,
    n257,
    n316,
    n466,
    n255
  );


  xnor
  g994
  (
    n975,
    n304,
    n258,
    n417,
    n467
  );


  nand
  g995
  (
    n817,
    n444,
    n368,
    n289,
    n570
  );


  nor
  g996
  (
    n771,
    n551,
    n265,
    n364,
    n401
  );


  or
  g997
  (
    n991,
    n241,
    n501,
    n352,
    n361
  );


  and
  g998
  (
    n905,
    n192,
    n436,
    n211,
    n391
  );


  xor
  g999
  (
    n839,
    n269,
    n330,
    n258,
    n278
  );


  xor
  g1000
  (
    n686,
    n173,
    n294,
    n526,
    n383
  );


  and
  g1001
  (
    n974,
    n263,
    n152,
    n158,
    n270
  );


  nor
  g1002
  (
    n803,
    n334,
    n308,
    n178,
    n457
  );


  and
  g1003
  (
    n873,
    n394,
    n250,
    n498,
    n472
  );


  and
  g1004
  (
    n1005,
    n439,
    n469,
    n350,
    n407
  );


  nor
  g1005
  (
    n698,
    n428,
    n229,
    n191,
    n351
  );


  nand
  g1006
  (
    n704,
    n440,
    n480,
    n268,
    n456
  );


  nand
  g1007
  (
    n992,
    n212,
    n534,
    n308,
    n327
  );


  or
  g1008
  (
    n651,
    n518,
    n578,
    n579,
    n497
  );


  and
  g1009
  (
    n979,
    n548,
    n440,
    n386,
    n204
  );


  or
  g1010
  (
    n784,
    n508,
    n543,
    n413,
    n485
  );


  nand
  g1011
  (
    n956,
    n552,
    n420,
    n419,
    n285
  );


  or
  g1012
  (
    n673,
    n198,
    n186,
    n235,
    n462
  );


  nor
  g1013
  (
    n769,
    n571,
    n530,
    n244,
    n389
  );


  nor
  g1014
  (
    n1006,
    n265,
    n348,
    n345,
    n347
  );


  nor
  g1015
  (
    n738,
    n432,
    n282,
    n177,
    n306
  );


  nand
  g1016
  (
    n1159,
    n222,
    n190,
    n557,
    n484
  );


  nand
  g1017
  (
    n1155,
    n572,
    n395,
    n269,
    n260
  );


  or
  g1018
  (
    n1103,
    n182,
    n530,
    n538,
    n190
  );


  nand
  g1019
  (
    n1032,
    n437,
    n482,
    n216,
    n566
  );


  or
  g1020
  (
    n762,
    n292,
    n408,
    n372,
    n349
  );


  nand
  g1021
  (
    n887,
    n317,
    n500,
    n511,
    n347
  );


  and
  g1022
  (
    n660,
    n585,
    n407,
    n265,
    n193
  );


  and
  g1023
  (
    n924,
    n505,
    n239,
    n174,
    n267
  );


  xnor
  g1024
  (
    n692,
    n477,
    n428,
    n547,
    n342
  );


  xnor
  g1025
  (
    n910,
    n455,
    n385,
    n326,
    n343
  );


  xor
  g1026
  (
    n1174,
    n172,
    n545,
    n460,
    n348
  );


  xor
  g1027
  (
    n1117,
    n308,
    n154,
    n541,
    n254
  );


  xnor
  g1028
  (
    n953,
    n155,
    n199,
    n458,
    n525
  );


  xnor
  g1029
  (
    n908,
    n413,
    n193,
    n321,
    n412
  );


  xor
  g1030
  (
    n674,
    n362,
    n543,
    n320,
    n386
  );


  xor
  g1031
  (
    n1183,
    n154,
    n316,
    n342,
    n445
  );


  xnor
  g1032
  (
    n652,
    n465,
    n401,
    n556,
    n183
  );


  or
  g1033
  (
    n1023,
    n517,
    n346,
    n400,
    n261
  );


  xor
  g1034
  (
    n906,
    n486,
    n220,
    n308,
    n340
  );


  or
  g1035
  (
    n697,
    n409,
    n504,
    n364,
    n341
  );


  xor
  g1036
  (
    n645,
    n464,
    n527,
    n190,
    n327
  );


  and
  g1037
  (
    n961,
    n218,
    n335,
    n180,
    n555
  );


  nand
  g1038
  (
    n781,
    n378,
    n392,
    n275,
    n309
  );


  or
  g1039
  (
    n768,
    n171,
    n450,
    n168,
    n270
  );


  xnor
  g1040
  (
    n859,
    n336,
    n291,
    n328,
    n241
  );


  xnor
  g1041
  (
    n740,
    n443,
    n388,
    n246,
    n378
  );


  xor
  g1042
  (
    n775,
    n204,
    n573,
    n449,
    n234
  );


  or
  g1043
  (
    n897,
    n370,
    n328,
    n511,
    n228
  );


  and
  g1044
  (
    n641,
    n302,
    n330,
    n306,
    n211
  );


  xnor
  g1045
  (
    n970,
    n478,
    n553,
    n388,
    n387
  );


  nand
  g1046
  (
    n795,
    n394,
    n493,
    n230,
    n174
  );


  nor
  g1047
  (
    n644,
    n165,
    n535,
    n341,
    n554
  );


  and
  g1048
  (
    n1205,
    n323,
    n404,
    n326,
    n169
  );


  nor
  g1049
  (
    n922,
    n283,
    n222,
    n325,
    n277
  );


  xor
  g1050
  (
    KeyWire_0_18,
    n261,
    n564,
    n325,
    n377
  );


  nand
  g1051
  (
    n971,
    n301,
    n397,
    n511,
    n262
  );


  nor
  g1052
  (
    n850,
    n254,
    n215,
    n267,
    n585
  );


  or
  g1053
  (
    n1116,
    n275,
    n233,
    n161,
    n493
  );


  and
  g1054
  (
    n666,
    n445,
    n387,
    n502,
    n378
  );


  xor
  g1055
  (
    n739,
    n572,
    n496,
    n456,
    n170
  );


  or
  g1056
  (
    n730,
    n276,
    n291,
    n213,
    n198
  );


  nor
  g1057
  (
    n669,
    n570,
    n546,
    n585,
    n388
  );


  xor
  g1058
  (
    n884,
    n223,
    n253,
    n425,
    n188
  );


  nand
  g1059
  (
    n967,
    n563,
    n348,
    n391
  );


  xnor
  g1060
  (
    n745,
    n241,
    n289,
    n540,
    n207
  );


  or
  g1061
  (
    n1053,
    n167,
    n440,
    n346,
    n539
  );


  xor
  g1062
  (
    n948,
    n177,
    n296,
    n488,
    n411
  );


  or
  g1063
  (
    n885,
    n170,
    n436,
    n458,
    n267
  );


  nand
  g1064
  (
    n926,
    n221,
    n497,
    n490,
    n165
  );


  or
  g1065
  (
    n1185,
    n562,
    n467,
    n274,
    n414
  );


  nand
  g1066
  (
    n1133,
    n301,
    n201,
    n184,
    n338
  );


  nand
  g1067
  (
    n990,
    n363,
    n523,
    n393,
    n379
  );


  and
  g1068
  (
    n1096,
    n452,
    n499,
    n588,
    n545
  );


  and
  g1069
  (
    n978,
    n576,
    n315,
    n379,
    n219
  );


  xor
  g1070
  (
    n1004,
    n519,
    n157,
    n359,
    n321
  );


  nor
  g1071
  (
    n670,
    n490,
    n565,
    n171,
    n314
  );


  xnor
  g1072
  (
    n916,
    n296,
    n494,
    n333,
    n197
  );


  nor
  g1073
  (
    n1059,
    n402,
    n378,
    n310,
    n538
  );


  and
  g1074
  (
    n705,
    n457,
    n429,
    n419,
    n427
  );


  xor
  g1075
  (
    n1052,
    n517,
    n424,
    n215,
    n481
  );


  nand
  g1076
  (
    n1033,
    n195,
    n313,
    n503,
    n512
  );


  xnor
  g1077
  (
    n802,
    n222,
    n536,
    n224,
    n399
  );


  xor
  g1078
  (
    n809,
    n464,
    n166,
    n275,
    n382
  );


  or
  g1079
  (
    n640,
    n285,
    n237,
    n167,
    n205
  );


  nor
  g1080
  (
    n678,
    n158,
    n185,
    n547,
    n475
  );


  xnor
  g1081
  (
    n706,
    n554,
    n455,
    n443,
    n242
  );


  xnor
  g1082
  (
    n987,
    n398,
    n546,
    n243,
    n171
  );


  xnor
  g1083
  (
    n635,
    n345,
    n211,
    n266,
    n297
  );


  and
  g1084
  (
    n1010,
    n570,
    n159,
    n182,
    n264
  );


  nand
  g1085
  (
    n870,
    n273,
    n264,
    n360,
    n206
  );


  xnor
  g1086
  (
    n995,
    n332,
    n516,
    n525,
    n556
  );


  or
  g1087
  (
    n1040,
    n240,
    n528,
    n329,
    n247
  );


  xor
  g1088
  (
    n907,
    n337,
    n436,
    n444,
    n360
  );


  nand
  g1089
  (
    n1101,
    n410,
    n433,
    n549,
    n460
  );


  nand
  g1090
  (
    n1178,
    n153,
    n445,
    n579,
    n572
  );


  nand
  g1091
  (
    n1203,
    n292,
    n156,
    n279,
    n447
  );


  nor
  g1092
  (
    n619,
    n290,
    n394,
    n302,
    n551
  );


  nor
  g1093
  (
    n847,
    n386,
    n174,
    n424,
    n262
  );


  xor
  g1094
  (
    n1036,
    n219,
    n318,
    n411,
    n163
  );


  xor
  g1095
  (
    n1177,
    n583,
    n411,
    n192,
    n435
  );


  nor
  g1096
  (
    n1113,
    n407,
    n551,
    n588,
    n347
  );


  and
  g1097
  (
    n767,
    n175,
    n232,
    n200,
    n371
  );


  xnor
  g1098
  (
    n821,
    n273,
    n532,
    n466,
    n392
  );


  nand
  g1099
  (
    n999,
    n428,
    n390,
    n317,
    n355
  );


  and
  g1100
  (
    n1188,
    n374,
    n557,
    n380,
    n443
  );


  nor
  g1101
  (
    n685,
    n535,
    n435,
    n206,
    n324
  );


  and
  g1102
  (
    n1048,
    n355,
    n534,
    n513,
    n209
  );


  xor
  g1103
  (
    n1184,
    n589,
    n521,
    n320,
    n475
  );


  nor
  g1104
  (
    n720,
    n440,
    n275,
    n561,
    n213
  );


  nor
  g1105
  (
    n750,
    n361,
    n568,
    n183,
    n403
  );


  nor
  g1106
  (
    n964,
    n312,
    n369,
    n448,
    n587
  );


  nor
  g1107
  (
    n1060,
    n469,
    n182,
    n184,
    n268
  );


  or
  g1108
  (
    n946,
    n218,
    n160,
    n163,
    n446
  );


  or
  g1109
  (
    n976,
    n179,
    n550,
    n367,
    n496
  );


  or
  g1110
  (
    n1149,
    n489,
    n162,
    n553,
    n325
  );


  xnor
  g1111
  (
    n798,
    n545,
    n181,
    n341,
    n372
  );


  or
  g1112
  (
    n1049,
    n170,
    n322,
    n346,
    n289
  );


  nor
  g1113
  (
    KeyWire_0_28,
    n354,
    n235,
    n208
  );


  nand
  g1114
  (
    n858,
    n339,
    n307,
    n178,
    n568
  );


  nand
  g1115
  (
    n997,
    n255,
    n403,
    n448,
    n460
  );


  xor
  g1116
  (
    n1167,
    n188,
    n166,
    n305,
    n186
  );


  or
  g1117
  (
    n1108,
    n421,
    n478,
    n230
  );


  nor
  g1118
  (
    n1038,
    n441,
    n162,
    n167,
    n218
  );


  or
  g1119
  (
    n621,
    n177,
    n387,
    n300,
    n516
  );


  nand
  g1120
  (
    n1011,
    n398,
    n451,
    n287,
    n432
  );


  xor
  g1121
  (
    n959,
    n301,
    n510,
    n496,
    n489
  );


  nor
  g1122
  (
    n1064,
    n342,
    n247,
    n310,
    n201
  );


  xor
  g1123
  (
    n1109,
    n552,
    n253,
    n243,
    n396
  );


  or
  g1124
  (
    n616,
    n322,
    n403,
    n576,
    n352
  );


  xnor
  g1125
  (
    n950,
    n261,
    n256,
    n223,
    n337
  );


  xnor
  g1126
  (
    n631,
    n159,
    n331,
    n526,
    n245
  );


  xor
  g1127
  (
    n1172,
    n575,
    n163,
    n504,
    n331
  );


  nor
  g1128
  (
    n749,
    n350,
    n179,
    n372,
    n324
  );


  nand
  g1129
  (
    n1137,
    n487,
    n499,
    n427,
    n262
  );


  and
  g1130
  (
    n1028,
    n514,
    n590,
    n248,
    n169
  );


  nand
  g1131
  (
    KeyWire_0_0,
    n510,
    n429,
    n547,
    n563
  );


  xnor
  g1132
  (
    n732,
    n360,
    n368,
    n424,
    n587
  );


  and
  g1133
  (
    n988,
    n217,
    n185,
    n397,
    n157
  );


  xor
  g1134
  (
    n636,
    n449,
    n312,
    n576,
    n472
  );


  xor
  g1135
  (
    n708,
    n284,
    n304,
    n373,
    n211
  );


  xnor
  g1136
  (
    n1022,
    n348,
    n172,
    n459,
    n418
  );


  nand
  g1137
  (
    n861,
    n373,
    n537,
    n166,
    n495
  );


  or
  g1138
  (
    n627,
    n317,
    n334,
    n411,
    n276
  );


  nand
  g1139
  (
    n761,
    n284,
    n447,
    n163,
    n536
  );


  nor
  g1140
  (
    n937,
    n382,
    n390,
    n329,
    n454
  );


  or
  g1141
  (
    n646,
    n493,
    n537,
    n441,
    n173
  );


  xor
  g1142
  (
    n679,
    n250,
    n482,
    n441,
    n590
  );


  xor
  g1143
  (
    n824,
    n574,
    n553,
    n280,
    n488
  );


  and
  g1144
  (
    n925,
    n560,
    n268,
    n558
  );


  and
  g1145
  (
    n663,
    n154,
    n302,
    n187,
    n312
  );


  nand
  g1146
  (
    n675,
    n477,
    n237,
    n368,
    n159
  );


  xor
  g1147
  (
    n757,
    n356,
    n167,
    n436,
    n442
  );


  and
  g1148
  (
    n632,
    n197,
    n507,
    n573,
    n371
  );


  xor
  g1149
  (
    n1055,
    n285,
    n303,
    n221,
    n226
  );


  nand
  g1150
  (
    n778,
    n353,
    n311,
    n215,
    n442
  );


  and
  g1151
  (
    n827,
    n388,
    n366,
    n546,
    n310
  );


  and
  g1152
  (
    n876,
    n514,
    n459,
    n381,
    n454
  );


  xor
  g1153
  (
    n642,
    n303,
    n384,
    n571,
    n449
  );


  xnor
  g1154
  (
    n751,
    n533,
    n201,
    n309,
    n209
  );


  xor
  g1155
  (
    n797,
    n260,
    n578,
    n227,
    n588
  );


  nor
  g1156
  (
    n1099,
    n351,
    n350,
    n535,
    n550
  );


  xnor
  g1157
  (
    n676,
    n221,
    n212,
    n162,
    n225
  );


  xnor
  g1158
  (
    n814,
    n309,
    n255,
    n269,
    n507
  );


  xnor
  g1159
  (
    n855,
    n298,
    n344,
    n531,
    n391
  );


  nor
  g1160
  (
    n620,
    n486,
    n476,
    n575,
    n187
  );


  nand
  g1161
  (
    n851,
    n165,
    n172,
    n370,
    n214
  );


  xnor
  g1162
  (
    n932,
    n480,
    n212,
    n235,
    n495
  );


  and
  g1163
  (
    n841,
    n473,
    n461,
    n266,
    n238
  );


  nor
  g1164
  (
    n688,
    n396,
    n317,
    n506,
    n321
  );


  nor
  g1165
  (
    n849,
    n295,
    n471,
    n339,
    n490
  );


  and
  g1166
  (
    n748,
    n501,
    n385,
    n168,
    n232
  );


  and
  g1167
  (
    n816,
    n173,
    n415,
    n576,
    n245
  );


  xnor
  g1168
  (
    n1071,
    n257,
    n487,
    n258,
    n274
  );


  nand
  g1169
  (
    n608,
    n193,
    n393,
    n503,
    n539
  );


  or
  g1170
  (
    n957,
    n169,
    n474,
    n327,
    n421
  );


  nor
  g1171
  (
    n1138,
    n320,
    n236,
    n372,
    n401
  );


  xor
  g1172
  (
    n753,
    n226,
    n384,
    n516,
    n421
  );


  xnor
  g1173
  (
    n1201,
    n152,
    n368,
    n203,
    n418
  );


  xnor
  g1174
  (
    n869,
    n313,
    n403,
    n303,
    n577
  );


  and
  g1175
  (
    n653,
    n384,
    n259,
    n295,
    n313
  );


  and
  g1176
  (
    n826,
    n438,
    n392,
    n337,
    n418
  );


  and
  g1177
  (
    n783,
    n535,
    n566,
    n390,
    n326
  );


  or
  g1178
  (
    n684,
    n502,
    n299,
    n530,
    n254
  );


  nor
  g1179
  (
    n1245,
    n745,
    n777,
    n716,
    n781
  );


  nand
  g1180
  (
    n1258,
    n763,
    n687,
    n718,
    n779
  );


  or
  g1181
  (
    n1257,
    n650,
    n695,
    n667,
    n608
  );


  and
  g1182
  (
    n1248,
    n646,
    n788,
    n797,
    n616
  );


  xnor
  g1183
  (
    n1246,
    n720,
    n782,
    n723,
    n800
  );


  xor
  g1184
  (
    n1237,
    n652,
    n784,
    n742,
    n673
  );


  nand
  g1185
  (
    n1213,
    n620,
    n713,
    n755,
    n666
  );


  nor
  g1186
  (
    n1252,
    n758,
    n632,
    n672,
    n705
  );


  xnor
  g1187
  (
    n1219,
    n661,
    n728,
    n792,
    n798
  );


  xnor
  g1188
  (
    n1253,
    n764,
    n760,
    n730,
    n736
  );


  or
  g1189
  (
    n1230,
    n765,
    n682,
    n756,
    n677
  );


  nand
  g1190
  (
    n1235,
    n701,
    n740,
    n729,
    n754
  );


  or
  g1191
  (
    n1211,
    n631,
    n702,
    n766,
    n612
  );


  nand
  g1192
  (
    n1215,
    n786,
    n645,
    n739,
    n611
  );


  nand
  g1193
  (
    n1225,
    n640,
    n649,
    n787,
    n796
  );


  nand
  g1194
  (
    n1254,
    n634,
    n618,
    n683,
    n783
  );


  and
  g1195
  (
    n1232,
    n628,
    n747,
    n735,
    n647
  );


  and
  g1196
  (
    n1249,
    n769,
    n700,
    n711,
    n717
  );


  xnor
  g1197
  (
    n1247,
    n746,
    n734,
    n703,
    n750
  );


  and
  g1198
  (
    n1231,
    n768,
    n693,
    n773,
    n657
  );


  nand
  g1199
  (
    n1227,
    n727,
    n725,
    n741,
    n653
  );


  and
  g1200
  (
    n1250,
    n708,
    n662,
    n780,
    n609
  );


  and
  g1201
  (
    n1241,
    n795,
    n655,
    n668,
    n676
  );


  nor
  g1202
  (
    n1214,
    n665,
    n675,
    n712,
    n680
  );


  nor
  g1203
  (
    n1210,
    n663,
    n791,
    n626,
    n644
  );


  xor
  g1204
  (
    n1242,
    n669,
    n651,
    n767,
    n721
  );


  nor
  g1205
  (
    n1223,
    n761,
    n733,
    n732,
    n776
  );


  nand
  g1206
  (
    n1212,
    n698,
    n689,
    n681,
    n793
  );


  nor
  g1207
  (
    n1236,
    n710,
    n694,
    n670,
    n751
  );


  xnor
  g1208
  (
    n1238,
    n629,
    n801,
    n744,
    n674
  );


  nor
  g1209
  (
    n1224,
    n759,
    n775,
    n637,
    n738
  );


  and
  g1210
  (
    n1259,
    n778,
    n656,
    n770,
    n774
  );


  and
  g1211
  (
    n1239,
    n762,
    n706,
    n686,
    n664
  );


  nand
  g1212
  (
    n1234,
    n639,
    n679,
    n642,
    n623
  );


  xor
  g1213
  (
    n1240,
    n684,
    n719,
    n614,
    n622
  );


  nand
  g1214
  (
    n1233,
    n799,
    n724,
    n749,
    n627
  );


  and
  g1215
  (
    n1244,
    n648,
    n804,
    n619,
    n621
  );


  nand
  g1216
  (
    n1218,
    n696,
    n633,
    n748,
    n726
  );


  xor
  g1217
  (
    n1243,
    n625,
    n707,
    n641,
    n722
  );


  nand
  g1218
  (
    n1222,
    n785,
    n636,
    n643,
    n638
  );


  xor
  g1219
  (
    n1216,
    n671,
    n803,
    n753,
    n692
  );


  nand
  g1220
  (
    n1220,
    n610,
    n624,
    n697,
    n678
  );


  xor
  g1221
  (
    n1255,
    n699,
    n772,
    n752,
    n607
  );


  xor
  g1222
  (
    n1226,
    n790,
    n660,
    n737,
    n613
  );


  and
  g1223
  (
    n1256,
    n794,
    n606,
    n743,
    n690
  );


  and
  g1224
  (
    n1217,
    n789,
    n617,
    n659,
    n658
  );


  xor
  g1225
  (
    n1229,
    n715,
    n654,
    n704,
    n802
  );


  nand
  g1226
  (
    n1251,
    n709,
    n771,
    n688,
    n691
  );


  xor
  g1227
  (
    n1228,
    n805,
    n685,
    n731,
    n757
  );


  xor
  g1228
  (
    n1221,
    n714,
    n635,
    n615,
    n630
  );


  and
  g1229
  (
    n1303,
    n1231,
    n811,
    n1240,
    n852
  );


  nor
  g1230
  (
    n1291,
    n819,
    n860,
    n854,
    n874
  );


  and
  g1231
  (
    n1298,
    n827,
    n930,
    n1232,
    n1229
  );


  and
  g1232
  (
    n1277,
    n917,
    n929,
    n833,
    n1247
  );


  xnor
  g1233
  (
    n1261,
    n935,
    n911,
    n1250,
    n876
  );


  nor
  g1234
  (
    n1294,
    n906,
    n1227,
    n925,
    n1222
  );


  nor
  g1235
  (
    n1283,
    n1246,
    n931,
    n888,
    n913
  );


  nand
  g1236
  (
    n1282,
    n864,
    n1235,
    n894,
    n812
  );


  nand
  g1237
  (
    n1295,
    n847,
    n937,
    n1217,
    n840
  );


  nand
  g1238
  (
    n1271,
    n901,
    n871,
    n845,
    n900
  );


  nor
  g1239
  (
    n1263,
    n1252,
    n1239,
    n869,
    n1244
  );


  nor
  g1240
  (
    n1262,
    n936,
    n934,
    n824,
    n835
  );


  xnor
  g1241
  (
    n1296,
    n1251,
    n831,
    n825,
    n868
  );


  or
  g1242
  (
    n1292,
    n870,
    n1221,
    n893,
    n1212
  );


  xor
  g1243
  (
    n1279,
    n928,
    n880,
    n818,
    n829
  );


  nor
  g1244
  (
    n1290,
    n909,
    n920,
    n883,
    n905
  );


  xor
  g1245
  (
    n1276,
    n821,
    n1218,
    n1233,
    n865
  );


  and
  g1246
  (
    KeyWire_0_31,
    n808,
    n866,
    n1228,
    n932
  );


  or
  g1247
  (
    n1260,
    n851,
    n927,
    n815,
    n806
  );


  and
  g1248
  (
    n1278,
    n1226,
    n907,
    n914,
    n918
  );


  xor
  g1249
  (
    n1281,
    n1249,
    n1236,
    n809,
    n841
  );


  xnor
  g1250
  (
    n1287,
    n890,
    n902,
    n889,
    n839
  );


  and
  g1251
  (
    n1266,
    n1211,
    n924,
    n842,
    n903
  );


  nand
  g1252
  (
    n1293,
    n910,
    n877,
    n887,
    n891
  );


  and
  g1253
  (
    n1289,
    n1253,
    n843,
    n1230,
    n850
  );


  xnor
  g1254
  (
    n1272,
    n861,
    n922,
    n1219,
    n1238
  );


  nand
  g1255
  (
    n1264,
    n892,
    n810,
    n1248,
    n1241
  );


  or
  g1256
  (
    n1270,
    n1242,
    n1213,
    n816,
    n830
  );


  nand
  g1257
  (
    n1267,
    n1210,
    n855,
    n933,
    n820
  );


  nor
  g1258
  (
    n1297,
    n838,
    n886,
    n1216,
    n919
  );


  and
  g1259
  (
    n1284,
    n828,
    n882,
    n858,
    n1215
  );


  and
  g1260
  (
    n1286,
    n875,
    n879,
    n898,
    n848
  );


  and
  g1261
  (
    n1300,
    n1214,
    n857,
    n896,
    n844
  );


  xnor
  g1262
  (
    n1274,
    n1234,
    n846,
    n859,
    n1225
  );


  xor
  g1263
  (
    n1302,
    n904,
    n908,
    n895,
    n834
  );


  nand
  g1264
  (
    n1301,
    n873,
    n826,
    n923,
    n817
  );


  nor
  g1265
  (
    n1280,
    n1237,
    n849,
    n823,
    n1220
  );


  or
  g1266
  (
    KeyWire_0_11,
    n1223,
    n807,
    n867,
    n814
  );


  and
  g1267
  (
    n1275,
    n862,
    n822,
    n832,
    n856
  );


  xnor
  g1268
  (
    n1265,
    n863,
    n884,
    n881,
    n1224
  );


  xor
  g1269
  (
    n1268,
    n921,
    n916,
    n878,
    n836
  );


  or
  g1270
  (
    n1299,
    n1243,
    n915,
    n912,
    n853
  );


  and
  g1271
  (
    n1288,
    n813,
    n872,
    n837,
    n885
  );


  or
  g1272
  (
    KeyWire_0_29,
    n897,
    n1245,
    n899,
    n926
  );


  xnor
  g1273
  (
    n1305,
    n938,
    n946,
    n1288
  );


  xnor
  g1274
  (
    n1307,
    n947,
    n1256,
    n941
  );


  and
  g1275
  (
    n1304,
    n1259,
    n945,
    n1255,
    n1290
  );


  nand
  g1276
  (
    n1308,
    n939,
    n940,
    n1287,
    n943
  );


  xnor
  g1277
  (
    n1306,
    n1258,
    n1257,
    n1291,
    n1286
  );


  xnor
  g1278
  (
    n1309,
    n942,
    n944,
    n1289,
    n1254
  );


  nand
  g1279
  (
    n1314,
    n952,
    n1309,
    n957,
    n1307
  );


  xnor
  g1280
  (
    n1316,
    n948,
    n1308,
    n959,
    n591
  );


  nand
  g1281
  (
    n1312,
    n960,
    n950,
    n1306,
    n1308
  );


  and
  g1282
  (
    n1317,
    n591,
    n953,
    n955,
    n961
  );


  or
  g1283
  (
    n1310,
    n1305,
    n591,
    n951,
    n592
  );


  xnor
  g1284
  (
    n1311,
    n1306,
    n1304,
    n954,
    n1309
  );


  and
  g1285
  (
    n1315,
    n591,
    n958,
    n949,
    n592
  );


  or
  g1286
  (
    n1313,
    n592,
    n956,
    n962,
    n1307
  );


  not
  g1287
  (
    n1325,
    n1317
  );


  not
  g1288
  (
    n1319,
    n1315
  );


  buf
  g1289
  (
    n1323,
    n1312
  );


  not
  g1290
  (
    n1320,
    n1314
  );


  not
  g1291
  (
    n1322,
    n1315
  );


  buf
  g1292
  (
    n1333,
    n1316
  );


  not
  g1293
  (
    n1330,
    n1315
  );


  not
  g1294
  (
    n1321,
    n1316
  );


  buf
  g1295
  (
    n1331,
    n1313
  );


  not
  g1296
  (
    n1326,
    n1314
  );


  not
  g1297
  (
    n1327,
    n1314
  );


  not
  g1298
  (
    n1332,
    n1316
  );


  not
  g1299
  (
    n1329,
    n1317
  );


  not
  g1300
  (
    n1328,
    n1311
  );


  not
  g1301
  (
    n1324,
    n1310
  );


  buf
  g1302
  (
    n1318,
    n1317
  );


  buf
  g1303
  (
    n1339,
    n1329
  );


  buf
  g1304
  (
    n1345,
    n593
  );


  not
  g1305
  (
    n1347,
    n1326
  );


  buf
  g1306
  (
    n1334,
    n146
  );


  nor
  g1307
  (
    n1335,
    n146,
    n1325,
    n596,
    n1322
  );


  xnor
  g1308
  (
    n1338,
    n595,
    n594,
    n147
  );


  or
  g1309
  (
    n1344,
    n144,
    n593,
    n1327
  );


  nand
  g1310
  (
    n1337,
    n963,
    n596,
    n595
  );


  xnor
  g1311
  (
    n1348,
    n1323,
    n145,
    n146,
    n148
  );


  nand
  g1312
  (
    n1349,
    n147,
    n1332,
    n964,
    n1328
  );


  xnor
  g1313
  (
    n1340,
    n594,
    n1330,
    n147,
    n1319
  );


  nor
  g1314
  (
    n1336,
    n1318,
    n146,
    n1333,
    n595
  );


  or
  g1315
  (
    n1342,
    n596,
    n597,
    n593,
    n1324
  );


  nor
  g1316
  (
    n1343,
    n147,
    n1320,
    n594,
    n965
  );


  and
  g1317
  (
    n1346,
    n148,
    n592,
    n145,
    n1321
  );


  xor
  g1318
  (
    n1341,
    n596,
    n145,
    n1331
  );


  not
  g1319
  (
    n1363,
    n1335
  );


  buf
  g1320
  (
    n1350,
    n1334
  );


  not
  g1321
  (
    n1351,
    n1336
  );


  not
  g1322
  (
    n1353,
    n1337
  );


  not
  g1323
  (
    n1356,
    n1334
  );


  not
  g1324
  (
    n1355,
    n1336
  );


  buf
  g1325
  (
    n1359,
    n1337
  );


  buf
  g1326
  (
    n1361,
    n1337
  );


  not
  g1327
  (
    n1360,
    n1334
  );


  not
  g1328
  (
    n1358,
    n1335
  );


  buf
  g1329
  (
    n1354,
    n1335
  );


  buf
  g1330
  (
    n1357,
    n1334
  );


  buf
  g1331
  (
    n1362,
    n1336
  );


  not
  g1332
  (
    n1352,
    n1335
  );


  buf
  g1333
  (
    n1364,
    n1336
  );


  xnor
  g1334
  (
    n1375,
    n1338,
    n1346,
    n1340,
    n1342
  );


  nand
  g1335
  (
    n1373,
    n1358,
    n1340,
    n1346,
    n1352
  );


  or
  g1336
  (
    n1368,
    n1349,
    n1358,
    n1359
  );


  xnor
  g1337
  (
    n1374,
    n1356,
    n1338,
    n1343,
    n1341
  );


  or
  g1338
  (
    n1382,
    n1356,
    n1348,
    n1354,
    n1343
  );


  nand
  g1339
  (
    n1381,
    n1342,
    n966,
    n1339,
    n1358
  );


  xor
  g1340
  (
    n1369,
    n1355,
    n1345,
    n1337
  );


  and
  g1341
  (
    n1377,
    n1348,
    n1357,
    n1342
  );


  xnor
  g1342
  (
    n1384,
    n1356,
    n1339,
    n1344,
    n1345
  );


  nor
  g1343
  (
    n1371,
    n1356,
    n1351,
    n1344,
    n1352
  );


  xnor
  g1344
  (
    n1366,
    n1349,
    n1345,
    n1358,
    n1340
  );


  xnor
  g1345
  (
    n1372,
    n1359,
    n1339,
    n1348,
    n1355
  );


  nor
  g1346
  (
    n1365,
    n1354,
    n1359,
    n1341,
    n1347
  );


  nand
  g1347
  (
    n1378,
    n1347,
    n1357,
    n1344,
    n1355
  );


  xnor
  g1348
  (
    n1380,
    n1341,
    n1353,
    n1338,
    n1349
  );


  and
  g1349
  (
    n1383,
    n1349,
    n1343,
    n1357,
    n1351
  );


  xor
  g1350
  (
    n1379,
    n1346,
    n1339,
    n1357,
    n1341
  );


  nor
  g1351
  (
    n1376,
    n1355,
    n1346,
    n1347,
    n1344
  );


  nor
  g1352
  (
    n1370,
    n1350,
    n1343,
    n1348,
    n1340
  );


  nor
  g1353
  (
    n1367,
    n1350,
    n1347,
    n1338,
    n1353
  );


  or
  g1354
  (
    n1393,
    n1361,
    n979,
    n983,
    n981
  );


  nand
  g1355
  (
    n1389,
    n970,
    n1374,
    n1360,
    n1384
  );


  xor
  g1356
  (
    n1395,
    n1363,
    n1376,
    n980,
    n969
  );


  or
  g1357
  (
    n1388,
    n984,
    n972,
    n974,
    n1361
  );


  nor
  g1358
  (
    n1392,
    n1360,
    n1360,
    n971,
    n1380
  );


  xnor
  g1359
  (
    n1386,
    n975,
    n1362,
    n1378,
    n982
  );


  nand
  g1360
  (
    n1390,
    n1382,
    n1381,
    n1361,
    n977
  );


  or
  g1361
  (
    n1391,
    n1361,
    n1360,
    n1375,
    n1363
  );


  and
  g1362
  (
    n1387,
    n973,
    n1362,
    n976
  );


  xnor
  g1363
  (
    n1394,
    n1377,
    n1362,
    n1363,
    n978
  );


  and
  g1364
  (
    n1385,
    n968,
    n967,
    n1383,
    n1379
  );


  not
  g1365
  (
    n1416,
    n987
  );


  not
  g1366
  (
    n1403,
    n1387
  );


  not
  g1367
  (
    n1433,
    n1390
  );


  buf
  g1368
  (
    n1432,
    n1389
  );


  not
  g1369
  (
    n1420,
    n150
  );


  not
  g1370
  (
    n1425,
    n1393
  );


  buf
  g1371
  (
    n1406,
    n1395
  );


  buf
  g1372
  (
    n1437,
    n1387
  );


  not
  g1373
  (
    n1428,
    n600
  );


  buf
  g1374
  (
    n1417,
    n1387
  );


  buf
  g1375
  (
    n1426,
    n1385
  );


  not
  g1376
  (
    n1411,
    n1389
  );


  not
  g1377
  (
    n1439,
    n601
  );


  buf
  g1378
  (
    n1402,
    n1391
  );


  buf
  g1379
  (
    n1418,
    n598
  );


  not
  g1380
  (
    n1401,
    n992
  );


  not
  g1381
  (
    n1438,
    n1386
  );


  buf
  g1382
  (
    n1404,
    n1364
  );


  buf
  g1383
  (
    n1427,
    n603
  );


  buf
  g1384
  (
    n1409,
    n601
  );


  buf
  g1385
  (
    n1423,
    n1395
  );


  and
  g1386
  (
    n1414,
    n149,
    n985,
    n150
  );


  and
  g1387
  (
    n1413,
    n1390,
    n1393,
    n1391
  );


  or
  g1388
  (
    n1399,
    n1393,
    n1388,
    n602
  );


  and
  g1389
  (
    n1407,
    n600,
    n986,
    n148
  );


  xor
  g1390
  (
    n1410,
    n1388,
    n1386,
    n1385
  );


  xor
  g1391
  (
    n1400,
    n601,
    n1385,
    n149
  );


  xnor
  g1392
  (
    n1436,
    n602,
    n1390,
    n1386
  );


  or
  g1393
  (
    n1398,
    n989,
    n600,
    n1394
  );


  xnor
  g1394
  (
    n1434,
    n601,
    n991,
    n990
  );


  xnor
  g1395
  (
    n1412,
    n599,
    n1394,
    n988
  );


  nor
  g1396
  (
    n1435,
    n598,
    n1388,
    n1393
  );


  xor
  g1397
  (
    n1421,
    n602,
    n1364,
    n1389
  );


  xnor
  g1398
  (
    n1419,
    n1387,
    n1392,
    n600
  );


  or
  g1399
  (
    n1429,
    n150,
    n599,
    n1363
  );


  and
  g1400
  (
    n1422,
    n1391,
    n1392
  );


  xor
  g1401
  (
    n1405,
    n603,
    n1392,
    n599
  );


  xnor
  g1402
  (
    n1430,
    n597,
    n1395
  );


  and
  g1403
  (
    n1408,
    n1385,
    n598,
    n1394
  );


  xnor
  g1404
  (
    n1424,
    n1391,
    n149
  );


  xor
  g1405
  (
    n1431,
    n1386,
    n597,
    n598
  );


  xor
  g1406
  (
    n1396,
    n597,
    n148,
    n1390
  );


  xnor
  g1407
  (
    n1397,
    n1388,
    n1389,
    n150
  );


  nor
  g1408
  (
    n1415,
    n1394,
    n599,
    n602
  );


  and
  g1409
  (
    n1440,
    n1439,
    n1422,
    n1419,
    n1431
  );


  or
  g1410
  (
    n1441,
    n1398,
    n1437,
    n1426,
    n1408
  );


  xor
  g1411
  (
    n1447,
    n1436,
    n1432,
    n1414,
    n1413
  );


  xor
  g1412
  (
    n1448,
    n1439,
    n1407,
    n1410
  );


  xor
  g1413
  (
    n1459,
    n1424,
    n1404,
    n1416,
    n1409
  );


  or
  g1414
  (
    n1445,
    n1414,
    n1430,
    n1416,
    n1411
  );


  and
  g1415
  (
    n1444,
    n1396,
    n1431,
    n1425,
    n1430
  );


  nor
  g1416
  (
    n1452,
    n1436,
    n1435,
    n1420
  );


  nand
  g1417
  (
    n1450,
    n1415,
    n1421,
    n1411
  );


  nor
  g1418
  (
    n1449,
    n1420,
    n1401,
    n1402,
    n1423
  );


  nand
  g1419
  (
    n1457,
    n1397,
    n1434,
    n1399,
    n1437
  );


  or
  g1420
  (
    n1451,
    n1433,
    n1429,
    n1406,
    n1427
  );


  xor
  g1421
  (
    n1446,
    n1438,
    n1418,
    n1429,
    n1412
  );


  xor
  g1422
  (
    n1455,
    n1409,
    n1428,
    n1427,
    n1417
  );


  xor
  g1423
  (
    n1454,
    n1425,
    n1405,
    n1403,
    n1428
  );


  xor
  g1424
  (
    n1442,
    n1424,
    n1417,
    n1438,
    n1410
  );


  xnor
  g1425
  (
    n1458,
    n1422,
    n1432,
    n1418,
    n1434
  );


  or
  g1426
  (
    n1453,
    n1415,
    n1400,
    n1419,
    n1408
  );


  xor
  g1427
  (
    n1456,
    n1412,
    n1433,
    n1426,
    n1406
  );


  and
  g1428
  (
    n1443,
    n1423,
    n1404,
    n1413,
    n1405
  );


  not
  g1429
  (
    n1463,
    n1440
  );


  not
  g1430
  (
    n1461,
    n1443
  );


  buf
  g1431
  (
    n1460,
    n1441
  );


  buf
  g1432
  (
    n1462,
    n1442
  );


  not
  g1433
  (
    n1464,
    n1463
  );


  buf
  g1434
  (
    n1466,
    n1462
  );


  and
  g1435
  (
    n1467,
    n1461,
    n604,
    n1460
  );


  and
  g1436
  (
    n1465,
    n605,
    n605,
    n603,
    n604
  );


  or
  g1437
  (
    n1468,
    n603,
    n1463,
    n605,
    n604
  );


  not
  g1438
  (
    n1474,
    n1465
  );


  not
  g1439
  (
    n1472,
    n1466
  );


  buf
  g1440
  (
    n1485,
    n1466
  );


  not
  g1441
  (
    n1477,
    n1468
  );


  buf
  g1442
  (
    n1469,
    n1467
  );


  not
  g1443
  (
    n1484,
    n1464
  );


  not
  g1444
  (
    n1486,
    n1467
  );


  not
  g1445
  (
    n1480,
    n1464
  );


  not
  g1446
  (
    n1479,
    n1466
  );


  not
  g1447
  (
    n1470,
    n1467
  );


  not
  g1448
  (
    n1475,
    n1468
  );


  buf
  g1449
  (
    n1478,
    n1468
  );


  not
  g1450
  (
    n1481,
    n1465
  );


  buf
  g1451
  (
    n1483,
    n1466
  );


  not
  g1452
  (
    n1482,
    n1465
  );


  not
  g1453
  (
    n1471,
    n1467
  );


  buf
  g1454
  (
    n1476,
    n1465
  );


  not
  g1455
  (
    n1473,
    n1468
  );


  or
  g1456
  (
    n1539,
    n1018,
    n1116,
    n1061,
    n1484
  );


  xnor
  g1457
  (
    n1525,
    n1043,
    n1084,
    n1135,
    n1005
  );


  and
  g1458
  (
    n1537,
    n1121,
    n1017,
    n1032,
    n1041
  );


  and
  g1459
  (
    n1494,
    n1030,
    n1206,
    n1022,
    n1031
  );


  xor
  g1460
  (
    n1551,
    n1002,
    n1015,
    n1062,
    n1474
  );


  and
  g1461
  (
    n1501,
    n1028,
    n1033,
    n1196,
    n1184
  );


  nor
  g1462
  (
    n1515,
    n1167,
    n1097,
    n1042,
    n1081
  );


  xor
  g1463
  (
    n1498,
    n1472,
    n1153,
    n1078,
    n1474
  );


  nor
  g1464
  (
    n1542,
    n1070,
    n1485,
    n1191,
    n1103
  );


  xor
  g1465
  (
    n1541,
    n1140,
    n1478,
    n1483,
    n1187
  );


  nor
  g1466
  (
    n1507,
    n1166,
    n1127,
    n1170,
    n1204
  );


  nand
  g1467
  (
    n1505,
    n1474,
    n1006,
    n1181,
    n1069
  );


  nand
  g1468
  (
    n1511,
    n1024,
    n1105,
    n1208,
    n1067
  );


  nor
  g1469
  (
    n1506,
    n1016,
    n1056,
    n1100,
    n1025
  );


  nor
  g1470
  (
    n1540,
    n1035,
    n1151,
    n1085,
    n1478
  );


  xnor
  g1471
  (
    n1513,
    n1480,
    n1484,
    n1045,
    n1066
  );


  xor
  g1472
  (
    n1528,
    n1125,
    n1161,
    n1478,
    n1149
  );


  and
  g1473
  (
    n1492,
    n1198,
    n1119,
    n1021,
    n1477
  );


  nand
  g1474
  (
    n1530,
    n1472,
    n1169,
    n1142,
    n1471
  );


  nand
  g1475
  (
    n1548,
    n1019,
    n1063,
    n1476,
    n1004
  );


  and
  g1476
  (
    n1523,
    n1136,
    n1177,
    n1477,
    n1160
  );


  nand
  g1477
  (
    n1538,
    n1171,
    n1026,
    n1088,
    n1175
  );


  and
  g1478
  (
    n1536,
    n1207,
    n1120,
    n1101,
    n1051
  );


  xnor
  g1479
  (
    n1547,
    n1172,
    n1165,
    n1481,
    n994
  );


  nor
  g1480
  (
    n1532,
    n1474,
    n1047,
    n1037,
    n1111
  );


  nand
  g1481
  (
    n1489,
    n1150,
    n1182,
    n1481,
    n1471
  );


  nor
  g1482
  (
    n1550,
    n996,
    n1482,
    n1193,
    n1057
  );


  xnor
  g1483
  (
    n1517,
    n1046,
    n1202,
    n1068,
    n1110
  );


  xor
  g1484
  (
    n1544,
    n1134,
    n1072,
    n1118,
    n1485
  );


  and
  g1485
  (
    n1491,
    n1090,
    n1020,
    n1482,
    n1479
  );


  and
  g1486
  (
    n1553,
    n1131,
    n1477,
    n1096,
    n1203
  );


  nand
  g1487
  (
    n1524,
    n1054,
    n1092,
    n1044,
    n1205
  );


  xor
  g1488
  (
    n1554,
    n1195,
    n1469,
    n1486,
    n1040
  );


  xnor
  g1489
  (
    n1512,
    n1077,
    n1122,
    n1098,
    n1174
  );


  nor
  g1490
  (
    n1503,
    n1094,
    n1477,
    n1482,
    n1117
  );


  xor
  g1491
  (
    n1545,
    n1476,
    n995,
    n1036,
    n1079
  );


  xnor
  g1492
  (
    n1499,
    n1129,
    n1139,
    n1470,
    n1186
  );


  xor
  g1493
  (
    n1497,
    n1055,
    n1093,
    n999,
    n1152
  );


  nor
  g1494
  (
    n1510,
    n1190,
    n1102,
    n1049,
    n1486
  );


  nor
  g1495
  (
    n1518,
    n1071,
    n1027,
    n1104,
    n1074
  );


  nand
  g1496
  (
    n1488,
    n1475,
    n1469,
    n1010,
    n1014
  );


  and
  g1497
  (
    n1520,
    n1180,
    n1107,
    n1179,
    n1008
  );


  xor
  g1498
  (
    n1555,
    n1178,
    n1173,
    n1475,
    n1194
  );


  xor
  g1499
  (
    n1556,
    n993,
    n1483,
    n1485,
    n1106
  );


  or
  g1500
  (
    n1549,
    n1145,
    n1000,
    n1130,
    n1483
  );


  xnor
  g1501
  (
    n1496,
    n1073,
    n1080,
    n1157,
    n1144
  );


  nand
  g1502
  (
    n1514,
    n1064,
    n1481,
    n1486,
    n1470
  );


  xor
  g1503
  (
    n1557,
    n1065,
    n1148,
    n1162,
    n1076
  );


  nand
  g1504
  (
    n1500,
    n1483,
    n1115,
    n1163,
    n1083
  );


  xor
  g1505
  (
    n1487,
    n1128,
    n1124,
    n1001,
    n1003
  );


  or
  g1506
  (
    n1502,
    n1075,
    n1479,
    n1470,
    n1473
  );


  xor
  g1507
  (
    n1521,
    n1472,
    n1137,
    n1486,
    n1053
  );


  nor
  g1508
  (
    n1558,
    n1199,
    n1086,
    n1479,
    n1082
  );


  xnor
  g1509
  (
    n1533,
    n1126,
    n1099,
    n1012,
    n1475
  );


  xor
  g1510
  (
    n1546,
    n1481,
    n1133,
    n1471,
    n1470
  );


  or
  g1511
  (
    n1529,
    n1011,
    n1478,
    n1473,
    n1485
  );


  xor
  g1512
  (
    n1490,
    n1197,
    n1060,
    n1113,
    n1038
  );


  and
  g1513
  (
    n1493,
    n1168,
    n1188,
    n1475,
    n1183
  );


  nand
  g1514
  (
    n1516,
    n1087,
    n1479,
    n1469,
    n998
  );


  nand
  g1515
  (
    n1526,
    n1192,
    n1108,
    n1480,
    n1473
  );


  xor
  g1516
  (
    n1535,
    n1156,
    n1039,
    n1007,
    n1123
  );


  xor
  g1517
  (
    n1495,
    n1058,
    n1048,
    n1089,
    n1138
  );


  nor
  g1518
  (
    n1543,
    n1476,
    n1472,
    n1484,
    n1009
  );


  and
  g1519
  (
    n1504,
    n1112,
    n1023,
    n1201,
    n1176
  );


  and
  g1520
  (
    n1522,
    n1200,
    n1469,
    n1109,
    n1480
  );


  nor
  g1521
  (
    n1508,
    n1034,
    n1471,
    n1484,
    n1480
  );


  xnor
  g1522
  (
    n1552,
    n1141,
    n1052,
    n1159,
    n1164
  );


  xor
  g1523
  (
    n1519,
    n1154,
    n1132,
    n1476,
    n1189
  );


  xnor
  g1524
  (
    n1527,
    n1473,
    n1029,
    n1059,
    n1185
  );


  nor
  g1525
  (
    n1509,
    n1114,
    n1095,
    n1091,
    n1158
  );


  nand
  g1526
  (
    n1534,
    n1155,
    n1482,
    n997,
    n1146
  );


  xor
  g1527
  (
    n1531,
    n1050,
    n1143,
    n1147,
    n1013
  );


  buf
  g1528
  (
    n1812,
    n1554
  );


  not
  g1529
  (
    n1588,
    n1494
  );


  not
  g1530
  (
    n1703,
    n1505
  );


  buf
  g1531
  (
    n1809,
    n1503
  );


  buf
  g1532
  (
    n1583,
    n1518
  );


  buf
  g1533
  (
    n1793,
    n1494
  );


  buf
  g1534
  (
    n1752,
    n1531
  );


  buf
  g1535
  (
    n1741,
    n1519
  );


  not
  g1536
  (
    n1842,
    n1539
  );


  not
  g1537
  (
    n1751,
    n1504
  );


  buf
  g1538
  (
    n1563,
    n1491
  );


  not
  g1539
  (
    n1660,
    n1526
  );


  buf
  g1540
  (
    n1621,
    n1506
  );


  buf
  g1541
  (
    n1726,
    n1539
  );


  buf
  g1542
  (
    n1608,
    n1492
  );


  buf
  g1543
  (
    n1845,
    n1556
  );


  buf
  g1544
  (
    n1780,
    n1551
  );


  buf
  g1545
  (
    n1828,
    n1519
  );


  buf
  g1546
  (
    n1843,
    n1489
  );


  buf
  g1547
  (
    n1618,
    n1536
  );


  not
  g1548
  (
    n1705,
    n1446
  );


  buf
  g1549
  (
    n1816,
    n1533
  );


  not
  g1550
  (
    n1821,
    n1543
  );


  not
  g1551
  (
    n1803,
    n1521
  );


  buf
  g1552
  (
    n1584,
    n1532
  );


  not
  g1553
  (
    n1657,
    n1549
  );


  not
  g1554
  (
    n1661,
    n1536
  );


  not
  g1555
  (
    n1593,
    n1517
  );


  not
  g1556
  (
    n1652,
    n1534
  );


  buf
  g1557
  (
    n1818,
    n1454
  );


  not
  g1558
  (
    n1770,
    n1551
  );


  not
  g1559
  (
    n1674,
    n1491
  );


  not
  g1560
  (
    n1586,
    n1551
  );


  not
  g1561
  (
    n1736,
    n1497
  );


  not
  g1562
  (
    n1638,
    n1523
  );


  not
  g1563
  (
    n1749,
    n1557
  );


  buf
  g1564
  (
    n1682,
    n1503
  );


  buf
  g1565
  (
    n1683,
    n1518
  );


  not
  g1566
  (
    n1701,
    n1453
  );


  not
  g1567
  (
    n1560,
    n1504
  );


  not
  g1568
  (
    n1822,
    n1540
  );


  not
  g1569
  (
    n1595,
    n1528
  );


  not
  g1570
  (
    n1704,
    n1552
  );


  buf
  g1571
  (
    n1581,
    n1530
  );


  buf
  g1572
  (
    n1727,
    n1524
  );


  not
  g1573
  (
    n1696,
    n1536
  );


  not
  g1574
  (
    n1624,
    n1491
  );


  buf
  g1575
  (
    n1656,
    n1540
  );


  not
  g1576
  (
    n1600,
    n1529
  );


  not
  g1577
  (
    n1790,
    n1512
  );


  not
  g1578
  (
    n1647,
    n1529
  );


  buf
  g1579
  (
    n1758,
    n1527
  );


  buf
  g1580
  (
    n1626,
    n1509
  );


  buf
  g1581
  (
    n1672,
    n1556
  );


  buf
  g1582
  (
    n1562,
    n1495
  );


  not
  g1583
  (
    n1761,
    n1492
  );


  not
  g1584
  (
    n1802,
    n1516
  );


  buf
  g1585
  (
    n1838,
    n1525
  );


  buf
  g1586
  (
    n1836,
    n1512
  );


  buf
  g1587
  (
    n1680,
    n1526
  );


  not
  g1588
  (
    n1671,
    n1538
  );


  buf
  g1589
  (
    n1561,
    n1452
  );


  not
  g1590
  (
    KeyWire_0_25,
    n1494
  );


  buf
  g1591
  (
    KeyWire_0_24,
    n1521
  );


  buf
  g1592
  (
    n1730,
    n1532
  );


  buf
  g1593
  (
    n1789,
    n1529
  );


  buf
  g1594
  (
    n1753,
    n1537
  );


  not
  g1595
  (
    n1635,
    n1487
  );


  not
  g1596
  (
    n1580,
    n1507
  );


  not
  g1597
  (
    n1788,
    n1545
  );


  buf
  g1598
  (
    n1759,
    n1549
  );


  not
  g1599
  (
    n1694,
    n1515
  );


  buf
  g1600
  (
    n1798,
    n1520
  );


  not
  g1601
  (
    n1605,
    n1558
  );


  not
  g1602
  (
    n1628,
    n1524
  );


  not
  g1603
  (
    n1817,
    n1495
  );


  buf
  g1604
  (
    n1659,
    n1510
  );


  buf
  g1605
  (
    n1718,
    n1501
  );


  not
  g1606
  (
    n1737,
    n1543
  );


  buf
  g1607
  (
    n1796,
    n1555
  );


  buf
  g1608
  (
    n1739,
    n1558
  );


  not
  g1609
  (
    n1766,
    n1499
  );


  not
  g1610
  (
    n1653,
    n1523
  );


  not
  g1611
  (
    n1702,
    n1540
  );


  buf
  g1612
  (
    n1754,
    n1293
  );


  not
  g1613
  (
    n1695,
    n1507
  );


  buf
  g1614
  (
    n1573,
    n1526
  );


  not
  g1615
  (
    n1716,
    n1507
  );


  buf
  g1616
  (
    n1643,
    n1490
  );


  not
  g1617
  (
    n1668,
    n1499
  );


  not
  g1618
  (
    KeyWire_0_3,
    n1538
  );


  buf
  g1619
  (
    n1797,
    n1545
  );


  not
  g1620
  (
    n1594,
    n1496
  );


  not
  g1621
  (
    n1642,
    n1512
  );


  buf
  g1622
  (
    n1575,
    n1502
  );


  not
  g1623
  (
    n1596,
    n1488
  );


  not
  g1624
  (
    n1662,
    n1554
  );


  not
  g1625
  (
    n1639,
    n1296
  );


  buf
  g1626
  (
    n1729,
    n1497
  );


  buf
  g1627
  (
    n1645,
    n1509
  );


  buf
  g1628
  (
    n1731,
    n1520
  );


  buf
  g1629
  (
    n1782,
    n1513
  );


  buf
  g1630
  (
    n1697,
    n1503
  );


  buf
  g1631
  (
    n1805,
    n1300
  );


  buf
  g1632
  (
    n1744,
    n1530
  );


  not
  g1633
  (
    n1792,
    n1552
  );


  not
  g1634
  (
    n1743,
    n1542
  );


  not
  g1635
  (
    n1801,
    n1521
  );


  not
  g1636
  (
    n1578,
    n1488
  );


  buf
  g1637
  (
    n1732,
    n1518
  );


  buf
  g1638
  (
    n1633,
    n1549
  );


  not
  g1639
  (
    n1786,
    n1455
  );


  not
  g1640
  (
    n1756,
    n1541
  );


  buf
  g1641
  (
    n1811,
    n1493
  );


  not
  g1642
  (
    n1712,
    n1551
  );


  not
  g1643
  (
    KeyWire_0_7,
    n1491
  );


  not
  g1644
  (
    n1623,
    n1543
  );


  not
  g1645
  (
    n1746,
    n1535
  );


  not
  g1646
  (
    n1677,
    n1543
  );


  not
  g1647
  (
    n1587,
    n1515
  );


  buf
  g1648
  (
    n1625,
    n1511
  );


  not
  g1649
  (
    n1781,
    n1498
  );


  buf
  g1650
  (
    n1765,
    n1557
  );


  not
  g1651
  (
    KeyWire_0_6,
    n1509
  );


  buf
  g1652
  (
    n1615,
    n1553
  );


  not
  g1653
  (
    n1776,
    n1549
  );


  buf
  g1654
  (
    n1709,
    n1528
  );


  not
  g1655
  (
    n1649,
    n1503
  );


  not
  g1656
  (
    n1655,
    n1548
  );


  buf
  g1657
  (
    n1827,
    n1548
  );


  buf
  g1658
  (
    n1693,
    n1302
  );


  buf
  g1659
  (
    n1666,
    n1554
  );


  buf
  g1660
  (
    n1819,
    n1487
  );


  buf
  g1661
  (
    n1571,
    n1297
  );


  buf
  g1662
  (
    n1764,
    n1525
  );


  not
  g1663
  (
    n1747,
    n1554
  );


  not
  g1664
  (
    n1582,
    n1299
  );


  not
  g1665
  (
    n1585,
    n1555
  );


  buf
  g1666
  (
    n1640,
    n1294
  );


  buf
  g1667
  (
    n1748,
    n1539
  );


  not
  g1668
  (
    n1733,
    n1516
  );


  buf
  g1669
  (
    n1734,
    n1507
  );


  buf
  g1670
  (
    n1698,
    n1492
  );


  not
  g1671
  (
    n1599,
    n1497
  );


  buf
  g1672
  (
    n1772,
    n1533
  );


  not
  g1673
  (
    n1665,
    n1301
  );


  buf
  g1674
  (
    n1823,
    n1550
  );


  buf
  g1675
  (
    n1681,
    n1303
  );


  not
  g1676
  (
    n1807,
    n1448
  );


  buf
  g1677
  (
    n1576,
    n1451
  );


  buf
  g1678
  (
    n1728,
    n1558
  );


  not
  g1679
  (
    n1837,
    n1508
  );


  buf
  g1680
  (
    n1641,
    n1537
  );


  buf
  g1681
  (
    n1745,
    n1494
  );


  buf
  g1682
  (
    n1713,
    n1502
  );


  not
  g1683
  (
    n1829,
    n1544
  );


  buf
  g1684
  (
    n1715,
    n1529
  );


  buf
  g1685
  (
    n1634,
    n1532
  );


  not
  g1686
  (
    n1572,
    n1541
  );


  buf
  g1687
  (
    n1835,
    n1364
  );


  buf
  g1688
  (
    n1688,
    n1517
  );


  buf
  g1689
  (
    n1650,
    n1528
  );


  not
  g1690
  (
    n1676,
    n1525
  );


  not
  g1691
  (
    n1717,
    n1546
  );


  buf
  g1692
  (
    n1791,
    n1557
  );


  not
  g1693
  (
    n1841,
    n1547
  );


  buf
  g1694
  (
    n1604,
    n1445
  );


  buf
  g1695
  (
    n1714,
    n1506
  );


  not
  g1696
  (
    n1566,
    n1546
  );


  buf
  g1697
  (
    n1654,
    n1498
  );


  not
  g1698
  (
    n1719,
    n1501
  );


  not
  g1699
  (
    n1799,
    n1508
  );


  buf
  g1700
  (
    n1710,
    n1499
  );


  not
  g1701
  (
    n1773,
    n1514
  );


  buf
  g1702
  (
    n1777,
    n1530
  );


  not
  g1703
  (
    n1775,
    n1488
  );


  buf
  g1704
  (
    n1720,
    n1493
  );


  buf
  g1705
  (
    n1601,
    n1501
  );


  buf
  g1706
  (
    n1738,
    n1534
  );


  not
  g1707
  (
    n1840,
    n1488
  );


  buf
  g1708
  (
    n1606,
    n1522
  );


  buf
  g1709
  (
    n1774,
    n1535
  );


  not
  g1710
  (
    n1627,
    n1499
  );


  not
  g1711
  (
    n1826,
    n1509
  );


  not
  g1712
  (
    n1844,
    n1520
  );


  buf
  g1713
  (
    KeyWire_0_23,
    n1519
  );


  not
  g1714
  (
    n1778,
    n1527
  );


  buf
  g1715
  (
    n1607,
    n1298
  );


  not
  g1716
  (
    n1569,
    n1511
  );


  not
  g1717
  (
    n1636,
    n1517
  );


  buf
  g1718
  (
    n1846,
    n1547
  );


  buf
  g1719
  (
    n1574,
    n1540
  );


  buf
  g1720
  (
    n1691,
    n1490
  );


  buf
  g1721
  (
    n1824,
    n1510
  );


  not
  g1722
  (
    n1577,
    n1492
  );


  buf
  g1723
  (
    n1757,
    n1538
  );


  buf
  g1724
  (
    n1663,
    n1521
  );


  not
  g1725
  (
    n1637,
    n1292
  );


  buf
  g1726
  (
    n1644,
    n1515
  );


  not
  g1727
  (
    n1687,
    n1531
  );


  buf
  g1728
  (
    n1567,
    n1525
  );


  not
  g1729
  (
    n1783,
    n1489
  );


  not
  g1730
  (
    n1830,
    n1533
  );


  not
  g1731
  (
    n1616,
    n1547
  );


  not
  g1732
  (
    n1564,
    n1542
  );


  buf
  g1733
  (
    n1675,
    n1496
  );


  not
  g1734
  (
    n1742,
    n1555
  );


  buf
  g1735
  (
    n1724,
    n1537
  );


  not
  g1736
  (
    n1609,
    n1531
  );


  buf
  g1737
  (
    n1667,
    n1511
  );


  buf
  g1738
  (
    n1814,
    n1548
  );


  buf
  g1739
  (
    n1690,
    n1505
  );


  buf
  g1740
  (
    n1568,
    n1545
  );


  buf
  g1741
  (
    n1686,
    n1496
  );


  not
  g1742
  (
    n1833,
    n1534
  );


  buf
  g1743
  (
    n1684,
    n1502
  );


  buf
  g1744
  (
    n1629,
    n1520
  );


  not
  g1745
  (
    n1612,
    n1209
  );


  not
  g1746
  (
    n1559,
    n1541
  );


  not
  g1747
  (
    n1750,
    n1495
  );


  buf
  g1748
  (
    n1631,
    n1545
  );


  not
  g1749
  (
    n1760,
    n1555
  );


  not
  g1750
  (
    n1815,
    n1487
  );


  not
  g1751
  (
    n1787,
    n1546
  );


  not
  g1752
  (
    n1679,
    n1496
  );


  not
  g1753
  (
    n1706,
    n1513
  );


  not
  g1754
  (
    n1755,
    n1515
  );


  buf
  g1755
  (
    n1685,
    n1553
  );


  buf
  g1756
  (
    n1602,
    n1517
  );


  buf
  g1757
  (
    n1813,
    n1514
  );


  buf
  g1758
  (
    n1579,
    n1552
  );


  not
  g1759
  (
    n1721,
    n1553
  );


  not
  g1760
  (
    n1610,
    n1500
  );


  not
  g1761
  (
    n1630,
    n1523
  );


  not
  g1762
  (
    n1808,
    n1505
  );


  buf
  g1763
  (
    n1785,
    n1490
  );


  not
  g1764
  (
    n1768,
    n1513
  );


  not
  g1765
  (
    n1651,
    n1489
  );


  buf
  g1766
  (
    n1603,
    n1505
  );


  buf
  g1767
  (
    n1771,
    n1506
  );


  not
  g1768
  (
    n1806,
    n1514
  );


  not
  g1769
  (
    n1598,
    n1522
  );


  not
  g1770
  (
    n1722,
    n1500
  );


  buf
  g1771
  (
    n1839,
    n1364
  );


  buf
  g1772
  (
    n1664,
    n1557
  );


  not
  g1773
  (
    n1834,
    n1504
  );


  not
  g1774
  (
    n1795,
    n1550
  );


  not
  g1775
  (
    n1810,
    n1532
  );


  not
  g1776
  (
    n1622,
    n1556
  );


  buf
  g1777
  (
    n1617,
    n1544
  );


  not
  g1778
  (
    n1794,
    n1510
  );


  not
  g1779
  (
    n1707,
    n1498
  );


  buf
  g1780
  (
    n1597,
    n1528
  );


  not
  g1781
  (
    n1592,
    n1524
  );


  buf
  g1782
  (
    n1831,
    n1539
  );


  buf
  g1783
  (
    n1825,
    n1490
  );


  not
  g1784
  (
    n1800,
    n1493
  );


  not
  g1785
  (
    n1820,
    n1295
  );


  buf
  g1786
  (
    n1769,
    n1541
  );


  buf
  g1787
  (
    n1614,
    n1512
  );


  not
  g1788
  (
    n1832,
    n1553
  );


  buf
  g1789
  (
    n1613,
    n1514
  );


  not
  g1790
  (
    n1763,
    n1487
  );


  buf
  g1791
  (
    n1570,
    n1537
  );


  buf
  g1792
  (
    n1632,
    n1519
  );


  not
  g1793
  (
    n1804,
    n1449
  );


  not
  g1794
  (
    n1723,
    n1516
  );


  buf
  g1795
  (
    n1658,
    n1544
  );


  buf
  g1796
  (
    n1678,
    n1531
  );


  not
  g1797
  (
    n1692,
    n1513
  );


  buf
  g1798
  (
    n1620,
    n1527
  );


  buf
  g1799
  (
    n1646,
    n1501
  );


  not
  g1800
  (
    n1689,
    n1450
  );


  not
  g1801
  (
    n1648,
    n1506
  );


  nor
  g1802
  (
    n1590,
    n1535,
    n1523,
    n1498
  );


  or
  g1803
  (
    n1670,
    n1518,
    n1444,
    n1546
  );


  nor
  g1804
  (
    n1762,
    n1530,
    n1522,
    n1510
  );


  or
  g1805
  (
    n1619,
    n1535,
    n1493,
    n1556
  );


  nand
  g1806
  (
    n1591,
    n1550,
    n1552,
    n1511
  );


  nor
  g1807
  (
    n1669,
    n1508,
    n1500,
    n1516
  );


  nor
  g1808
  (
    n1700,
    n1538,
    n1542,
    n1508
  );


  xor
  g1809
  (
    n1740,
    n1500,
    n1456,
    n1497
  );


  xor
  g1810
  (
    n1779,
    n1536,
    n1504,
    n1447
  );


  nand
  g1811
  (
    n1611,
    n1522,
    n1558,
    n1495
  );


  xor
  g1812
  (
    n1735,
    n1550,
    n1547,
    n1524
  );


  nor
  g1813
  (
    n1767,
    n1542,
    n1534,
    n1544
  );


  and
  g1814
  (
    n1699,
    n1489,
    n1526,
    n1533
  );


  and
  g1815
  (
    n1784,
    n1502,
    n1548,
    n1527
  );


  nor
  g1816
  (
    n2032,
    n1833,
    n1698,
    n1836,
    n1775
  );


  nor
  g1817
  (
    n2001,
    n1819,
    n1840,
    n1761,
    n1737
  );


  nand
  g1818
  (
    n1991,
    n1712,
    n1838,
    n1581,
    n1708
  );


  nand
  g1819
  (
    n1847,
    n1700,
    n1794,
    n1715,
    n1831
  );


  nor
  g1820
  (
    n1994,
    n1815,
    n1599,
    n1647,
    n1843
  );


  xor
  g1821
  (
    n1861,
    n1587,
    n1772,
    n1670,
    n1781
  );


  xnor
  g1822
  (
    n1920,
    n1603,
    n1714,
    n1728,
    n1563
  );


  nor
  g1823
  (
    n1891,
    n1814,
    n1787,
    n1846,
    n1607
  );


  xnor
  g1824
  (
    n2018,
    n1725,
    n1802,
    n1695,
    n1832
  );


  xnor
  g1825
  (
    n1928,
    n1812,
    n1781,
    n1840,
    n1751
  );


  and
  g1826
  (
    n2038,
    n1688,
    n1778,
    n1704,
    n1824
  );


  xor
  g1827
  (
    n1865,
    n1458,
    n1835,
    n1679,
    n1838
  );


  xnor
  g1828
  (
    n1848,
    n1831,
    n1708,
    n1709,
    n1668
  );


  nor
  g1829
  (
    n2034,
    n1715,
    n1744,
    n1565,
    n1765
  );


  xor
  g1830
  (
    n2027,
    n1725,
    n1594,
    n1692,
    n1635
  );


  xor
  g1831
  (
    n2026,
    n1730,
    n1713,
    n1795,
    n1845
  );


  nand
  g1832
  (
    n1988,
    n1782,
    n1786,
    n1711,
    n1730
  );


  and
  g1833
  (
    n2008,
    n1810,
    n1769,
    n1801,
    n1731
  );


  nor
  g1834
  (
    n1915,
    n1667,
    n1567,
    n1753,
    n1807
  );


  or
  g1835
  (
    n1996,
    n1780,
    n1459,
    n1645,
    n1758
  );


  nand
  g1836
  (
    n1881,
    n1826,
    n1693,
    n1756,
    n1721
  );


  and
  g1837
  (
    n2023,
    n1839,
    n1712,
    n1702,
    n1723
  );


  nor
  g1838
  (
    n1883,
    n1777,
    n1663,
    n1792,
    n1833
  );


  nand
  g1839
  (
    n1975,
    n1694,
    n1753,
    n1616,
    n1826
  );


  xor
  g1840
  (
    n1893,
    n1723,
    n1724,
    n1765,
    n1756
  );


  or
  g1841
  (
    n2015,
    n1838,
    n1670,
    n1778,
    n1752
  );


  nor
  g1842
  (
    n1856,
    n1648,
    n1726,
    n1773,
    n1628
  );


  and
  g1843
  (
    n1917,
    n1624,
    n1754,
    n1650,
    n1590
  );


  and
  g1844
  (
    n1936,
    n1737,
    n1813,
    n1748,
    n1819
  );


  xor
  g1845
  (
    n1860,
    n1814,
    n1606,
    n1780,
    n1810
  );


  and
  g1846
  (
    n1958,
    n1816,
    n1807,
    n1841,
    n1760
  );


  xnor
  g1847
  (
    n1877,
    n1737,
    n1830,
    n1677,
    n1785
  );


  nand
  g1848
  (
    n2009,
    n1705,
    n1844,
    n1727,
    n1611
  );


  nand
  g1849
  (
    n1954,
    n1651,
    n1731,
    n1714,
    n1688
  );


  or
  g1850
  (
    n1962,
    n1789,
    n1806,
    n1676,
    n1693
  );


  or
  g1851
  (
    n1898,
    n1716,
    n1826,
    n1798,
    n1790
  );


  xor
  g1852
  (
    n1873,
    n1811,
    n1726,
    n1814,
    n1620
  );


  nor
  g1853
  (
    KeyWire_0_27,
    n1717,
    n1800,
    n1747,
    n1709
  );


  and
  g1854
  (
    n2037,
    n1788,
    n1738,
    n1843,
    n1786
  );


  nand
  g1855
  (
    n1885,
    n1673,
    n1759,
    n1569,
    n1757
  );


  xnor
  g1856
  (
    n1867,
    n1784,
    n1828,
    n1792,
    n1788
  );


  xnor
  g1857
  (
    n1943,
    n1617,
    n1815,
    n1800,
    n1786
  );


  xor
  g1858
  (
    n1869,
    n1777,
    n1707,
    n1818,
    n1693
  );


  nor
  g1859
  (
    n1987,
    n1824,
    n1742,
    n1560,
    n1706
  );


  and
  g1860
  (
    n2024,
    n1691,
    n1686,
    n1830,
    n1820
  );


  nand
  g1861
  (
    n2002,
    n1827,
    n1752,
    n1694,
    n1811
  );


  xor
  g1862
  (
    n2014,
    n1799,
    n1707,
    n1614,
    n1715
  );


  or
  g1863
  (
    n2004,
    n1740,
    n1797,
    n1818,
    n1653
  );


  xnor
  g1864
  (
    n1849,
    n1830,
    n1738,
    n1775,
    n1843
  );


  xor
  g1865
  (
    n1929,
    n1724,
    n1829,
    n1739,
    n1791
  );


  xnor
  g1866
  (
    n1990,
    n1716,
    n1597,
    n1808,
    n1610
  );


  xnor
  g1867
  (
    n1910,
    n1812,
    n1750,
    n1804,
    n1793
  );


  xnor
  g1868
  (
    n1961,
    n1809,
    n1753,
    n1754,
    n1808
  );


  xor
  g1869
  (
    n1934,
    n1718,
    n1604,
    n1733,
    n1827
  );


  and
  g1870
  (
    n1982,
    n1740,
    n1584,
    n1844,
    n1643
  );


  and
  g1871
  (
    n1956,
    n1741,
    n1800,
    n1613,
    n1457
  );


  xor
  g1872
  (
    n2007,
    n1819,
    n1631,
    n1705,
    n1589
  );


  xor
  g1873
  (
    n1901,
    n1837,
    n1766,
    n1769,
    n1652
  );


  xnor
  g1874
  (
    n1974,
    n1741,
    n1699,
    n1739,
    n1736
  );


  xnor
  g1875
  (
    n1963,
    n1767,
    n1801,
    n1820,
    n1621
  );


  xor
  g1876
  (
    n1926,
    n1797,
    n1772,
    n1811,
    n1760
  );


  nand
  g1877
  (
    n1960,
    n1820,
    n1681,
    n1739,
    n1776
  );


  or
  g1878
  (
    n2011,
    n1761,
    n1784,
    n1672,
    n1828
  );


  nand
  g1879
  (
    n1892,
    n1839,
    n1839,
    n1666,
    n1811
  );


  or
  g1880
  (
    n2031,
    n1730,
    n1783,
    n1809,
    n1798
  );


  or
  g1881
  (
    n1935,
    n1703,
    n1780,
    n1712,
    n1698
  );


  nand
  g1882
  (
    n1980,
    n1817,
    n1762,
    n1803,
    n1683
  );


  or
  g1883
  (
    n2021,
    n1727,
    n1744,
    n1696,
    n1755
  );


  or
  g1884
  (
    n1932,
    n1723,
    n1732,
    n1742,
    n1796
  );


  and
  g1885
  (
    n1977,
    n1679,
    n1773,
    n1774,
    n1649
  );


  xor
  g1886
  (
    n2036,
    n1784,
    n1812,
    n1741,
    n1626
  );


  and
  g1887
  (
    n1937,
    n1790,
    n1736,
    n1575,
    n1729
  );


  xnor
  g1888
  (
    n1886,
    n1755,
    n1783,
    n1719,
    n1787
  );


  nand
  g1889
  (
    n1889,
    n1802,
    n1778,
    n1699,
    n1795
  );


  nor
  g1890
  (
    n1850,
    n1789,
    n1769,
    n1574,
    n1823
  );


  or
  g1891
  (
    n2006,
    n1734,
    n1826,
    n1803,
    n1632
  );


  and
  g1892
  (
    n1964,
    n1780,
    n1766,
    n1627,
    n1763
  );


  nand
  g1893
  (
    n2010,
    n1605,
    n1825,
    n1783,
    n1735
  );


  xor
  g1894
  (
    n1945,
    n1837,
    n1661,
    n1794,
    n1750
  );


  or
  g1895
  (
    n1950,
    n1803,
    n1692,
    n1608,
    n1781
  );


  xor
  g1896
  (
    n2005,
    n1736,
    n1846,
    n1709,
    n1671
  );


  nand
  g1897
  (
    n1955,
    n1805,
    n1825,
    n1745,
    n1725
  );


  xnor
  g1898
  (
    n1947,
    n1596,
    n1674,
    n1746,
    n1754
  );


  or
  g1899
  (
    n2028,
    n1699,
    n1771,
    n1720,
    n1571
  );


  xor
  g1900
  (
    n1938,
    n1782,
    n1568,
    n1808,
    n1664
  );


  nor
  g1901
  (
    n2033,
    n1816,
    n1772,
    n1842,
    n1776
  );


  nor
  g1902
  (
    n1925,
    n1798,
    n1751,
    n1703,
    n1582
  );


  nand
  g1903
  (
    n1909,
    n1722,
    n1709,
    n1659,
    n1833
  );


  nand
  g1904
  (
    n1905,
    n1646,
    n1706,
    n1799,
    n1822
  );


  xnor
  g1905
  (
    n1986,
    n1680,
    n1767,
    n1711,
    n1675
  );


  xnor
  g1906
  (
    n1983,
    n1676,
    n1838,
    n1815,
    n1779
  );


  nand
  g1907
  (
    n1957,
    n1598,
    n1717,
    n1702,
    n1749
  );


  or
  g1908
  (
    n1916,
    n1834,
    n1809,
    n1763,
    n1713
  );


  xor
  g1909
  (
    n1908,
    n1768,
    n1710,
    n1743,
    n1717
  );


  or
  g1910
  (
    n1953,
    n1701,
    n1718,
    n1745,
    n1682
  );


  nand
  g1911
  (
    n1874,
    n1573,
    n1562,
    n1743,
    n1726
  );


  nand
  g1912
  (
    n1911,
    n1841,
    n1685,
    n1821,
    n1751
  );


  nor
  g1913
  (
    n1882,
    n1757,
    n1823,
    n1791,
    n1712
  );


  xor
  g1914
  (
    n2029,
    n1706,
    n1720,
    n1668,
    n1830
  );


  nor
  g1915
  (
    n1875,
    n1766,
    n1764,
    n1696,
    n1771
  );


  or
  g1916
  (
    n1949,
    n1721,
    n1829,
    n1719,
    n1786
  );


  xor
  g1917
  (
    n1946,
    n1714,
    n1619,
    n1734,
    n1723
  );


  nand
  g1918
  (
    n1912,
    n1821,
    n1586,
    n1593,
    n1768
  );


  xor
  g1919
  (
    n1914,
    n1743,
    n1797,
    n1795,
    n1730
  );


  or
  g1920
  (
    n1866,
    n1687,
    n1718,
    n1708,
    n1686
  );


  xor
  g1921
  (
    n1863,
    n1680,
    n1790,
    n1817,
    n1800
  );


  or
  g1922
  (
    n2019,
    n1771,
    n1749,
    n1841,
    n1804
  );


  xnor
  g1923
  (
    n1862,
    n1739,
    n1656,
    n1733,
    n1640
  );


  xor
  g1924
  (
    n1997,
    n1720,
    n1774,
    n1576,
    n1633
  );


  nor
  g1925
  (
    n1995,
    n1776,
    n1638,
    n1803,
    n1761
  );


  nor
  g1926
  (
    n1923,
    n1825,
    n1726,
    n1705,
    n1756
  );


  or
  g1927
  (
    n1979,
    n1623,
    n1667,
    n1728,
    n1745
  );


  nand
  g1928
  (
    n1871,
    n1787,
    n1669,
    n1700,
    n1824
  );


  nor
  g1929
  (
    n1857,
    n1765,
    n1724,
    n1818,
    n1703
  );


  xor
  g1930
  (
    n1896,
    n1685,
    n1728,
    n1758,
    n1732
  );


  and
  g1931
  (
    n1927,
    n1700,
    n1791,
    n1843,
    n1583
  );


  nand
  g1932
  (
    n1904,
    n1840,
    n1779,
    n1828,
    n1689
  );


  and
  g1933
  (
    n1993,
    n1695,
    n1773,
    n1836,
    n1715
  );


  xor
  g1934
  (
    n1854,
    n1662,
    n1736,
    n1766,
    n1810
  );


  xor
  g1935
  (
    n1870,
    n1711,
    n1729,
    n1837,
    n1775
  );


  or
  g1936
  (
    n1998,
    n1823,
    n1694,
    n1717,
    n1822
  );


  nor
  g1937
  (
    n1976,
    n1718,
    n1745,
    n1806,
    n1769
  );


  nor
  g1938
  (
    n1852,
    n1759,
    n1772,
    n1600,
    n1819
  );


  nand
  g1939
  (
    n1864,
    n1559,
    n1823,
    n1763,
    n1810
  );


  or
  g1940
  (
    n1967,
    n1764,
    n1822,
    n1789,
    n1829
  );


  nand
  g1941
  (
    n1989,
    n1746,
    n1655,
    n1735,
    n1713
  );


  nor
  g1942
  (
    n1984,
    n1724,
    n1816,
    n1641
  );


  or
  g1943
  (
    n1884,
    n1636,
    n1578,
    n1710,
    n1601
  );


  xor
  g1944
  (
    n2003,
    n1697,
    n1666,
    n1732,
    n1728
  );


  xnor
  g1945
  (
    n1970,
    n1825,
    n1764,
    n1763,
    n1708
  );


  xor
  g1946
  (
    n1952,
    n1733,
    n1682,
    n1760,
    n1697
  );


  xor
  g1947
  (
    n1894,
    n1770,
    n1591,
    n1776,
    n1764
  );


  or
  g1948
  (
    n1922,
    n1832,
    n1561,
    n1767,
    n1625
  );


  and
  g1949
  (
    n1899,
    n1774,
    n1612,
    n1794,
    n1770
  );


  nor
  g1950
  (
    n1851,
    n1722,
    n1765,
    n1802,
    n1658
  );


  nor
  g1951
  (
    n1907,
    n1793,
    n1796,
    n1812,
    n1846
  );


  xor
  g1952
  (
    n2030,
    n1762,
    n1609,
    n1585,
    n1748
  );


  xor
  g1953
  (
    n1951,
    n1807,
    n1753,
    n1796,
    n1592
  );


  nand
  g1954
  (
    n2013,
    n1639,
    n1749,
    n1721,
    n1821
  );


  xnor
  g1955
  (
    n1913,
    n1704,
    n1644,
    n1828,
    n1714
  );


  nand
  g1956
  (
    n1876,
    n1757,
    n1744,
    n605,
    n1720
  );


  nand
  g1957
  (
    n1868,
    n1750,
    n1748,
    n1704,
    n1792
  );


  and
  g1958
  (
    n1903,
    n1701,
    n1831,
    n1707,
    n1752
  );


  nand
  g1959
  (
    n1858,
    n1750,
    n1683,
    n1813,
    n1827
  );


  and
  g1960
  (
    n1965,
    n1657,
    n1806,
    n1827,
    n1642
  );


  nor
  g1961
  (
    n1919,
    n1707,
    n1793,
    n1674,
    n1837
  );


  or
  g1962
  (
    n1902,
    n1768,
    n1839,
    n1799,
    n1665
  );


  or
  g1963
  (
    n1880,
    n1787,
    n1721,
    n1727,
    n1805
  );


  or
  g1964
  (
    n1906,
    n1801,
    n1842,
    n1564,
    n1687
  );


  nand
  g1965
  (
    n1992,
    n1570,
    n1701,
    n1790,
    n1795
  );


  xor
  g1966
  (
    n1966,
    n1654,
    n1813,
    n1735,
    n1738
  );


  xnor
  g1967
  (
    n2000,
    n1835,
    n1684,
    n1588,
    n1779
  );


  and
  g1968
  (
    n1939,
    n1722,
    n1807,
    n1775,
    n1822
  );


  nor
  g1969
  (
    n1973,
    n1779,
    n1774,
    n1660,
    n1729
  );


  nand
  g1970
  (
    n1878,
    n1759,
    n1762,
    n1665,
    n1833
  );


  nor
  g1971
  (
    n1853,
    n1782,
    n1831,
    n1845,
    n1622
  );


  xor
  g1972
  (
    n1942,
    n1777,
    n1727,
    n1615,
    n1781
  );


  nand
  g1973
  (
    n1941,
    n1758,
    n1634,
    n1711,
    n1834
  );


  xnor
  g1974
  (
    n1931,
    n1747,
    n1681,
    n1618,
    n1684
  );


  nand
  g1975
  (
    n1933,
    n1671,
    n1777,
    n1842,
    n1579
  );


  nand
  g1976
  (
    n1855,
    n1690,
    n1752,
    n1804,
    n1815
  );


  nand
  g1977
  (
    n1944,
    n1757,
    n1758,
    n1580,
    n1771
  );


  and
  g1978
  (
    n1959,
    n1768,
    n1572,
    n1788,
    n1629
  );


  nand
  g1979
  (
    n1897,
    n1836,
    n1778,
    n1824,
    n1595
  );


  nand
  g1980
  (
    n1924,
    n1829,
    n1740,
    n1735,
    n1844
  );


  nor
  g1981
  (
    n2020,
    n1832,
    n1817,
    n1835,
    n1793
  );


  and
  g1982
  (
    n1981,
    n1630,
    n1760,
    n1716,
    n1740
  );


  nor
  g1983
  (
    n1978,
    n1805,
    n1731,
    n1749,
    n1566
  );


  and
  g1984
  (
    n1921,
    n1741,
    n1840,
    n1842,
    n1782
  );


  and
  g1985
  (
    n1999,
    n1841,
    n1754,
    n1577,
    n1698
  );


  nand
  g1986
  (
    n2022,
    n1696,
    n1719,
    n1785,
    n1798
  );


  xor
  g1987
  (
    n1859,
    n1719,
    n1844,
    n1743,
    n1818
  );


  or
  g1988
  (
    n1940,
    n1773,
    n1761,
    n1702,
    n1748
  );


  xor
  g1989
  (
    n2016,
    n1799,
    n1729,
    n1678,
    n1689
  );


  or
  g1990
  (
    n1888,
    n1738,
    n1809,
    n1846,
    n1836
  );


  and
  g1991
  (
    n1900,
    n1746,
    n1733,
    n1734,
    n1806
  );


  or
  g1992
  (
    n1985,
    n1751,
    n1805,
    n1797,
    n1637
  );


  and
  g1993
  (
    n2025,
    n1792,
    n1731,
    n1801,
    n1835
  );


  nor
  g1994
  (
    KeyWire_0_16,
    n1767,
    n1695,
    n1817,
    n1690
  );


  xnor
  g1995
  (
    KeyWire_0_17,
    n1742,
    n1716,
    n1770,
    n1834
  );


  xor
  g1996
  (
    n1930,
    n1722,
    n1755,
    n1794,
    n1796
  );


  nand
  g1997
  (
    n1969,
    n1783,
    n1725,
    n1744,
    n1697
  );


  nand
  g1998
  (
    n1890,
    n1791,
    n1802,
    n1845,
    n1770
  );


  nor
  g1999
  (
    n1879,
    n1669,
    n1820,
    n1834,
    n1759
  );


  nand
  g2000
  (
    n1887,
    n1673,
    n1677,
    n1713,
    n1808
  );


  nor
  g2001
  (
    n2035,
    n1675,
    n1747,
    n1821,
    n1742
  );


  or
  g2002
  (
    n1968,
    n1832,
    n1691,
    n1804,
    n1788
  );


  nand
  g2003
  (
    n2017,
    n1602,
    n1672,
    n1678,
    n1755
  );


  xnor
  g2004
  (
    n1918,
    n1845,
    n1784,
    n1813,
    n1737
  );


  xnor
  g2005
  (
    n1948,
    n1762,
    n1746,
    n1785
  );


  and
  g2006
  (
    n1872,
    n1747,
    n1814,
    n1710,
    n1732
  );


  nand
  g2007
  (
    n1895,
    n1734,
    n1789,
    n1710,
    n1756
  );


  or
  g2008
  (
    n2082,
    n1849,
    n1922,
    n2028,
    n1911
  );


  nand
  g2009
  (
    n2062,
    n1951,
    n1933,
    n1909,
    n1955
  );


  or
  g2010
  (
    n2043,
    n1857,
    n1937,
    n2029,
    n1938
  );


  nand
  g2011
  (
    n2047,
    n1917,
    n1956,
    n1866,
    n2032
  );


  nor
  g2012
  (
    n2080,
    n2022,
    n2026,
    n1981,
    n1993
  );


  nor
  g2013
  (
    n2045,
    n2015,
    n2018,
    n1996,
    n1847
  );


  or
  g2014
  (
    n2070,
    n1998,
    n1930,
    n1855,
    n1876
  );


  nor
  g2015
  (
    n2063,
    n2021,
    n1910,
    n1905,
    n1990
  );


  and
  g2016
  (
    n2064,
    n1897,
    n1851,
    n2008,
    n1874
  );


  xor
  g2017
  (
    n2054,
    n1952,
    n1870,
    n1880,
    n1900
  );


  xor
  g2018
  (
    n2059,
    n1966,
    n1853,
    n2009,
    n1946
  );


  nor
  g2019
  (
    n2069,
    n1976,
    n1877,
    n1878,
    n2030
  );


  and
  g2020
  (
    n2056,
    n1929,
    n1901,
    n1924,
    n1859
  );


  and
  g2021
  (
    n2068,
    n1919,
    n1983,
    n1931,
    n1899
  );


  xnor
  g2022
  (
    n2049,
    n1989,
    n1982,
    n1960,
    n1967
  );


  and
  g2023
  (
    n2042,
    n1949,
    n1892,
    n1872,
    n1973
  );


  and
  g2024
  (
    n2084,
    n1896,
    n1894,
    n1945,
    n1913
  );


  nor
  g2025
  (
    n2057,
    n1860,
    n1869,
    n2000,
    n1898
  );


  or
  g2026
  (
    n2053,
    n1974,
    n1939,
    n2016,
    n1915
  );


  nor
  g2027
  (
    n2065,
    n1965,
    n1882,
    n2038,
    n1959
  );


  or
  g2028
  (
    n2071,
    n1902,
    n2013,
    n1958,
    n1980
  );


  and
  g2029
  (
    n2081,
    n1884,
    n2020,
    n1888,
    n2014
  );


  and
  g2030
  (
    n2076,
    n2036,
    n1883,
    n1927,
    n1948
  );


  xnor
  g2031
  (
    n2061,
    n1963,
    n1991,
    n2023,
    n1947
  );


  and
  g2032
  (
    n2039,
    n2034,
    n2027,
    n1992,
    n2033
  );


  nor
  g2033
  (
    n2085,
    n1848,
    n1916,
    n1932,
    n1925
  );


  nor
  g2034
  (
    n2051,
    n1968,
    n1864,
    n1923,
    n1986
  );


  nor
  g2035
  (
    KeyWire_0_12,
    n1858,
    n2019,
    n1904,
    n1926
  );


  xor
  g2036
  (
    n2074,
    n1865,
    n1994,
    n1850,
    n1940
  );


  or
  g2037
  (
    n2078,
    n1962,
    n2024,
    n2002,
    n1891
  );


  or
  g2038
  (
    n2040,
    n1914,
    n1988,
    n2037,
    n1997
  );


  or
  g2039
  (
    n2055,
    n1912,
    n2010,
    n1979,
    n2005
  );


  xor
  g2040
  (
    n2050,
    n1887,
    n1935,
    n1999,
    n1920
  );


  xor
  g2041
  (
    n2083,
    n1985,
    n1953,
    n1944,
    n1928
  );


  nand
  g2042
  (
    n2067,
    n2001,
    n1995,
    n1954,
    n1941
  );


  nor
  g2043
  (
    n2041,
    n2011,
    n1881,
    n1868,
    n1978
  );


  nand
  g2044
  (
    n2066,
    n1971,
    n1936,
    n1934,
    n1903
  );


  nand
  g2045
  (
    n2046,
    n1889,
    n1918,
    n1984,
    n1852
  );


  nor
  g2046
  (
    n2077,
    n1969,
    n1908,
    n1921,
    n1890
  );


  xnor
  g2047
  (
    n2075,
    n1871,
    n1975,
    n1893,
    n1907
  );


  xor
  g2048
  (
    n2058,
    n1862,
    n1863,
    n1970,
    n2035
  );


  xor
  g2049
  (
    n2072,
    n2025,
    n1856,
    n2004,
    n1964
  );


  nor
  g2050
  (
    n2086,
    n1987,
    n1943,
    n1875,
    n1885
  );


  nand
  g2051
  (
    n2060,
    n1972,
    n2017,
    n2007,
    n2031
  );


  or
  g2052
  (
    n2044,
    n2012,
    n1879,
    n1950,
    n1942
  );


  or
  g2053
  (
    n2052,
    n1961,
    n1854,
    n1861,
    n1895
  );


  nand
  g2054
  (
    n2048,
    n1873,
    n1977,
    n2003,
    n1906
  );


  or
  g2055
  (
    n2073,
    n1886,
    n1867,
    n1957,
    n2006
  );


  nor
  g2056
  (
    n2095,
    n2052,
    n2049,
    n2068,
    n2054
  );


  xor
  g2057
  (
    n2089,
    n2070,
    n2060,
    n2083,
    n2074
  );


  or
  g2058
  (
    n2093,
    n2045,
    n2085,
    n2081,
    n2067
  );


  nor
  g2059
  (
    n2094,
    n2069,
    n2039,
    n2061,
    n2077
  );


  nand
  g2060
  (
    n2091,
    n2062,
    n2056,
    n2058,
    n2053
  );


  xnor
  g2061
  (
    n2098,
    n2047,
    n2059,
    n2046,
    n2066
  );


  xnor
  g2062
  (
    n2088,
    n2065,
    n2073,
    n2048,
    n2044
  );


  or
  g2063
  (
    n2096,
    n2076,
    n2086,
    n2043,
    n2078
  );


  nand
  g2064
  (
    n2092,
    n2084,
    n2051,
    n2050,
    n2072
  );


  nor
  g2065
  (
    n2087,
    n2041,
    n2082,
    n2055,
    n2080
  );


  xor
  g2066
  (
    n2090,
    n2064,
    n2075,
    n2063,
    n2079
  );


  xor
  g2067
  (
    n2097,
    n2057,
    n2042,
    n2071,
    n2040
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1160,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n756,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n48,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1565,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n269,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n613,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1673,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1589,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n339,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n347,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n947,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1273,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n2079,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1105,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1168,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n82,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n1972,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n2012,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n634,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n351,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n968,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n40,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n105,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n1725,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n1708,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1711,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n410,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1971,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n918,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1269,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n235,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1285,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

