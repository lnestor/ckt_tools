

module Stat_277_639
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n298,
  n293,
  n286,
  n291,
  n282,
  n294,
  n283,
  n296,
  n278,
  n287,
  n288,
  n279,
  n280,
  n276,
  n295,
  n277,
  n290,
  n281,
  n284,
  n285,
  n275,
  n289,
  n292,
  n297
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n298;output n293;output n286;output n291;output n282;output n294;output n283;output n296;output n278;output n287;output n288;output n279;output n280;output n276;output n295;output n277;output n290;output n281;output n284;output n285;output n275;output n289;output n292;output n297;
  wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    n22,
    n5
  );


  buf
  g1
  (
    n24,
    n2
  );


  not
  g2
  (
    n25,
    n1
  );


  not
  g3
  (
    n26,
    n4
  );


  not
  g4
  (
    n23,
    n3
  );


  not
  g5
  (
    n38,
    n25
  );


  not
  g6
  (
    KeyWire_0_59,
    n24
  );


  not
  g7
  (
    n43,
    n23
  );


  not
  g8
  (
    n37,
    n25
  );


  buf
  g9
  (
    n32,
    n23
  );


  buf
  g10
  (
    n36,
    n26
  );


  not
  g11
  (
    n33,
    n26
  );


  buf
  g12
  (
    n30,
    n24
  );


  buf
  g13
  (
    KeyWire_0_44,
    n23
  );


  buf
  g14
  (
    n42,
    n26
  );


  not
  g15
  (
    n29,
    n26
  );


  buf
  g16
  (
    n35,
    n24
  );


  not
  g17
  (
    n40,
    n25
  );


  not
  g18
  (
    n28,
    n24
  );


  not
  g19
  (
    n31,
    n23
  );


  buf
  g20
  (
    KeyWire_0_24,
    n25
  );


  buf
  g21
  (
    KeyWire_0_54,
    n22
  );


  not
  g22
  (
    n62,
    n30
  );


  not
  g23
  (
    n86,
    n32
  );


  buf
  g24
  (
    n57,
    n39
  );


  not
  g25
  (
    n88,
    n31
  );


  buf
  g26
  (
    n69,
    n43
  );


  buf
  g27
  (
    n102,
    n28
  );


  buf
  g28
  (
    n50,
    n36
  );


  buf
  g29
  (
    n96,
    n41
  );


  buf
  g30
  (
    n58,
    n33
  );


  not
  g31
  (
    n56,
    n42
  );


  buf
  g32
  (
    n71,
    n39
  );


  not
  g33
  (
    n98,
    n33
  );


  not
  g34
  (
    n45,
    n29
  );


  buf
  g35
  (
    n59,
    n42
  );


  buf
  g36
  (
    n55,
    n28
  );


  not
  g37
  (
    n68,
    n30
  );


  buf
  g38
  (
    n66,
    n30
  );


  buf
  g39
  (
    n78,
    n37
  );


  not
  g40
  (
    KeyWire_0_28,
    n43
  );


  buf
  g41
  (
    n99,
    n43
  );


  not
  g42
  (
    n95,
    n37
  );


  not
  g43
  (
    n87,
    n33
  );


  not
  g44
  (
    n63,
    n27
  );


  buf
  g45
  (
    n67,
    n38
  );


  buf
  g46
  (
    n80,
    n39
  );


  buf
  g47
  (
    KeyWire_0_2,
    n31
  );


  not
  g48
  (
    n74,
    n29
  );


  buf
  g49
  (
    n54,
    n33
  );


  buf
  g50
  (
    n49,
    n38
  );


  not
  g51
  (
    n64,
    n40
  );


  not
  g52
  (
    n79,
    n32
  );


  not
  g53
  (
    KeyWire_0_20,
    n41
  );


  not
  g54
  (
    n103,
    n35
  );


  not
  g55
  (
    n92,
    n37
  );


  not
  g56
  (
    n46,
    n38
  );


  buf
  g57
  (
    KeyWire_0_62,
    n37
  );


  not
  g58
  (
    n82,
    n29
  );


  buf
  g59
  (
    n97,
    n28
  );


  not
  g60
  (
    KeyWire_0_30,
    n34
  );


  buf
  g61
  (
    n109,
    n41
  );


  not
  g62
  (
    KeyWire_0_55,
    n32
  );


  buf
  g63
  (
    n51,
    n42
  );


  buf
  g64
  (
    n85,
    n40
  );


  not
  g65
  (
    n81,
    n34
  );


  not
  g66
  (
    n72,
    n38
  );


  not
  g67
  (
    n110,
    n39
  );


  buf
  g68
  (
    n111,
    n34
  );


  buf
  g69
  (
    n108,
    n27
  );


  not
  g70
  (
    KeyWire_0_43,
    n31
  );


  not
  g71
  (
    KeyWire_0_21,
    n28
  );


  not
  g72
  (
    n100,
    n34
  );


  buf
  g73
  (
    n89,
    n27
  );


  not
  g74
  (
    n77,
    n40
  );


  buf
  g75
  (
    n47,
    n35
  );


  buf
  g76
  (
    n93,
    n30
  );


  buf
  g77
  (
    n75,
    n29
  );


  not
  g78
  (
    n83,
    n43
  );


  buf
  g79
  (
    n52,
    n27
  );


  buf
  g80
  (
    n73,
    n36
  );


  not
  g81
  (
    KeyWire_0_18,
    n41
  );


  buf
  g82
  (
    n61,
    n35
  );


  not
  g83
  (
    KeyWire_0_13,
    n35
  );


  not
  g84
  (
    KeyWire_0_46,
    n40
  );


  not
  g85
  (
    KeyWire_0_15,
    n42
  );


  buf
  g86
  (
    n106,
    n31
  );


  buf
  g87
  (
    KeyWire_0_38,
    n36
  );


  not
  g88
  (
    KeyWire_0_6,
    n32
  );


  buf
  g89
  (
    n91,
    n36
  );


  not
  g90
  (
    KeyWire_0_57,
    n95
  );


  buf
  g91
  (
    n189,
    n60
  );


  buf
  g92
  (
    n180,
    n68
  );


  not
  g93
  (
    n163,
    n76
  );


  not
  g94
  (
    n178,
    n84
  );


  not
  g95
  (
    n123,
    n65
  );


  not
  g96
  (
    n187,
    n84
  );


  buf
  g97
  (
    n193,
    n73
  );


  buf
  g98
  (
    n179,
    n100
  );


  buf
  g99
  (
    KeyWire_0_16,
    n74
  );


  not
  g100
  (
    n143,
    n19
  );


  buf
  g101
  (
    KeyWire_0_37,
    n10
  );


  not
  g102
  (
    n167,
    n67
  );


  nor
  g103
  (
    n130,
    n18,
    n51,
    n48
  );


  and
  g104
  (
    n171,
    n82,
    n81,
    n51,
    n52
  );


  nand
  g105
  (
    n185,
    n67,
    n73,
    n106,
    n89
  );


  and
  g106
  (
    n138,
    n17,
    n99,
    n60,
    n104
  );


  nand
  g107
  (
    n151,
    n87,
    n110,
    n55,
    n109
  );


  and
  g108
  (
    n141,
    n56,
    n61,
    n82,
    n90
  );


  nand
  g109
  (
    n118,
    n101,
    n51,
    n61,
    n106
  );


  nor
  g110
  (
    n152,
    n109,
    n75,
    n100
  );


  xor
  g111
  (
    n160,
    n74,
    n111,
    n96
  );


  xor
  g112
  (
    n135,
    n49,
    n56,
    n91,
    n97
  );


  or
  g113
  (
    n186,
    n93,
    n84,
    n65,
    n85
  );


  xor
  g114
  (
    n168,
    n46,
    n63,
    n75,
    n99
  );


  and
  g115
  (
    n117,
    n102,
    n59,
    n64,
    n65
  );


  or
  g116
  (
    n121,
    n83,
    n54,
    n76,
    n71
  );


  and
  g117
  (
    n166,
    n106,
    n81,
    n104,
    n108
  );


  xor
  g118
  (
    KeyWire_0_10,
    n108,
    n53,
    n16,
    n11
  );


  and
  g119
  (
    n164,
    n77,
    n54,
    n68,
    n21
  );


  xnor
  g120
  (
    n173,
    n45,
    n57,
    n44,
    n95
  );


  and
  g121
  (
    n176,
    n82,
    n47,
    n44,
    n85
  );


  nor
  g122
  (
    n153,
    n53,
    n69,
    n107,
    n68
  );


  xor
  g123
  (
    n139,
    n58,
    n108,
    n52,
    n103
  );


  and
  g124
  (
    n137,
    n51,
    n67,
    n110,
    n54
  );


  and
  g125
  (
    KeyWire_0_34,
    n80,
    n59,
    n53,
    n96
  );


  xor
  g126
  (
    n128,
    n103,
    n93,
    n72,
    n84
  );


  nand
  g127
  (
    n155,
    n94,
    n55,
    n79,
    n49
  );


  and
  g128
  (
    KeyWire_0_50,
    n95,
    n57,
    n99,
    n105
  );


  or
  g129
  (
    n142,
    n57,
    n89,
    n101,
    n88
  );


  xnor
  g130
  (
    n149,
    n94,
    n87,
    n95,
    n91
  );


  xnor
  g131
  (
    n182,
    n69,
    n66,
    n93,
    n92
  );


  or
  g132
  (
    n136,
    n64,
    n100,
    n13,
    n54
  );


  nand
  g133
  (
    n114,
    n71,
    n111,
    n62,
    n58
  );


  xnor
  g134
  (
    n133,
    n97,
    n48,
    n109,
    n90
  );


  and
  g135
  (
    n165,
    n64,
    n111,
    n50,
    n62
  );


  xnor
  g136
  (
    n190,
    n46,
    n75,
    n63,
    n66
  );


  nand
  g137
  (
    n144,
    n91,
    n49,
    n69,
    n87
  );


  xnor
  g138
  (
    n156,
    n62,
    n80,
    n73,
    n74
  );


  nand
  g139
  (
    n112,
    n98,
    n7,
    n105,
    n89
  );


  or
  g140
  (
    n159,
    n109,
    n50,
    n70,
    n90
  );


  and
  g141
  (
    n140,
    n102,
    n92,
    n48,
    n104
  );


  xor
  g142
  (
    n175,
    n61,
    n68,
    n70,
    n97
  );


  nand
  g143
  (
    KeyWire_0_60,
    n50,
    n98,
    n77,
    n96
  );


  or
  g144
  (
    n177,
    n98,
    n107,
    n87,
    n81
  );


  nand
  g145
  (
    n131,
    n58,
    n79,
    n103,
    n45
  );


  nand
  g146
  (
    n174,
    n63,
    n8,
    n110,
    n60
  );


  xnor
  g147
  (
    n169,
    n88,
    n45,
    n102,
    n97
  );


  or
  g148
  (
    KeyWire_0_41,
    n103,
    n104,
    n83,
    n88
  );


  or
  g149
  (
    n146,
    n46,
    n49,
    n71,
    n59
  );


  xnor
  g150
  (
    KeyWire_0_11,
    n101,
    n12,
    n71,
    n85
  );


  nand
  g151
  (
    n129,
    n89,
    n60,
    n83,
    n86
  );


  xnor
  g152
  (
    n116,
    n52,
    n45,
    n98,
    n66
  );


  xor
  g153
  (
    n192,
    n99,
    n44,
    n80,
    n77
  );


  xor
  g154
  (
    KeyWire_0_39,
    n70,
    n79,
    n107,
    n72
  );


  nor
  g155
  (
    n191,
    n61,
    n108,
    n96,
    n107
  );


  xor
  g156
  (
    n134,
    n56,
    n86,
    n64,
    n79
  );


  xnor
  g157
  (
    n158,
    n110,
    n105,
    n70,
    n48
  );


  nor
  g158
  (
    KeyWire_0_7,
    n6,
    n58,
    n102,
    n59
  );


  or
  g159
  (
    n127,
    n77,
    n57,
    n55,
    n80
  );


  nor
  g160
  (
    n148,
    n74,
    n56,
    n72,
    n50
  );


  or
  g161
  (
    n172,
    n85,
    n55,
    n72,
    n106
  );


  xnor
  g162
  (
    KeyWire_0_35,
    n78,
    n67,
    n47,
    n92
  );


  and
  g163
  (
    KeyWire_0_36,
    n78,
    n91,
    n92,
    n65
  );


  xor
  g164
  (
    n113,
    n52,
    n82,
    n101,
    n90
  );


  and
  g165
  (
    n183,
    n66,
    n86,
    n46,
    n76
  );


  nand
  g166
  (
    n188,
    n83,
    n9,
    n20,
    n47
  );


  and
  g167
  (
    KeyWire_0_23,
    n76,
    n44,
    n53,
    n78
  );


  nand
  g168
  (
    n115,
    n94,
    n78,
    n93,
    n62
  );


  and
  g169
  (
    KeyWire_0_52,
    n100,
    n105,
    n47,
    n94
  );


  and
  g170
  (
    KeyWire_0_58,
    n69,
    n15,
    n63,
    n81
  );


  and
  g171
  (
    KeyWire_0_8,
    n88,
    n86,
    n73,
    n14
  );


  xor
  g172
  (
    KeyWire_0_33,
    n134,
    n179,
    n148,
    n144
  );


  nor
  g173
  (
    KeyWire_0_5,
    n126,
    n124,
    n150,
    n136
  );


  or
  g174
  (
    KeyWire_0_32,
    n180,
    n112,
    n146,
    n182
  );


  nand
  g175
  (
    n258,
    n145,
    n123,
    n133
  );


  and
  g176
  (
    KeyWire_0_47,
    n129,
    n154,
    n190,
    n146
  );


  nand
  g177
  (
    n210,
    n114,
    n157,
    n128,
    n178
  );


  and
  g178
  (
    KeyWire_0_9,
    n182,
    n173,
    n162,
    n141
  );


  xnor
  g179
  (
    n268,
    n163,
    n166,
    n158,
    n134
  );


  nand
  g180
  (
    KeyWire_0_14,
    n193,
    n172,
    n158,
    n177
  );


  xnor
  g181
  (
    n255,
    n174,
    n188,
    n159,
    n138
  );


  xnor
  g182
  (
    n260,
    n123,
    n168,
    n169
  );


  or
  g183
  (
    n274,
    n168,
    n151,
    n164,
    n130
  );


  and
  g184
  (
    n197,
    n156,
    n178,
    n190,
    n159
  );


  nor
  g185
  (
    KeyWire_0_49,
    n173,
    n152,
    n135,
    n141
  );


  xor
  g186
  (
    n254,
    n126,
    n113,
    n130,
    n158
  );


  or
  g187
  (
    n236,
    n141,
    n165,
    n183,
    n137
  );


  xnor
  g188
  (
    KeyWire_0_56,
    n192,
    n124,
    n166,
    n119
  );


  xor
  g189
  (
    n219,
    n120,
    n152,
    n142,
    n155
  );


  and
  g190
  (
    n223,
    n170,
    n167,
    n136,
    n187
  );


  xnor
  g191
  (
    KeyWire_0_42,
    n184,
    n118,
    n153,
    n120
  );


  nand
  g192
  (
    n246,
    n177,
    n188,
    n131,
    n141
  );


  xor
  g193
  (
    n238,
    n176,
    n157,
    n114,
    n190
  );


  nor
  g194
  (
    n213,
    n138,
    n127,
    n120,
    n152
  );


  nor
  g195
  (
    KeyWire_0_17,
    n176,
    n140,
    n118,
    n189
  );


  nand
  g196
  (
    KeyWire_0_45,
    n185,
    n155,
    n179,
    n118
  );


  nand
  g197
  (
    KeyWire_0_22,
    n155,
    n123,
    n163,
    n149
  );


  and
  g198
  (
    n257,
    n191,
    n124,
    n116,
    n164
  );


  and
  g199
  (
    n270,
    n174,
    n179,
    n125
  );


  nor
  g200
  (
    n198,
    n161,
    n139,
    n174,
    n175
  );


  or
  g201
  (
    n202,
    n192,
    n139,
    n134,
    n115
  );


  or
  g202
  (
    KeyWire_0_48,
    n177,
    n165,
    n147,
    n128
  );


  xnor
  g203
  (
    KeyWire_0_3,
    n186,
    n164,
    n122,
    n157
  );


  nand
  g204
  (
    n229,
    n132,
    n186,
    n176,
    n169
  );


  nor
  g205
  (
    n200,
    n177,
    n150,
    n162,
    n185
  );


  nor
  g206
  (
    n206,
    n130,
    n136,
    n173,
    n134
  );


  xnor
  g207
  (
    n269,
    n116,
    n131,
    n150,
    n187
  );


  xnor
  g208
  (
    n194,
    n186,
    n183,
    n163,
    n148
  );


  nand
  g209
  (
    KeyWire_0_53,
    n140,
    n138,
    n178,
    n121
  );


  nand
  g210
  (
    n195,
    n185,
    n140,
    n168,
    n143
  );


  and
  g211
  (
    n271,
    n173,
    n132,
    n191,
    n167
  );


  xnor
  g212
  (
    n240,
    n135,
    n162,
    n159,
    n164
  );


  and
  g213
  (
    n272,
    n147,
    n122,
    n145,
    n139
  );


  xnor
  g214
  (
    n261,
    n138,
    n157,
    n137,
    n156
  );


  nor
  g215
  (
    n273,
    n151,
    n175,
    n149,
    n126
  );


  and
  g216
  (
    n263,
    n137,
    n171,
    n121,
    n182
  );


  xnor
  g217
  (
    n211,
    n158,
    n130,
    n190,
    n170
  );


  nor
  g218
  (
    n199,
    n113,
    n115,
    n125,
    n117
  );


  or
  g219
  (
    KeyWire_0_26,
    n142,
    n175,
    n181,
    n131
  );


  nor
  g220
  (
    KeyWire_0_31,
    n156,
    n128,
    n115,
    n132
  );


  xor
  g221
  (
    n247,
    n153,
    n118,
    n182,
    n167
  );


  and
  g222
  (
    n244,
    n115,
    n116,
    n117,
    n163
  );


  or
  g223
  (
    n208,
    n144,
    n180,
    n187,
    n148
  );


  or
  g224
  (
    n231,
    n161,
    n184,
    n127,
    n135
  );


  and
  g225
  (
    KeyWire_0_0,
    n125,
    n170,
    n127,
    n168
  );


  xor
  g226
  (
    n265,
    n122,
    n181,
    n136,
    n189
  );


  or
  g227
  (
    n242,
    n161,
    n176,
    n147,
    n124
  );


  xnor
  g228
  (
    n221,
    n191,
    n183,
    n154,
    n178
  );


  nor
  g229
  (
    n256,
    n119,
    n133,
    n151,
    n117
  );


  xor
  g230
  (
    n205,
    n171,
    n172,
    n142
  );


  nor
  g231
  (
    KeyWire_0_51,
    n160,
    n148,
    n152,
    n156
  );


  xnor
  g232
  (
    n204,
    n160,
    n169,
    n143,
    n180
  );


  or
  g233
  (
    n226,
    n112,
    n189,
    n193,
    n174
  );


  or
  g234
  (
    KeyWire_0_19,
    n123,
    n145,
    n181,
    n140
  );


  nand
  g235
  (
    n214,
    n160,
    n116,
    n165,
    n143
  );


  or
  g236
  (
    n232,
    n131,
    n150,
    n146,
    n132
  );


  nor
  g237
  (
    n234,
    n129,
    n167,
    n153,
    n149
  );


  nor
  g238
  (
    n245,
    n185,
    n137,
    n145,
    n192
  );


  xnor
  g239
  (
    n267,
    n122,
    n128,
    n184,
    n188
  );


  nor
  g240
  (
    n230,
    n126,
    n186,
    n188,
    n159
  );


  and
  g241
  (
    n222,
    n192,
    n135,
    n147,
    n149
  );


  xnor
  g242
  (
    n209,
    n144,
    n129,
    n121,
    n191
  );


  xnor
  g243
  (
    KeyWire_0_27,
    n139,
    n143,
    n161,
    n119
  );


  or
  g244
  (
    n259,
    n153,
    n187,
    n183,
    n142
  );


  nor
  g245
  (
    n264,
    n184,
    n189,
    n170,
    n144
  );


  nor
  g246
  (
    n228,
    n165,
    n119,
    n151,
    n114
  );


  or
  g247
  (
    n237,
    n180,
    n146,
    n155,
    n166
  );


  nor
  g248
  (
    n225,
    n162,
    n175,
    n121,
    n193
  );


  xnor
  g249
  (
    n207,
    n127,
    n171,
    n129,
    n133
  );


  xnor
  g250
  (
    n243,
    n193,
    n120,
    n154,
    n114
  );


  and
  g251
  (
    n201,
    n181,
    n172,
    n171,
    n166
  );


  xor
  g252
  (
    n216,
    n117,
    n160,
    n154,
    n125
  );


  nand
  g253
  (
    n289,
    n197,
    n245,
    n216,
    n223
  );


  and
  g254
  (
    n276,
    n244,
    n208,
    n227,
    n273
  );


  nand
  g255
  (
    n293,
    n221,
    n203,
    n268,
    n194
  );


  or
  g256
  (
    KeyWire_0_12,
    n259,
    n254,
    n260,
    n246
  );


  xor
  g257
  (
    n278,
    n226,
    n261,
    n270,
    n235
  );


  xnor
  g258
  (
    n294,
    n272,
    n270,
    n266,
    n198
  );


  or
  g259
  (
    KeyWire_0_61,
    n204,
    n220,
    n217,
    n239
  );


  nor
  g260
  (
    n295,
    n222,
    n236,
    n256,
    n196
  );


  xnor
  g261
  (
    n290,
    n257,
    n232,
    n247,
    n274
  );


  nand
  g262
  (
    n286,
    n215,
    n274,
    n266,
    n269
  );


  xnor
  g263
  (
    KeyWire_0_1,
    n234,
    n201,
    n274,
    n233
  );


  xnor
  g264
  (
    KeyWire_0_29,
    n241,
    n264,
    n250,
    n253
  );


  and
  g265
  (
    n285,
    n212,
    n238,
    n224,
    n248
  );


  nor
  g266
  (
    KeyWire_0_40,
    n249,
    n252,
    n210,
    n265
  );


  xor
  g267
  (
    KeyWire_0_4,
    n195,
    n240,
    n225,
    n205
  );


  xor
  g268
  (
    n284,
    n264,
    n262,
    n219,
    n206
  );


  xor
  g269
  (
    n287,
    n267,
    n237,
    n200,
    n271
  );


  or
  g270
  (
    n288,
    n262,
    n230,
    n213,
    n263
  );


  nor
  g271
  (
    KeyWire_0_25,
    n229,
    n218,
    n265,
    n211
  );


  xor
  g272
  (
    n280,
    n272,
    n268,
    n274,
    n271
  );


  nand
  g273
  (
    n281,
    n251,
    n202,
    n269,
    n267
  );


  or
  g274
  (
    KeyWire_0_63,
    n207,
    n228,
    n209,
    n214
  );


  xnor
  g275
  (
    n279,
    n255,
    n263,
    n258,
    n242
  );


  and
  g276
  (
    n297,
    n199,
    n243,
    n231,
    n273
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n203,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n275,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n101,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n249,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n296,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n212,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n105,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n150,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n122,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n252,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n124,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n154,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n298,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n65,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n220,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n48,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n125,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n241,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n76,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n224,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n44,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n107,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n235,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n145,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n27,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n277,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n196,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n251,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n60,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n291,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n94,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n248,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n218,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n217,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n147,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n126,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n161,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n120,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n90,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n157,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n292,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n119,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n239,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n104,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n34,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n253,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n70,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n215,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n250,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n233,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n184,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n262,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n162,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n266,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n41,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n53,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n227,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n181,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n170,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n39,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n132,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n282,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n84,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n283,
    KeyNOTWire_0_63
  );


endmodule


