

module Stat_1000_156
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1023,
  n1025,
  n1006,
  n1013,
  n1030,
  n1002,
  n1016,
  n1011,
  n1022,
  n1014,
  n1027,
  n1019,
  n1018,
  n1004,
  n1028,
  n1005,
  n1008,
  n1026,
  n1001,
  n1021,
  n1029,
  n1012,
  n1032,
  n1031,
  n1003,
  n1017,
  n1010,
  n1007,
  n1024,
  n1015,
  n1009,
  n1020,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1023;output n1025;output n1006;output n1013;output n1030;output n1002;output n1016;output n1011;output n1022;output n1014;output n1027;output n1019;output n1018;output n1004;output n1028;output n1005;output n1008;output n1026;output n1001;output n1021;output n1029;output n1012;output n1032;output n1031;output n1003;output n1017;output n1010;output n1007;output n1024;output n1015;output n1009;output n1020;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n68,
    n1
  );


  not
  g1
  (
    n109,
    n4
  );


  not
  g2
  (
    n95,
    n8
  );


  not
  g3
  (
    n89,
    n17
  );


  buf
  g4
  (
    n111,
    n13
  );


  not
  g5
  (
    n74,
    n18
  );


  not
  g6
  (
    n110,
    n18
  );


  not
  g7
  (
    n49,
    n13
  );


  not
  g8
  (
    n57,
    n16
  );


  buf
  g9
  (
    n54,
    n7
  );


  not
  g10
  (
    n35,
    n24
  );


  buf
  g11
  (
    n102,
    n5
  );


  not
  g12
  (
    n71,
    n4
  );


  buf
  g13
  (
    n59,
    n20
  );


  not
  g14
  (
    n77,
    n16
  );


  not
  g15
  (
    n56,
    n23
  );


  not
  g16
  (
    n86,
    n26
  );


  not
  g17
  (
    n70,
    n7
  );


  not
  g18
  (
    n94,
    n10
  );


  buf
  g19
  (
    n48,
    n8
  );


  not
  g20
  (
    n63,
    n12
  );


  not
  g21
  (
    n60,
    n6
  );


  buf
  g22
  (
    n55,
    n4
  );


  buf
  g23
  (
    n88,
    n3
  );


  buf
  g24
  (
    n38,
    n13
  );


  not
  g25
  (
    n87,
    n9
  );


  not
  g26
  (
    n66,
    n26
  );


  not
  g27
  (
    n42,
    n11
  );


  buf
  g28
  (
    n84,
    n4
  );


  not
  g29
  (
    n79,
    n8
  );


  not
  g30
  (
    n81,
    n25
  );


  buf
  g31
  (
    n46,
    n9
  );


  buf
  g32
  (
    n58,
    n1
  );


  not
  g33
  (
    n34,
    n24
  );


  buf
  g34
  (
    n96,
    n18
  );


  buf
  g35
  (
    n33,
    n25
  );


  not
  g36
  (
    n51,
    n14
  );


  not
  g37
  (
    n104,
    n3
  );


  buf
  g38
  (
    n98,
    n12
  );


  buf
  g39
  (
    n40,
    n24
  );


  buf
  g40
  (
    n52,
    n16
  );


  not
  g41
  (
    n80,
    n11
  );


  not
  g42
  (
    n108,
    n25
  );


  buf
  g43
  (
    n75,
    n15
  );


  buf
  g44
  (
    n103,
    n6
  );


  buf
  g45
  (
    n39,
    n15
  );


  buf
  g46
  (
    n72,
    n26
  );


  not
  g47
  (
    n61,
    n7
  );


  buf
  g48
  (
    n100,
    n19
  );


  buf
  g49
  (
    n36,
    n16
  );


  buf
  g50
  (
    n83,
    n20
  );


  buf
  g51
  (
    n97,
    n21
  );


  buf
  g52
  (
    n90,
    n17
  );


  buf
  g53
  (
    n99,
    n22
  );


  not
  g54
  (
    n45,
    n13
  );


  buf
  g55
  (
    n44,
    n22
  );


  buf
  g56
  (
    n43,
    n27
  );


  buf
  g57
  (
    n64,
    n12
  );


  buf
  g58
  (
    n41,
    n12
  );


  not
  g59
  (
    n93,
    n6
  );


  buf
  g60
  (
    n47,
    n6
  );


  not
  g61
  (
    n53,
    n23
  );


  not
  g62
  (
    n106,
    n9
  );


  not
  g63
  (
    n91,
    n5
  );


  buf
  g64
  (
    n76,
    n1
  );


  not
  g65
  (
    n85,
    n3
  );


  not
  g66
  (
    n73,
    n2
  );


  buf
  g67
  (
    n37,
    n11
  );


  buf
  g68
  (
    n62,
    n9
  );


  buf
  g69
  (
    n78,
    n3
  );


  not
  g70
  (
    n65,
    n24
  );


  xnor
  g71
  (
    n107,
    n1,
    n23,
    n11
  );


  and
  g72
  (
    n101,
    n5,
    n15,
    n23
  );


  nor
  g73
  (
    n105,
    n21,
    n27,
    n19
  );


  or
  g74
  (
    n67,
    n21,
    n8,
    n10,
    n14
  );


  xnor
  g75
  (
    n82,
    n25,
    n20,
    n14,
    n17
  );


  xor
  g76
  (
    n50,
    n10,
    n18,
    n2,
    n21
  );


  or
  g77
  (
    n92,
    n19,
    n26,
    n14,
    n22
  );


  xor
  g78
  (
    n69,
    n2,
    n10,
    n5,
    n17
  );


  xor
  g79
  (
    n112,
    n22,
    n2,
    n20,
    n7
  );


  buf
  g80
  (
    n238,
    n48
  );


  not
  g81
  (
    n161,
    n68
  );


  buf
  g82
  (
    n145,
    n37
  );


  buf
  g83
  (
    n226,
    n93
  );


  not
  g84
  (
    n119,
    n107
  );


  not
  g85
  (
    n183,
    n53
  );


  buf
  g86
  (
    n160,
    n56
  );


  buf
  g87
  (
    n202,
    n95
  );


  buf
  g88
  (
    n115,
    n51
  );


  buf
  g89
  (
    n212,
    n38
  );


  not
  g90
  (
    n125,
    n104
  );


  not
  g91
  (
    n219,
    n85
  );


  buf
  g92
  (
    n193,
    n41
  );


  not
  g93
  (
    n120,
    n33
  );


  buf
  g94
  (
    n234,
    n104
  );


  not
  g95
  (
    n171,
    n76
  );


  buf
  g96
  (
    n124,
    n94
  );


  buf
  g97
  (
    n213,
    n87
  );


  not
  g98
  (
    n140,
    n49
  );


  not
  g99
  (
    n233,
    n110
  );


  buf
  g100
  (
    n116,
    n62
  );


  buf
  g101
  (
    n200,
    n54
  );


  not
  g102
  (
    n228,
    n47
  );


  buf
  g103
  (
    n205,
    n75
  );


  buf
  g104
  (
    n242,
    n102
  );


  buf
  g105
  (
    n169,
    n78
  );


  buf
  g106
  (
    n209,
    n96
  );


  buf
  g107
  (
    n184,
    n52
  );


  buf
  g108
  (
    n144,
    n89
  );


  buf
  g109
  (
    n166,
    n109
  );


  buf
  g110
  (
    n173,
    n47
  );


  buf
  g111
  (
    n240,
    n65
  );


  buf
  g112
  (
    n231,
    n73
  );


  not
  g113
  (
    n186,
    n40
  );


  not
  g114
  (
    n117,
    n51
  );


  buf
  g115
  (
    n187,
    n76
  );


  not
  g116
  (
    n154,
    n95
  );


  buf
  g117
  (
    n182,
    n64
  );


  not
  g118
  (
    n135,
    n87
  );


  buf
  g119
  (
    n156,
    n56
  );


  nor
  g120
  (
    n235,
    n35,
    n106,
    n100
  );


  xor
  g121
  (
    n153,
    n39,
    n86,
    n105
  );


  nor
  g122
  (
    n129,
    n59,
    n35,
    n60
  );


  xnor
  g123
  (
    n151,
    n72,
    n85,
    n74
  );


  nor
  g124
  (
    n114,
    n41,
    n35,
    n79
  );


  xnor
  g125
  (
    n163,
    n78,
    n52,
    n90
  );


  xor
  g126
  (
    n195,
    n60,
    n44,
    n103
  );


  nor
  g127
  (
    n147,
    n51,
    n101,
    n34
  );


  or
  g128
  (
    n152,
    n47,
    n105,
    n101
  );


  nor
  g129
  (
    n241,
    n58,
    n65,
    n92
  );


  nand
  g130
  (
    n201,
    n98,
    n108,
    n45
  );


  xnor
  g131
  (
    n220,
    n59,
    n80,
    n108
  );


  nand
  g132
  (
    n211,
    n54,
    n61,
    n83
  );


  and
  g133
  (
    n198,
    n58,
    n111,
    n63
  );


  and
  g134
  (
    n139,
    n97,
    n109,
    n53
  );


  nor
  g135
  (
    n142,
    n81,
    n73,
    n76
  );


  and
  g136
  (
    n168,
    n46,
    n52,
    n77
  );


  nor
  g137
  (
    n199,
    n84,
    n91,
    n72
  );


  nor
  g138
  (
    n237,
    n94,
    n83,
    n79
  );


  nand
  g139
  (
    n218,
    n55,
    n94,
    n44
  );


  nor
  g140
  (
    n123,
    n55,
    n99,
    n41
  );


  nand
  g141
  (
    n143,
    n80,
    n49,
    n33
  );


  and
  g142
  (
    n207,
    n71,
    n43,
    n35
  );


  or
  g143
  (
    n131,
    n60,
    n107,
    n98
  );


  nor
  g144
  (
    n172,
    n86,
    n68,
    n56
  );


  and
  g145
  (
    n224,
    n42,
    n98,
    n78
  );


  nand
  g146
  (
    n197,
    n81,
    n101,
    n69
  );


  nand
  g147
  (
    n146,
    n90,
    n105,
    n38
  );


  xnor
  g148
  (
    n157,
    n72,
    n99,
    n50
  );


  nor
  g149
  (
    n179,
    n57,
    n43,
    n91
  );


  nor
  g150
  (
    n150,
    n40,
    n75,
    n87
  );


  nor
  g151
  (
    n138,
    n82,
    n106,
    n54
  );


  nand
  g152
  (
    n158,
    n93,
    n81,
    n94
  );


  xor
  g153
  (
    n221,
    n103,
    n71,
    n72
  );


  xor
  g154
  (
    n181,
    n38,
    n89,
    n85
  );


  nor
  g155
  (
    n164,
    n65,
    n89,
    n109
  );


  or
  g156
  (
    n127,
    n62,
    n46,
    n42
  );


  or
  g157
  (
    n128,
    n33,
    n63,
    n40
  );


  nor
  g158
  (
    n149,
    n97,
    n39,
    n106
  );


  nor
  g159
  (
    n180,
    n66,
    n75,
    n83
  );


  and
  g160
  (
    n177,
    n62,
    n49,
    n45
  );


  nand
  g161
  (
    n133,
    n45,
    n100,
    n54
  );


  xnor
  g162
  (
    n239,
    n61,
    n36,
    n58
  );


  xor
  g163
  (
    n203,
    n55,
    n57,
    n41
  );


  xnor
  g164
  (
    n136,
    n104,
    n82,
    n101
  );


  nand
  g165
  (
    n204,
    n82,
    n80
  );


  xor
  g166
  (
    n122,
    n88,
    n40,
    n104
  );


  xnor
  g167
  (
    n196,
    n36,
    n34,
    n52
  );


  xor
  g168
  (
    n194,
    n76,
    n93
  );


  xor
  g169
  (
    n191,
    n62,
    n86,
    n49
  );


  nand
  g170
  (
    n225,
    n55,
    n64,
    n84
  );


  xnor
  g171
  (
    n165,
    n78,
    n77,
    n84
  );


  and
  g172
  (
    n227,
    n66,
    n88,
    n64
  );


  xnor
  g173
  (
    n132,
    n88,
    n71,
    n39
  );


  nand
  g174
  (
    n190,
    n60,
    n43,
    n103
  );


  nor
  g175
  (
    n170,
    n58,
    n33,
    n57
  );


  or
  g176
  (
    n230,
    n46,
    n103,
    n96
  );


  nand
  g177
  (
    n236,
    n57,
    n96,
    n48
  );


  xor
  g178
  (
    n175,
    n108,
    n107,
    n84
  );


  xor
  g179
  (
    n223,
    n81,
    n91,
    n70
  );


  xor
  g180
  (
    n141,
    n97,
    n110,
    n108
  );


  and
  g181
  (
    n134,
    n50,
    n102,
    n74
  );


  nor
  g182
  (
    n188,
    n53,
    n90,
    n64
  );


  nor
  g183
  (
    n206,
    n110,
    n96,
    n107
  );


  xor
  g184
  (
    n214,
    n39,
    n36,
    n67
  );


  nand
  g185
  (
    n118,
    n100,
    n51,
    n38
  );


  xnor
  g186
  (
    n189,
    n44,
    n110,
    n65
  );


  nand
  g187
  (
    n232,
    n66,
    n70,
    n73
  );


  or
  g188
  (
    n229,
    n53,
    n46,
    n61
  );


  xnor
  g189
  (
    n210,
    n36,
    n42,
    n69
  );


  and
  g190
  (
    n137,
    n92,
    n45,
    n88
  );


  nor
  g191
  (
    n243,
    n82,
    n86,
    n100
  );


  and
  g192
  (
    n222,
    n98,
    n77
  );


  xnor
  g193
  (
    n148,
    n67,
    n37,
    n63
  );


  nand
  g194
  (
    n217,
    n90,
    n70,
    n47
  );


  or
  g195
  (
    n121,
    n95,
    n105,
    n92
  );


  xor
  g196
  (
    n215,
    n102,
    n42,
    n106
  );


  xnor
  g197
  (
    n174,
    n75,
    n79,
    n85
  );


  and
  g198
  (
    n126,
    n59,
    n67
  );


  xor
  g199
  (
    n216,
    n56,
    n73,
    n66
  );


  nand
  g200
  (
    n167,
    n43,
    n63,
    n102
  );


  xor
  g201
  (
    n185,
    n48,
    n79,
    n71
  );


  or
  g202
  (
    n113,
    n99,
    n61,
    n74
  );


  nand
  g203
  (
    n192,
    n70,
    n95,
    n69
  );


  nand
  g204
  (
    n130,
    n92,
    n68,
    n34
  );


  xor
  g205
  (
    n178,
    n69,
    n50
  );


  nand
  g206
  (
    n176,
    n34,
    n59,
    n91
  );


  and
  g207
  (
    n162,
    n87,
    n37,
    n48
  );


  nand
  g208
  (
    n208,
    n68,
    n89,
    n99
  );


  xnor
  g209
  (
    n155,
    n83,
    n74,
    n97
  );


  nand
  g210
  (
    n159,
    n37,
    n44,
    n109
  );


  not
  g211
  (
    n300,
    n127
  );


  buf
  g212
  (
    n339,
    n113
  );


  buf
  g213
  (
    n315,
    n127
  );


  not
  g214
  (
    n245,
    n125
  );


  buf
  g215
  (
    n348,
    n115
  );


  buf
  g216
  (
    n316,
    n123
  );


  not
  g217
  (
    n354,
    n128
  );


  not
  g218
  (
    n318,
    n142
  );


  buf
  g219
  (
    n351,
    n123
  );


  buf
  g220
  (
    n273,
    n120
  );


  not
  g221
  (
    n319,
    n120
  );


  not
  g222
  (
    n272,
    n121
  );


  not
  g223
  (
    n337,
    n121
  );


  not
  g224
  (
    n249,
    n141
  );


  not
  g225
  (
    n342,
    n133
  );


  not
  g226
  (
    n280,
    n126
  );


  buf
  g227
  (
    n266,
    n133
  );


  buf
  g228
  (
    n358,
    n115
  );


  not
  g229
  (
    n327,
    n118
  );


  not
  g230
  (
    n289,
    n125
  );


  not
  g231
  (
    n331,
    n117
  );


  not
  g232
  (
    n244,
    n135
  );


  buf
  g233
  (
    n290,
    n135
  );


  buf
  g234
  (
    n279,
    n129
  );


  buf
  g235
  (
    n341,
    n130
  );


  not
  g236
  (
    n326,
    n114
  );


  not
  g237
  (
    n284,
    n138
  );


  not
  g238
  (
    n323,
    n127
  );


  buf
  g239
  (
    n340,
    n127
  );


  not
  g240
  (
    n302,
    n130
  );


  not
  g241
  (
    n260,
    n141
  );


  buf
  g242
  (
    n322,
    n115
  );


  buf
  g243
  (
    n275,
    n132
  );


  not
  g244
  (
    n285,
    n123
  );


  buf
  g245
  (
    n254,
    n126
  );


  not
  g246
  (
    n291,
    n139
  );


  buf
  g247
  (
    n248,
    n128
  );


  not
  g248
  (
    n335,
    n119
  );


  buf
  g249
  (
    n287,
    n134
  );


  not
  g250
  (
    n252,
    n132
  );


  buf
  g251
  (
    n309,
    n131
  );


  not
  g252
  (
    n265,
    n118
  );


  not
  g253
  (
    n256,
    n117
  );


  not
  g254
  (
    n262,
    n128
  );


  not
  g255
  (
    n310,
    n137
  );


  buf
  g256
  (
    n277,
    n130
  );


  not
  g257
  (
    n333,
    n119
  );


  buf
  g258
  (
    n283,
    n137
  );


  buf
  g259
  (
    n274,
    n129
  );


  buf
  g260
  (
    n336,
    n134
  );


  not
  g261
  (
    n301,
    n136
  );


  not
  g262
  (
    n347,
    n121
  );


  buf
  g263
  (
    n320,
    n119
  );


  not
  g264
  (
    n250,
    n131
  );


  not
  g265
  (
    n294,
    n119
  );


  not
  g266
  (
    n356,
    n136
  );


  not
  g267
  (
    n346,
    n122
  );


  buf
  g268
  (
    n355,
    n138
  );


  buf
  g269
  (
    n324,
    n133
  );


  buf
  g270
  (
    n271,
    n124
  );


  not
  g271
  (
    n267,
    n139
  );


  not
  g272
  (
    n314,
    n117
  );


  buf
  g273
  (
    n334,
    n139
  );


  buf
  g274
  (
    n286,
    n123
  );


  not
  g275
  (
    n247,
    n125
  );


  buf
  g276
  (
    n345,
    n114
  );


  not
  g277
  (
    n352,
    n135
  );


  not
  g278
  (
    n292,
    n124
  );


  not
  g279
  (
    n312,
    n120
  );


  not
  g280
  (
    n255,
    n114
  );


  buf
  g281
  (
    n305,
    n122
  );


  buf
  g282
  (
    n321,
    n117
  );


  not
  g283
  (
    n353,
    n140
  );


  not
  g284
  (
    n257,
    n128
  );


  buf
  g285
  (
    n343,
    n129
  );


  buf
  g286
  (
    n357,
    n118
  );


  not
  g287
  (
    n264,
    n140
  );


  not
  g288
  (
    n303,
    n131
  );


  not
  g289
  (
    n278,
    n137
  );


  buf
  g290
  (
    n253,
    n124
  );


  buf
  g291
  (
    n270,
    n130
  );


  not
  g292
  (
    n295,
    n116
  );


  not
  g293
  (
    n293,
    n132
  );


  buf
  g294
  (
    n299,
    n138
  );


  buf
  g295
  (
    n344,
    n138
  );


  buf
  g296
  (
    n311,
    n121
  );


  buf
  g297
  (
    n308,
    n126
  );


  not
  g298
  (
    n349,
    n120
  );


  not
  g299
  (
    n251,
    n134
  );


  not
  g300
  (
    n269,
    n113
  );


  buf
  g301
  (
    n329,
    n140
  );


  not
  g302
  (
    n261,
    n139
  );


  buf
  g303
  (
    n328,
    n142
  );


  buf
  g304
  (
    n313,
    n113
  );


  buf
  g305
  (
    n282,
    n125
  );


  not
  g306
  (
    n276,
    n124
  );


  not
  g307
  (
    n258,
    n141
  );


  buf
  g308
  (
    n246,
    n122
  );


  buf
  g309
  (
    n268,
    n131
  );


  buf
  g310
  (
    n317,
    n115
  );


  buf
  g311
  (
    n263,
    n140
  );


  buf
  g312
  (
    n281,
    n135
  );


  not
  g313
  (
    n259,
    n116
  );


  buf
  g314
  (
    n338,
    n137
  );


  not
  g315
  (
    n296,
    n136
  );


  buf
  g316
  (
    n298,
    n134
  );


  buf
  g317
  (
    n332,
    n126
  );


  buf
  g318
  (
    n304,
    n136
  );


  buf
  g319
  (
    n325,
    n113
  );


  buf
  g320
  (
    n350,
    n114
  );


  buf
  g321
  (
    n288,
    n141
  );


  buf
  g322
  (
    n297,
    n129
  );


  buf
  g323
  (
    n330,
    n118
  );


  buf
  g324
  (
    n306,
    n122
  );


  nand
  g325
  (
    n307,
    n116,
    n116,
    n133,
    n132
  );


  buf
  g326
  (
    n365,
    n320
  );


  buf
  g327
  (
    n441,
    n152
  );


  buf
  g328
  (
    n436,
    n156
  );


  not
  g329
  (
    n407,
    n150
  );


  not
  g330
  (
    n375,
    n142
  );


  not
  g331
  (
    n404,
    n255
  );


  buf
  g332
  (
    n382,
    n307
  );


  buf
  g333
  (
    n389,
    n152
  );


  buf
  g334
  (
    n438,
    n144
  );


  not
  g335
  (
    n414,
    n111
  );


  not
  g336
  (
    n384,
    n276
  );


  buf
  g337
  (
    n437,
    n315
  );


  buf
  g338
  (
    n403,
    n295
  );


  buf
  g339
  (
    n413,
    n149
  );


  buf
  g340
  (
    n385,
    n287
  );


  buf
  g341
  (
    n387,
    n259
  );


  buf
  g342
  (
    n439,
    n149
  );


  not
  g343
  (
    n425,
    n155
  );


  buf
  g344
  (
    n405,
    n291
  );


  buf
  g345
  (
    n372,
    n286
  );


  buf
  g346
  (
    n399,
    n268
  );


  not
  g347
  (
    n411,
    n278
  );


  not
  g348
  (
    n377,
    n152
  );


  not
  g349
  (
    n381,
    n153
  );


  not
  g350
  (
    n431,
    n145
  );


  buf
  g351
  (
    n435,
    n252
  );


  buf
  g352
  (
    n363,
    n303
  );


  buf
  g353
  (
    n434,
    n287
  );


  buf
  g354
  (
    n364,
    n112
  );


  not
  g355
  (
    n417,
    n151
  );


  not
  g356
  (
    n400,
    n270
  );


  not
  g357
  (
    n402,
    n313
  );


  not
  g358
  (
    n374,
    n312
  );


  not
  g359
  (
    n409,
    n301
  );


  buf
  g360
  (
    n392,
    n265
  );


  not
  g361
  (
    n420,
    n146
  );


  not
  g362
  (
    n408,
    n260
  );


  buf
  g363
  (
    n433,
    n245
  );


  not
  g364
  (
    n360,
    n294
  );


  buf
  g365
  (
    n366,
    n154
  );


  buf
  g366
  (
    n376,
    n253
  );


  buf
  g367
  (
    n398,
    n300
  );


  not
  g368
  (
    n421,
    n157
  );


  not
  g369
  (
    n371,
    n294
  );


  nor
  g370
  (
    n361,
    n289,
    n276,
    n302,
    n292
  );


  nor
  g371
  (
    n370,
    n248,
    n144,
    n151,
    n282
  );


  and
  g372
  (
    n419,
    n302,
    n151,
    n305,
    n268
  );


  and
  g373
  (
    n367,
    n152,
    n295,
    n111,
    n246
  );


  or
  g374
  (
    n390,
    n149,
    n275,
    n254,
    n306
  );


  xnor
  g375
  (
    n388,
    n278,
    n310,
    n155
  );


  xnor
  g376
  (
    n396,
    n272,
    n156,
    n308,
    n304
  );


  nand
  g377
  (
    n380,
    n281,
    n313,
    n298,
    n150
  );


  xor
  g378
  (
    n429,
    n153,
    n301,
    n154,
    n277
  );


  nor
  g379
  (
    n394,
    n311,
    n112,
    n269,
    n148
  );


  nand
  g380
  (
    n418,
    n290,
    n147,
    n143,
    n251
  );


  xnor
  g381
  (
    n415,
    n285,
    n284,
    n257,
    n308
  );


  nand
  g382
  (
    n359,
    n155,
    n27,
    n320,
    n280
  );


  xor
  g383
  (
    n424,
    n305,
    n304,
    n286,
    n150
  );


  xor
  g384
  (
    n410,
    n153,
    n307,
    n275,
    n266
  );


  nand
  g385
  (
    n426,
    n296,
    n154,
    n146,
    n148
  );


  nor
  g386
  (
    n373,
    n145,
    n279,
    n281,
    n288
  );


  nor
  g387
  (
    n427,
    n146,
    n144,
    n317,
    n258
  );


  and
  g388
  (
    n369,
    n277,
    n309,
    n315,
    n297
  );


  nor
  g389
  (
    n379,
    n292,
    n155,
    n148,
    n143
  );


  nor
  g390
  (
    n395,
    n145,
    n306,
    n314,
    n267
  );


  nor
  g391
  (
    n391,
    n273,
    n290,
    n112,
    n144
  );


  xor
  g392
  (
    n386,
    n291,
    n256,
    n269,
    n264
  );


  xnor
  g393
  (
    n378,
    n319,
    n293,
    n303,
    n148
  );


  xor
  g394
  (
    n401,
    n271,
    n274,
    n316,
    n288
  );


  and
  g395
  (
    n406,
    n143,
    n311,
    n314,
    n284
  );


  and
  g396
  (
    n393,
    n282,
    n147,
    n289,
    n299
  );


  xnor
  g397
  (
    n397,
    n147,
    n111,
    n280,
    n142
  );


  or
  g398
  (
    n432,
    n312,
    n293,
    n154,
    n271
  );


  and
  g399
  (
    n412,
    n262,
    n272,
    n298,
    n299
  );


  xor
  g400
  (
    n362,
    n244,
    n151,
    n112,
    n285
  );


  or
  g401
  (
    n416,
    n318,
    n267,
    n27,
    n283
  );


  and
  g402
  (
    n422,
    n274,
    n143,
    n283,
    n146
  );


  nor
  g403
  (
    n428,
    n156,
    n249,
    n296,
    n316
  );


  and
  g404
  (
    n368,
    n270,
    n317,
    n263,
    n319
  );


  or
  g405
  (
    n430,
    n145,
    n318,
    n273,
    n149
  );


  and
  g406
  (
    n440,
    n153,
    n266,
    n147,
    n156
  );


  and
  g407
  (
    n383,
    n279,
    n309,
    n247,
    n250
  );


  xnor
  g408
  (
    n423,
    n300,
    n150,
    n297,
    n261
  );


  xnor
  g409
  (
    n445,
    n362,
    n364,
    n363
  );


  xnor
  g410
  (
    n448,
    n364,
    n360
  );


  and
  g411
  (
    n447,
    n361,
    n360,
    n363
  );


  or
  g412
  (
    n444,
    n360,
    n361,
    n366,
    n362
  );


  xnor
  g413
  (
    n442,
    n362,
    n361,
    n366,
    n364
  );


  xnor
  g414
  (
    n443,
    n362,
    n366,
    n365
  );


  nor
  g415
  (
    n446,
    n364,
    n365
  );


  xnor
  g416
  (
    n449,
    n359,
    n363,
    n361,
    n367
  );


  nor
  g417
  (
    n452,
    n157,
    n28,
    n158
  );


  xnor
  g418
  (
    n451,
    n443,
    n445,
    n157,
    n29
  );


  nand
  g419
  (
    n450,
    n28,
    n158,
    n157
  );


  xor
  g420
  (
    n453,
    n158,
    n28,
    n444,
    n442
  );


  nor
  g421
  (
    n463,
    n450,
    n369,
    n453,
    n373
  );


  or
  g422
  (
    n461,
    n371,
    n372,
    n367
  );


  nor
  g423
  (
    n456,
    n370,
    n373,
    n368
  );


  nand
  g424
  (
    n460,
    n374,
    n371,
    n452,
    n369
  );


  nand
  g425
  (
    n458,
    n370,
    n369,
    n452
  );


  nor
  g426
  (
    n454,
    n453,
    n453,
    n374,
    n371
  );


  or
  g427
  (
    n455,
    n368,
    n372,
    n451,
    n369
  );


  xnor
  g428
  (
    n457,
    n368,
    n453,
    n372,
    n367
  );


  or
  g429
  (
    n462,
    n370,
    n372,
    n373,
    n374
  );


  nand
  g430
  (
    n459,
    n452,
    n370,
    n373,
    n371
  );


  or
  g431
  (
    n497,
    n160,
    n463,
    n383,
    n461
  );


  xnor
  g432
  (
    n498,
    n167,
    n159,
    n171,
    n166
  );


  xor
  g433
  (
    n489,
    n160,
    n164,
    n460,
    n457
  );


  xor
  g434
  (
    n483,
    n381,
    n170,
    n456,
    n175
  );


  xnor
  g435
  (
    n468,
    n384,
    n177,
    n168,
    n383
  );


  and
  g436
  (
    n492,
    n459,
    n163,
    n171,
    n461
  );


  xnor
  g437
  (
    n501,
    n159,
    n457,
    n379,
    n177
  );


  nand
  g438
  (
    n465,
    n164,
    n383,
    n173,
    n163
  );


  nand
  g439
  (
    n485,
    n164,
    n456,
    n378,
    n376
  );


  xnor
  g440
  (
    n477,
    n178,
    n457,
    n162
  );


  nand
  g441
  (
    n491,
    n379,
    n173,
    n459,
    n381
  );


  nand
  g442
  (
    n499,
    n455,
    n174,
    n159,
    n171
  );


  or
  g443
  (
    n480,
    n461,
    n455,
    n462,
    n169
  );


  and
  g444
  (
    n500,
    n455,
    n177,
    n174
  );


  nand
  g445
  (
    n478,
    n161,
    n461,
    n380,
    n383
  );


  nor
  g446
  (
    n479,
    n378,
    n379,
    n377,
    n165
  );


  xor
  g447
  (
    n503,
    n460,
    n160,
    n169,
    n378
  );


  xor
  g448
  (
    n482,
    n172,
    n169,
    n375,
    n161
  );


  xor
  g449
  (
    n487,
    n172,
    n169,
    n380,
    n170
  );


  nand
  g450
  (
    n502,
    n454,
    n382,
    n168,
    n375
  );


  and
  g451
  (
    n488,
    n175,
    n454,
    n163,
    n166
  );


  nor
  g452
  (
    n495,
    n160,
    n377,
    n176,
    n167
  );


  nor
  g453
  (
    n496,
    n176,
    n458,
    n384,
    n382
  );


  and
  g454
  (
    n466,
    n455,
    n172,
    n457,
    n463
  );


  nor
  g455
  (
    n486,
    n379,
    n175,
    n459,
    n162
  );


  or
  g456
  (
    n494,
    n463,
    n376,
    n176,
    n166
  );


  nor
  g457
  (
    n472,
    n460,
    n165,
    n458,
    n175
  );


  nand
  g458
  (
    n470,
    n458,
    n170,
    n163,
    n167
  );


  nor
  g459
  (
    n471,
    n172,
    n381,
    n173,
    n376
  );


  xnor
  g460
  (
    n481,
    n456,
    n384,
    n377,
    n176
  );


  and
  g461
  (
    n490,
    n382,
    n380,
    n454,
    n462
  );


  xor
  g462
  (
    n469,
    n374,
    n178,
    n168,
    n161
  );


  xnor
  g463
  (
    n484,
    n463,
    n159,
    n460,
    n173
  );


  or
  g464
  (
    n467,
    n165,
    n462,
    n381,
    n161
  );


  xnor
  g465
  (
    n475,
    n384,
    n166,
    n459,
    n375
  );


  or
  g466
  (
    n473,
    n454,
    n382,
    n168,
    n380
  );


  xnor
  g467
  (
    n476,
    n376,
    n378,
    n462,
    n174
  );


  xnor
  g468
  (
    n474,
    n377,
    n170,
    n456,
    n177
  );


  nand
  g469
  (
    n464,
    n162,
    n375,
    n171,
    n164
  );


  or
  g470
  (
    n493,
    n167,
    n458,
    n165,
    n178
  );


  and
  g471
  (
    n554,
    n343,
    n345,
    n391,
    n470
  );


  xnor
  g472
  (
    n551,
    n399,
    n397,
    n343,
    n478
  );


  nand
  g473
  (
    n530,
    n332,
    n350,
    n487,
    n347
  );


  nor
  g474
  (
    n574,
    n467,
    n396,
    n464,
    n332
  );


  xor
  g475
  (
    n508,
    n346,
    n358,
    n405,
    n487
  );


  xnor
  g476
  (
    n525,
    n349,
    n350,
    n386,
    n329
  );


  nand
  g477
  (
    n571,
    n483,
    n390,
    n485,
    n400
  );


  xnor
  g478
  (
    n548,
    n339,
    n327,
    n335,
    n386
  );


  nor
  g479
  (
    n519,
    n397,
    n486,
    n475,
    n471
  );


  xnor
  g480
  (
    n512,
    n474,
    n393,
    n466,
    n355
  );


  xnor
  g481
  (
    n547,
    n487,
    n331,
    n330
  );


  nor
  g482
  (
    n568,
    n354,
    n336,
    n346,
    n491
  );


  xnor
  g483
  (
    n572,
    n343,
    n345,
    n327,
    n349
  );


  or
  g484
  (
    n529,
    n480,
    n355,
    n392,
    n485
  );


  xor
  g485
  (
    n523,
    n355,
    n336,
    n348,
    n393
  );


  or
  g486
  (
    n544,
    n321,
    n326,
    n332,
    n395
  );


  xor
  g487
  (
    n567,
    n489,
    n404,
    n399,
    n391
  );


  xor
  g488
  (
    n520,
    n385,
    n398,
    n395,
    n490
  );


  xnor
  g489
  (
    n504,
    n325,
    n388,
    n394,
    n341
  );


  nand
  g490
  (
    n536,
    n484,
    n488,
    n340,
    n321
  );


  xor
  g491
  (
    n560,
    n484,
    n337,
    n396,
    n467
  );


  or
  g492
  (
    n531,
    n400,
    n334,
    n335,
    n491
  );


  xor
  g493
  (
    n527,
    n404,
    n348,
    n351,
    n388
  );


  xor
  g494
  (
    n553,
    n482,
    n339,
    n328,
    n485
  );


  xnor
  g495
  (
    n555,
    n474,
    n336,
    n397,
    n485
  );


  xnor
  g496
  (
    n521,
    n401,
    n396,
    n358,
    n354
  );


  xnor
  g497
  (
    n549,
    n352,
    n387,
    n326,
    n338
  );


  nand
  g498
  (
    n558,
    n490,
    n489,
    n400,
    n335
  );


  xor
  g499
  (
    n522,
    n357,
    n352,
    n472,
    n405
  );


  or
  g500
  (
    n576,
    n464,
    n338,
    n337,
    n331
  );


  and
  g501
  (
    n524,
    n338,
    n332,
    n385,
    n478
  );


  nor
  g502
  (
    n575,
    n394,
    n352,
    n339,
    n403
  );


  or
  g503
  (
    n557,
    n334,
    n385,
    n386,
    n477
  );


  or
  g504
  (
    n569,
    n395,
    n353,
    n484,
    n487
  );


  nand
  g505
  (
    n528,
    n401,
    n390,
    n354,
    n490
  );


  or
  g506
  (
    n518,
    n393,
    n483,
    n336,
    n356
  );


  or
  g507
  (
    n507,
    n347,
    n340,
    n398,
    n472
  );


  nand
  g508
  (
    n566,
    n347,
    n339,
    n351,
    n398
  );


  nor
  g509
  (
    n517,
    n356,
    n350,
    n387,
    n395
  );


  xnor
  g510
  (
    n573,
    n388,
    n324,
    n325,
    n391
  );


  xor
  g511
  (
    n526,
    n335,
    n387,
    n340,
    n483
  );


  nand
  g512
  (
    n511,
    n466,
    n329,
    n405,
    n354
  );


  nand
  g513
  (
    n564,
    n473,
    n386,
    n398,
    n404
  );


  xor
  g514
  (
    n546,
    n469,
    n331,
    n403,
    n481
  );


  xor
  g515
  (
    n514,
    n337,
    n396,
    n394,
    n352
  );


  nor
  g516
  (
    n539,
    n341,
    n390,
    n323,
    n322
  );


  xor
  g517
  (
    n545,
    n402,
    n480,
    n330,
    n353
  );


  xor
  g518
  (
    n550,
    n490,
    n402,
    n477,
    n355
  );


  or
  g519
  (
    n542,
    n349,
    n330,
    n333,
    n358
  );


  and
  g520
  (
    n537,
    n406,
    n337,
    n402,
    n342
  );


  xor
  g521
  (
    n505,
    n473,
    n479,
    n322,
    n393
  );


  nor
  g522
  (
    n562,
    n471,
    n402,
    n397,
    n481
  );


  and
  g523
  (
    n535,
    n476,
    n333,
    n389,
    n486
  );


  nor
  g524
  (
    n552,
    n331,
    n345,
    n399,
    n357
  );


  nand
  g525
  (
    n540,
    n479,
    n358,
    n392,
    n356
  );


  xor
  g526
  (
    n509,
    n491,
    n344,
    n399,
    n400
  );


  xor
  g527
  (
    n515,
    n324,
    n343,
    n338,
    n357
  );


  and
  g528
  (
    n563,
    n465,
    n385,
    n486,
    n341
  );


  nor
  g529
  (
    n559,
    n488,
    n475,
    n389,
    n333
  );


  or
  g530
  (
    n543,
    n347,
    n353,
    n392,
    n334
  );


  nand
  g531
  (
    n534,
    n488,
    n345,
    n391,
    n390
  );


  and
  g532
  (
    n570,
    n488,
    n340,
    n482,
    n468
  );


  xor
  g533
  (
    n533,
    n489,
    n470,
    n476,
    n348
  );


  nand
  g534
  (
    n565,
    n394,
    n344,
    n349,
    n401
  );


  xnor
  g535
  (
    n516,
    n333,
    n484,
    n323,
    n357
  );


  nand
  g536
  (
    n532,
    n465,
    n403,
    n344,
    n405
  );


  xor
  g537
  (
    n506,
    n334,
    n483,
    n401,
    n351
  );


  or
  g538
  (
    n541,
    n342,
    n328,
    n387,
    n348
  );


  nand
  g539
  (
    n538,
    n342,
    n342,
    n350,
    n344
  );


  nor
  g540
  (
    n561,
    n351,
    n468,
    n469,
    n403
  );


  nor
  g541
  (
    n513,
    n486,
    n341,
    n392,
    n346
  );


  or
  g542
  (
    n556,
    n404,
    n353,
    n389
  );


  xnor
  g543
  (
    n510,
    n388,
    n346,
    n489,
    n356
  );


  xor
  g544
  (
    n584,
    n407,
    n510
  );


  nor
  g545
  (
    n580,
    n406,
    n508
  );


  nand
  g546
  (
    n579,
    n504,
    n506
  );


  xor
  g547
  (
    n582,
    n507,
    n505
  );


  and
  g548
  (
    n578,
    n511,
    n408
  );


  or
  g549
  (
    n583,
    n509,
    n406
  );


  not
  g550
  (
    n581,
    n407
  );


  xnor
  g551
  (
    n577,
    n407,
    n406
  );


  xnor
  g552
  (
    n608,
    n411,
    n522,
    n448,
    n180
  );


  xnor
  g553
  (
    n603,
    n183,
    n583,
    n521,
    n578
  );


  xnor
  g554
  (
    n606,
    n409,
    n409,
    n551,
    n579
  );


  and
  g555
  (
    n595,
    n525,
    n584,
    n526,
    n181
  );


  or
  g556
  (
    n602,
    n183,
    n577,
    n181,
    n411
  );


  and
  g557
  (
    n613,
    n578,
    n512,
    n534,
    n543
  );


  nor
  g558
  (
    n607,
    n582,
    n180,
    n181,
    n579
  );


  or
  g559
  (
    n612,
    n181,
    n179,
    n581
  );


  nand
  g560
  (
    n611,
    n449,
    n179,
    n580,
    n531
  );


  nand
  g561
  (
    n610,
    n532,
    n178,
    n411,
    n582
  );


  xnor
  g562
  (
    n609,
    n514,
    n446,
    n538,
    n410
  );


  xnor
  g563
  (
    n596,
    n180,
    n516,
    n581,
    n527
  );


  nor
  g564
  (
    n592,
    n580,
    n523,
    n518,
    n515
  );


  or
  g565
  (
    n588,
    n179,
    n408,
    n579,
    n183
  );


  nor
  g566
  (
    n591,
    n546,
    n182,
    n410,
    n582
  );


  xnor
  g567
  (
    n587,
    n579,
    n547,
    n541,
    n580
  );


  nand
  g568
  (
    n604,
    n409,
    n550,
    n583,
    n517
  );


  or
  g569
  (
    n593,
    n540,
    n533,
    n548,
    n182
  );


  nand
  g570
  (
    n599,
    n539,
    n583,
    n182,
    n584
  );


  xnor
  g571
  (
    n601,
    n410,
    n448,
    n449
  );


  nand
  g572
  (
    n594,
    n513,
    n583,
    n447,
    n520
  );


  nand
  g573
  (
    n600,
    n578,
    n524,
    n580,
    n544
  );


  and
  g574
  (
    n589,
    n449,
    n581,
    n549
  );


  or
  g575
  (
    n605,
    n447,
    n182,
    n578,
    n446
  );


  nand
  g576
  (
    n598,
    n582,
    n584,
    n408,
    n535
  );


  and
  g577
  (
    n586,
    n584,
    n448,
    n491,
    n537
  );


  xnor
  g578
  (
    n597,
    n545,
    n409,
    n529,
    n542
  );


  or
  g579
  (
    n585,
    n449,
    n536,
    n519,
    n180
  );


  or
  g580
  (
    n590,
    n408,
    n528,
    n530,
    n410
  );


  not
  g581
  (
    n658,
    n429
  );


  buf
  g582
  (
    n665,
    n608
  );


  not
  g583
  (
    n638,
    n610
  );


  not
  g584
  (
    n620,
    n593
  );


  not
  g585
  (
    n625,
    n596
  );


  buf
  g586
  (
    n656,
    n592
  );


  buf
  g587
  (
    n621,
    n594
  );


  buf
  g588
  (
    n701,
    n590
  );


  buf
  g589
  (
    n615,
    n594
  );


  buf
  g590
  (
    n671,
    n599
  );


  buf
  g591
  (
    n618,
    n591
  );


  buf
  g592
  (
    n691,
    n418
  );


  not
  g593
  (
    n666,
    n593
  );


  not
  g594
  (
    n630,
    n603
  );


  buf
  g595
  (
    n708,
    n613
  );


  buf
  g596
  (
    n676,
    n417
  );


  buf
  g597
  (
    n644,
    n589
  );


  buf
  g598
  (
    n640,
    n595
  );


  not
  g599
  (
    n672,
    n603
  );


  buf
  g600
  (
    n633,
    n418
  );


  not
  g601
  (
    n704,
    n606
  );


  buf
  g602
  (
    n702,
    n608
  );


  not
  g603
  (
    n614,
    n606
  );


  not
  g604
  (
    n646,
    n590
  );


  buf
  g605
  (
    n634,
    n604
  );


  buf
  g606
  (
    n693,
    n600
  );


  not
  g607
  (
    n684,
    n421
  );


  not
  g608
  (
    n668,
    n598
  );


  buf
  g609
  (
    n639,
    n564
  );


  buf
  g610
  (
    n631,
    n432
  );


  buf
  g611
  (
    n685,
    n436
  );


  not
  g612
  (
    n653,
    n596
  );


  not
  g613
  (
    n632,
    n613
  );


  buf
  g614
  (
    n663,
    n593
  );


  not
  g615
  (
    n675,
    n422
  );


  buf
  g616
  (
    n679,
    n596
  );


  not
  g617
  (
    n689,
    n607
  );


  not
  g618
  (
    n623,
    n595
  );


  not
  g619
  (
    n682,
    n604
  );


  buf
  g620
  (
    n619,
    n594
  );


  not
  g621
  (
    n698,
    n586
  );


  not
  g622
  (
    n700,
    n554
  );


  buf
  g623
  (
    n617,
    n592
  );


  buf
  g624
  (
    n686,
    n415
  );


  not
  g625
  (
    n648,
    n589
  );


  buf
  g626
  (
    n664,
    n417
  );


  buf
  g627
  (
    n667,
    n597
  );


  not
  g628
  (
    n699,
    n607
  );


  not
  g629
  (
    n641,
    n612
  );


  xnor
  g630
  (
    n705,
    n421,
    n493,
    n604
  );


  nand
  g631
  (
    n624,
    n420,
    n413,
    n434,
    n585
  );


  nand
  g632
  (
    n627,
    n420,
    n563,
    n492,
    n428
  );


  nor
  g633
  (
    n637,
    n607,
    n426,
    n430,
    n417
  );


  nor
  g634
  (
    n695,
    n587,
    n425,
    n424,
    n599
  );


  xor
  g635
  (
    n661,
    n592,
    n426,
    n585,
    n588
  );


  and
  g636
  (
    n696,
    n588,
    n428,
    n604,
    n559
  );


  xor
  g637
  (
    n669,
    n412,
    n589,
    n429,
    n601
  );


  xor
  g638
  (
    n642,
    n414,
    n435,
    n597,
    n436
  );


  nand
  g639
  (
    n655,
    n608,
    n595,
    n601,
    n416
  );


  and
  g640
  (
    n673,
    n422,
    n594,
    n418,
    n600
  );


  xnor
  g641
  (
    n659,
    n424,
    n419,
    n602,
    n586
  );


  and
  g642
  (
    n654,
    n601,
    n419,
    n608,
    n416
  );


  nand
  g643
  (
    n680,
    n609,
    n605,
    n420
  );


  xnor
  g644
  (
    n662,
    n427,
    n603,
    n426,
    n434
  );


  xor
  g645
  (
    n690,
    n431,
    n599,
    n412,
    n585
  );


  or
  g646
  (
    n687,
    n586,
    n427,
    n428,
    n588
  );


  nor
  g647
  (
    n692,
    n597,
    n427,
    n416,
    n561
  );


  nor
  g648
  (
    n651,
    n610,
    n613,
    n612,
    n598
  );


  and
  g649
  (
    n706,
    n553,
    n432,
    n611,
    n590
  );


  nand
  g650
  (
    n626,
    n431,
    n415,
    n423
  );


  xor
  g651
  (
    n678,
    n434,
    n492,
    n600,
    n423
  );


  and
  g652
  (
    n703,
    n432,
    n421,
    n605,
    n593
  );


  xor
  g653
  (
    n652,
    n430,
    n599,
    n421,
    n436
  );


  nor
  g654
  (
    n694,
    n585,
    n592,
    n417,
    n425
  );


  and
  g655
  (
    n709,
    n595,
    n414,
    n412,
    n424
  );


  or
  g656
  (
    n677,
    n436,
    n590,
    n610,
    n557
  );


  or
  g657
  (
    n636,
    n610,
    n435,
    n430,
    n429
  );


  and
  g658
  (
    n616,
    n611,
    n596,
    n492,
    n430
  );


  nor
  g659
  (
    n649,
    n415,
    n419,
    n432
  );


  nor
  g660
  (
    n657,
    n612,
    n435,
    n414,
    n420
  );


  or
  g661
  (
    n628,
    n556,
    n598,
    n413,
    n424
  );


  or
  g662
  (
    n629,
    n586,
    n434,
    n611,
    n603
  );


  xnor
  g663
  (
    n660,
    n492,
    n598,
    n602,
    n425
  );


  nor
  g664
  (
    n683,
    n429,
    n413,
    n613,
    n411
  );


  and
  g665
  (
    n647,
    n428,
    n607,
    n609,
    n422
  );


  nand
  g666
  (
    n697,
    n431,
    n558,
    n433,
    n435
  );


  or
  g667
  (
    n707,
    n560,
    n588,
    n605,
    n426
  );


  nor
  g668
  (
    n674,
    n433,
    n587,
    n611,
    n600
  );


  and
  g669
  (
    n645,
    n437,
    n602,
    n606,
    n601
  );


  and
  g670
  (
    n670,
    n425,
    n589,
    n418,
    n609
  );


  nor
  g671
  (
    n688,
    n552,
    n609,
    n591,
    n423
  );


  nand
  g672
  (
    n643,
    n597,
    n612,
    n427,
    n433
  );


  nor
  g673
  (
    n681,
    n422,
    n555,
    n416,
    n602
  );


  xnor
  g674
  (
    n650,
    n414,
    n591,
    n413,
    n412
  );


  and
  g675
  (
    n635,
    n606,
    n591,
    n587,
    n415
  );


  xnor
  g676
  (
    n622,
    n562,
    n587,
    n431,
    n433
  );


  xor
  g677
  (
    n769,
    n184,
    n225,
    n706,
    n238
  );


  nand
  g678
  (
    n778,
    n198,
    n570,
    n188,
    n201
  );


  nand
  g679
  (
    n741,
    n617,
    n625,
    n643,
    n187
  );


  nand
  g680
  (
    n714,
    n189,
    n665,
    n623,
    n199
  );


  xnor
  g681
  (
    n755,
    n664,
    n672,
    n197,
    n627
  );


  nor
  g682
  (
    n798,
    n681,
    n651,
    n668,
    n623
  );


  or
  g683
  (
    n760,
    n686,
    n202,
    n661,
    n230
  );


  or
  g684
  (
    n870,
    n238,
    n232,
    n672,
    n660
  );


  and
  g685
  (
    n869,
    n241,
    n202,
    n679,
    n628
  );


  or
  g686
  (
    n810,
    n688,
    n183,
    n208,
    n684
  );


  and
  g687
  (
    n752,
    n690,
    n669,
    n682,
    n200
  );


  nor
  g688
  (
    n751,
    n662,
    n663,
    n231,
    n614
  );


  and
  g689
  (
    n802,
    n239,
    n186,
    n222,
    n194
  );


  xor
  g690
  (
    n759,
    n217,
    n666,
    n243,
    n657
  );


  and
  g691
  (
    n816,
    n619,
    n661,
    n683,
    n185
  );


  nor
  g692
  (
    n844,
    n650,
    n683,
    n208,
    n673
  );


  xnor
  g693
  (
    n849,
    n677,
    n630,
    n642,
    n676
  );


  or
  g694
  (
    n744,
    n224,
    n698,
    n628,
    n208
  );


  xnor
  g695
  (
    n713,
    n695,
    n635,
    n234,
    n216
  );


  xor
  g696
  (
    n806,
    n196,
    n29,
    n630,
    n658
  );


  nor
  g697
  (
    n753,
    n692,
    n617,
    n651,
    n622
  );


  or
  g698
  (
    n850,
    n619,
    n203,
    n236,
    n211
  );


  nand
  g699
  (
    n848,
    n692,
    n237,
    n645,
    n243
  );


  nand
  g700
  (
    n818,
    n615,
    n235,
    n32,
    n625
  );


  or
  g701
  (
    n854,
    n224,
    n646,
    n621,
    n620
  );


  xnor
  g702
  (
    n780,
    n653,
    n665,
    n631,
    n614
  );


  xor
  g703
  (
    n735,
    n186,
    n209,
    n31,
    n236
  );


  xnor
  g704
  (
    n772,
    n701,
    n188,
    n689,
    n695
  );


  xnor
  g705
  (
    n811,
    n32,
    n232,
    n229,
    n646
  );


  nand
  g706
  (
    n716,
    n238,
    n654,
    n636,
    n632
  );


  or
  g707
  (
    n732,
    n619,
    n666,
    n199,
    n639
  );


  xor
  g708
  (
    n862,
    n659,
    n239,
    n706,
    n648
  );


  nand
  g709
  (
    n825,
    n659,
    n624,
    n184,
    n206
  );


  xnor
  g710
  (
    n787,
    n615,
    n652,
    n677,
    n223
  );


  xnor
  g711
  (
    n842,
    n694,
    n631,
    n30,
    n681
  );


  nor
  g712
  (
    n796,
    n685,
    n187,
    n200,
    n680
  );


  nand
  g713
  (
    n710,
    n690,
    n650,
    n32,
    n693
  );


  or
  g714
  (
    n853,
    n678,
    n702,
    n687,
    n654
  );


  nand
  g715
  (
    n805,
    n229,
    n228,
    n668,
    n618
  );


  xor
  g716
  (
    n717,
    n184,
    n697,
    n632,
    n676
  );


  nand
  g717
  (
    n828,
    n214,
    n687,
    n194,
    n235
  );


  and
  g718
  (
    n726,
    n653,
    n692,
    n626,
    n651
  );


  or
  g719
  (
    n777,
    n213,
    n657,
    n696,
    n214
  );


  and
  g720
  (
    n747,
    n226,
    n681,
    n682,
    n204
  );


  nand
  g721
  (
    n843,
    n635,
    n650,
    n693,
    n653
  );


  and
  g722
  (
    n739,
    n189,
    n660,
    n215
  );


  xnor
  g723
  (
    n773,
    n218,
    n198,
    n695,
    n615
  );


  and
  g724
  (
    n761,
    n703,
    n630,
    n203,
    n657
  );


  xnor
  g725
  (
    n856,
    n674,
    n677,
    n649,
    n234
  );


  and
  g726
  (
    n768,
    n220,
    n678,
    n701,
    n615
  );


  and
  g727
  (
    n738,
    n700,
    n185,
    n216,
    n637
  );


  nor
  g728
  (
    n799,
    n237,
    n664,
    n201,
    n658
  );


  nor
  g729
  (
    n861,
    n29,
    n231,
    n640,
    n652
  );


  or
  g730
  (
    n840,
    n207,
    n184,
    n705,
    n627
  );


  nor
  g731
  (
    n823,
    n239,
    n637,
    n221,
    n231
  );


  or
  g732
  (
    n779,
    n617,
    n229,
    n678,
    n675
  );


  xnor
  g733
  (
    n871,
    n31,
    n618,
    n709,
    n191
  );


  xnor
  g734
  (
    n785,
    n699,
    n192,
    n220,
    n189
  );


  or
  g735
  (
    n792,
    n201,
    n207,
    n645,
    n668
  );


  xor
  g736
  (
    n794,
    n656,
    n679,
    n708,
    n698
  );


  nor
  g737
  (
    n724,
    n669,
    n199,
    n639,
    n242
  );


  or
  g738
  (
    n764,
    n225,
    n210,
    n204,
    n205
  );


  xnor
  g739
  (
    n733,
    n567,
    n193,
    n212,
    n655
  );


  and
  g740
  (
    n743,
    n684,
    n190,
    n680,
    n212
  );


  nor
  g741
  (
    n809,
    n650,
    n654,
    n236,
    n234
  );


  nand
  g742
  (
    n784,
    n242,
    n230,
    n31,
    n685
  );


  or
  g743
  (
    n866,
    n235,
    n640,
    n656,
    n694
  );


  xor
  g744
  (
    n837,
    n571,
    n689,
    n697,
    n645
  );


  nor
  g745
  (
    n841,
    n206,
    n672,
    n212,
    n691
  );


  or
  g746
  (
    n770,
    n675,
    n621,
    n620,
    n667
  );


  or
  g747
  (
    n774,
    n572,
    n209,
    n236,
    n219
  );


  xor
  g748
  (
    n807,
    n223,
    n233,
    n195,
    n621
  );


  nand
  g749
  (
    n725,
    n680,
    n696,
    n668,
    n624
  );


  nand
  g750
  (
    n762,
    n679,
    n639,
    n673,
    n235
  );


  xnor
  g751
  (
    n728,
    n691,
    n622,
    n687,
    n631
  );


  or
  g752
  (
    n852,
    n654,
    n699,
    n671,
    n709
  );


  nor
  g753
  (
    n833,
    n243,
    n689,
    n634,
    n209
  );


  nand
  g754
  (
    n808,
    n658,
    n662,
    n664,
    n240
  );


  xor
  g755
  (
    n771,
    n200,
    n633,
    n241,
    n217
  );


  xor
  g756
  (
    n832,
    n237,
    n706,
    n691,
    n651
  );


  nor
  g757
  (
    n788,
    n194,
    n225,
    n709,
    n704
  );


  or
  g758
  (
    n789,
    n704,
    n222,
    n210,
    n241
  );


  nor
  g759
  (
    n863,
    n228,
    n189,
    n227,
    n637
  );


  xor
  g760
  (
    n839,
    n217,
    n30,
    n240,
    n196
  );


  xor
  g761
  (
    n814,
    n242,
    n221,
    n645,
    n614
  );


  and
  g762
  (
    n845,
    n197,
    n697,
    n662,
    n660
  );


  or
  g763
  (
    n864,
    n617,
    n618,
    n671,
    n679
  );


  and
  g764
  (
    n781,
    n192,
    n633,
    n675,
    n569
  );


  xor
  g765
  (
    n765,
    n202,
    n205,
    n627,
    n223
  );


  and
  g766
  (
    n775,
    n216,
    n622,
    n638,
    n620
  );


  nand
  g767
  (
    n859,
    n694,
    n211,
    n648,
    n616
  );


  nand
  g768
  (
    n829,
    n206,
    n683,
    n700,
    n669
  );


  nand
  g769
  (
    n855,
    n641,
    n191,
    n672
  );


  and
  g770
  (
    n860,
    n663,
    n685,
    n652,
    n618
  );


  nor
  g771
  (
    n748,
    n698,
    n195,
    n691,
    n207
  );


  and
  g772
  (
    n718,
    n629,
    n655,
    n215,
    n692
  );


  or
  g773
  (
    n783,
    n662,
    n671,
    n218,
    n211
  );


  xnor
  g774
  (
    n750,
    n210,
    n212,
    n648,
    n702
  );


  nand
  g775
  (
    n820,
    n628,
    n242,
    n185,
    n674
  );


  xnor
  g776
  (
    n793,
    n690,
    n186,
    n667,
    n657
  );


  nand
  g777
  (
    n812,
    n576,
    n203,
    n688,
    n638
  );


  xor
  g778
  (
    n831,
    n193,
    n211,
    n705,
    n641
  );


  nand
  g779
  (
    n786,
    n209,
    n226,
    n217,
    n31
  );


  xnor
  g780
  (
    n819,
    n222,
    n203,
    n221,
    n202
  );


  and
  g781
  (
    n737,
    n233,
    n670,
    n683,
    n197
  );


  nor
  g782
  (
    n740,
    n630,
    n204,
    n636,
    n656
  );


  nor
  g783
  (
    n867,
    n634,
    n663,
    n701,
    n647
  );


  or
  g784
  (
    n817,
    n685,
    n702,
    n616,
    n629
  );


  nand
  g785
  (
    n711,
    n195,
    n625,
    n640,
    n226
  );


  and
  g786
  (
    n746,
    n695,
    n661,
    n636,
    n233
  );


  xor
  g787
  (
    n797,
    n207,
    n208,
    n190
  );


  nor
  g788
  (
    n834,
    n677,
    n638,
    n637,
    n204
  );


  xnor
  g789
  (
    n804,
    n642,
    n218,
    n641,
    n188
  );


  or
  g790
  (
    n846,
    n214,
    n199,
    n633,
    n213
  );


  nor
  g791
  (
    n721,
    n619,
    n644,
    n675,
    n655
  );


  nor
  g792
  (
    n835,
    n648,
    n231,
    n193,
    n232
  );


  nand
  g793
  (
    n865,
    n703,
    n693,
    n700,
    n225
  );


  xor
  g794
  (
    n715,
    n661,
    n214,
    n680,
    n684
  );


  nand
  g795
  (
    n857,
    n708,
    n671,
    n240,
    n647
  );


  nand
  g796
  (
    n749,
    n638,
    n227,
    n215,
    n224
  );


  or
  g797
  (
    n754,
    n626,
    n566,
    n565,
    n240
  );


  xor
  g798
  (
    n868,
    n674,
    n646,
    n206,
    n219
  );


  and
  g799
  (
    n830,
    n660,
    n643,
    n190,
    n658
  );


  nor
  g800
  (
    n791,
    n201,
    n699,
    n674,
    n633
  );


  xor
  g801
  (
    n722,
    n186,
    n187,
    n655
  );


  nor
  g802
  (
    n790,
    n29,
    n640,
    n621,
    n670
  );


  or
  g803
  (
    n763,
    n676,
    n690,
    n688,
    n639
  );


  nor
  g804
  (
    n742,
    n652,
    n686,
    n193,
    n626
  );


  xor
  g805
  (
    n782,
    n620,
    n205,
    n644,
    n32
  );


  and
  g806
  (
    n824,
    n684,
    n643,
    n234,
    n649
  );


  xor
  g807
  (
    n858,
    n665,
    n229,
    n624,
    n641
  );


  xnor
  g808
  (
    n821,
    n699,
    n625,
    n669,
    n632
  );


  and
  g809
  (
    n734,
    n227,
    n205,
    n707,
    n197
  );


  xnor
  g810
  (
    n723,
    n697,
    n708,
    n649,
    n30
  );


  or
  g811
  (
    n801,
    n702,
    n696,
    n230,
    n653
  );


  nor
  g812
  (
    n827,
    n705,
    n200,
    n701,
    n673
  );


  and
  g813
  (
    n730,
    n647,
    n659,
    n670,
    n693
  );


  xnor
  g814
  (
    n712,
    n227,
    n196,
    n213,
    n707
  );


  or
  g815
  (
    n795,
    n614,
    n195,
    n629,
    n704
  );


  xor
  g816
  (
    n776,
    n664,
    n241,
    n646,
    n673
  );


  nor
  g817
  (
    n847,
    n222,
    n676,
    n624,
    n686
  );


  xnor
  g818
  (
    n822,
    n192,
    n682,
    n191,
    n196
  );


  xor
  g819
  (
    n758,
    n623,
    n221,
    n243,
    n696
  );


  or
  g820
  (
    n836,
    n228,
    n198,
    n659,
    n213
  );


  xnor
  g821
  (
    n736,
    n670,
    n681,
    n708,
    n642
  );


  or
  g822
  (
    n803,
    n705,
    n686,
    n706,
    n574
  );


  xor
  g823
  (
    n800,
    n698,
    n220,
    n30,
    n623
  );


  or
  g824
  (
    n851,
    n223,
    n704,
    n228,
    n649
  );


  xor
  g825
  (
    n767,
    n634,
    n636,
    n707,
    n666
  );


  nand
  g826
  (
    n766,
    n682,
    n628,
    n631,
    n629
  );


  and
  g827
  (
    n756,
    n687,
    n573,
    n233,
    n689
  );


  nand
  g828
  (
    n719,
    n627,
    n194,
    n703,
    n666
  );


  nand
  g829
  (
    n727,
    n694,
    n220,
    n622,
    n568
  );


  xnor
  g830
  (
    n720,
    n575,
    n700,
    n626,
    n678
  );


  xnor
  g831
  (
    n838,
    n616,
    n219,
    n218,
    n188
  );


  nand
  g832
  (
    n731,
    n667,
    n198,
    n185,
    n665
  );


  xnor
  g833
  (
    n745,
    n239,
    n709,
    n667,
    n226
  );


  xnor
  g834
  (
    n872,
    n688,
    n656,
    n644,
    n237
  );


  xor
  g835
  (
    n826,
    n230,
    n224,
    n232,
    n703
  );


  and
  g836
  (
    n813,
    n644,
    n219,
    n238,
    n616
  );


  and
  g837
  (
    n757,
    n643,
    n192,
    n647,
    n635
  );


  or
  g838
  (
    n729,
    n216,
    n635,
    n634,
    n632
  );


  nand
  g839
  (
    n815,
    n663,
    n642,
    n707,
    n210
  );


  nand
  g840
  (
    n873,
    n840,
    n813,
    n499,
    n860
  );


  xnor
  g841
  (
    n874,
    n754,
    n846,
    n815,
    n729
  );


  xor
  g842
  (
    n907,
    n744,
    n755,
    n772,
    n831
  );


  xor
  g843
  (
    n994,
    n503,
    n813,
    n869,
    n860
  );


  xor
  g844
  (
    n990,
    n500,
    n867,
    n857,
    n777
  );


  nor
  g845
  (
    n977,
    n712,
    n720,
    n779,
    n732
  );


  or
  g846
  (
    n922,
    n765,
    n501,
    n819,
    n759
  );


  or
  g847
  (
    n902,
    n791,
    n839,
    n726,
    n725
  );


  nand
  g848
  (
    n976,
    n749,
    n719,
    n751,
    n780
  );


  and
  g849
  (
    n894,
    n748,
    n845,
    n820,
    n730
  );


  xnor
  g850
  (
    n941,
    n735,
    n764,
    n852,
    n503
  );


  xnor
  g851
  (
    n964,
    n843,
    n771,
    n441,
    n830
  );


  nand
  g852
  (
    n933,
    n827,
    n715,
    n870,
    n844
  );


  nor
  g853
  (
    n958,
    n502,
    n822,
    n838,
    n438
  );


  nor
  g854
  (
    n961,
    n821,
    n824,
    n865,
    n807
  );


  or
  g855
  (
    n997,
    n857,
    n716,
    n765,
    n757
  );


  nand
  g856
  (
    n978,
    n762,
    n864,
    n816,
    n739
  );


  and
  g857
  (
    n885,
    n734,
    n745,
    n728,
    n768
  );


  xor
  g858
  (
    n955,
    n871,
    n828,
    n439,
    n494
  );


  xor
  g859
  (
    n896,
    n499,
    n819,
    n835,
    n501
  );


  nor
  g860
  (
    n965,
    n837,
    n806,
    n860,
    n856
  );


  or
  g861
  (
    n995,
    n764,
    n761,
    n782,
    n824
  );


  xor
  g862
  (
    n884,
    n800,
    n857,
    n774,
    n799
  );


  or
  g863
  (
    n917,
    n835,
    n809,
    n743,
    n758
  );


  xor
  g864
  (
    n932,
    n830,
    n864,
    n797,
    n847
  );


  nor
  g865
  (
    n929,
    n718,
    n859,
    n823,
    n867
  );


  and
  g866
  (
    n935,
    n752,
    n866,
    n857,
    n724
  );


  xnor
  g867
  (
    n892,
    n803,
    n786,
    n750,
    n837
  );


  and
  g868
  (
    n943,
    n439,
    n803,
    n870,
    n817
  );


  nand
  g869
  (
    n887,
    n737,
    n871,
    n805,
    n786
  );


  xnor
  g870
  (
    n938,
    n727,
    n866,
    n710,
    n844
  );


  xor
  g871
  (
    n942,
    n785,
    n806,
    n822,
    n790
  );


  and
  g872
  (
    n973,
    n872,
    n823,
    n438,
    n862
  );


  xnor
  g873
  (
    n970,
    n828,
    n869,
    n836,
    n816
  );


  xnor
  g874
  (
    n881,
    n812,
    n805,
    n712,
    n822
  );


  xor
  g875
  (
    n975,
    n866,
    n868,
    n842,
    n858
  );


  xor
  g876
  (
    n918,
    n710,
    n812,
    n498,
    n865
  );


  nand
  g877
  (
    n927,
    n851,
    n494,
    n835,
    n804
  );


  xnor
  g878
  (
    n882,
    n437,
    n821,
    n841,
    n767
  );


  or
  g879
  (
    n948,
    n830,
    n787,
    n441,
    n789
  );


  nor
  g880
  (
    n987,
    n838,
    n440,
    n758,
    n794
  );


  nand
  g881
  (
    n969,
    n772,
    n747,
    n727,
    n501
  );


  nand
  g882
  (
    n924,
    n716,
    n856,
    n865,
    n736
  );


  and
  g883
  (
    n891,
    n811,
    n755,
    n812,
    n852
  );


  nor
  g884
  (
    n951,
    n776,
    n843,
    n761,
    n852
  );


  and
  g885
  (
    n899,
    n719,
    n859,
    n814,
    n834
  );


  xor
  g886
  (
    n993,
    n840,
    n869,
    n827,
    n731
  );


  nand
  g887
  (
    n926,
    n815,
    n833,
    n808,
    n438
  );


  xor
  g888
  (
    n998,
    n815,
    n863,
    n853,
    n725
  );


  xor
  g889
  (
    n963,
    n437,
    n802,
    n729,
    n438
  );


  and
  g890
  (
    n999,
    n818,
    n849,
    n836,
    n824
  );


  nand
  g891
  (
    n931,
    n773,
    n868,
    n778,
    n825
  );


  xnor
  g892
  (
    n984,
    n770,
    n739,
    n763,
    n734
  );


  xor
  g893
  (
    n880,
    n868,
    n793,
    n816,
    n503
  );


  or
  g894
  (
    n986,
    n497,
    n495,
    n503,
    n861
  );


  xnor
  g895
  (
    n879,
    n846,
    n809,
    n850,
    n751
  );


  nor
  g896
  (
    n979,
    n826,
    n733,
    n834,
    n441
  );


  xnor
  g897
  (
    n903,
    n826,
    n831,
    n847,
    n759
  );


  and
  g898
  (
    n966,
    n849,
    n831,
    n722,
    n795
  );


  or
  g899
  (
    n962,
    n753,
    n863,
    n495,
    n829
  );


  xnor
  g900
  (
    n991,
    n810,
    n818,
    n717,
    n842
  );


  nand
  g901
  (
    n901,
    n860,
    n837,
    n717,
    n825
  );


  nor
  g902
  (
    n906,
    n754,
    n730,
    n791,
    n781
  );


  nand
  g903
  (
    n960,
    n796,
    n437,
    n836,
    n841
  );


  xnor
  g904
  (
    n928,
    n867,
    n496,
    n820,
    n846
  );


  nand
  g905
  (
    n980,
    n817,
    n845,
    n784,
    n833
  );


  nand
  g906
  (
    n919,
    n798,
    n496,
    n840,
    n807
  );


  nor
  g907
  (
    n972,
    n748,
    n861,
    n817,
    n823
  );


  xor
  g908
  (
    n936,
    n778,
    n871,
    n851,
    n753
  );


  xnor
  g909
  (
    n920,
    n866,
    n854,
    n711,
    n439
  );


  or
  g910
  (
    n953,
    n721,
    n827,
    n845,
    n499
  );


  nor
  g911
  (
    n944,
    n811,
    n855,
    n835,
    n856
  );


  xnor
  g912
  (
    n921,
    n850,
    n752,
    n496,
    n771
  );


  nand
  g913
  (
    n949,
    n819,
    n830,
    n840,
    n861
  );


  xor
  g914
  (
    n908,
    n826,
    n818,
    n870,
    n781
  );


  and
  g915
  (
    n952,
    n841,
    n834,
    n728,
    n863
  );


  nand
  g916
  (
    n1000,
    n726,
    n847,
    n797,
    n826
  );


  and
  g917
  (
    n945,
    n747,
    n494,
    n824,
    n838
  );


  or
  g918
  (
    n915,
    n849,
    n777,
    n762,
    n838
  );


  nor
  g919
  (
    n897,
    n812,
    n832,
    n766,
    n825
  );


  nand
  g920
  (
    n946,
    n837,
    n774,
    n839,
    n871
  );


  nand
  g921
  (
    n937,
    n740,
    n862,
    n813,
    n497
  );


  xor
  g922
  (
    n959,
    n832,
    n502,
    n831,
    n796
  );


  xor
  g923
  (
    n895,
    n861,
    n802,
    n746,
    n864
  );


  xnor
  g924
  (
    n940,
    n440,
    n801,
    n843,
    n821
  );


  or
  g925
  (
    n878,
    n800,
    n783,
    n855,
    n769
  );


  or
  g926
  (
    n883,
    n849,
    n844,
    n848,
    n845
  );


  nor
  g927
  (
    n890,
    n848,
    n767,
    n850,
    n822
  );


  xnor
  g928
  (
    n898,
    n779,
    n872,
    n495,
    n783
  );


  nor
  g929
  (
    n983,
    n500,
    n869,
    n713,
    n497
  );


  xnor
  g930
  (
    n981,
    n742,
    n868,
    n821,
    n862
  );


  xor
  g931
  (
    n914,
    n780,
    n763,
    n801,
    n858
  );


  nand
  g932
  (
    n925,
    n834,
    n808,
    n851,
    n493
  );


  xor
  g933
  (
    n947,
    n863,
    n833,
    n740,
    n746
  );


  and
  g934
  (
    n886,
    n804,
    n832,
    n792,
    n776
  );


  xnor
  g935
  (
    n877,
    n789,
    n718,
    n501,
    n724
  );


  nor
  g936
  (
    n889,
    n735,
    n440,
    n496,
    n741
  );


  nand
  g937
  (
    n888,
    n825,
    n768,
    n766,
    n815
  );


  xnor
  g938
  (
    n909,
    n757,
    n814,
    n775,
    n817
  );


  or
  g939
  (
    n996,
    n723,
    n811,
    n502,
    n848
  );


  xor
  g940
  (
    n930,
    n798,
    n738,
    n852,
    n745
  );


  or
  g941
  (
    n971,
    n441,
    n782,
    n714,
    n721
  );


  and
  g942
  (
    n934,
    n722,
    n744,
    n858,
    n788
  );


  and
  g943
  (
    n904,
    n720,
    n736,
    n827,
    n829
  );


  or
  g944
  (
    n893,
    n864,
    n855,
    n499,
    n738
  );


  and
  g945
  (
    n985,
    n823,
    n500,
    n756,
    n819
  );


  nor
  g946
  (
    n900,
    n836,
    n498,
    n872,
    n795
  );


  or
  g947
  (
    n875,
    n829,
    n775,
    n498,
    n847
  );


  xnor
  g948
  (
    n967,
    n853,
    n816,
    n750,
    n713
  );


  xnor
  g949
  (
    n905,
    n440,
    n756,
    n493,
    n799
  );


  xor
  g950
  (
    n956,
    n813,
    n714,
    n853,
    n787
  );


  and
  g951
  (
    n968,
    n867,
    n773,
    n865,
    n828
  );


  nand
  g952
  (
    n923,
    n832,
    n493,
    n870,
    n502
  );


  and
  g953
  (
    n910,
    n810,
    n732,
    n770,
    n829
  );


  xnor
  g954
  (
    n950,
    n828,
    n731,
    n737,
    n858
  );


  and
  g955
  (
    n954,
    n872,
    n498,
    n814,
    n497
  );


  nor
  g956
  (
    n916,
    n794,
    n842,
    n741,
    n495
  );


  nor
  g957
  (
    n939,
    n859,
    n711,
    n855,
    n833
  );


  and
  g958
  (
    n989,
    n818,
    n844,
    n839,
    n854
  );


  nor
  g959
  (
    n913,
    n792,
    n854,
    n760,
    n715
  );


  nor
  g960
  (
    n992,
    n851,
    n856,
    n788,
    n500
  );


  nor
  g961
  (
    n911,
    n793,
    n841,
    n846,
    n814
  );


  or
  g962
  (
    n982,
    n843,
    n862,
    n854,
    n784
  );


  or
  g963
  (
    n974,
    n743,
    n494,
    n853,
    n439
  );


  or
  g964
  (
    n912,
    n760,
    n769,
    n842,
    n820
  );


  nand
  g965
  (
    n876,
    n749,
    n848,
    n790,
    n742
  );


  nand
  g966
  (
    n988,
    n811,
    n850,
    n733,
    n820
  );


  nor
  g967
  (
    n957,
    n785,
    n859,
    n839,
    n723
  );


  xnor
  g968
  (
    n1004,
    n878,
    n920,
    n958,
    n953
  );


  nor
  g969
  (
    n1008,
    n996,
    n905,
    n992,
    n933
  );


  or
  g970
  (
    n1021,
    n894,
    n909,
    n961,
    n918
  );


  nand
  g971
  (
    n1012,
    n881,
    n998,
    n934,
    n962
  );


  xnor
  g972
  (
    n1005,
    n883,
    n923,
    n874,
    n989
  );


  nor
  g973
  (
    n1029,
    n939,
    n899,
    n926,
    n1000
  );


  xor
  g974
  (
    n1023,
    n877,
    n959,
    n990,
    n936
  );


  or
  g975
  (
    n1003,
    n982,
    n978,
    n882,
    n980
  );


  nor
  g976
  (
    n1026,
    n949,
    n965,
    n979,
    n976
  );


  nand
  g977
  (
    n1013,
    n937,
    n960,
    n928,
    n999
  );


  and
  g978
  (
    n1025,
    n985,
    n925,
    n890,
    n993
  );


  and
  g979
  (
    n1010,
    n893,
    n900,
    n930,
    n895
  );


  xor
  g980
  (
    n1011,
    n947,
    n903,
    n889,
    n946
  );


  xnor
  g981
  (
    n1015,
    n885,
    n897,
    n932,
    n983
  );


  and
  g982
  (
    AntiSAT_key_wire,
    n986,
    n921,
    n951,
    n945
  );


  xor
  g983
  (
    n1019,
    n964,
    n922,
    n896,
    n944
  );


  nand
  g984
  (
    n1027,
    n876,
    n888,
    n913,
    n910
  );


  xnor
  g985
  (
    n1009,
    n919,
    n972,
    n943,
    n935
  );


  xnor
  g986
  (
    n1028,
    n908,
    n954,
    n955,
    n880
  );


  and
  g987
  (
    n1017,
    n940,
    n884,
    n929,
    n892
  );


  xor
  g988
  (
    n1024,
    n995,
    n912,
    n991,
    n963
  );


  nand
  g989
  (
    n1030,
    n974,
    n952,
    n956,
    n970
  );


  nor
  g990
  (
    n1016,
    n975,
    n948,
    n994,
    n927
  );


  nand
  g991
  (
    n1032,
    n906,
    n988,
    n931,
    n969
  );


  xnor
  g992
  (
    n1014,
    n981,
    n917,
    n987,
    n967
  );


  nor
  g993
  (
    n1002,
    n957,
    n941,
    n875,
    n942
  );


  xnor
  g994
  (
    n1020,
    n911,
    n916,
    n887,
    n915
  );


  xnor
  g995
  (
    n1007,
    n977,
    n886,
    n966,
    n984
  );


  nor
  g996
  (
    n1006,
    n898,
    n907,
    n971,
    n968
  );


  and
  g997
  (
    n1022,
    n873,
    n904,
    n902,
    n924
  );


  xor
  g998
  (
    n1001,
    n938,
    n950,
    n891,
    n914
  );


  nand
  g999
  (
    n1031,
    n997,
    n901,
    n973,
    n879
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n1018,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

