

module Stat_100_55
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n98,
  n103,
  n107,
  n109,
  n104,
  n112,
  n131,
  n117,
  n113,
  n126,
  n116,
  n120,
  n114,
  n115,
  n132,
  n108,
  n127,
  n121,
  n122,
  n128,
  n111,
  n106,
  n125,
  n123,
  n102,
  n118,
  n105,
  n129,
  n110,
  n119,
  n130,
  n124
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n98;output n103;output n107;output n109;output n104;output n112;output n131;output n117;output n113;output n126;output n116;output n120;output n114;output n115;output n132;output n108;output n127;output n121;output n122;output n128;output n111;output n106;output n125;output n123;output n102;output n118;output n105;output n129;output n110;output n119;output n130;output n124;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n99;wire n100;wire n101;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  not
  g0
  (
    n33,
    n9
  );


  buf
  g1
  (
    n37,
    n4
  );


  buf
  g2
  (
    n42,
    n6
  );


  buf
  g3
  (
    KeyWire_0_4,
    n10
  );


  buf
  g4
  (
    KeyWire_0_58,
    n3
  );


  buf
  g5
  (
    KeyWire_0_3,
    n2
  );


  buf
  g6
  (
    KeyWire_0_43,
    n5
  );


  buf
  g7
  (
    KeyWire_0_59,
    n1
  );


  buf
  g8
  (
    KeyWire_0_17,
    n8
  );


  not
  g9
  (
    n35,
    n7
  );


  buf
  g10
  (
    KeyWire_0_29,
    n36
  );


  not
  g11
  (
    KeyWire_0_32,
    n35
  );


  not
  g12
  (
    KeyWire_0_0,
    n36
  );


  not
  g13
  (
    n61,
    n34
  );


  buf
  g14
  (
    KeyWire_0_46,
    n38
  );


  buf
  g15
  (
    KeyWire_0_16,
    n12
  );


  not
  g16
  (
    n62,
    n37
  );


  buf
  g17
  (
    n52,
    n38
  );


  buf
  g18
  (
    KeyWire_0_30,
    n37
  );


  not
  g19
  (
    KeyWire_0_15,
    n40
  );


  not
  g20
  (
    KeyWire_0_19,
    n35
  );


  not
  g21
  (
    KeyWire_0_26,
    n38
  );


  buf
  g22
  (
    n60,
    n11
  );


  buf
  g23
  (
    KeyWire_0_9,
    n38
  );


  buf
  g24
  (
    KeyWire_0_1,
    n34
  );


  buf
  g25
  (
    KeyWire_0_31,
    n37
  );


  buf
  g26
  (
    KeyWire_0_54,
    n39
  );


  not
  g27
  (
    KeyWire_0_49,
    n40
  );


  not
  g28
  (
    n76,
    n13
  );


  not
  g29
  (
    KeyWire_0_48,
    n39
  );


  buf
  g30
  (
    n56,
    n33
  );


  not
  g31
  (
    KeyWire_0_52,
    n36
  );


  not
  g32
  (
    n58,
    n33
  );


  buf
  g33
  (
    n53,
    n41
  );


  not
  g34
  (
    KeyWire_0_11,
    n35
  );


  not
  g35
  (
    KeyWire_0_53,
    n33
  );


  buf
  g36
  (
    n71,
    n34
  );


  not
  g37
  (
    KeyWire_0_33,
    n35
  );


  buf
  g38
  (
    KeyWire_0_25,
    n33
  );


  not
  g39
  (
    KeyWire_0_50,
    n37
  );


  buf
  g40
  (
    KeyWire_0_36,
    n39
  );


  not
  g41
  (
    KeyWire_0_14,
    n40
  );


  buf
  g42
  (
    KeyWire_0_51,
    n39
  );


  buf
  g43
  (
    KeyWire_0_2,
    n36
  );


  or
  g44
  (
    KeyWire_0_60,
    n40,
    n34,
    n41
  );


  nor
  g45
  (
    KeyWire_0_24,
    n22,
    n46,
    n24,
    n32
  );


  nor
  g46
  (
    n80,
    n32,
    n32,
    n16,
    n31
  );


  nand
  g47
  (
    n81,
    n43,
    n29,
    n47,
    n23
  );


  and
  g48
  (
    n79,
    n18,
    n45,
    n20,
    n21
  );


  nand
  g49
  (
    n82,
    n30,
    n30,
    n44,
    n14
  );


  or
  g50
  (
    n85,
    n28,
    n19,
    n25,
    n50
  );


  or
  g51
  (
    KeyWire_0_35,
    n51,
    n49,
    n17,
    n27
  );


  nor
  g52
  (
    KeyWire_0_28,
    n26,
    n31,
    n48,
    n15
  );


  buf
  g53
  (
    KeyWire_0_42,
    n80
  );


  not
  g54
  (
    KeyWire_0_62,
    n83
  );


  not
  g55
  (
    n86,
    n53
  );


  not
  g56
  (
    KeyWire_0_37,
    n42
  );


  not
  g57
  (
    n94,
    n42
  );


  not
  g58
  (
    n91,
    n83
  );


  buf
  g59
  (
    n88,
    n32
  );


  buf
  g60
  (
    KeyWire_0_20,
    n55
  );


  buf
  g61
  (
    n99,
    n55
  );


  buf
  g62
  (
    KeyWire_0_18,
    n83
  );


  xor
  g63
  (
    KeyWire_0_57,
    n54,
    n82
  );


  and
  g64
  (
    KeyWire_0_44,
    n79,
    n85,
    n41,
    n84
  );


  or
  g65
  (
    KeyWire_0_41,
    n52,
    n84,
    n82
  );


  and
  g66
  (
    n93,
    n82,
    n54,
    n42
  );


  and
  g67
  (
    KeyWire_0_27,
    n84,
    n53,
    n54,
    n83
  );


  xor
  g68
  (
    KeyWire_0_45,
    n84,
    n42,
    n81,
    n78
  );


  and
  g69
  (
    KeyWire_0_7,
    n58,
    n73,
    n65,
    n62
  );


  or
  g70
  (
    KeyWire_0_38,
    n68,
    n70,
    n61,
    n69
  );


  nand
  g71
  (
    n106,
    n59,
    n61,
    n56,
    n100
  );


  or
  g72
  (
    n128,
    n74,
    n66,
    n72,
    n62
  );


  xnor
  g73
  (
    KeyWire_0_23,
    n55,
    n70,
    n63,
    n92
  );


  xnor
  g74
  (
    KeyWire_0_63,
    n87,
    n56,
    n64,
    n95
  );


  nor
  g75
  (
    KeyWire_0_40,
    n67,
    n88,
    n61,
    n60
  );


  xor
  g76
  (
    KeyWire_0_22,
    n68,
    n77,
    n74,
    n64
  );


  nor
  g77
  (
    n110,
    n75,
    n101,
    n55,
    n67
  );


  or
  g78
  (
    KeyWire_0_21,
    n65,
    n97,
    n71,
    n60
  );


  xor
  g79
  (
    KeyWire_0_61,
    n56,
    n62,
    n99,
    n100
  );


  xor
  g80
  (
    n111,
    n100,
    n62,
    n74,
    n91
  );


  xnor
  g81
  (
    KeyWire_0_10,
    n96,
    n58,
    n67,
    n90
  );


  nand
  g82
  (
    n121,
    n57,
    n66,
    n99,
    n69
  );


  nor
  g83
  (
    n116,
    n75,
    n69,
    n59,
    n94
  );


  xnor
  g84
  (
    n118,
    n72,
    n97,
    n61,
    n98
  );


  nand
  g85
  (
    n112,
    n75,
    n59,
    n57,
    n100
  );


  and
  g86
  (
    KeyWire_0_12,
    n64,
    n85,
    n58,
    n77
  );


  and
  g87
  (
    n103,
    n69,
    n98,
    n65
  );


  xnor
  g88
  (
    n102,
    n56,
    n76,
    n73
  );


  xnor
  g89
  (
    n130,
    n89,
    n59,
    n97,
    n74
  );


  nand
  g90
  (
    KeyWire_0_55,
    n101,
    n66,
    n71
  );


  nor
  g91
  (
    KeyWire_0_56,
    n76,
    n97,
    n71,
    n86
  );


  xnor
  g92
  (
    KeyWire_0_34,
    n63,
    n63,
    n99,
    n75
  );


  xnor
  g93
  (
    KeyWire_0_47,
    n60,
    n76,
    n85,
    n101
  );


  and
  g94
  (
    n105,
    n77,
    n73,
    n72,
    n68
  );


  and
  g95
  (
    KeyWire_0_39,
    n57,
    n70,
    n66,
    n85
  );


  xor
  g96
  (
    KeyWire_0_6,
    n99,
    n68,
    n73,
    n58
  );


  nand
  g97
  (
    KeyWire_0_8,
    n64,
    n98,
    n101,
    n70
  );


  nand
  g98
  (
    KeyWire_0_5,
    n93,
    n63,
    n65,
    n67
  );


  and
  g99
  (
    KeyWire_0_13,
    n72,
    n57,
    n60,
    n77
  );


  xor
  KeyGate_0_0
  (
    n59,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n63,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n51,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n36,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n41,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n129,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n117,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n132,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n119,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n50,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n126,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n54,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n107,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n131,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n73,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n49,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n57,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n40,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n101,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n69,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n87,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n125,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n114,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n108,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n78,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n45,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n77,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n95,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n84,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n74,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n67,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n70,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n46,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n66,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n124,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n83,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n75,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n100,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n115,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n127,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n104,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n90,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n92,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n34,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n96,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n98,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n44,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n113,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n68,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n65,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n55,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n72,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n64,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n43,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n47,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n109,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n122,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n89,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n38,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n39,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n48,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n120,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n97,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n123,
    KeyNOTWire_0_63
  );


endmodule


