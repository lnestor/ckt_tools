

module Stat_100_43
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n108,
  n118,
  n127,
  n131,
  n124,
  n115,
  n125,
  n116,
  n101,
  n126,
  n129,
  n111,
  n112,
  n110,
  n120,
  n123,
  n104,
  n130,
  n113,
  n132,
  n128,
  n102,
  n114,
  n119,
  n109,
  n121,
  n122,
  n105,
  n106,
  n107,
  n117,
  n103,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n108;
  output n118;
  output n127;
  output n131;
  output n124;
  output n115;
  output n125;
  output n116;
  output n101;
  output n126;
  output n129;
  output n111;
  output n112;
  output n110;
  output n120;
  output n123;
  output n104;
  output n130;
  output n113;
  output n132;
  output n128;
  output n102;
  output n114;
  output n119;
  output n109;
  output n121;
  output n122;
  output n105;
  output n106;
  output n107;
  output n117;
  output n103;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    KeyWire_0_27,
    n3
  );


  not
  g1
  (
    n46,
    n4
  );


  not
  g2
  (
    KeyWire_0_20,
    n2
  );


  buf
  g3
  (
    KeyWire_0_13,
    n2
  );


  not
  g4
  (
    KeyWire_0_48,
    n2
  );


  not
  g5
  (
    n47,
    n1
  );


  not
  g6
  (
    KeyWire_0_14,
    n1
  );


  not
  g7
  (
    KeyWire_0_46,
    n3
  );


  not
  g8
  (
    KeyWire_0_8,
    n3
  );


  not
  g9
  (
    n37,
    n3
  );


  not
  g10
  (
    n40,
    n4
  );


  not
  g11
  (
    KeyWire_0_41,
    n1
  );


  buf
  g12
  (
    n34,
    n4
  );


  not
  g13
  (
    n41,
    n1
  );


  buf
  g14
  (
    n42,
    n2
  );


  buf
  g15
  (
    n55,
    n7
  );


  not
  g16
  (
    KeyWire_0_42,
    n44
  );


  not
  g17
  (
    KeyWire_0_11,
    n24
  );


  not
  g18
  (
    KeyWire_0_16,
    n27
  );


  not
  g19
  (
    KeyWire_0_33,
    n38
  );


  buf
  g20
  (
    KeyWire_0_60,
    n35
  );


  or
  g21
  (
    KeyWire_0_21,
    n12,
    n9,
    n13
  );


  xnor
  g22
  (
    KeyWire_0_40,
    n34,
    n24,
    n8,
    n7
  );


  nand
  g23
  (
    n88,
    n38,
    n5,
    n22,
    n21
  );


  xor
  g24
  (
    KeyWire_0_34,
    n29,
    n11,
    n31,
    n39
  );


  xor
  g25
  (
    KeyWire_0_52,
    n37,
    n30,
    n20,
    n43
  );


  and
  g26
  (
    KeyWire_0_24,
    n23,
    n20,
    n14,
    n44
  );


  xnor
  g27
  (
    KeyWire_0_17,
    n27,
    n10,
    n34,
    n15
  );


  nand
  g28
  (
    KeyWire_0_57,
    n39,
    n19,
    n17,
    n37
  );


  nand
  g29
  (
    n72,
    n34,
    n15,
    n29,
    n31
  );


  xnor
  g30
  (
    n64,
    n41,
    n37,
    n6,
    n26
  );


  nor
  g31
  (
    n75,
    n22,
    n22,
    n30,
    n35
  );


  nand
  g32
  (
    KeyWire_0_2,
    n29,
    n44,
    n18,
    n17
  );


  nand
  g33
  (
    n56,
    n33,
    n29,
    n10,
    n17
  );


  xor
  g34
  (
    KeyWire_0_19,
    n43,
    n28,
    n41,
    n14
  );


  or
  g35
  (
    n81,
    n32,
    n21,
    n42,
    n26
  );


  or
  g36
  (
    KeyWire_0_18,
    n17,
    n12,
    n30,
    n26
  );


  nand
  g37
  (
    KeyWire_0_63,
    n16,
    n9,
    n26,
    n43
  );


  xor
  g38
  (
    KeyWire_0_44,
    n31,
    n42,
    n20,
    n30
  );


  xnor
  g39
  (
    n82,
    n21,
    n19,
    n6,
    n5
  );


  and
  g40
  (
    KeyWire_0_6,
    n45,
    n16,
    n9,
    n23
  );


  xor
  g41
  (
    n86,
    n18,
    n18,
    n24,
    n36
  );


  xor
  g42
  (
    KeyWire_0_32,
    n44,
    n11,
    n5,
    n25
  );


  nor
  g43
  (
    n67,
    n45,
    n40,
    n19,
    n42
  );


  and
  g44
  (
    KeyWire_0_23,
    n25,
    n12,
    n38,
    n22
  );


  xor
  g45
  (
    KeyWire_0_43,
    n32,
    n42,
    n8,
    n35
  );


  nor
  g46
  (
    KeyWire_0_38,
    n40,
    n14,
    n15,
    n7
  );


  and
  g47
  (
    n66,
    n23,
    n15,
    n37,
    n32
  );


  and
  g48
  (
    KeyWire_0_53,
    n28,
    n5,
    n25,
    n41
  );


  nand
  g49
  (
    KeyWire_0_50,
    n16,
    n23,
    n31,
    n34
  );


  and
  g50
  (
    KeyWire_0_61,
    n16,
    n45,
    n6,
    n10
  );


  or
  g51
  (
    KeyWire_0_29,
    n39,
    n9,
    n25,
    n7
  );


  nor
  g52
  (
    n60,
    n36,
    n40,
    n35,
    n38
  );


  xor
  g53
  (
    KeyWire_0_36,
    n14,
    n28,
    n36
  );


  nor
  g54
  (
    n58,
    n21,
    n40,
    n27,
    n43
  );


  nand
  g55
  (
    KeyWire_0_45,
    n41,
    n8,
    n28
  );


  nand
  g56
  (
    KeyWire_0_31,
    n18,
    n27,
    n11
  );


  xnor
  g57
  (
    n65,
    n12,
    n13,
    n24
  );


  nand
  g58
  (
    KeyWire_0_51,
    n39,
    n4,
    n10,
    n6
  );


  and
  g59
  (
    KeyWire_0_5,
    n20,
    n45,
    n19,
    n32
  );


  buf
  g60
  (
    KeyWire_0_59,
    n51
  );


  not
  g61
  (
    KeyWire_0_26,
    n47
  );


  not
  g62
  (
    KeyWire_0_35,
    n48
  );


  not
  g63
  (
    KeyWire_0_30,
    n50
  );


  xor
  g64
  (
    KeyWire_0_15,
    n47,
    n58,
    n46
  );


  nand
  g65
  (
    n93,
    n47,
    n49,
    n57,
    n53
  );


  xnor
  g66
  (
    n94,
    n56,
    n46,
    n52
  );


  nor
  g67
  (
    n98,
    n47,
    n59,
    n54,
    n55
  );


  or
  g68
  (
    KeyWire_0_22,
    n90,
    n75,
    n87,
    n83
  );


  xor
  g69
  (
    n104,
    n96,
    n90,
    n79,
    n89
  );


  xnor
  g70
  (
    n106,
    n67,
    n72,
    n60,
    n90
  );


  nand
  g71
  (
    KeyWire_0_1,
    n81,
    n61,
    n84,
    n93
  );


  nor
  g72
  (
    n113,
    n85,
    n73,
    n77,
    n93
  );


  xnor
  g73
  (
    KeyWire_0_3,
    n97,
    n80,
    n83,
    n89
  );


  xor
  g74
  (
    KeyWire_0_9,
    n85,
    n95,
    n99,
    n90
  );


  xor
  g75
  (
    KeyWire_0_25,
    n99,
    n89,
    n77,
    n68
  );


  or
  g76
  (
    n117,
    n75,
    n74,
    n78,
    n92
  );


  xnor
  g77
  (
    KeyWire_0_7,
    n81,
    n76,
    n72,
    n85
  );


  nor
  g78
  (
    n123,
    n85,
    n77,
    n82,
    n92
  );


  nor
  g79
  (
    KeyWire_0_39,
    n89,
    n76,
    n70,
    n64
  );


  nand
  g80
  (
    KeyWire_0_47,
    n100,
    n74,
    n96,
    n95
  );


  xnor
  g81
  (
    KeyWire_0_58,
    n83,
    n75,
    n93,
    n73
  );


  xnor
  g82
  (
    KeyWire_0_56,
    n96,
    n88,
    n95,
    n79
  );


  xnor
  g83
  (
    KeyWire_0_37,
    n80,
    n65,
    n81,
    n73
  );


  xor
  g84
  (
    n112,
    n86,
    n87,
    n91,
    n97
  );


  or
  g85
  (
    n111,
    n100,
    n82,
    n66,
    n72
  );


  nor
  g86
  (
    KeyWire_0_54,
    n100,
    n96,
    n93,
    n92
  );


  xnor
  g87
  (
    KeyWire_0_62,
    n94,
    n95,
    n62,
    n86
  );


  or
  g88
  (
    KeyWire_0_10,
    n79,
    n78,
    n98,
    n81
  );


  nand
  g89
  (
    n101,
    n84,
    n94,
    n72,
    n88
  );


  xor
  g90
  (
    n105,
    n91,
    n77,
    n97,
    n71
  );


  xnor
  g91
  (
    n110,
    n98,
    n86,
    n99,
    n97
  );


  xor
  g92
  (
    n124,
    n91,
    n82,
    n74,
    n76
  );


  or
  g93
  (
    KeyWire_0_28,
    n94,
    n94,
    n87,
    n76
  );


  xnor
  g94
  (
    KeyWire_0_0,
    n86,
    n88,
    n78,
    n82
  );


  nand
  g95
  (
    KeyWire_0_55,
    n63,
    n73,
    n99,
    n80
  );


  and
  g96
  (
    n103,
    n74,
    n79,
    n84,
    n91
  );


  nand
  g97
  (
    KeyWire_0_4,
    n92,
    n88,
    n80,
    n98
  );


  and
  g98
  (
    KeyWire_0_49,
    n87,
    n75,
    n100,
    n69
  );


  or
  g99
  (
    KeyWire_0_12,
    n83,
    n84,
    n98,
    n78
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n115,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n130,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n77,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n122,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n119,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n74,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n84,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n125,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n36,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n109,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n131,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n49,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n120,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n39,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n38,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n96,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n57,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n48,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n91,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n53,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n33,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n79,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n102,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n62,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n92,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n118,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n100,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n43,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n132,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n59,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n99,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n70,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n80,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n63,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n78,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n95,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n54,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n127,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n83,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n114,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n89,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n45,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n76,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n87,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n52,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n69,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n35,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n128,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n44,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n121,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n68,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n85,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n51,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n90,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n126,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n108,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n107,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n71,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n129,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n97,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n73,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n50,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n116,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n61,
    KeyNOTWire_0_63
  );


endmodule

