// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_114_49 written by SynthGen on 2021/05/24 19:42:17
module Stat_114_49( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17,
 n130, n118, n131, n123, n115, n117, n114, n120,
 n128, n121, n119, n126, n129, n124, n116, n125,
 n127, n122, n113);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17;

output n130, n118, n131, n123, n115, n117, n114, n120,
 n128, n121, n119, n126, n129, n124, n116, n125,
 n127, n122, n113;

wire n18, n19, n20, n21, n22, n23, n24, n25,
 n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112;

buf  g0 (n32, n17);
buf  g1 (n26, n7);
buf  g2 (n20, n11);
not  g3 (n24, n6);
not  g4 (n18, n9);
buf  g5 (n25, n17);
buf  g6 (n23, n12);
buf  g7 (n28, n15);
buf  g8 (n30, n14);
not  g9 (n35, n13);
buf  g10 (n27, n10);
not  g11 (n22, n16);
buf  g12 (n34, n5);
not  g13 (n33, n3);
buf  g14 (n21, n1);
buf  g15 (n19, n4);
buf  g16 (n31, n2);
buf  g17 (n29, n8);
not  g18 (n41, n31);
buf  g19 (n63, n34);
not  g20 (n43, n24);
not  g21 (n65, n20);
buf  g22 (n52, n27);
not  g23 (n39, n35);
not  g24 (n64, n19);
buf  g25 (n49, n26);
not  g26 (n42, n24);
buf  g27 (n45, n35);
not  g28 (n36, n27);
not  g29 (n48, n29);
not  g30 (n72, n30);
buf  g31 (n50, n35);
not  g32 (n60, n31);
not  g33 (n70, n33);
buf  g34 (n55, n22);
not  g35 (n44, n18);
not  g36 (n66, n29);
not  g37 (n61, n23);
not  g38 (n37, n22);
buf  g39 (n68, n18);
not  g40 (n40, n34);
not  g41 (n47, n28);
not  g42 (n56, n34);
buf  g43 (n69, n25);
not  g44 (n38, n30);
buf  g45 (n58, n20);
buf  g46 (n51, n19);
buf  g47 (n57, n33);
buf  g48 (n73, n28);
buf  g49 (n62, n23);
buf  g50 (n54, n32);
not  g51 (n46, n21);
not  g52 (n67, n26);
not  g53 (n71, n21);
buf  g54 (n53, n32);
not  g55 (n59, n25);
not  g56 (n76, n49);
not  g57 (n104, n68);
buf  g58 (n100, n39);
buf  g59 (n107, n38);
buf  g60 (n74, n55);
buf  g61 (n106, n43);
not  g62 (n94, n37);
buf  g63 (n92, n42);
buf  g64 (n90, n51);
not  g65 (n75, n65);
buf  g66 (n83, n66);
not  g67 (n112, n60);
not  g68 (n103, n64);
buf  g69 (n91, n53);
buf  g70 (n78, n69);
not  g71 (n93, n40);
buf  g72 (n97, n72);
not  g73 (n96, n36);
buf  g74 (n85, n46);
buf  g75 (n98, n48);
not  g76 (n79, n71);
buf  g77 (n88, n57);
buf  g78 (n105, n73);
buf  g79 (n89, n58);
not  g80 (n99, n61);
buf  g81 (n101, n41);
buf  g82 (n102, n54);
not  g83 (n86, n59);
not  g84 (n77, n52);
not  g85 (n84, n67);
not  g86 (n110, n73);
not  g87 (n80, n63);
buf  g88 (n87, n62);
buf  g89 (n109, n56);
buf  g90 (n82, n50);
not  g91 (n111, n70);
not  g92 (n108, n44);
buf  g93 (n81, n45);
not  g94 (n95, n47);
not  g95 (n115, n88);
buf  g96 (n123, n108);
not  g97 (n129, n107);
buf  g98 (n124, n106);
buf  g99 (n119, n75);
buf  g100 (n128, n100);
buf  g101 (n126, n98);
buf  g102 (n131, n78);
not  g103 (n125, n82);
not  g104 (n120, n93);
not  g105 (n127, n110);
not  g106 (n121, n94);
xnor g107 (n116, n105, n101, n92);
xor  g108 (n130, n102, n109, n87, n96);
and  g109 (n118, n91, n97, n77, n99);
xor  g110 (n114, n80, n90, n76, n79);
nor  g111 (n117, n74, n111, n95, n83);
nand g112 (n113, n81, n104, n112, n86);
or   g113 (n122, n84, n103, n89, n85);
endmodule
