

module Stat_1000_155
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n225,
  n588,
  n589,
  n597,
  n596,
  n602,
  n585,
  n600,
  n592,
  n581,
  n595,
  n593,
  n616,
  n619,
  n622,
  n1032,
  n1016,
  n1029,
  n1020,
  n1031,
  n1021,
  n1022,
  n1023,
  n1027,
  n1026,
  n1024,
  n1018,
  n1028,
  n1017,
  n1019,
  n1030,
  n1025,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n225;output n588;output n589;output n597;output n596;output n602;output n585;output n600;output n592;output n581;output n595;output n593;output n616;output n619;output n622;output n1032;output n1016;output n1029;output n1020;output n1031;output n1021;output n1022;output n1023;output n1027;output n1026;output n1024;output n1018;output n1028;output n1017;output n1019;output n1030;output n1025;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n582;wire n583;wire n584;wire n586;wire n587;wire n590;wire n591;wire n594;wire n598;wire n599;wire n601;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n617;wire n618;wire n620;wire n621;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  buf
  g0
  (
    n37,
    n2
  );


  buf
  g1
  (
    n54,
    n1
  );


  buf
  g2
  (
    n53,
    n4
  );


  buf
  g3
  (
    n38,
    n3
  );


  buf
  g4
  (
    n56,
    n3
  );


  buf
  g5
  (
    n40,
    n2
  );


  not
  g6
  (
    n51,
    n6
  );


  not
  g7
  (
    n57,
    n3
  );


  buf
  g8
  (
    n43,
    n4
  );


  not
  g9
  (
    n41,
    n6
  );


  buf
  g10
  (
    n35,
    n1
  );


  not
  g11
  (
    n47,
    n5
  );


  not
  g12
  (
    n55,
    n5
  );


  buf
  g13
  (
    n36,
    n2
  );


  buf
  g14
  (
    n58,
    n5
  );


  not
  g15
  (
    n52,
    n7
  );


  not
  g16
  (
    n44,
    n2
  );


  buf
  g17
  (
    n46,
    n1
  );


  not
  g18
  (
    n59,
    n6
  );


  not
  g19
  (
    n50,
    n1
  );


  not
  g20
  (
    n49,
    n7
  );


  buf
  g21
  (
    n34,
    n6
  );


  buf
  g22
  (
    n48,
    n4
  );


  buf
  g23
  (
    n45,
    n7
  );


  buf
  g24
  (
    n33,
    n3
  );


  buf
  g25
  (
    n42,
    n4
  );


  buf
  g26
  (
    n39,
    n5
  );


  not
  g27
  (
    n88,
    n36
  );


  buf
  g28
  (
    n60,
    n34
  );


  buf
  g29
  (
    n64,
    n36
  );


  not
  g30
  (
    n69,
    n38
  );


  not
  g31
  (
    n67,
    n43
  );


  not
  g32
  (
    n76,
    n43
  );


  buf
  g33
  (
    n63,
    n34
  );


  buf
  g34
  (
    n79,
    n35
  );


  not
  g35
  (
    n86,
    n38
  );


  buf
  g36
  (
    n61,
    n39
  );


  buf
  g37
  (
    n62,
    n42
  );


  not
  g38
  (
    n83,
    n43
  );


  not
  g39
  (
    n66,
    n41
  );


  not
  g40
  (
    n70,
    n40
  );


  not
  g41
  (
    n77,
    n42
  );


  not
  g42
  (
    n75,
    n41
  );


  not
  g43
  (
    n78,
    n42
  );


  buf
  g44
  (
    n65,
    n43
  );


  buf
  g45
  (
    KeyWire_0_26,
    n37
  );


  buf
  g46
  (
    n71,
    n41
  );


  not
  g47
  (
    n85,
    n42
  );


  buf
  g48
  (
    n74,
    n36
  );


  buf
  g49
  (
    n90,
    n33
  );


  buf
  g50
  (
    n80,
    n40
  );


  not
  g51
  (
    n68,
    n40
  );


  not
  g52
  (
    n87,
    n41
  );


  buf
  g53
  (
    n89,
    n35
  );


  buf
  g54
  (
    n82,
    n37
  );


  not
  g55
  (
    n72,
    n37
  );


  buf
  g56
  (
    n84,
    n40
  );


  xor
  g57
  (
    n81,
    n33,
    n38,
    n44,
    n39
  );


  and
  g58
  (
    n91,
    n33,
    n34,
    n35,
    n39
  );


  not
  g59
  (
    n161,
    n76
  );


  buf
  g60
  (
    KeyWire_0_21,
    n87
  );


  buf
  g61
  (
    n183,
    n64
  );


  buf
  g62
  (
    n172,
    n63
  );


  not
  g63
  (
    n177,
    n64
  );


  not
  g64
  (
    n135,
    n65
  );


  buf
  g65
  (
    n189,
    n66
  );


  buf
  g66
  (
    n120,
    n72
  );


  buf
  g67
  (
    n192,
    n84
  );


  buf
  g68
  (
    n153,
    n63
  );


  not
  g69
  (
    n190,
    n65
  );


  not
  g70
  (
    n111,
    n82
  );


  not
  g71
  (
    n100,
    n76
  );


  not
  g72
  (
    n103,
    n44
  );


  not
  g73
  (
    n152,
    n72
  );


  buf
  g74
  (
    n169,
    n73
  );


  not
  g75
  (
    n159,
    n79
  );


  buf
  g76
  (
    n147,
    n61
  );


  not
  g77
  (
    n197,
    n84
  );


  buf
  g78
  (
    n99,
    n7
  );


  buf
  g79
  (
    n92,
    n67
  );


  buf
  g80
  (
    n155,
    n60
  );


  buf
  g81
  (
    n146,
    n81
  );


  buf
  g82
  (
    n173,
    n78
  );


  buf
  g83
  (
    n141,
    n79
  );


  not
  g84
  (
    n105,
    n81
  );


  buf
  g85
  (
    n127,
    n63
  );


  buf
  g86
  (
    n138,
    n60
  );


  not
  g87
  (
    n193,
    n75
  );


  buf
  g88
  (
    n96,
    n70
  );


  not
  g89
  (
    n196,
    n69
  );


  buf
  g90
  (
    n191,
    n81
  );


  buf
  g91
  (
    n98,
    n85
  );


  buf
  g92
  (
    n118,
    n80
  );


  not
  g93
  (
    n206,
    n75
  );


  buf
  g94
  (
    n200,
    n84
  );


  not
  g95
  (
    n150,
    n85
  );


  not
  g96
  (
    n93,
    n68
  );


  not
  g97
  (
    KeyWire_0_6,
    n71
  );


  not
  g98
  (
    n195,
    n80
  );


  not
  g99
  (
    n95,
    n76
  );


  buf
  g100
  (
    n182,
    n87
  );


  buf
  g101
  (
    n198,
    n65
  );


  not
  g102
  (
    n139,
    n44
  );


  buf
  g103
  (
    n106,
    n61
  );


  buf
  g104
  (
    n125,
    n66
  );


  buf
  g105
  (
    n115,
    n60
  );


  buf
  g106
  (
    n174,
    n79
  );


  buf
  g107
  (
    n123,
    n78
  );


  buf
  g108
  (
    n122,
    n85
  );


  buf
  g109
  (
    n107,
    n74
  );


  buf
  g110
  (
    n187,
    n86
  );


  not
  g111
  (
    n124,
    n67
  );


  not
  g112
  (
    n188,
    n65
  );


  not
  g113
  (
    n149,
    n80
  );


  buf
  g114
  (
    n205,
    n86
  );


  not
  g115
  (
    n128,
    n64
  );


  not
  g116
  (
    n143,
    n71
  );


  not
  g117
  (
    n94,
    n77
  );


  buf
  g118
  (
    n130,
    n70
  );


  not
  g119
  (
    n112,
    n86
  );


  not
  g120
  (
    n151,
    n77
  );


  buf
  g121
  (
    n126,
    n83
  );


  not
  g122
  (
    n181,
    n71
  );


  not
  g123
  (
    n204,
    n81
  );


  not
  g124
  (
    n102,
    n87
  );


  not
  g125
  (
    n170,
    n73
  );


  not
  g126
  (
    n108,
    n67
  );


  buf
  g127
  (
    n160,
    n88
  );


  buf
  g128
  (
    n158,
    n73
  );


  buf
  g129
  (
    KeyWire_0_2,
    n66
  );


  not
  g130
  (
    n201,
    n72
  );


  buf
  g131
  (
    n113,
    n88
  );


  not
  g132
  (
    n176,
    n63
  );


  buf
  g133
  (
    n144,
    n69
  );


  not
  g134
  (
    n110,
    n75
  );


  not
  g135
  (
    n154,
    n74
  );


  not
  g136
  (
    n142,
    n61
  );


  buf
  g137
  (
    n186,
    n68
  );


  not
  g138
  (
    n185,
    n85
  );


  not
  g139
  (
    n202,
    n82
  );


  buf
  g140
  (
    n180,
    n72
  );


  not
  g141
  (
    n148,
    n74
  );


  buf
  g142
  (
    KeyWire_0_16,
    n75
  );


  not
  g143
  (
    n136,
    n77
  );


  buf
  g144
  (
    n101,
    n78
  );


  not
  g145
  (
    n166,
    n77
  );


  buf
  g146
  (
    n175,
    n79
  );


  buf
  g147
  (
    n145,
    n69
  );


  buf
  g148
  (
    n164,
    n68
  );


  not
  g149
  (
    n116,
    n61
  );


  buf
  g150
  (
    n131,
    n68
  );


  not
  g151
  (
    n117,
    n62
  );


  buf
  g152
  (
    n129,
    n66
  );


  buf
  g153
  (
    n163,
    n88
  );


  buf
  g154
  (
    n171,
    n86
  );


  buf
  g155
  (
    n97,
    n74
  );


  not
  g156
  (
    n184,
    n71
  );


  buf
  g157
  (
    n121,
    n62
  );


  not
  g158
  (
    n179,
    n67
  );


  buf
  g159
  (
    n114,
    n78
  );


  not
  g160
  (
    n137,
    n83
  );


  not
  g161
  (
    n178,
    n64
  );


  not
  g162
  (
    n134,
    n60
  );


  buf
  g163
  (
    n157,
    n69
  );


  not
  g164
  (
    n119,
    n82
  );


  not
  g165
  (
    n104,
    n83
  );


  not
  g166
  (
    n168,
    n70
  );


  buf
  g167
  (
    n156,
    n70
  );


  not
  g168
  (
    n203,
    n84
  );


  not
  g169
  (
    n140,
    n73
  );


  not
  g170
  (
    n194,
    n87
  );


  buf
  g171
  (
    n132,
    n76
  );


  not
  g172
  (
    n133,
    n83
  );


  nand
  g173
  (
    n109,
    n80,
    n82,
    n62
  );


  buf
  g174
  (
    n248,
    n182
  );


  buf
  g175
  (
    n285,
    n162
  );


  not
  g176
  (
    n307,
    n160
  );


  buf
  g177
  (
    n211,
    n100
  );


  not
  g178
  (
    n231,
    n158
  );


  buf
  g179
  (
    n215,
    n183
  );


  not
  g180
  (
    n322,
    n152
  );


  buf
  g181
  (
    n247,
    n124
  );


  buf
  g182
  (
    n348,
    n178
  );


  not
  g183
  (
    n359,
    n155
  );


  buf
  g184
  (
    n213,
    n120
  );


  not
  g185
  (
    n281,
    n179
  );


  not
  g186
  (
    n237,
    n151
  );


  buf
  g187
  (
    n309,
    n176
  );


  not
  g188
  (
    n297,
    n185
  );


  not
  g189
  (
    n350,
    n101
  );


  not
  g190
  (
    n391,
    n150
  );


  buf
  g191
  (
    n409,
    n159
  );


  buf
  g192
  (
    n361,
    n180
  );


  buf
  g193
  (
    n216,
    n108
  );


  buf
  g194
  (
    n218,
    n140
  );


  buf
  g195
  (
    n209,
    n181
  );


  buf
  g196
  (
    n384,
    n127
  );


  buf
  g197
  (
    n267,
    n99
  );


  not
  g198
  (
    n400,
    n156
  );


  not
  g199
  (
    n303,
    n138
  );


  buf
  g200
  (
    n355,
    n191
  );


  not
  g201
  (
    n336,
    n171
  );


  not
  g202
  (
    n395,
    n193
  );


  buf
  g203
  (
    n383,
    n170
  );


  not
  g204
  (
    n379,
    n148
  );


  buf
  g205
  (
    n230,
    n119
  );


  buf
  g206
  (
    n214,
    n157
  );


  buf
  g207
  (
    n257,
    n167
  );


  not
  g208
  (
    n408,
    n172
  );


  buf
  g209
  (
    n427,
    n109
  );


  buf
  g210
  (
    n420,
    n110
  );


  buf
  g211
  (
    n325,
    n159
  );


  buf
  g212
  (
    n426,
    n182
  );


  not
  g213
  (
    n329,
    n140
  );


  not
  g214
  (
    n376,
    n145
  );


  buf
  g215
  (
    n212,
    n146
  );


  not
  g216
  (
    n282,
    n174
  );


  not
  g217
  (
    n287,
    n167
  );


  not
  g218
  (
    n269,
    n146
  );


  buf
  g219
  (
    n291,
    n173
  );


  not
  g220
  (
    KeyWire_0_29,
    n100
  );


  not
  g221
  (
    n254,
    n126
  );


  not
  g222
  (
    n260,
    n133
  );


  not
  g223
  (
    n241,
    n187
  );


  not
  g224
  (
    n338,
    n133
  );


  not
  g225
  (
    n378,
    n186
  );


  buf
  g226
  (
    n334,
    n115
  );


  not
  g227
  (
    n380,
    n153
  );


  not
  g228
  (
    n347,
    n134
  );


  not
  g229
  (
    n377,
    n187
  );


  not
  g230
  (
    n403,
    n149
  );


  buf
  g231
  (
    n227,
    n147
  );


  not
  g232
  (
    n299,
    n154
  );


  buf
  g233
  (
    n341,
    n128
  );


  not
  g234
  (
    n394,
    n174
  );


  buf
  g235
  (
    n351,
    n108
  );


  not
  g236
  (
    n327,
    n143
  );


  buf
  g237
  (
    n259,
    n147
  );


  not
  g238
  (
    n245,
    n134
  );


  buf
  g239
  (
    KeyWire_0_10,
    n188
  );


  buf
  g240
  (
    n393,
    n173
  );


  not
  g241
  (
    n273,
    n120
  );


  buf
  g242
  (
    n265,
    n155
  );


  not
  g243
  (
    n272,
    n103
  );


  not
  g244
  (
    n318,
    n135
  );


  buf
  g245
  (
    n210,
    n152
  );


  not
  g246
  (
    n387,
    n177
  );


  not
  g247
  (
    n219,
    n144
  );


  not
  g248
  (
    n279,
    n109
  );


  buf
  g249
  (
    n238,
    n181
  );


  not
  g250
  (
    n239,
    n176
  );


  buf
  g251
  (
    KeyWire_0_12,
    n116
  );


  buf
  g252
  (
    n372,
    n172
  );


  not
  g253
  (
    n366,
    n184
  );


  buf
  g254
  (
    n405,
    n178
  );


  buf
  g255
  (
    n305,
    n121
  );


  not
  g256
  (
    n319,
    n110
  );


  not
  g257
  (
    n345,
    n145
  );


  buf
  g258
  (
    n392,
    n116
  );


  not
  g259
  (
    n386,
    n180
  );


  not
  g260
  (
    n222,
    n144
  );


  not
  g261
  (
    n242,
    n169
  );


  not
  g262
  (
    n417,
    n158
  );


  not
  g263
  (
    n311,
    n148
  );


  not
  g264
  (
    n258,
    n158
  );


  buf
  g265
  (
    n410,
    n136
  );


  not
  g266
  (
    n293,
    n190
  );


  buf
  g267
  (
    n277,
    n160
  );


  buf
  g268
  (
    n407,
    n168
  );


  not
  g269
  (
    n294,
    n132
  );


  buf
  g270
  (
    n292,
    n118
  );


  buf
  g271
  (
    n340,
    n150
  );


  buf
  g272
  (
    n250,
    n124
  );


  buf
  g273
  (
    n360,
    n163
  );


  not
  g274
  (
    n264,
    n157
  );


  buf
  g275
  (
    n317,
    n177
  );


  buf
  g276
  (
    n276,
    n188
  );


  buf
  g277
  (
    n418,
    n104
  );


  buf
  g278
  (
    n304,
    n181
  );


  not
  g279
  (
    n251,
    n143
  );


  buf
  g280
  (
    n308,
    n135
  );


  not
  g281
  (
    n321,
    n149
  );


  not
  g282
  (
    n320,
    n92
  );


  buf
  g283
  (
    n411,
    n126
  );


  buf
  g284
  (
    n406,
    n145
  );


  not
  g285
  (
    n220,
    n159
  );


  not
  g286
  (
    n223,
    n136
  );


  buf
  g287
  (
    n289,
    n143
  );


  not
  g288
  (
    n396,
    n177
  );


  not
  g289
  (
    KeyWire_0_15,
    n167
  );


  buf
  g290
  (
    n208,
    n123
  );


  not
  g291
  (
    n349,
    n185
  );


  not
  g292
  (
    n367,
    n156
  );


  buf
  g293
  (
    n424,
    n136
  );


  not
  g294
  (
    n226,
    n149
  );


  buf
  g295
  (
    n382,
    n114
  );


  buf
  g296
  (
    n255,
    n173
  );


  not
  g297
  (
    n316,
    n178
  );


  buf
  g298
  (
    n261,
    n156
  );


  buf
  g299
  (
    n333,
    n139
  );


  not
  g300
  (
    n271,
    n153
  );


  buf
  g301
  (
    n310,
    n175
  );


  not
  g302
  (
    n404,
    n123
  );


  not
  g303
  (
    n354,
    n180
  );


  not
  g304
  (
    n296,
    n146
  );


  not
  g305
  (
    n425,
    n126
  );


  buf
  g306
  (
    n368,
    n179
  );


  buf
  g307
  (
    n234,
    n169
  );


  buf
  g308
  (
    n381,
    n177
  );


  not
  g309
  (
    n286,
    n150
  );


  buf
  g310
  (
    n399,
    n188
  );


  not
  g311
  (
    n328,
    n182
  );


  buf
  g312
  (
    n335,
    n164
  );


  buf
  g313
  (
    n371,
    n139
  );


  buf
  g314
  (
    n415,
    n131
  );


  buf
  g315
  (
    n295,
    n192
  );


  buf
  g316
  (
    n290,
    n137
  );


  not
  g317
  (
    n362,
    n111
  );


  buf
  g318
  (
    n375,
    n112
  );


  not
  g319
  (
    n306,
    n192
  );


  buf
  g320
  (
    n357,
    n117
  );


  buf
  g321
  (
    n249,
    n122
  );


  buf
  g322
  (
    n365,
    n152
  );


  not
  g323
  (
    n275,
    n175
  );


  not
  g324
  (
    n385,
    n156
  );


  not
  g325
  (
    n419,
    n151
  );


  buf
  g326
  (
    n412,
    n173
  );


  not
  g327
  (
    n314,
    n105
  );


  buf
  g328
  (
    n326,
    n164
  );


  not
  g329
  (
    n313,
    n191
  );


  not
  g330
  (
    n225,
    n141
  );


  buf
  g331
  (
    n401,
    n165
  );


  not
  g332
  (
    n246,
    n117
  );


  not
  g333
  (
    KeyWire_0_11,
    n149
  );


  buf
  g334
  (
    n339,
    n111
  );


  not
  g335
  (
    n302,
    n162
  );


  not
  g336
  (
    n374,
    n183
  );


  buf
  g337
  (
    n278,
    n154
  );


  buf
  g338
  (
    n342,
    n164
  );


  buf
  g339
  (
    KeyWire_0_30,
    n179
  );


  not
  g340
  (
    n244,
    n136
  );


  buf
  g341
  (
    n363,
    n113
  );


  buf
  g342
  (
    n240,
    n181
  );


  not
  g343
  (
    n232,
    n140
  );


  not
  g344
  (
    KeyWire_0_23,
    n122
  );


  buf
  g345
  (
    n332,
    n147
  );


  not
  g346
  (
    n217,
    n98
  );


  buf
  g347
  (
    n343,
    n107
  );


  buf
  g348
  (
    n352,
    n93
  );


  buf
  g349
  (
    n421,
    n165
  );


  not
  g350
  (
    n284,
    n138
  );


  buf
  g351
  (
    n252,
    n125
  );


  buf
  g352
  (
    n270,
    n154
  );


  nand
  g353
  (
    n364,
    n192,
    n159,
    n168,
    n132
  );


  xnor
  g354
  (
    n236,
    n150,
    n168,
    n131,
    n182
  );


  or
  g355
  (
    n283,
    n166,
    n106,
    n127,
    n185
  );


  xnor
  g356
  (
    n414,
    n106,
    n157,
    n130,
    n161
  );


  nor
  g357
  (
    n268,
    n105,
    n148,
    n160,
    n178
  );


  or
  g358
  (
    n373,
    n162,
    n171,
    n174,
    n176
  );


  or
  g359
  (
    n331,
    n110,
    n141,
    n115,
    n184
  );


  or
  g360
  (
    n228,
    n187,
    n101,
    n122,
    n118
  );


  nand
  g361
  (
    n207,
    n186,
    n142,
    n165,
    n144
  );


  or
  g362
  (
    n229,
    n106,
    n101,
    n143,
    n152
  );


  nor
  g363
  (
    n274,
    n114,
    n128,
    n165,
    n112
  );


  nor
  g364
  (
    n324,
    n189,
    n167,
    n184,
    n161
  );


  or
  g365
  (
    n330,
    n164,
    n186,
    n147,
    n137
  );


  nor
  g366
  (
    n280,
    n175,
    n108,
    n160,
    n102
  );


  nor
  g367
  (
    n422,
    n113,
    n112,
    n117,
    n172
  );


  nand
  g368
  (
    n369,
    n138,
    n174,
    n107,
    n103
  );


  nand
  g369
  (
    n288,
    n141,
    n183,
    n134,
    n170
  );


  nor
  g370
  (
    n256,
    n118,
    n135,
    n188,
    n109
  );


  nor
  g371
  (
    n346,
    n134,
    n125,
    n163,
    n138
  );


  or
  g372
  (
    n312,
    n142,
    n161,
    n102,
    n104
  );


  nand
  g373
  (
    n402,
    n158,
    n135,
    n189,
    n113
  );


  xor
  g374
  (
    n353,
    n137,
    n153,
    n116,
    n111
  );


  or
  g375
  (
    n337,
    n121,
    n189,
    n180,
    n94
  );


  xnor
  g376
  (
    n298,
    n168,
    n151,
    n171,
    n120
  );


  nor
  g377
  (
    n397,
    n161,
    n189,
    n104,
    n155
  );


  xnor
  g378
  (
    n388,
    n132,
    n151,
    n170,
    n103
  );


  and
  g379
  (
    n370,
    n169,
    n131,
    n137,
    n146
  );


  or
  g380
  (
    n423,
    n129,
    n130,
    n114,
    n187
  );


  xnor
  g381
  (
    n233,
    n171,
    n183,
    n125,
    n96
  );


  nand
  g382
  (
    n224,
    n157,
    n141,
    n124,
    n123
  );


  or
  g383
  (
    n262,
    n121,
    n184,
    n163,
    n129
  );


  xor
  g384
  (
    n356,
    n133,
    n142,
    n176,
    n166
  );


  or
  g385
  (
    n300,
    n119,
    n142,
    n127,
    n163
  );


  and
  g386
  (
    n221,
    n186,
    n155,
    n153,
    n119
  );


  nand
  g387
  (
    n315,
    n140,
    n133,
    n128,
    n190
  );


  xor
  g388
  (
    n390,
    n139,
    n192,
    n170,
    n144
  );


  xor
  g389
  (
    n358,
    n105,
    n169,
    n166,
    n102
  );


  and
  g390
  (
    n413,
    n166,
    n97,
    n154,
    n115
  );


  xnor
  g391
  (
    n253,
    n190,
    n130,
    n129,
    n145
  );


  nand
  g392
  (
    n263,
    n162,
    n139,
    n175,
    n191
  );


  nand
  g393
  (
    n398,
    n185,
    n148,
    n107,
    n179
  );


  nor
  g394
  (
    n416,
    n191,
    n95,
    n172,
    n190
  );


  not
  g395
  (
    KeyWire_0_5,
    n13
  );


  not
  g396
  (
    n510,
    n270
  );


  not
  g397
  (
    n432,
    n266
  );


  buf
  g398
  (
    n440,
    n274
  );


  not
  g399
  (
    n489,
    n277
  );


  not
  g400
  (
    n438,
    n287
  );


  buf
  g401
  (
    n443,
    n349
  );


  buf
  g402
  (
    n467,
    n250
  );


  not
  g403
  (
    n504,
    n340
  );


  buf
  g404
  (
    n484,
    n344
  );


  not
  g405
  (
    n458,
    n303
  );


  buf
  g406
  (
    n495,
    n254
  );


  not
  g407
  (
    n450,
    n285
  );


  not
  g408
  (
    n511,
    n350
  );


  buf
  g409
  (
    n490,
    n331
  );


  buf
  g410
  (
    n501,
    n233
  );


  not
  g411
  (
    n508,
    n263
  );


  buf
  g412
  (
    n524,
    n242
  );


  not
  g413
  (
    n428,
    n221
  );


  not
  g414
  (
    n519,
    n10
  );


  buf
  g415
  (
    n499,
    n231
  );


  buf
  g416
  (
    n478,
    n302
  );


  buf
  g417
  (
    n472,
    n304
  );


  buf
  g418
  (
    n480,
    n280
  );


  buf
  g419
  (
    n464,
    n260
  );


  buf
  g420
  (
    n470,
    n333
  );


  not
  g421
  (
    n498,
    n11
  );


  buf
  g422
  (
    n515,
    n246
  );


  not
  g423
  (
    n505,
    n307
  );


  not
  g424
  (
    n460,
    n44
  );


  not
  g425
  (
    n500,
    n352
  );


  not
  g426
  (
    n463,
    n306
  );


  buf
  g427
  (
    n456,
    n332
  );


  not
  g428
  (
    KeyWire_0_1,
    n343
  );


  not
  g429
  (
    n468,
    n251
  );


  buf
  g430
  (
    n448,
    n318
  );


  buf
  g431
  (
    n477,
    n224
  );


  buf
  g432
  (
    n449,
    n334
  );


  buf
  g433
  (
    n494,
    n244
  );


  buf
  g434
  (
    n469,
    n346
  );


  not
  g435
  (
    n466,
    n9
  );


  not
  g436
  (
    n527,
    n12
  );


  not
  g437
  (
    n444,
    n226
  );


  not
  g438
  (
    n506,
    n223
  );


  buf
  g439
  (
    n526,
    n267
  );


  not
  g440
  (
    n513,
    n220
  );


  not
  g441
  (
    n461,
    n294
  );


  buf
  g442
  (
    n485,
    n290
  );


  buf
  g443
  (
    n521,
    n8
  );


  buf
  g444
  (
    n471,
    n241
  );


  not
  g445
  (
    n514,
    n243
  );


  buf
  g446
  (
    n433,
    n12
  );


  buf
  g447
  (
    n525,
    n269
  );


  buf
  g448
  (
    n509,
    n299
  );


  not
  g449
  (
    n447,
    n315
  );


  buf
  g450
  (
    n497,
    n10
  );


  buf
  g451
  (
    n429,
    n300
  );


  buf
  g452
  (
    n487,
    n292
  );


  buf
  g453
  (
    n441,
    n248
  );


  buf
  g454
  (
    n491,
    n298
  );


  buf
  g455
  (
    n507,
    n222
  );


  not
  g456
  (
    n522,
    n335
  );


  not
  g457
  (
    n481,
    n308
  );


  not
  g458
  (
    n516,
    n13
  );


  buf
  g459
  (
    n518,
    n234
  );


  buf
  g460
  (
    n431,
    n289
  );


  not
  g461
  (
    n517,
    n193
  );


  buf
  g462
  (
    n473,
    n230
  );


  buf
  g463
  (
    n486,
    n261
  );


  buf
  g464
  (
    n454,
    n229
  );


  not
  g465
  (
    n520,
    n239
  );


  buf
  g466
  (
    n493,
    n211
  );


  buf
  g467
  (
    n452,
    n253
  );


  buf
  g468
  (
    n512,
    n272
  );


  not
  g469
  (
    n459,
    n245
  );


  not
  g470
  (
    n483,
    n193
  );


  and
  g471
  (
    n475,
    n323,
    n219
  );


  nor
  g472
  (
    n502,
    n227,
    n193,
    n12
  );


  nor
  g473
  (
    n476,
    n11,
    n8,
    n311,
    n218
  );


  nand
  g474
  (
    n482,
    n295,
    n271,
    n296,
    n9
  );


  xnor
  g475
  (
    n451,
    n207,
    n264,
    n273,
    n310
  );


  nor
  g476
  (
    n453,
    n324,
    n9,
    n212,
    n314
  );


  xor
  g477
  (
    n455,
    n237,
    n240,
    n325,
    n208
  );


  and
  g478
  (
    n465,
    n336,
    n347,
    n13,
    n348
  );


  or
  g479
  (
    n523,
    n339,
    n328,
    n213,
    n238
  );


  xor
  g480
  (
    n492,
    n209,
    n252,
    n278,
    n9
  );


  and
  g481
  (
    n457,
    n284,
    n301,
    n293,
    n309
  );


  or
  g482
  (
    n474,
    n281,
    n255,
    n312,
    n279
  );


  nor
  g483
  (
    n496,
    n341,
    n286,
    n258,
    n235
  );


  nor
  g484
  (
    n430,
    n338,
    n317,
    n11,
    n288
  );


  nand
  g485
  (
    n479,
    n11,
    n313,
    n216,
    n321
  );


  or
  g486
  (
    n445,
    n329,
    n215,
    n8,
    n228
  );


  and
  g487
  (
    n442,
    n283,
    n249,
    n10,
    n282
  );


  xor
  g488
  (
    n434,
    n342,
    n275,
    n268,
    n316
  );


  xor
  g489
  (
    n439,
    n259,
    n214,
    n326,
    n330
  );


  xor
  g490
  (
    n437,
    n327,
    n210,
    n13,
    n305
  );


  nand
  g491
  (
    n446,
    n247,
    n297,
    n232,
    n8
  );


  xor
  g492
  (
    n436,
    n225,
    n217,
    n256,
    n345
  );


  and
  g493
  (
    KeyWire_0_8,
    n257,
    n351,
    n291,
    n236
  );


  xnor
  g494
  (
    n435,
    n322,
    n337,
    n276,
    n10
  );


  nor
  g495
  (
    n488,
    n265,
    n319,
    n320,
    n262
  );


  buf
  g496
  (
    n577,
    n14
  );


  not
  g497
  (
    n552,
    n19
  );


  not
  g498
  (
    n571,
    n31
  );


  not
  g499
  (
    n546,
    n459
  );


  not
  g500
  (
    n548,
    n475
  );


  buf
  g501
  (
    n567,
    n31
  );


  not
  g502
  (
    n535,
    n456
  );


  not
  g503
  (
    n556,
    n24
  );


  not
  g504
  (
    n543,
    n29
  );


  not
  g505
  (
    n561,
    n23
  );


  buf
  g506
  (
    n550,
    n466
  );


  not
  g507
  (
    n570,
    n17
  );


  xor
  g508
  (
    n547,
    n18,
    n21,
    n446
  );


  nor
  g509
  (
    n557,
    n469,
    n16,
    n22
  );


  or
  g510
  (
    n559,
    n24,
    n471,
    n432
  );


  nor
  g511
  (
    n562,
    n26,
    n15,
    n439
  );


  nor
  g512
  (
    n538,
    n23,
    n443,
    n452
  );


  xnor
  g513
  (
    n566,
    n430,
    n473,
    n436
  );


  or
  g514
  (
    n531,
    n20,
    n32,
    n435
  );


  xor
  g515
  (
    n564,
    n431,
    n460,
    n18
  );


  and
  g516
  (
    n553,
    n462,
    n19,
    n470
  );


  xnor
  g517
  (
    n569,
    n26,
    n20,
    n434
  );


  xor
  g518
  (
    n534,
    n450,
    n440,
    n18
  );


  or
  g519
  (
    n555,
    n31,
    n477,
    n448
  );


  and
  g520
  (
    n542,
    n476,
    n25,
    n18
  );


  xor
  g521
  (
    n530,
    n428,
    n27,
    n447
  );


  and
  g522
  (
    n536,
    n15,
    n463,
    n474
  );


  nor
  g523
  (
    n549,
    n19,
    n453,
    n30
  );


  xnor
  g524
  (
    n554,
    n16,
    n21,
    n27
  );


  nand
  g525
  (
    n545,
    n17,
    n472,
    n465
  );


  nor
  g526
  (
    n563,
    n457,
    n445,
    n22
  );


  xnor
  g527
  (
    n551,
    n30,
    n24
  );


  nand
  g528
  (
    n532,
    n429,
    n17,
    n21
  );


  nand
  g529
  (
    n533,
    n449,
    n21,
    n29
  );


  nor
  g530
  (
    n537,
    n29,
    n28,
    n19
  );


  and
  g531
  (
    n529,
    n14,
    n451,
    n28
  );


  and
  g532
  (
    n574,
    n26,
    n454,
    n32
  );


  xor
  g533
  (
    n560,
    n23,
    n437,
    n30
  );


  xnor
  g534
  (
    n541,
    n15,
    n455,
    n20
  );


  xnor
  g535
  (
    n565,
    n31,
    n26,
    n458
  );


  xnor
  g536
  (
    n544,
    n15,
    n16
  );


  xnor
  g537
  (
    n572,
    n433,
    n28,
    n22
  );


  or
  g538
  (
    n540,
    n27,
    n25
  );


  nand
  g539
  (
    n575,
    n461,
    n28,
    n464
  );


  nor
  g540
  (
    n578,
    n30,
    n20,
    n14
  );


  xor
  g541
  (
    n576,
    n441,
    n442,
    n467
  );


  xor
  g542
  (
    n568,
    n32,
    n25,
    n23
  );


  nand
  g543
  (
    n573,
    n14,
    n17,
    n22
  );


  xor
  g544
  (
    n558,
    n27,
    n32,
    n444
  );


  and
  g545
  (
    n539,
    n438,
    n468,
    n29
  );


  buf
  g546
  (
    n596,
    n534
  );


  not
  g547
  (
    n597,
    n529
  );


  not
  g548
  (
    n595,
    n535
  );


  not
  g549
  (
    n587,
    n534
  );


  buf
  g550
  (
    n586,
    n534
  );


  not
  g551
  (
    n588,
    n535
  );


  not
  g552
  (
    n581,
    n529
  );


  buf
  g553
  (
    n584,
    n46
  );


  not
  g554
  (
    n580,
    n533
  );


  not
  g555
  (
    n590,
    n536
  );


  buf
  g556
  (
    n601,
    n530
  );


  buf
  g557
  (
    n605,
    n532
  );


  buf
  g558
  (
    n599,
    n532
  );


  buf
  g559
  (
    n592,
    n529
  );


  not
  g560
  (
    n604,
    n531
  );


  not
  g561
  (
    n582,
    n534
  );


  buf
  g562
  (
    n591,
    n536
  );


  not
  g563
  (
    n602,
    n533
  );


  buf
  g564
  (
    n603,
    n535
  );


  not
  g565
  (
    n598,
    n45
  );


  not
  g566
  (
    n585,
    n530
  );


  buf
  g567
  (
    n594,
    n531
  );


  buf
  g568
  (
    n579,
    n45
  );


  not
  g569
  (
    n593,
    n45
  );


  and
  g570
  (
    n589,
    n532,
    n530
  );


  or
  g571
  (
    KeyWire_0_24,
    n531,
    n533,
    n535
  );


  and
  g572
  (
    n583,
    n45,
    n532,
    n533
  );


  xnor
  g573
  (
    KeyWire_0_9,
    n46,
    n53
  );


  and
  g574
  (
    n606,
    n51,
    n50,
    n52
  );


  and
  g575
  (
    n610,
    n598,
    n49,
    n593,
    n91
  );


  and
  g576
  (
    n613,
    n47,
    n590,
    n90,
    n46
  );


  xor
  g577
  (
    n615,
    n49,
    n51,
    n602,
    n48
  );


  or
  g578
  (
    n618,
    n50,
    n592,
    n48
  );


  xor
  g579
  (
    n612,
    n90,
    n591,
    n52,
    n91
  );


  nor
  g580
  (
    n614,
    n89,
    n89,
    n91,
    n49
  );


  nor
  g581
  (
    n616,
    n603,
    n604,
    n47,
    n50
  );


  xor
  g582
  (
    n607,
    n595,
    n53,
    n49,
    n89
  );


  nand
  g583
  (
    n611,
    n47,
    n48,
    n51,
    n90
  );


  or
  g584
  (
    n608,
    n89,
    n47,
    n52,
    n597
  );


  nand
  g585
  (
    n617,
    n91,
    n594,
    n53,
    n601
  );


  nor
  g586
  (
    n620,
    n599,
    n46,
    n51,
    n596
  );


  nand
  g587
  (
    n619,
    n90,
    n52,
    n600,
    n88
  );


  and
  g588
  (
    n627,
    n609,
    n198
  );


  xor
  g589
  (
    n628,
    n194,
    n196,
    n201
  );


  nand
  g590
  (
    n635,
    n616,
    n199,
    n194
  );


  or
  g591
  (
    n632,
    n197,
    n196,
    n608
  );


  xnor
  g592
  (
    n636,
    n197,
    n200
  );


  and
  g593
  (
    n622,
    n195,
    n201,
    n619
  );


  and
  g594
  (
    n623,
    n198,
    n197,
    n195
  );


  xnor
  g595
  (
    n626,
    n201,
    n199,
    n613
  );


  xor
  g596
  (
    n625,
    n195,
    n615,
    n196
  );


  xor
  g597
  (
    n629,
    n620,
    n610,
    n607
  );


  xnor
  g598
  (
    n633,
    n202,
    n200,
    n194
  );


  xor
  g599
  (
    n631,
    n195,
    n614,
    n200
  );


  nand
  g600
  (
    n621,
    n606,
    n199
  );


  or
  g601
  (
    n624,
    n197,
    n611,
    n194
  );


  and
  g602
  (
    n630,
    n620,
    n618,
    n196,
    n612
  );


  xnor
  g603
  (
    n634,
    n617,
    n201,
    n202,
    n198
  );


  buf
  g604
  (
    n660,
    n381
  );


  not
  g605
  (
    n641,
    n365
  );


  not
  g606
  (
    n639,
    n54
  );


  buf
  g607
  (
    n638,
    n56
  );


  buf
  g608
  (
    n644,
    n58
  );


  nor
  g609
  (
    n661,
    n625,
    n357,
    n622
  );


  xor
  g610
  (
    n643,
    n373,
    n424,
    n624,
    n426
  );


  xnor
  g611
  (
    n647,
    n398,
    n627,
    n391,
    n425
  );


  and
  g612
  (
    n665,
    n405,
    n406,
    n366,
    n58
  );


  xnor
  g613
  (
    n658,
    n383,
    n630,
    n625,
    n629
  );


  or
  g614
  (
    n663,
    n392,
    n394,
    n390,
    n55
  );


  or
  g615
  (
    n669,
    n629,
    n413,
    n627,
    n389
  );


  xnor
  g616
  (
    n668,
    n625,
    n418,
    n54,
    n417
  );


  xnor
  g617
  (
    KeyWire_0_13,
    n393,
    n403,
    n53,
    n625
  );


  nor
  g618
  (
    n666,
    n415,
    n362,
    n627,
    n621
  );


  and
  g619
  (
    n653,
    n380,
    n423,
    n626,
    n421
  );


  nor
  g620
  (
    n648,
    n623,
    n414,
    n408,
    n374
  );


  xnor
  g621
  (
    n642,
    n57,
    n400,
    n621,
    n626
  );


  xnor
  g622
  (
    n673,
    n623,
    n376,
    n626,
    n427
  );


  xor
  g623
  (
    n671,
    n55,
    n56,
    n364,
    n399
  );


  nand
  g624
  (
    n672,
    n355,
    n56,
    n371,
    n358
  );


  xor
  g625
  (
    n651,
    n382,
    n57,
    n626
  );


  nor
  g626
  (
    n655,
    n623,
    n412,
    n353,
    n370
  );


  nor
  g627
  (
    n646,
    n377,
    n54,
    n387
  );


  xnor
  g628
  (
    n645,
    n57,
    n629,
    n404
  );


  xnor
  g629
  (
    n670,
    n628,
    n56,
    n622,
    n372
  );


  xor
  g630
  (
    n652,
    n422,
    n369,
    n419,
    n388
  );


  and
  g631
  (
    KeyWire_0_25,
    n411,
    n354,
    n386,
    n622
  );


  and
  g632
  (
    n640,
    n409,
    n624,
    n410,
    n630
  );


  xor
  g633
  (
    n662,
    n375,
    n395,
    n628,
    n396
  );


  nand
  g634
  (
    n637,
    n623,
    n397,
    n624,
    n361
  );


  xor
  g635
  (
    n656,
    n628,
    n385,
    n55,
    n621
  );


  nand
  g636
  (
    n667,
    n401,
    n624,
    n420,
    n407
  );


  nor
  g637
  (
    n654,
    n363,
    n360,
    n378,
    n58
  );


  xnor
  g638
  (
    n650,
    n416,
    n359,
    n368,
    n628
  );


  nand
  g639
  (
    n664,
    n55,
    n384,
    n367,
    n622
  );


  xor
  g640
  (
    n657,
    n356,
    n627,
    n379,
    n402
  );


  nor
  g641
  (
    n674,
    n483,
    n672,
    n513,
    n59
  );


  xor
  g642
  (
    n688,
    n662,
    n666,
    n518,
    n481
  );


  or
  g643
  (
    n683,
    n512,
    n491,
    n649,
    n669
  );


  nand
  g644
  (
    n681,
    n654,
    n523,
    n526,
    n643
  );


  xnor
  g645
  (
    n675,
    n668,
    n652,
    n525,
    n659
  );


  xnor
  g646
  (
    n692,
    n669,
    n59,
    n668,
    n653
  );


  xnor
  g647
  (
    n696,
    n519,
    n670,
    n58,
    n486
  );


  and
  g648
  (
    n694,
    n663,
    n639,
    n664,
    n527
  );


  and
  g649
  (
    n701,
    n59,
    n638,
    n480,
    n662
  );


  xnor
  g650
  (
    n695,
    n660,
    n637,
    n500,
    n504
  );


  nor
  g651
  (
    n685,
    n511,
    n655,
    n494,
    n507
  );


  xnor
  g652
  (
    n687,
    n672,
    n654,
    n665,
    n650
  );


  xor
  g653
  (
    n689,
    n671,
    n658,
    n515,
    n495
  );


  and
  g654
  (
    n697,
    n671,
    n478,
    n508,
    n59
  );


  xnor
  g655
  (
    n698,
    n487,
    n484,
    n498,
    n652
  );


  nand
  g656
  (
    n678,
    n647,
    n490,
    n653,
    n488
  );


  xor
  g657
  (
    n682,
    n482,
    n516,
    n501,
    n502
  );


  or
  g658
  (
    n699,
    n665,
    n645,
    n499,
    n505
  );


  and
  g659
  (
    n679,
    n664,
    n521,
    n661,
    n479
  );


  xnor
  g660
  (
    n680,
    n655,
    n640,
    n509,
    n517
  );


  nor
  g661
  (
    n686,
    n666,
    n524,
    n661,
    n489
  );


  or
  g662
  (
    n690,
    n503,
    n485,
    n656,
    n659
  );


  nand
  g663
  (
    n677,
    n642,
    n651,
    n522,
    n658
  );


  xnor
  g664
  (
    n676,
    n644,
    n497,
    n496,
    n667
  );


  nor
  g665
  (
    n693,
    n673,
    n646,
    n510,
    n506
  );


  xnor
  g666
  (
    KeyWire_0_0,
    n493,
    n514,
    n660,
    n657
  );


  xnor
  g667
  (
    n691,
    n648,
    n673,
    n520,
    n656
  );


  nand
  g668
  (
    n702,
    n670,
    n663,
    n528,
    n667
  );


  nand
  g669
  (
    n684,
    n657,
    n492,
    n641,
    n651
  );


  buf
  g670
  (
    n766,
    n685
  );


  not
  g671
  (
    n717,
    n696
  );


  buf
  g672
  (
    n761,
    n680
  );


  buf
  g673
  (
    n741,
    n678
  );


  not
  g674
  (
    n794,
    n694
  );


  not
  g675
  (
    n723,
    n674
  );


  not
  g676
  (
    n810,
    n698
  );


  buf
  g677
  (
    n729,
    n681
  );


  buf
  g678
  (
    n769,
    n674
  );


  not
  g679
  (
    n798,
    n691
  );


  buf
  g680
  (
    n796,
    n682
  );


  not
  g681
  (
    n774,
    n686
  );


  not
  g682
  (
    n773,
    n690
  );


  buf
  g683
  (
    n726,
    n697
  );


  buf
  g684
  (
    n714,
    n687
  );


  buf
  g685
  (
    n763,
    n677
  );


  not
  g686
  (
    n768,
    n675
  );


  not
  g687
  (
    n805,
    n691
  );


  not
  g688
  (
    n720,
    n698
  );


  not
  g689
  (
    KeyWire_0_17,
    n680
  );


  not
  g690
  (
    n713,
    n684
  );


  buf
  g691
  (
    n781,
    n674
  );


  buf
  g692
  (
    n748,
    n695
  );


  not
  g693
  (
    n733,
    n692
  );


  buf
  g694
  (
    n750,
    n683
  );


  buf
  g695
  (
    KeyWire_0_27,
    n683
  );


  not
  g696
  (
    n737,
    n696
  );


  not
  g697
  (
    n724,
    n686
  );


  buf
  g698
  (
    KeyWire_0_14,
    n676
  );


  not
  g699
  (
    n706,
    n681
  );


  buf
  g700
  (
    n749,
    n682
  );


  buf
  g701
  (
    n765,
    n694
  );


  buf
  g702
  (
    n747,
    n686
  );


  buf
  g703
  (
    n716,
    n698
  );


  not
  g704
  (
    n771,
    n691
  );


  not
  g705
  (
    n705,
    n693
  );


  buf
  g706
  (
    n734,
    n681
  );


  buf
  g707
  (
    KeyWire_0_28,
    n700
  );


  buf
  g708
  (
    n806,
    n699
  );


  buf
  g709
  (
    n753,
    n690
  );


  buf
  g710
  (
    n809,
    n675
  );


  not
  g711
  (
    n772,
    n679
  );


  not
  g712
  (
    n715,
    n676
  );


  buf
  g713
  (
    n784,
    n682
  );


  buf
  g714
  (
    n745,
    n678
  );


  buf
  g715
  (
    KeyWire_0_3,
    n689
  );


  not
  g716
  (
    n703,
    n700
  );


  not
  g717
  (
    n791,
    n676
  );


  not
  g718
  (
    n709,
    n696
  );


  not
  g719
  (
    n792,
    n685
  );


  buf
  g720
  (
    n719,
    n700
  );


  not
  g721
  (
    n802,
    n679
  );


  not
  g722
  (
    n731,
    n680
  );


  not
  g723
  (
    n752,
    n677
  );


  buf
  g724
  (
    KeyWire_0_31,
    n677
  );


  buf
  g725
  (
    n808,
    n675
  );


  buf
  g726
  (
    n762,
    n682
  );


  buf
  g727
  (
    n718,
    n687
  );


  not
  g728
  (
    n758,
    n692
  );


  not
  g729
  (
    n740,
    n692
  );


  buf
  g730
  (
    n770,
    n687
  );


  buf
  g731
  (
    n760,
    n685
  );


  not
  g732
  (
    n776,
    n695
  );


  buf
  g733
  (
    n754,
    n684
  );


  buf
  g734
  (
    n803,
    n678
  );


  buf
  g735
  (
    n795,
    n700
  );


  buf
  g736
  (
    n712,
    n681
  );


  not
  g737
  (
    n744,
    n694
  );


  not
  g738
  (
    n783,
    n699
  );


  not
  g739
  (
    n725,
    n675
  );


  not
  g740
  (
    n778,
    n687
  );


  buf
  g741
  (
    n730,
    n699
  );


  buf
  g742
  (
    n777,
    n695
  );


  not
  g743
  (
    n767,
    n689
  );


  buf
  g744
  (
    n797,
    n691
  );


  not
  g745
  (
    n735,
    n693
  );


  buf
  g746
  (
    n782,
    n697
  );


  not
  g747
  (
    n751,
    n686
  );


  not
  g748
  (
    n722,
    n698
  );


  not
  g749
  (
    n728,
    n680
  );


  buf
  g750
  (
    n790,
    n694
  );


  buf
  g751
  (
    n727,
    n695
  );


  not
  g752
  (
    n756,
    n697
  );


  not
  g753
  (
    n787,
    n676
  );


  not
  g754
  (
    n764,
    n690
  );


  buf
  g755
  (
    n736,
    n693
  );


  not
  g756
  (
    n707,
    n679
  );


  buf
  g757
  (
    n708,
    n683
  );


  buf
  g758
  (
    n721,
    n689
  );


  not
  g759
  (
    n710,
    n679
  );


  buf
  g760
  (
    n757,
    n677
  );


  not
  g761
  (
    n799,
    n684
  );


  buf
  g762
  (
    n779,
    n690
  );


  buf
  g763
  (
    n800,
    n697
  );


  not
  g764
  (
    KeyWire_0_19,
    n692
  );


  buf
  g765
  (
    n793,
    n674
  );


  not
  g766
  (
    n742,
    n688
  );


  buf
  g767
  (
    n732,
    n688
  );


  not
  g768
  (
    n788,
    n678
  );


  buf
  g769
  (
    n746,
    n688
  );


  not
  g770
  (
    n780,
    n683
  );


  buf
  g771
  (
    n804,
    n696
  );


  not
  g772
  (
    n739,
    n685
  );


  buf
  g773
  (
    n755,
    n689
  );


  buf
  g774
  (
    n738,
    n699
  );


  buf
  g775
  (
    n785,
    n688
  );


  not
  g776
  (
    n775,
    n684
  );


  buf
  g777
  (
    n786,
    n693
  );


  nand
  g778
  (
    n926,
    n794,
    n761,
    n759
  );


  and
  g779
  (
    n930,
    n708,
    n578,
    n569
  );


  nand
  g780
  (
    n901,
    n709,
    n555,
    n553
  );


  nand
  g781
  (
    n843,
    n722,
    n204,
    n802
  );


  and
  g782
  (
    n871,
    n569,
    n778,
    n564
  );


  nor
  g783
  (
    n878,
    n551,
    n806,
    n750
  );


  and
  g784
  (
    n842,
    n787,
    n739,
    n723
  );


  xnor
  g785
  (
    n956,
    n784,
    n546,
    n705
  );


  xor
  g786
  (
    KeyWire_0_20,
    n564,
    n559,
    n561
  );


  or
  g787
  (
    n826,
    n753,
    n740,
    n754
  );


  nor
  g788
  (
    n834,
    n704,
    n743,
    n776
  );


  xor
  g789
  (
    n873,
    n537,
    n764,
    n710
  );


  nand
  g790
  (
    n865,
    n555,
    n701,
    n745
  );


  nor
  g791
  (
    n909,
    n777,
    n726,
    n779
  );


  xor
  g792
  (
    n933,
    n543,
    n783,
    n605
  );


  xor
  g793
  (
    n898,
    n718,
    n805,
    n804
  );


  nor
  g794
  (
    n812,
    n780,
    n722,
    n782
  );


  or
  g795
  (
    n846,
    n765,
    n543,
    n548
  );


  xor
  g796
  (
    n876,
    n575,
    n771,
    n547
  );


  xnor
  g797
  (
    n914,
    n576,
    n731,
    n577
  );


  or
  g798
  (
    n932,
    n742,
    n807,
    n574
  );


  nor
  g799
  (
    n913,
    n547,
    n205,
    n566
  );


  nand
  g800
  (
    n897,
    n785,
    n738,
    n792
  );


  xnor
  g801
  (
    n820,
    n770,
    n789,
    n753
  );


  nand
  g802
  (
    n858,
    n729,
    n706,
    n578
  );


  nand
  g803
  (
    n825,
    n776,
    n728,
    n205
  );


  and
  g804
  (
    n867,
    n554,
    n794,
    n727
  );


  xor
  g805
  (
    n823,
    n545,
    n784,
    n577
  );


  or
  g806
  (
    n813,
    n557,
    n767,
    n788
  );


  nand
  g807
  (
    n963,
    n769,
    n741,
    n783
  );


  nor
  g808
  (
    n855,
    n707,
    n801,
    n550
  );


  xnor
  g809
  (
    n817,
    n791,
    n551,
    n720
  );


  xor
  g810
  (
    n881,
    n749,
    n540,
    n559
  );


  nor
  g811
  (
    n877,
    n547,
    n563,
    n559
  );


  xnor
  g812
  (
    n952,
    n745,
    n727,
    n787
  );


  and
  g813
  (
    n936,
    n704,
    n770,
    n572
  );


  nor
  g814
  (
    n973,
    n567,
    n804,
    n756
  );


  xnor
  g815
  (
    n951,
    n714,
    n809,
    n724
  );


  nor
  g816
  (
    n905,
    n204,
    n559,
    n568
  );


  xor
  g817
  (
    n864,
    n551,
    n544,
    n761
  );


  xnor
  g818
  (
    n838,
    n544,
    n806,
    n549
  );


  and
  g819
  (
    n893,
    n766,
    n740,
    n571
  );


  nand
  g820
  (
    n844,
    n550,
    n726,
    n740
  );


  nor
  g821
  (
    n852,
    n563,
    n805,
    n742
  );


  nor
  g822
  (
    n859,
    n721,
    n567,
    n800
  );


  nand
  g823
  (
    n957,
    n767,
    n736,
    n798
  );


  nand
  g824
  (
    n971,
    n759,
    n727,
    n541
  );


  xor
  g825
  (
    n872,
    n541,
    n786,
    n778
  );


  nand
  g826
  (
    n961,
    n725,
    n711,
    n784
  );


  xnor
  g827
  (
    n960,
    n722,
    n763,
    n536
  );


  xor
  g828
  (
    n937,
    n745,
    n577,
    n756
  );


  xor
  g829
  (
    n887,
    n786,
    n792,
    n735
  );


  xor
  g830
  (
    n839,
    n786,
    n555,
    n709
  );


  xor
  g831
  (
    n869,
    n763,
    n565,
    n749
  );


  nor
  g832
  (
    n943,
    n747,
    n546,
    n202
  );


  nand
  g833
  (
    n964,
    n752,
    n554,
    n725
  );


  xnor
  g834
  (
    n962,
    n573,
    n772,
    n769
  );


  nand
  g835
  (
    n811,
    n772,
    n574,
    n810
  );


  or
  g836
  (
    n860,
    n539,
    n557,
    n711
  );


  and
  g837
  (
    n922,
    n737,
    n736,
    n728
  );


  and
  g838
  (
    n832,
    n574,
    n773,
    n565
  );


  and
  g839
  (
    n885,
    n569,
    n576,
    n571
  );


  and
  g840
  (
    n892,
    n558,
    n575,
    n710
  );


  nor
  g841
  (
    n924,
    n780,
    n801,
    n556
  );


  nor
  g842
  (
    n907,
    n567,
    n765,
    n560
  );


  nand
  g843
  (
    n947,
    n751,
    n717,
    n733
  );


  xor
  g844
  (
    n889,
    n781,
    n793,
    n575
  );


  xor
  g845
  (
    n840,
    n755,
    n540,
    n720
  );


  and
  g846
  (
    n875,
    n542,
    n545,
    n802
  );


  xor
  g847
  (
    n849,
    n541,
    n539,
    n548
  );


  or
  g848
  (
    n950,
    n805,
    n576,
    n809
  );


  xor
  g849
  (
    n828,
    n798,
    n748,
    n715
  );


  and
  g850
  (
    n814,
    n721,
    n747,
    n703
  );


  xnor
  g851
  (
    n853,
    n552,
    n716,
    n558
  );


  or
  g852
  (
    n856,
    n204,
    n541,
    n571
  );


  or
  g853
  (
    n967,
    n789,
    n800,
    n741
  );


  nand
  g854
  (
    n906,
    n542,
    n751,
    n701
  );


  nand
  g855
  (
    n946,
    n765,
    n744,
    n734
  );


  and
  g856
  (
    n866,
    n538,
    n782,
    n557
  );


  nand
  g857
  (
    n847,
    n566,
    n561,
    n558
  );


  xor
  g858
  (
    n845,
    n773,
    n573,
    n542
  );


  or
  g859
  (
    n827,
    n746,
    n719,
    n712
  );


  and
  g860
  (
    n925,
    n570,
    n734,
    n790
  );


  xor
  g861
  (
    n970,
    n787,
    n789,
    n552
  );


  xnor
  g862
  (
    n819,
    n803,
    n556,
    n545
  );


  nand
  g863
  (
    n919,
    n567,
    n205,
    n546
  );


  xor
  g864
  (
    n942,
    n795,
    n799,
    n730
  );


  xor
  g865
  (
    n861,
    n205,
    n762,
    n757
  );


  nor
  g866
  (
    n923,
    n744,
    n768,
    n562
  );


  and
  g867
  (
    n822,
    n552,
    n569,
    n565
  );


  xor
  g868
  (
    n831,
    n573,
    n578,
    n719
  );


  or
  g869
  (
    n958,
    n777,
    n737,
    n756
  );


  xor
  g870
  (
    n833,
    n775,
    n571,
    n785
  );


  and
  g871
  (
    n848,
    n780,
    n701,
    n538
  );


  xnor
  g872
  (
    n880,
    n755,
    n796,
    n773
  );


  xor
  g873
  (
    n910,
    n714,
    n560,
    n538
  );


  xnor
  g874
  (
    n954,
    n796,
    n563,
    n770
  );


  and
  g875
  (
    n928,
    n752,
    n575,
    n726
  );


  nor
  g876
  (
    n816,
    n790,
    n743,
    n750
  );


  or
  g877
  (
    n841,
    n809,
    n748,
    n540
  );


  nor
  g878
  (
    n931,
    n545,
    n753,
    n720
  );


  and
  g879
  (
    n915,
    n702,
    n810,
    n570
  );


  xnor
  g880
  (
    n948,
    n739,
    n554,
    n731
  );


  or
  g881
  (
    n938,
    n762,
    n754,
    n721
  );


  xor
  g882
  (
    n916,
    n563,
    n803,
    n783
  );


  nor
  g883
  (
    n953,
    n793,
    n556,
    n735
  );


  and
  g884
  (
    n870,
    n548,
    n807,
    n778
  );


  and
  g885
  (
    KeyWire_0_22,
    n543,
    n707,
    n768
  );


  and
  g886
  (
    n851,
    n747,
    n754,
    n748
  );


  xnor
  g887
  (
    n955,
    n764,
    n774,
    n750
  );


  or
  g888
  (
    n900,
    n738,
    n549,
    n795
  );


  and
  g889
  (
    n911,
    n576,
    n801,
    n731
  );


  xnor
  g890
  (
    n836,
    n807,
    n775,
    n718
  );


  xnor
  g891
  (
    n959,
    n724,
    n788,
    n562
  );


  nand
  g892
  (
    n934,
    n539,
    n702,
    n566
  );


  xor
  g893
  (
    n927,
    n774,
    n782,
    n204
  );


  nand
  g894
  (
    n857,
    n570,
    n565,
    n806
  );


  xnor
  g895
  (
    n835,
    n732,
    n556,
    n203
  );


  xnor
  g896
  (
    n908,
    n794,
    n553,
    n549
  );


  and
  g897
  (
    n884,
    n749,
    n791,
    n568
  );


  xor
  g898
  (
    n968,
    n759,
    n561,
    n560
  );


  or
  g899
  (
    n904,
    n746,
    n752,
    n539
  );


  nand
  g900
  (
    n821,
    n572,
    n554,
    n758
  );


  and
  g901
  (
    n972,
    n555,
    n203,
    n547
  );


  xnor
  g902
  (
    n912,
    n732,
    n562,
    n779
  );


  xor
  g903
  (
    n879,
    n792,
    n742,
    n713
  );


  nand
  g904
  (
    n886,
    n757,
    n716,
    n706
  );


  xor
  g905
  (
    n890,
    n548,
    n537,
    n774
  );


  nor
  g906
  (
    n815,
    n540,
    n549,
    n791
  );


  and
  g907
  (
    n824,
    n776,
    n800,
    n553
  );


  xnor
  g908
  (
    n945,
    n544,
    n572,
    n771
  );


  xnor
  g909
  (
    n895,
    n708,
    n542,
    n769
  );


  and
  g910
  (
    n891,
    n730,
    n578,
    n766
  );


  or
  g911
  (
    n829,
    n790,
    n741,
    n715
  );


  nor
  g912
  (
    n939,
    n723,
    n568,
    n560
  );


  nor
  g913
  (
    n940,
    n763,
    n557,
    n802
  );


  nand
  g914
  (
    n874,
    n546,
    n758,
    n760
  );


  xor
  g915
  (
    n830,
    n712,
    n537,
    n755
  );


  or
  g916
  (
    n854,
    n733,
    n799,
    n724
  );


  or
  g917
  (
    n883,
    n730,
    n808,
    n572
  );


  xnor
  g918
  (
    n899,
    n766,
    n725,
    n797
  );


  or
  g919
  (
    n920,
    n797,
    n202,
    n758
  );


  nand
  g920
  (
    n917,
    n796,
    n734,
    n738
  );


  xor
  g921
  (
    n862,
    n788,
    n705,
    n739
  );


  or
  g922
  (
    n882,
    n732,
    n764,
    n203
  );


  xor
  g923
  (
    n888,
    n550,
    n768,
    n553
  );


  nand
  g924
  (
    n863,
    n544,
    n561,
    n543
  );


  nand
  g925
  (
    n894,
    n760,
    n803,
    n562
  );


  xnor
  g926
  (
    n837,
    n568,
    n723,
    n702
  );


  or
  g927
  (
    n966,
    n729,
    n808,
    n795
  );


  xor
  g928
  (
    n896,
    n736,
    n570,
    n573
  );


  xnor
  g929
  (
    n918,
    n733,
    n798,
    n762
  );


  xor
  g930
  (
    KeyWire_0_18,
    n779,
    n810,
    n558
  );


  xnor
  g931
  (
    n868,
    n701,
    n574,
    n799
  );


  and
  g932
  (
    n944,
    n577,
    n552,
    n744,
    n536
  );


  or
  g933
  (
    n969,
    n729,
    n737,
    n564,
    n743
  );


  xnor
  g934
  (
    n921,
    n797,
    n808,
    n771,
    n767
  );


  nor
  g935
  (
    n903,
    n203,
    n551,
    n728,
    n713
  );


  nand
  g936
  (
    n818,
    n781,
    n793,
    n760,
    n772
  );


  nor
  g937
  (
    n941,
    n735,
    n751,
    n781,
    n550
  );


  xnor
  g938
  (
    n850,
    n537,
    n757,
    n785,
    n746
  );


  nand
  g939
  (
    n949,
    n761,
    n777,
    n775,
    n717
  );


  xor
  g940
  (
    n929,
    n564,
    n538,
    n566,
    n804
  );


  and
  g941
  (
    n980,
    n836,
    n822,
    n878,
    n824
  );


  and
  g942
  (
    n981,
    n854,
    n970,
    n958,
    n888
  );


  nor
  g943
  (
    n978,
    n932,
    n889,
    n918,
    n960
  );


  or
  g944
  (
    n1013,
    n814,
    n901,
    n815,
    n895
  );


  xor
  g945
  (
    n1001,
    n881,
    n937,
    n933,
    n965
  );


  or
  g946
  (
    n977,
    n812,
    n906,
    n206,
    n828
  );


  nor
  g947
  (
    n1011,
    n839,
    n817,
    n873,
    n957
  );


  or
  g948
  (
    n990,
    n894,
    n206,
    n863,
    n853
  );


  xor
  g949
  (
    n1006,
    n944,
    n907,
    n930,
    n964
  );


  or
  g950
  (
    n989,
    n856,
    n949,
    n862,
    n953
  );


  nor
  g951
  (
    n1014,
    n880,
    n905,
    n869,
    n206
  );


  xor
  g952
  (
    n995,
    n830,
    n943,
    n831,
    n952
  );


  xnor
  g953
  (
    n1002,
    n946,
    n911,
    n842,
    n821
  );


  xor
  g954
  (
    n1007,
    n896,
    n940,
    n859,
    n904
  );


  nand
  g955
  (
    n982,
    n899,
    n811,
    n867,
    n835
  );


  xnor
  g956
  (
    n999,
    n858,
    n860,
    n887,
    n840
  );


  nor
  g957
  (
    n983,
    n947,
    n816,
    n913,
    n882
  );


  xor
  g958
  (
    n988,
    n865,
    n833,
    n838,
    n870
  );


  and
  g959
  (
    n1004,
    n855,
    n972,
    n900,
    n898
  );


  xnor
  g960
  (
    n1010,
    n866,
    n834,
    n928,
    n969
  );


  or
  g961
  (
    n996,
    n925,
    n868,
    n890,
    n850
  );


  xnor
  g962
  (
    n984,
    n916,
    n846,
    n915,
    n844
  );


  nand
  g963
  (
    n1008,
    n823,
    n921,
    n877,
    n891
  );


  nand
  g964
  (
    n987,
    n939,
    n938,
    n945,
    n852
  );


  and
  g965
  (
    n1005,
    n206,
    n825,
    n948,
    n902
  );


  xor
  g966
  (
    n1000,
    n886,
    n936,
    n885,
    n919
  );


  xnor
  g967
  (
    n976,
    n883,
    n962,
    n832,
    n874
  );


  or
  g968
  (
    n1015,
    n845,
    n954,
    n956,
    n909
  );


  and
  g969
  (
    n1003,
    n861,
    n820,
    n924,
    n827
  );


  xnor
  g970
  (
    n1012,
    n841,
    n950,
    n968,
    n847
  );


  xnor
  g971
  (
    n974,
    n864,
    n912,
    n871,
    n923
  );


  xor
  g972
  (
    KeyWire_0_4,
    n926,
    n963,
    n941,
    n897
  );


  nand
  g973
  (
    n992,
    n927,
    n843,
    n813,
    n917
  );


  nor
  g974
  (
    n998,
    n955,
    n884,
    n829,
    n922
  );


  or
  g975
  (
    n993,
    n931,
    n702,
    n935,
    n851
  );


  xor
  g976
  (
    n1009,
    n837,
    n819,
    n966,
    n910
  );


  xnor
  g977
  (
    n991,
    n920,
    n903,
    n942,
    n849
  );


  nand
  g978
  (
    n979,
    n875,
    n914,
    n967,
    n971
  );


  nor
  g979
  (
    n986,
    n892,
    n961,
    n951,
    n893
  );


  xnor
  g980
  (
    n985,
    n908,
    n934,
    n959,
    n848
  );


  nor
  g981
  (
    n975,
    n879,
    n826,
    n876,
    n818
  );


  and
  g982
  (
    n994,
    n857,
    n872,
    n973,
    n929
  );


  nand
  g983
  (
    n1021,
    n981,
    n630,
    n996,
    n1002
  );


  nor
  g984
  (
    n1017,
    n990,
    n1005,
    n631,
    n634
  );


  xnor
  g985
  (
    KeyWire_0_7,
    n1009,
    n636,
    n984,
    n1007
  );


  and
  g986
  (
    n1028,
    n631,
    n994,
    n632,
    n979
  );


  nand
  g987
  (
    n1027,
    n974,
    n1008,
    n998,
    n977
  );


  xnor
  g988
  (
    n1029,
    n633,
    n636,
    n985,
    n976
  );


  xnor
  g989
  (
    n1022,
    n635,
    n634,
    n995
  );


  xnor
  g990
  (
    n1020,
    n1013,
    n632,
    n631,
    n630
  );


  xnor
  g991
  (
    n1030,
    n631,
    n986,
    n635,
    n997
  );


  and
  g992
  (
    n1019,
    n1006,
    n987,
    n635,
    n1014
  );


  xnor
  g993
  (
    n1018,
    n1012,
    n1000,
    n992,
    n634
  );


  nor
  g994
  (
    n1025,
    n982,
    n636,
    n633
  );


  nand
  g995
  (
    n1026,
    n1001,
    n989,
    n999,
    n975
  );


  or
  g996
  (
    n1024,
    n993,
    n635,
    n1010,
    n991
  );


  xnor
  g997
  (
    n1023,
    n1004,
    n1011,
    n632
  );


  or
  g998
  (
    n1031,
    n1015,
    n633,
    n983,
    n988
  );


  nand
  g999
  (
    n1016,
    n980,
    n636,
    n1003,
    n978
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n700,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n503,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n165,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n801,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n997,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n528,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n167,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1032,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n462,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n609,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n266,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n301,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n389,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n659,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n807,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n235,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n199,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n704,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n902,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n743,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n965,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n162,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n935,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n243,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n600,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n649,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n73,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n711,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n759,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n323,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n344,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n789,
    KeyNOTWire_0_31
  );


endmodule

