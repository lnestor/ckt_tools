

module Stat_1352_44_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n986,
  n983,
  n979,
  n981,
  n974,
  n980,
  n987,
  n975,
  n978,
  n976,
  n1097,
  n1375,
  n1370,
  n1371,
  n1377,
  n1376,
  n1374,
  n1372,
  n1383
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n986;output n983;output n979;output n981;output n974;output n980;output n987;output n975;output n978;output n976;output n1097;output n1375;output n1370;output n1371;output n1377;output n1376;output n1374;output n1372;output n1383;
  wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n977;wire n982;wire n984;wire n985;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1373;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n36,
    n1
  );


  not
  g1
  (
    n126,
    n24
  );


  buf
  g2
  (
    n52,
    n27
  );


  not
  g3
  (
    n51,
    n25
  );


  buf
  g4
  (
    n80,
    n16
  );


  buf
  g5
  (
    n137,
    n31
  );


  not
  g6
  (
    n144,
    n29
  );


  buf
  g7
  (
    n141,
    n26
  );


  buf
  g8
  (
    n140,
    n12
  );


  not
  g9
  (
    n39,
    n20
  );


  not
  g10
  (
    n70,
    n6
  );


  not
  g11
  (
    n152,
    n16
  );


  buf
  g12
  (
    n101,
    n26
  );


  not
  g13
  (
    n65,
    n11
  );


  not
  g14
  (
    n143,
    n13
  );


  not
  g15
  (
    n132,
    n22
  );


  buf
  g16
  (
    n49,
    n15
  );


  buf
  g17
  (
    n63,
    n11
  );


  not
  g18
  (
    n35,
    n12
  );


  buf
  g19
  (
    n40,
    n12
  );


  not
  g20
  (
    n68,
    n30
  );


  not
  g21
  (
    n125,
    n20
  );


  not
  g22
  (
    n62,
    n18
  );


  buf
  g23
  (
    n103,
    n3
  );


  buf
  g24
  (
    n147,
    n1
  );


  not
  g25
  (
    n90,
    n8
  );


  not
  g26
  (
    n114,
    n21
  );


  not
  g27
  (
    n96,
    n24
  );


  not
  g28
  (
    n98,
    n13
  );


  buf
  g29
  (
    n86,
    n25
  );


  buf
  g30
  (
    n122,
    n4
  );


  not
  g31
  (
    n118,
    n6
  );


  not
  g32
  (
    n46,
    n16
  );


  buf
  g33
  (
    n131,
    n19
  );


  buf
  g34
  (
    n115,
    n30
  );


  not
  g35
  (
    n33,
    n26
  );


  buf
  g36
  (
    n151,
    n4
  );


  not
  g37
  (
    n111,
    n25
  );


  buf
  g38
  (
    n135,
    n23
  );


  not
  g39
  (
    n102,
    n22
  );


  not
  g40
  (
    n64,
    n21
  );


  buf
  g41
  (
    n83,
    n7
  );


  buf
  g42
  (
    n138,
    n5
  );


  not
  g43
  (
    n121,
    n9
  );


  buf
  g44
  (
    n85,
    n13
  );


  not
  g45
  (
    n55,
    n1
  );


  not
  g46
  (
    n44,
    n20
  );


  buf
  g47
  (
    n79,
    n30
  );


  buf
  g48
  (
    n155,
    n3
  );


  buf
  g49
  (
    n72,
    n24
  );


  not
  g50
  (
    n74,
    n4
  );


  buf
  g51
  (
    n104,
    n9
  );


  buf
  g52
  (
    n56,
    n29
  );


  buf
  g53
  (
    n117,
    n23
  );


  buf
  g54
  (
    n139,
    n2
  );


  not
  g55
  (
    n50,
    n23
  );


  buf
  g56
  (
    n76,
    n22
  );


  not
  g57
  (
    n53,
    n12
  );


  buf
  g58
  (
    n134,
    n3
  );


  not
  g59
  (
    n112,
    n19
  );


  not
  g60
  (
    n145,
    n2
  );


  not
  g61
  (
    n41,
    n5
  );


  buf
  g62
  (
    n82,
    n4
  );


  buf
  g63
  (
    n149,
    n7
  );


  not
  g64
  (
    n47,
    n22
  );


  buf
  g65
  (
    n123,
    n6
  );


  buf
  g66
  (
    n81,
    n15
  );


  not
  g67
  (
    n129,
    n11
  );


  buf
  g68
  (
    n107,
    n17
  );


  not
  g69
  (
    n95,
    n15
  );


  not
  g70
  (
    n88,
    n28
  );


  not
  g71
  (
    n154,
    n8
  );


  not
  g72
  (
    n59,
    n18
  );


  buf
  g73
  (
    n57,
    n1
  );


  not
  g74
  (
    n61,
    n10
  );


  buf
  g75
  (
    n128,
    n28
  );


  buf
  g76
  (
    n119,
    n27
  );


  not
  g77
  (
    n42,
    n20
  );


  buf
  g78
  (
    n73,
    n26
  );


  not
  g79
  (
    n37,
    n2
  );


  buf
  g80
  (
    n113,
    n7
  );


  not
  g81
  (
    n94,
    n14
  );


  buf
  g82
  (
    n69,
    n8
  );


  buf
  g83
  (
    n105,
    n19
  );


  buf
  g84
  (
    n77,
    n10
  );


  buf
  g85
  (
    n146,
    n11
  );


  buf
  g86
  (
    n84,
    n18
  );


  buf
  g87
  (
    n133,
    n31
  );


  buf
  g88
  (
    n67,
    n17
  );


  buf
  g89
  (
    n54,
    n10
  );


  not
  g90
  (
    n130,
    n31
  );


  buf
  g91
  (
    n58,
    n8
  );


  not
  g92
  (
    n110,
    n25
  );


  not
  g93
  (
    n109,
    n17
  );


  not
  g94
  (
    n108,
    n9
  );


  buf
  g95
  (
    n100,
    n19
  );


  not
  g96
  (
    n78,
    n31
  );


  buf
  g97
  (
    n34,
    n27
  );


  not
  g98
  (
    n66,
    n10
  );


  buf
  g99
  (
    n150,
    n5
  );


  not
  g100
  (
    n75,
    n17
  );


  buf
  g101
  (
    n148,
    n24
  );


  buf
  g102
  (
    n48,
    n14
  );


  not
  g103
  (
    n142,
    n9
  );


  not
  g104
  (
    n43,
    n3
  );


  buf
  g105
  (
    n71,
    n2
  );


  not
  g106
  (
    n136,
    n21
  );


  buf
  g107
  (
    n127,
    n16
  );


  not
  g108
  (
    n93,
    n27
  );


  buf
  g109
  (
    n87,
    n29
  );


  buf
  g110
  (
    n45,
    n15
  );


  buf
  g111
  (
    n106,
    n13
  );


  buf
  g112
  (
    n116,
    n30
  );


  not
  g113
  (
    KeyWire_0_25,
    n28
  );


  buf
  g114
  (
    n153,
    n7
  );


  not
  g115
  (
    n99,
    n28
  );


  buf
  g116
  (
    n60,
    n6
  );


  not
  g117
  (
    n32,
    n14
  );


  not
  g118
  (
    n91,
    n23
  );


  not
  g119
  (
    n120,
    n29
  );


  buf
  g120
  (
    n124,
    n14
  );


  not
  g121
  (
    n97,
    n18
  );


  buf
  g122
  (
    n92,
    n21
  );


  buf
  g123
  (
    n38,
    n5
  );


  not
  g124
  (
    n179,
    n113
  );


  buf
  g125
  (
    n291,
    n110
  );


  not
  g126
  (
    n203,
    n49
  );


  not
  g127
  (
    n185,
    n116
  );


  not
  g128
  (
    n400,
    n151
  );


  buf
  g129
  (
    n236,
    n100
  );


  not
  g130
  (
    KeyWire_0_21,
    n103
  );


  buf
  g131
  (
    n262,
    n94
  );


  buf
  g132
  (
    n201,
    n51
  );


  not
  g133
  (
    n274,
    n68
  );


  buf
  g134
  (
    n200,
    n49
  );


  buf
  g135
  (
    n250,
    n95
  );


  not
  g136
  (
    n269,
    n59
  );


  buf
  g137
  (
    n293,
    n153
  );


  not
  g138
  (
    n342,
    n68
  );


  buf
  g139
  (
    n268,
    n81
  );


  buf
  g140
  (
    n401,
    n96
  );


  not
  g141
  (
    n298,
    n138
  );


  buf
  g142
  (
    n156,
    n55
  );


  not
  g143
  (
    n176,
    n130
  );


  buf
  g144
  (
    n296,
    n149
  );


  buf
  g145
  (
    n260,
    n85
  );


  not
  g146
  (
    n227,
    n42
  );


  buf
  g147
  (
    n208,
    n154
  );


  not
  g148
  (
    n302,
    n147
  );


  buf
  g149
  (
    n390,
    n81
  );


  buf
  g150
  (
    n270,
    n140
  );


  not
  g151
  (
    n213,
    n137
  );


  not
  g152
  (
    n166,
    n63
  );


  not
  g153
  (
    n281,
    n97
  );


  not
  g154
  (
    KeyWire_0_15,
    n111
  );


  not
  g155
  (
    n228,
    n122
  );


  not
  g156
  (
    n277,
    n126
  );


  not
  g157
  (
    n170,
    n34
  );


  buf
  g158
  (
    n285,
    n93
  );


  buf
  g159
  (
    n244,
    n113
  );


  not
  g160
  (
    n326,
    n90
  );


  not
  g161
  (
    n346,
    n102
  );


  not
  g162
  (
    n340,
    n44
  );


  not
  g163
  (
    n252,
    n141
  );


  not
  g164
  (
    n239,
    n44
  );


  buf
  g165
  (
    n218,
    n39
  );


  not
  g166
  (
    n329,
    n122
  );


  not
  g167
  (
    n348,
    n102
  );


  not
  g168
  (
    n339,
    n35
  );


  not
  g169
  (
    n328,
    n76
  );


  buf
  g170
  (
    n362,
    n63
  );


  buf
  g171
  (
    n397,
    n115
  );


  not
  g172
  (
    n283,
    n45
  );


  not
  g173
  (
    KeyWire_0_14,
    n88
  );


  not
  g174
  (
    n160,
    n94
  );


  buf
  g175
  (
    n369,
    n132
  );


  not
  g176
  (
    n365,
    n117
  );


  not
  g177
  (
    n377,
    n48
  );


  buf
  g178
  (
    n187,
    n70
  );


  buf
  g179
  (
    KeyWire_0_28,
    n139
  );


  not
  g180
  (
    n199,
    n54
  );


  buf
  g181
  (
    n387,
    n35
  );


  buf
  g182
  (
    n210,
    n57
  );


  not
  g183
  (
    n163,
    n135
  );


  not
  g184
  (
    n168,
    n135
  );


  buf
  g185
  (
    n192,
    n144
  );


  buf
  g186
  (
    n261,
    n74
  );


  buf
  g187
  (
    n157,
    n65
  );


  buf
  g188
  (
    n247,
    n125
  );


  not
  g189
  (
    n374,
    n77
  );


  buf
  g190
  (
    n164,
    n74
  );


  buf
  g191
  (
    n386,
    n120
  );


  not
  g192
  (
    n195,
    n150
  );


  buf
  g193
  (
    n169,
    n63
  );


  not
  g194
  (
    n198,
    n53
  );


  buf
  g195
  (
    n307,
    n98
  );


  buf
  g196
  (
    n224,
    n151
  );


  buf
  g197
  (
    n321,
    n114
  );


  buf
  g198
  (
    n324,
    n96
  );


  not
  g199
  (
    n344,
    n75
  );


  buf
  g200
  (
    n354,
    n117
  );


  buf
  g201
  (
    n217,
    n91
  );


  buf
  g202
  (
    n193,
    n58
  );


  not
  g203
  (
    n197,
    n147
  );


  not
  g204
  (
    n189,
    n111
  );


  buf
  g205
  (
    n259,
    n71
  );


  not
  g206
  (
    n186,
    n70
  );


  buf
  g207
  (
    n212,
    n77
  );


  buf
  g208
  (
    n368,
    n77
  );


  not
  g209
  (
    n371,
    n148
  );


  not
  g210
  (
    n347,
    n33
  );


  not
  g211
  (
    KeyWire_0_6,
    n152
  );


  not
  g212
  (
    n367,
    n50
  );


  buf
  g213
  (
    n353,
    n103
  );


  buf
  g214
  (
    n319,
    n38
  );


  not
  g215
  (
    n209,
    n78
  );


  not
  g216
  (
    n318,
    n33
  );


  not
  g217
  (
    n309,
    n138
  );


  buf
  g218
  (
    n216,
    n70
  );


  not
  g219
  (
    n159,
    n37
  );


  buf
  g220
  (
    n240,
    n107
  );


  buf
  g221
  (
    n273,
    n60
  );


  buf
  g222
  (
    n337,
    n133
  );


  not
  g223
  (
    n297,
    n86
  );


  not
  g224
  (
    n161,
    n138
  );


  buf
  g225
  (
    n278,
    n64
  );


  not
  g226
  (
    n320,
    n142
  );


  buf
  g227
  (
    n359,
    n154
  );


  buf
  g228
  (
    n194,
    n55
  );


  not
  g229
  (
    n338,
    n54
  );


  buf
  g230
  (
    n233,
    n79
  );


  not
  g231
  (
    n178,
    n40
  );


  not
  g232
  (
    n222,
    n99
  );


  not
  g233
  (
    n280,
    n68
  );


  not
  g234
  (
    n290,
    n137
  );


  buf
  g235
  (
    n266,
    n83
  );


  not
  g236
  (
    n393,
    n131
  );


  not
  g237
  (
    n349,
    n106
  );


  buf
  g238
  (
    n196,
    n78
  );


  buf
  g239
  (
    n255,
    n61
  );


  not
  g240
  (
    KeyWire_0_16,
    n127
  );


  not
  g241
  (
    n295,
    n45
  );


  not
  g242
  (
    n288,
    n86
  );


  not
  g243
  (
    n287,
    n133
  );


  not
  g244
  (
    n330,
    n47
  );


  buf
  g245
  (
    n177,
    n100
  );


  not
  g246
  (
    n271,
    n56
  );


  buf
  g247
  (
    n165,
    n67
  );


  not
  g248
  (
    n301,
    n97
  );


  buf
  g249
  (
    n219,
    n151
  );


  buf
  g250
  (
    n305,
    n144
  );


  buf
  g251
  (
    n174,
    n80
  );


  not
  g252
  (
    n246,
    n41
  );


  not
  g253
  (
    n317,
    n101
  );


  buf
  g254
  (
    n292,
    n82
  );


  not
  g255
  (
    n171,
    n76
  );


  buf
  g256
  (
    n322,
    n42
  );


  not
  g257
  (
    n395,
    n46
  );


  not
  g258
  (
    n331,
    n91
  );


  not
  g259
  (
    n299,
    n123
  );


  not
  g260
  (
    n363,
    n61
  );


  buf
  g261
  (
    n207,
    n121
  );


  not
  g262
  (
    n223,
    n45
  );


  not
  g263
  (
    KeyWire_0_0,
    n142
  );


  buf
  g264
  (
    n383,
    n37
  );


  not
  g265
  (
    n300,
    n116
  );


  not
  g266
  (
    n180,
    n120
  );


  not
  g267
  (
    n308,
    n148
  );


  not
  g268
  (
    n242,
    n143
  );


  buf
  g269
  (
    n182,
    n143
  );


  not
  g270
  (
    n238,
    n51
  );


  buf
  g271
  (
    n241,
    n61
  );


  buf
  g272
  (
    n235,
    n75
  );


  buf
  g273
  (
    n230,
    n101
  );


  buf
  g274
  (
    n265,
    n149
  );


  not
  g275
  (
    n289,
    n119
  );


  buf
  g276
  (
    n398,
    n85
  );


  not
  g277
  (
    n335,
    n132
  );


  not
  g278
  (
    KeyWire_0_5,
    n58
  );


  not
  g279
  (
    n257,
    n52
  );


  buf
  g280
  (
    n181,
    n52
  );


  not
  g281
  (
    n336,
    n47
  );


  buf
  g282
  (
    n282,
    n133
  );


  buf
  g283
  (
    n345,
    n64
  );


  not
  g284
  (
    n284,
    n81
  );


  not
  g285
  (
    n378,
    n121
  );


  buf
  g286
  (
    n373,
    n109
  );


  not
  g287
  (
    n272,
    n43
  );


  xnor
  g288
  (
    n351,
    n144,
    n150
  );


  and
  g289
  (
    KeyWire_0_22,
    n136,
    n58,
    n69,
    n85
  );


  or
  g290
  (
    n229,
    n84,
    n129,
    n35,
    n120
  );


  xnor
  g291
  (
    n304,
    n66,
    n119,
    n80,
    n99
  );


  and
  g292
  (
    n343,
    n66,
    n114,
    n126,
    n37
  );


  xnor
  g293
  (
    n356,
    n127,
    n36,
    n146,
    n124
  );


  xnor
  g294
  (
    n358,
    n125,
    n69,
    n100
  );


  xnor
  g295
  (
    n364,
    n59,
    n34,
    n48,
    n124
  );


  xor
  g296
  (
    n352,
    n67,
    n75,
    n90,
    n41
  );


  xnor
  g297
  (
    n361,
    n54,
    n121,
    n83,
    n95
  );


  xor
  g298
  (
    n382,
    n78,
    n60,
    n101,
    n52
  );


  nor
  g299
  (
    n396,
    n126,
    n84,
    n88,
    n48
  );


  nor
  g300
  (
    n220,
    n123,
    n110,
    n32,
    n111
  );


  xor
  g301
  (
    n314,
    n104,
    n65,
    n34,
    n103
  );


  or
  g302
  (
    n245,
    n108,
    n147,
    n115,
    n91
  );


  xor
  g303
  (
    n276,
    n142,
    n80,
    n42,
    n107
  );


  nor
  g304
  (
    n311,
    n66,
    n43,
    n45,
    n130
  );


  nand
  g305
  (
    n184,
    n127,
    n101,
    n88,
    n59
  );


  nand
  g306
  (
    n399,
    n134,
    n76,
    n69,
    n96
  );


  and
  g307
  (
    n267,
    n77,
    n72,
    n107,
    n91
  );


  xnor
  g308
  (
    n375,
    n80,
    n83,
    n86,
    n110
  );


  nor
  g309
  (
    n323,
    n64,
    n93,
    n153,
    n109
  );


  or
  g310
  (
    n249,
    n132,
    n129,
    n38,
    n65
  );


  nand
  g311
  (
    n248,
    n126,
    n62,
    n128,
    n110
  );


  and
  g312
  (
    n384,
    n96,
    n112,
    n84,
    n94
  );


  or
  g313
  (
    n333,
    n62,
    n104,
    n40,
    n93
  );


  or
  g314
  (
    n350,
    n62,
    n88,
    n148,
    n49
  );


  xnor
  g315
  (
    n332,
    n129,
    n89,
    n98,
    n54
  );


  nand
  g316
  (
    n286,
    n36,
    n72,
    n47,
    n46
  );


  and
  g317
  (
    n232,
    n44,
    n151,
    n95,
    n102
  );


  and
  g318
  (
    n167,
    n122,
    n115,
    n132,
    n149
  );


  or
  g319
  (
    n264,
    n66,
    n108,
    n39,
    n128
  );


  nand
  g320
  (
    n388,
    n33,
    n67,
    n94,
    n113
  );


  and
  g321
  (
    n392,
    n58,
    n141,
    n139,
    n113
  );


  nor
  g322
  (
    n372,
    n71,
    n102,
    n72,
    n127
  );


  nand
  g323
  (
    n391,
    n141,
    n118,
    n130,
    n116
  );


  and
  g324
  (
    n226,
    n108,
    n52,
    n134,
    n128
  );


  or
  g325
  (
    n325,
    n150,
    n43,
    n147,
    n129
  );


  nor
  g326
  (
    n231,
    n56,
    n32,
    n143,
    n47
  );


  nand
  g327
  (
    n379,
    n146,
    n135,
    n84,
    n140
  );


  xnor
  g328
  (
    n256,
    n92,
    n152,
    n123,
    n61
  );


  xor
  g329
  (
    n205,
    n136,
    n98,
    n140,
    n139
  );


  nand
  g330
  (
    n370,
    n50,
    n90,
    n86,
    n145
  );


  nand
  g331
  (
    n360,
    n108,
    n57,
    n87,
    n89
  );


  nor
  g332
  (
    n310,
    n60,
    n36,
    n146,
    n49
  );


  or
  g333
  (
    n303,
    n55,
    n136,
    n140,
    n64
  );


  nand
  g334
  (
    n327,
    n124,
    n117,
    n130,
    n57
  );


  and
  g335
  (
    n190,
    n92,
    n81,
    n69,
    n79
  );


  xnor
  g336
  (
    n191,
    n149,
    n34,
    n63,
    n118
  );


  or
  g337
  (
    n234,
    n90,
    n97,
    n139,
    n60
  );


  nor
  g338
  (
    n279,
    n117,
    n134,
    n73,
    n121
  );


  nor
  g339
  (
    n306,
    n106,
    n145,
    n33,
    n89
  );


  nor
  g340
  (
    n204,
    n135,
    n53,
    n87
  );


  or
  g341
  (
    n263,
    n71,
    n105,
    n98,
    n32
  );


  or
  g342
  (
    n275,
    n103,
    n73,
    n74
  );


  xor
  g343
  (
    n183,
    n148,
    n114,
    n85,
    n107
  );


  nor
  g344
  (
    n315,
    n93,
    n134,
    n70,
    n50
  );


  xor
  g345
  (
    n389,
    n82,
    n131,
    n145,
    n153
  );


  and
  g346
  (
    n225,
    n41,
    n125,
    n111,
    n83
  );


  or
  g347
  (
    n172,
    n142,
    n141,
    n137,
    n125
  );


  xnor
  g348
  (
    KeyWire_0_24,
    n92,
    n78,
    n119,
    n118
  );


  nor
  g349
  (
    n258,
    n138,
    n79,
    n87,
    n42
  );


  xnor
  g350
  (
    n173,
    n116,
    n109,
    n137,
    n152
  );


  and
  g351
  (
    n215,
    n43,
    n73,
    n76,
    n44
  );


  nand
  g352
  (
    n316,
    n82,
    n152,
    n65,
    n75
  );


  or
  g353
  (
    n206,
    n82,
    n57,
    n109,
    n99
  );


  or
  g354
  (
    n334,
    n112,
    n99,
    n105,
    n119
  );


  xor
  g355
  (
    n341,
    n89,
    n36,
    n79,
    n46
  );


  or
  g356
  (
    n381,
    n56,
    n133,
    n46,
    n73
  );


  and
  g357
  (
    n202,
    n40,
    n118,
    n114,
    n146
  );


  xnor
  g358
  (
    n312,
    n51,
    n153,
    n50,
    n104
  );


  xor
  g359
  (
    n357,
    n112,
    n55,
    n32,
    n92
  );


  and
  g360
  (
    n158,
    n128,
    n106,
    n120,
    n131
  );


  xnor
  g361
  (
    n175,
    n56,
    n97,
    n105,
    n95
  );


  or
  g362
  (
    n385,
    n124,
    n144,
    n48,
    n112
  );


  nand
  g363
  (
    n243,
    n136,
    n115,
    n71,
    n39
  );


  nand
  g364
  (
    n394,
    n53,
    n40,
    n41,
    n123
  );


  xnor
  g365
  (
    n366,
    n62,
    n122,
    n67,
    n53
  );


  xnor
  g366
  (
    n254,
    n131,
    n38,
    n150,
    n104
  );


  nor
  g367
  (
    n188,
    n39,
    n105,
    n106,
    n38
  );


  xnor
  g368
  (
    n380,
    n72,
    n51,
    n68,
    n59
  );


  xor
  g369
  (
    n355,
    n35,
    n145,
    n37,
    n143
  );


  nand
  g370
  (
    n614,
    n231,
    n233,
    n250,
    n219
  );


  or
  g371
  (
    n473,
    n182,
    n288,
    n318,
    n210
  );


  and
  g372
  (
    n612,
    n324,
    n206,
    n267,
    n189
  );


  nand
  g373
  (
    n444,
    n234,
    n246,
    n157,
    n277
  );


  xnor
  g374
  (
    n565,
    n160,
    n271,
    n363,
    n199
  );


  nand
  g375
  (
    n531,
    n218,
    n257,
    n337,
    n295
  );


  or
  g376
  (
    n427,
    n206,
    n180,
    n353,
    n322
  );


  nor
  g377
  (
    n586,
    n191,
    n185,
    n275,
    n377
  );


  and
  g378
  (
    n410,
    n211,
    n215,
    n178,
    n337
  );


  and
  g379
  (
    n432,
    n242,
    n272,
    n350,
    n237
  );


  and
  g380
  (
    KeyWire_0_17,
    n357,
    n171,
    n311,
    n215
  );


  nor
  g381
  (
    n581,
    n346,
    n207,
    n221
  );


  xnor
  g382
  (
    n430,
    n298,
    n259,
    n339,
    n165
  );


  and
  g383
  (
    n541,
    n286,
    n304,
    n265,
    n226
  );


  xnor
  g384
  (
    n470,
    n247,
    n255,
    n240,
    n224
  );


  nor
  g385
  (
    n456,
    n181,
    n266,
    n184,
    n241
  );


  or
  g386
  (
    n551,
    n200,
    n190,
    n314,
    n222
  );


  xor
  g387
  (
    n591,
    n192,
    n376,
    n323,
    n346
  );


  nand
  g388
  (
    n461,
    n286,
    n213,
    n195,
    n167
  );


  or
  g389
  (
    n424,
    n335,
    n302,
    n311,
    n296
  );


  xor
  g390
  (
    n516,
    n220,
    n352,
    n244,
    n270
  );


  xor
  g391
  (
    n471,
    n347,
    n201,
    n179,
    n213
  );


  nand
  g392
  (
    n517,
    n231,
    n217,
    n375,
    n234
  );


  or
  g393
  (
    n404,
    n358,
    n230,
    n207,
    n355
  );


  xor
  g394
  (
    n537,
    n355,
    n156,
    n342,
    n191
  );


  or
  g395
  (
    n509,
    n374,
    n193,
    n290,
    n331
  );


  and
  g396
  (
    n577,
    n296,
    n287,
    n162,
    n240
  );


  xor
  g397
  (
    n536,
    n319,
    n270,
    n350,
    n251
  );


  nor
  g398
  (
    n447,
    n189,
    n334,
    n320,
    n364
  );


  and
  g399
  (
    n440,
    n165,
    n379,
    n310,
    n264
  );


  and
  g400
  (
    n532,
    n278,
    n219,
    n216,
    n263
  );


  nand
  g401
  (
    n535,
    n284,
    n179,
    n188,
    n264
  );


  nand
  g402
  (
    n479,
    n301,
    n348,
    n220,
    n346
  );


  xor
  g403
  (
    n606,
    n261,
    n239,
    n380,
    n303
  );


  xor
  g404
  (
    n467,
    n367,
    n252,
    n371,
    n381
  );


  and
  g405
  (
    n550,
    n351,
    n238,
    n166,
    n308
  );


  xnor
  g406
  (
    n623,
    n168,
    n316,
    n275,
    n297
  );


  nand
  g407
  (
    n522,
    n159,
    n236,
    n286,
    n282
  );


  or
  g408
  (
    n469,
    n211,
    n241,
    n281,
    n327
  );


  nor
  g409
  (
    n575,
    n336,
    n366,
    n310,
    n313
  );


  nand
  g410
  (
    n406,
    n201,
    n209,
    n292,
    n228
  );


  xnor
  g411
  (
    n482,
    n315,
    n284,
    n293,
    n338
  );


  xor
  g412
  (
    n553,
    n208,
    n159,
    n276,
    n356
  );


  xor
  g413
  (
    n474,
    n378,
    n331,
    n194,
    n376
  );


  xnor
  g414
  (
    n562,
    n170,
    n343,
    n282,
    n231
  );


  and
  g415
  (
    n620,
    n164,
    n381,
    n245,
    n312
  );


  nand
  g416
  (
    n428,
    n209,
    n285,
    n334,
    n300
  );


  xor
  g417
  (
    KeyWire_0_29,
    n337,
    n321,
    n299,
    n263
  );


  xnor
  g418
  (
    n403,
    n371,
    n360,
    n374,
    n187
  );


  xnor
  g419
  (
    n437,
    n288,
    n317,
    n297,
    n238
  );


  or
  g420
  (
    n411,
    n279,
    n309,
    n306,
    n333
  );


  and
  g421
  (
    n557,
    n232,
    n280,
    n372,
    n168
  );


  xor
  g422
  (
    n413,
    n257,
    n289,
    n266,
    n377
  );


  or
  g423
  (
    n602,
    n232,
    n289,
    n192,
    n322
  );


  nand
  g424
  (
    n506,
    n233,
    n343,
    n347,
    n176
  );


  xor
  g425
  (
    n483,
    n252,
    n208,
    n205,
    n228
  );


  and
  g426
  (
    n502,
    n191,
    n335,
    n206,
    n365
  );


  nand
  g427
  (
    n615,
    n244,
    n259,
    n334,
    n212
  );


  xor
  g428
  (
    n543,
    n367,
    n320,
    n301,
    n275
  );


  nand
  g429
  (
    n567,
    n270,
    n193,
    n178,
    n180
  );


  or
  g430
  (
    n464,
    n305,
    n262,
    n315,
    n269
  );


  xnor
  g431
  (
    n457,
    n309,
    n288,
    n262,
    n339
  );


  xor
  g432
  (
    n415,
    n226,
    n242,
    n295,
    n158
  );


  nand
  g433
  (
    n592,
    n266,
    n244,
    n280,
    n380
  );


  nor
  g434
  (
    n435,
    n275,
    n368,
    n382,
    n364
  );


  xor
  g435
  (
    n569,
    n354,
    n261,
    n163,
    n361
  );


  and
  g436
  (
    n465,
    n304,
    n376,
    n222,
    n347
  );


  or
  g437
  (
    n405,
    n181,
    n244,
    n370,
    n352
  );


  and
  g438
  (
    n547,
    n321,
    n249,
    n281,
    n221
  );


  nor
  g439
  (
    n618,
    n235,
    n299,
    n274,
    n358
  );


  xor
  g440
  (
    n625,
    n254,
    n261,
    n292,
    n367
  );


  or
  g441
  (
    n608,
    n303,
    n205,
    n167,
    n328
  );


  nand
  g442
  (
    n594,
    n223,
    n247,
    n378,
    n183
  );


  xor
  g443
  (
    n564,
    n382,
    n360,
    n330,
    n259
  );


  nor
  g444
  (
    n488,
    n189,
    n350,
    n278,
    n309
  );


  or
  g445
  (
    n610,
    n197,
    n246,
    n209,
    n375
  );


  xor
  g446
  (
    n554,
    n291,
    n373,
    n309,
    n274
  );


  nand
  g447
  (
    n490,
    n306,
    n369,
    n379,
    n203
  );


  nand
  g448
  (
    n500,
    n163,
    n317,
    n255,
    n264
  );


  and
  g449
  (
    n549,
    n203,
    n260,
    n374,
    n258
  );


  and
  g450
  (
    n595,
    n230,
    n213,
    n381,
    n258
  );


  nor
  g451
  (
    n556,
    n196,
    n305,
    n193,
    n366
  );


  or
  g452
  (
    n476,
    n292,
    n174,
    n283,
    n357
  );


  nand
  g453
  (
    n499,
    n258,
    n377,
    n333,
    n229
  );


  or
  g454
  (
    n438,
    n303,
    n185,
    n256,
    n194
  );


  xnor
  g455
  (
    n475,
    n181,
    n157,
    n324,
    n317
  );


  or
  g456
  (
    n421,
    n260,
    n310,
    n186,
    n211
  );


  nor
  g457
  (
    n582,
    n358,
    n362,
    n352,
    n341
  );


  or
  g458
  (
    n485,
    n285,
    n161,
    n326,
    n278
  );


  xor
  g459
  (
    n584,
    n370,
    n362,
    n280,
    n187
  );


  nor
  g460
  (
    n508,
    n365,
    n170,
    n324,
    n182
  );


  or
  g461
  (
    n628,
    n315,
    n268,
    n162,
    n182
  );


  xnor
  g462
  (
    n627,
    n227,
    n256,
    n157,
    n186
  );


  xnor
  g463
  (
    n420,
    n175,
    n321,
    n359,
    n190
  );


  nand
  g464
  (
    n548,
    n266,
    n180,
    n306,
    n161
  );


  and
  g465
  (
    n491,
    n248,
    n253,
    n370,
    n372
  );


  and
  g466
  (
    n605,
    n251,
    n217,
    n169,
    n284
  );


  nand
  g467
  (
    n559,
    n289,
    n222,
    n292,
    n302
  );


  xnor
  g468
  (
    n573,
    n239,
    n287,
    n280,
    n217
  );


  nand
  g469
  (
    n496,
    n223,
    n355,
    n327,
    n171
  );


  xor
  g470
  (
    n561,
    n190,
    n353,
    n215,
    n316
  );


  nand
  g471
  (
    n510,
    n314,
    n301,
    n237,
    n163
  );


  xnor
  g472
  (
    n617,
    n371,
    n248,
    n204,
    n353
  );


  or
  g473
  (
    n604,
    n381,
    n194,
    n326,
    n320
  );


  or
  g474
  (
    n505,
    n331,
    n295,
    n156,
    n351
  );


  and
  g475
  (
    n563,
    n205,
    n203,
    n315,
    n332
  );


  xor
  g476
  (
    n527,
    n380,
    n296,
    n310,
    n161
  );


  nand
  g477
  (
    n478,
    n335,
    n243,
    n246,
    n374
  );


  or
  g478
  (
    n619,
    n291,
    n300,
    n299,
    n200
  );


  or
  g479
  (
    n468,
    n261,
    n352,
    n361,
    n342
  );


  and
  g480
  (
    n472,
    n172,
    n255,
    n289,
    n225
  );


  xnor
  g481
  (
    n523,
    n156,
    n365,
    n363,
    n200
  );


  or
  g482
  (
    n626,
    n312,
    n224,
    n339,
    n202
  );


  xnor
  g483
  (
    n429,
    n358,
    n364,
    n198,
    n323
  );


  or
  g484
  (
    n451,
    n319,
    n282,
    n269,
    n316
  );


  xnor
  g485
  (
    n454,
    n277,
    n360,
    n159,
    n183
  );


  xor
  g486
  (
    n585,
    n186,
    n347,
    n201,
    n290
  );


  nand
  g487
  (
    n409,
    n171,
    n274,
    n242,
    n184
  );


  nor
  g488
  (
    n544,
    n329,
    n252,
    n322,
    n363
  );


  xnor
  g489
  (
    n449,
    n188,
    n219,
    n311,
    n225
  );


  nand
  g490
  (
    n542,
    n299,
    n227,
    n221,
    n354
  );


  xnor
  g491
  (
    n504,
    n160,
    n173,
    n240,
    n216
  );


  xor
  g492
  (
    n503,
    n276,
    n349,
    n203,
    n294
  );


  xnor
  g493
  (
    n560,
    n258,
    n334,
    n208,
    n165
  );


  nand
  g494
  (
    n446,
    n195,
    n342,
    n363,
    n168
  );


  nand
  g495
  (
    n486,
    n379,
    n345,
    n245,
    n298
  );


  nor
  g496
  (
    n622,
    n294,
    n284,
    n346,
    n212
  );


  xnor
  g497
  (
    n596,
    n173,
    n178,
    n325,
    n314
  );


  and
  g498
  (
    n515,
    n325,
    n257,
    n207,
    n342
  );


  or
  g499
  (
    n538,
    n368,
    n227,
    n196,
    n336
  );


  or
  g500
  (
    n603,
    n356,
    n234,
    n214,
    n286
  );


  xor
  g501
  (
    n607,
    n257,
    n167,
    n318,
    n164
  );


  xor
  g502
  (
    n416,
    n157,
    n220,
    n192,
    n364
  );


  and
  g503
  (
    n526,
    n336,
    n279,
    n169,
    n218
  );


  or
  g504
  (
    n419,
    n250,
    n187,
    n353,
    n182
  );


  xor
  g505
  (
    n579,
    n170,
    n362,
    n187,
    n311
  );


  xor
  g506
  (
    n583,
    n175,
    n229,
    n323,
    n294
  );


  and
  g507
  (
    n412,
    n225,
    n226,
    n190,
    n341
  );


  xor
  g508
  (
    n425,
    n236,
    n354,
    n376,
    n184
  );


  nor
  g509
  (
    n621,
    n262,
    n297,
    n168,
    n373
  );


  or
  g510
  (
    n558,
    n253,
    n343,
    n181,
    n349
  );


  and
  g511
  (
    n520,
    n192,
    n297,
    n166,
    n370
  );


  or
  g512
  (
    n588,
    n375,
    n326,
    n285,
    n161
  );


  xor
  g513
  (
    n576,
    n217,
    n287,
    n365,
    n366
  );


  nand
  g514
  (
    n484,
    n267,
    n273,
    n288,
    n176
  );


  nand
  g515
  (
    n418,
    n214,
    n291,
    n241,
    n232
  );


  nor
  g516
  (
    n601,
    n287,
    n274,
    n179,
    n279
  );


  xnor
  g517
  (
    n498,
    n158,
    n338,
    n223,
    n359
  );


  xnor
  g518
  (
    n452,
    n318,
    n172,
    n238,
    n184
  );


  xnor
  g519
  (
    n448,
    n254,
    n332,
    n209,
    n281
  );


  xnor
  g520
  (
    n546,
    n382,
    n204,
    n330,
    n216
  );


  nand
  g521
  (
    n528,
    n259,
    n177,
    n268,
    n378
  );


  and
  g522
  (
    n431,
    n233,
    n263,
    n178,
    n321
  );


  nand
  g523
  (
    n434,
    n369,
    n210,
    n324,
    n171
  );


  and
  g524
  (
    n402,
    n329,
    n198,
    n335,
    n298
  );


  nand
  g525
  (
    n459,
    n314,
    n262,
    n279,
    n307
  );


  nor
  g526
  (
    n519,
    n317,
    n298,
    n243,
    n237
  );


  or
  g527
  (
    n458,
    n271,
    n176,
    n201,
    n243
  );


  xor
  g528
  (
    n441,
    n272,
    n272,
    n349,
    n207
  );


  nand
  g529
  (
    n477,
    n162,
    n351,
    n158
  );


  nand
  g530
  (
    n507,
    n174,
    n328,
    n273,
    n340
  );


  or
  g531
  (
    n439,
    n382,
    n216,
    n338,
    n219
  );


  nor
  g532
  (
    n463,
    n350,
    n322,
    n197,
    n170
  );


  or
  g533
  (
    n407,
    n272,
    n340,
    n256,
    n231
  );


  or
  g534
  (
    n613,
    n238,
    n373,
    n380,
    n333
  );


  xor
  g535
  (
    n489,
    n235,
    n239,
    n211,
    n251
  );


  nand
  g536
  (
    n513,
    n248,
    n172,
    n176,
    n356
  );


  nor
  g537
  (
    n574,
    n225,
    n167,
    n263,
    n253
  );


  xnor
  g538
  (
    n501,
    n361,
    n372,
    n332,
    n189
  );


  nand
  g539
  (
    n443,
    n283,
    n196,
    n235,
    n331
  );


  and
  g540
  (
    n460,
    n333,
    n188,
    n304,
    n341
  );


  or
  g541
  (
    n455,
    n199,
    n173,
    n349,
    n177
  );


  nand
  g542
  (
    n590,
    n193,
    n233,
    n175,
    n226
  );


  xor
  g543
  (
    n518,
    n319,
    n328,
    n377,
    n269
  );


  nor
  g544
  (
    n533,
    n229,
    n247,
    n198,
    n276
  );


  xnor
  g545
  (
    n462,
    n268,
    n204,
    n249
  );


  xor
  g546
  (
    n530,
    n164,
    n336,
    n296,
    n351
  );


  nor
  g547
  (
    n487,
    n200,
    n308,
    n196,
    n294
  );


  xnor
  g548
  (
    n593,
    n267,
    n166,
    n245,
    n243
  );


  and
  g549
  (
    n426,
    n344,
    n359,
    n308,
    n210
  );


  and
  g550
  (
    n512,
    n254,
    n214,
    n195,
    n159
  );


  nand
  g551
  (
    n417,
    n345,
    n173,
    n227,
    n340
  );


  and
  g552
  (
    n525,
    n245,
    n162,
    n247,
    n362
  );


  xor
  g553
  (
    n481,
    n223,
    n301,
    n222,
    n337
  );


  nand
  g554
  (
    n514,
    n290,
    n273,
    n241,
    n237
  );


  and
  g555
  (
    n495,
    n312,
    n283,
    n368,
    n206
  );


  or
  g556
  (
    n466,
    n197,
    n308,
    n214,
    n185
  );


  nand
  g557
  (
    n571,
    n177,
    n293,
    n165,
    n260
  );


  or
  g558
  (
    KeyWire_0_12,
    n265,
    n252,
    n180,
    n371
  );


  nand
  g559
  (
    n568,
    n239,
    n319,
    n368,
    n305
  );


  nand
  g560
  (
    n600,
    n236,
    n345,
    n271,
    n235
  );


  xnor
  g561
  (
    n566,
    n188,
    n348,
    n295,
    n246
  );


  nor
  g562
  (
    n442,
    n185,
    n208,
    n341,
    n177
  );


  nor
  g563
  (
    n521,
    n205,
    n290,
    n199,
    n304
  );


  and
  g564
  (
    n545,
    n169,
    n202,
    n240,
    n218
  );


  and
  g565
  (
    n497,
    n174,
    n282,
    n344,
    n320
  );


  or
  g566
  (
    n570,
    n220,
    n267,
    n186,
    n372
  );


  nand
  g567
  (
    n589,
    n344,
    n234,
    n306,
    n348
  );


  nor
  g568
  (
    n453,
    n218,
    n338,
    n183,
    n242
  );


  nor
  g569
  (
    n511,
    n169,
    n302,
    n345,
    n340
  );


  nor
  g570
  (
    n524,
    n172,
    n307,
    n163,
    n313
  );


  xnor
  g571
  (
    n445,
    n326,
    n307,
    n379,
    n300
  );


  xnor
  g572
  (
    n611,
    n213,
    n260,
    n305,
    n291
  );


  nand
  g573
  (
    n422,
    n256,
    n360,
    n264,
    n354
  );


  xnor
  g574
  (
    n609,
    n361,
    n278,
    n164,
    n230
  );


  nand
  g575
  (
    n492,
    n198,
    n250,
    n344,
    n228
  );


  or
  g576
  (
    n534,
    n378,
    n202,
    n277,
    n199
  );


  xnor
  g577
  (
    n572,
    n375,
    n303,
    n212,
    n230
  );


  xor
  g578
  (
    n529,
    n293,
    n339,
    n327,
    n248
  );


  nor
  g579
  (
    n624,
    n224,
    n330,
    n232,
    n265
  );


  xor
  g580
  (
    n436,
    n328,
    n183,
    n160
  );


  nand
  g581
  (
    n580,
    n366,
    n194,
    n179,
    n269
  );


  nor
  g582
  (
    n494,
    n313,
    n293,
    n359,
    n202
  );


  or
  g583
  (
    n423,
    n329,
    n318,
    n325,
    n332
  );


  and
  g584
  (
    n552,
    n357,
    n197,
    n166,
    n224
  );


  xnor
  g585
  (
    n450,
    n268,
    n249,
    n357,
    n255
  );


  or
  g586
  (
    n598,
    n312,
    n316,
    n369,
    n343
  );


  xor
  g587
  (
    n539,
    n195,
    n228,
    n325,
    n356
  );


  nor
  g588
  (
    n587,
    n367,
    n254,
    n253,
    n300
  );


  nor
  g589
  (
    n555,
    n281,
    n277,
    n250,
    n265
  );


  and
  g590
  (
    n597,
    n307,
    n212,
    n229,
    n174
  );


  nor
  g591
  (
    n599,
    n373,
    n215,
    n283,
    n327
  );


  nor
  g592
  (
    n480,
    n236,
    n175,
    n323,
    n302
  );


  or
  g593
  (
    n414,
    n249,
    n313,
    n355,
    n276
  );


  xnor
  g594
  (
    n540,
    n270,
    n330,
    n273,
    n251
  );


  xor
  g595
  (
    n578,
    n329,
    n191,
    n369,
    n285
  );


  xor
  g596
  (
    KeyWire_0_26,
    n348,
    n271,
    n210,
    n156
  );


  nand
  g597
  (
    n663,
    n436,
    n544,
    n465,
    n415
  );


  xnor
  g598
  (
    n664,
    n623,
    n519,
    n515,
    n482
  );


  xnor
  g599
  (
    n631,
    n416,
    n518,
    n590,
    n539
  );


  or
  g600
  (
    n644,
    n597,
    n526,
    n452,
    n532
  );


  xnor
  g601
  (
    n630,
    n549,
    n506,
    n565,
    n466
  );


  xnor
  g602
  (
    n679,
    n592,
    n509,
    n445,
    n481
  );


  or
  g603
  (
    n676,
    n468,
    n496,
    n538,
    n475
  );


  xnor
  g604
  (
    n642,
    n479,
    n523,
    n494,
    n530
  );


  nand
  g605
  (
    n673,
    n531,
    n561,
    n507,
    n489
  );


  nor
  g606
  (
    n646,
    n424,
    n458,
    n497,
    n469
  );


  and
  g607
  (
    n669,
    n456,
    n533,
    n569,
    n484
  );


  xor
  g608
  (
    n668,
    n622,
    n541,
    n462,
    n520
  );


  or
  g609
  (
    n653,
    n624,
    n608,
    n459,
    n448
  );


  or
  g610
  (
    n651,
    n568,
    n614,
    n451,
    n610
  );


  nor
  g611
  (
    n677,
    n578,
    n609,
    n500,
    n429
  );


  xor
  g612
  (
    n635,
    n471,
    n557,
    n419,
    n405
  );


  and
  g613
  (
    n682,
    n583,
    n470,
    n463,
    n599
  );


  xor
  g614
  (
    n678,
    n612,
    n502,
    n461,
    n447
  );


  nor
  g615
  (
    n640,
    n426,
    n620,
    n553,
    n559
  );


  xor
  g616
  (
    n666,
    n534,
    n460,
    n488,
    n556
  );


  nor
  g617
  (
    n684,
    n495,
    n435,
    n499,
    n431
  );


  nor
  g618
  (
    n662,
    n472,
    n591,
    n414,
    n584
  );


  nor
  g619
  (
    n671,
    n564,
    n586,
    n453,
    n477
  );


  or
  g620
  (
    n649,
    n555,
    n404,
    n603,
    n483
  );


  xor
  g621
  (
    n661,
    n558,
    n587,
    n542,
    n487
  );


  or
  g622
  (
    n650,
    n516,
    n407,
    n574,
    n524
  );


  and
  g623
  (
    n629,
    n604,
    n464,
    n573,
    n449
  );


  xor
  g624
  (
    n638,
    n525,
    n517,
    n474,
    n430
  );


  xnor
  g625
  (
    KeyWire_0_3,
    n546,
    n606,
    n513,
    n601
  );


  nor
  g626
  (
    n659,
    n528,
    n594,
    n438,
    n563
  );


  nor
  g627
  (
    n665,
    n572,
    n410,
    n616,
    n476
  );


  nand
  g628
  (
    n658,
    n598,
    n444,
    n593,
    n570
  );


  xor
  g629
  (
    n674,
    n508,
    n403,
    n422,
    n537
  );


  and
  g630
  (
    n683,
    n413,
    n540,
    n440,
    n446
  );


  and
  g631
  (
    n634,
    n478,
    n432,
    n562,
    n560
  );


  or
  g632
  (
    n633,
    n535,
    n576,
    n600,
    n418
  );


  nor
  g633
  (
    n647,
    n441,
    n514,
    n579,
    n490
  );


  xor
  g634
  (
    n672,
    n433,
    n588,
    n437,
    n582
  );


  and
  g635
  (
    n645,
    n406,
    n420,
    n402,
    n522
  );


  xnor
  g636
  (
    n648,
    n617,
    n580,
    n485,
    n504
  );


  nor
  g637
  (
    n639,
    n548,
    n434,
    n411,
    n486
  );


  xnor
  g638
  (
    n660,
    n421,
    n552,
    n536,
    n625
  );


  xnor
  g639
  (
    n655,
    n501,
    n577,
    n529,
    n443
  );


  and
  g640
  (
    n632,
    n602,
    n605,
    n551,
    n595
  );


  nor
  g641
  (
    n654,
    n442,
    n457,
    n412,
    n427
  );


  xnor
  g642
  (
    n643,
    n521,
    n425,
    n511,
    n607
  );


  xnor
  g643
  (
    n657,
    n503,
    n547,
    n567,
    n512
  );


  or
  g644
  (
    n637,
    n543,
    n480,
    n423,
    n611
  );


  nand
  g645
  (
    n656,
    n571,
    n467,
    n498,
    n473
  );


  nand
  g646
  (
    n670,
    n505,
    n613,
    n596,
    n491
  );


  nor
  g647
  (
    n681,
    n409,
    n454,
    n408,
    n615
  );


  nor
  g648
  (
    n680,
    n618,
    n439,
    n589,
    n450
  );


  nand
  g649
  (
    n667,
    n545,
    n492,
    n510,
    n581
  );


  xnor
  g650
  (
    n675,
    n455,
    n575,
    n554,
    n493
  );


  nor
  g651
  (
    n652,
    n619,
    n527,
    n585,
    n566
  );


  xnor
  g652
  (
    n636,
    n621,
    n428,
    n417,
    n550
  );


  buf
  g653
  (
    n686,
    n631
  );


  buf
  g654
  (
    n688,
    n629
  );


  not
  g655
  (
    n692,
    n631
  );


  buf
  g656
  (
    n691,
    n629
  );


  nand
  g657
  (
    n685,
    n630,
    n633,
    n631
  );


  nand
  g658
  (
    n687,
    n630,
    n629,
    n633,
    n632
  );


  nand
  g659
  (
    n690,
    n630,
    n632,
    n633
  );


  xor
  g660
  (
    n689,
    n633,
    n629,
    n632,
    n630
  );


  buf
  g661
  (
    n693,
    n386
  );


  or
  g662
  (
    n695,
    n384,
    n686,
    n385,
    n383
  );


  xor
  g663
  (
    n702,
    n386,
    n384,
    n387
  );


  or
  g664
  (
    n699,
    n685,
    n388,
    n383,
    n385
  );


  nand
  g665
  (
    n700,
    n686,
    n386,
    n389
  );


  nand
  g666
  (
    n696,
    n687,
    n387,
    n388,
    n685
  );


  nand
  g667
  (
    n698,
    n383,
    n384,
    n686,
    n387
  );


  and
  g668
  (
    n701,
    n685,
    n686,
    n389,
    n383
  );


  xor
  g669
  (
    n694,
    n388,
    n385,
    n389
  );


  xor
  g670
  (
    n697,
    n388,
    n387,
    n685,
    n687
  );


  buf
  g671
  (
    n714,
    n694
  );


  buf
  g672
  (
    n705,
    n694
  );


  not
  g673
  (
    n703,
    n390
  );


  not
  g674
  (
    n712,
    n695
  );


  buf
  g675
  (
    n708,
    n693
  );


  buf
  g676
  (
    n707,
    n628
  );


  not
  g677
  (
    n706,
    n695
  );


  buf
  g678
  (
    n710,
    n390
  );


  xnor
  g679
  (
    n704,
    n626,
    n695,
    n390
  );


  and
  g680
  (
    n709,
    n695,
    n694,
    n693
  );


  or
  g681
  (
    n711,
    n627,
    n693
  );


  nor
  g682
  (
    n713,
    n694,
    n390,
    n389
  );


  nand
  g683
  (
    n715,
    n635,
    n703,
    n638
  );


  or
  g684
  (
    n720,
    n703,
    n640,
    n704
  );


  nor
  g685
  (
    n716,
    n704,
    n703,
    n639,
    n638
  );


  xnor
  g686
  (
    n721,
    n640,
    n636,
    n635,
    n634
  );


  xor
  g687
  (
    n717,
    n636,
    n635,
    n638,
    n639
  );


  nand
  g688
  (
    n723,
    n634,
    n637,
    n636,
    n635
  );


  or
  g689
  (
    n718,
    n639,
    n637,
    n634
  );


  nand
  g690
  (
    n722,
    n638,
    n637,
    n639,
    n705
  );


  or
  g691
  (
    n719,
    n634,
    n704,
    n636
  );


  and
  g692
  (
    n732,
    n715,
    n720,
    n689,
    n646
  );


  xor
  g693
  (
    n739,
    n718,
    n643,
    n691,
    n723
  );


  and
  g694
  (
    n728,
    n689,
    n645,
    n690
  );


  or
  g695
  (
    n727,
    n647,
    n647,
    n723,
    n687
  );


  or
  g696
  (
    n731,
    n644,
    n717,
    n648,
    n647
  );


  xor
  g697
  (
    n734,
    n722,
    n642,
    n690,
    n643
  );


  nand
  g698
  (
    KeyWire_0_30,
    n642,
    n716,
    n647,
    n721
  );


  xnor
  g699
  (
    n740,
    n642,
    n692,
    n691,
    n646
  );


  xnor
  g700
  (
    n736,
    n689,
    n723,
    n719,
    n687
  );


  xor
  g701
  (
    n730,
    n640,
    n646,
    n645,
    n648
  );


  xor
  g702
  (
    KeyWire_0_19,
    n689,
    n721,
    n643,
    n644
  );


  and
  g703
  (
    n726,
    n644,
    n648,
    n688
  );


  and
  g704
  (
    n725,
    n720,
    n722,
    n641,
    n691
  );


  xnor
  g705
  (
    n729,
    n648,
    n688,
    n646,
    n641
  );


  xor
  g706
  (
    n733,
    n642,
    n722,
    n645,
    n723
  );


  nand
  g707
  (
    n735,
    n690,
    n644,
    n722,
    n719
  );


  xor
  g708
  (
    n737,
    n641,
    n645,
    n643,
    n691
  );


  nor
  g709
  (
    n741,
    n649,
    n692,
    n688,
    n641
  );


  not
  g710
  (
    n806,
    n696
  );


  buf
  g711
  (
    n783,
    n740
  );


  buf
  g712
  (
    n755,
    n736
  );


  not
  g713
  (
    n793,
    n649
  );


  buf
  g714
  (
    n785,
    n735
  );


  not
  g715
  (
    n747,
    n697
  );


  not
  g716
  (
    n761,
    n393
  );


  buf
  g717
  (
    n805,
    n699
  );


  not
  g718
  (
    n762,
    n696
  );


  buf
  g719
  (
    n776,
    n650
  );


  buf
  g720
  (
    n787,
    n724
  );


  buf
  g721
  (
    n752,
    n701
  );


  buf
  g722
  (
    n758,
    n733
  );


  buf
  g723
  (
    n773,
    n702
  );


  buf
  g724
  (
    n763,
    n706
  );


  buf
  g725
  (
    n767,
    n692
  );


  buf
  g726
  (
    n743,
    n707
  );


  not
  g727
  (
    n750,
    n697
  );


  buf
  g728
  (
    n784,
    n727
  );


  buf
  g729
  (
    n742,
    n649
  );


  buf
  g730
  (
    n769,
    n697
  );


  not
  g731
  (
    n779,
    n730
  );


  not
  g732
  (
    n812,
    n739
  );


  not
  g733
  (
    n756,
    n707
  );


  buf
  g734
  (
    n789,
    n730
  );


  not
  g735
  (
    n780,
    n740
  );


  buf
  g736
  (
    n774,
    n727
  );


  buf
  g737
  (
    n775,
    n725
  );


  not
  g738
  (
    n777,
    n700
  );


  buf
  g739
  (
    n794,
    n730
  );


  not
  g740
  (
    n772,
    n698
  );


  buf
  g741
  (
    n749,
    n392
  );


  buf
  g742
  (
    n782,
    n729
  );


  buf
  g743
  (
    n791,
    n698
  );


  buf
  g744
  (
    n802,
    n732
  );


  buf
  g745
  (
    n803,
    n726
  );


  not
  g746
  (
    n801,
    n735
  );


  not
  g747
  (
    KeyWire_0_11,
    n698
  );


  buf
  g748
  (
    n744,
    n699
  );


  not
  g749
  (
    n766,
    n392
  );


  not
  g750
  (
    n808,
    n728
  );


  buf
  g751
  (
    n790,
    n737
  );


  not
  g752
  (
    n745,
    n729
  );


  not
  g753
  (
    n746,
    n740
  );


  buf
  g754
  (
    n811,
    n741
  );


  not
  g755
  (
    n813,
    n737
  );


  buf
  g756
  (
    n795,
    n705
  );


  not
  g757
  (
    n781,
    n731
  );


  buf
  g758
  (
    n748,
    n737
  );


  buf
  g759
  (
    n754,
    n728
  );


  buf
  g760
  (
    n798,
    n739
  );


  not
  g761
  (
    n753,
    n735
  );


  nor
  g762
  (
    n778,
    n734,
    n741,
    n729,
    n736
  );


  nand
  g763
  (
    n796,
    n726,
    n393,
    n706,
    n741
  );


  nand
  g764
  (
    n757,
    n731,
    n733,
    n707,
    n728
  );


  nor
  g765
  (
    n800,
    n725,
    n738,
    n727,
    n702
  );


  nor
  g766
  (
    n786,
    n649,
    n705,
    n734
  );


  xor
  g767
  (
    n770,
    n726,
    n725,
    n391
  );


  xnor
  g768
  (
    n799,
    n699,
    n739,
    n741,
    n738
  );


  nor
  g769
  (
    n751,
    n393,
    n392,
    n650,
    n701
  );


  nand
  g770
  (
    n760,
    n733,
    n733,
    n730,
    n728
  );


  nand
  g771
  (
    n759,
    n726,
    n724,
    n701,
    n727
  );


  xnor
  g772
  (
    n810,
    n391,
    n697,
    n707,
    n394
  );


  xnor
  g773
  (
    n804,
    n650,
    n732,
    n737,
    n740
  );


  xor
  g774
  (
    n792,
    n732,
    n700,
    n736,
    n701
  );


  xor
  g775
  (
    n807,
    n696,
    n698,
    n732,
    n393
  );


  xnor
  g776
  (
    n788,
    n734,
    n725,
    n731
  );


  xor
  g777
  (
    n797,
    n392,
    n699,
    n702,
    n692
  );


  xor
  g778
  (
    n764,
    n702,
    n706,
    n724
  );


  and
  g779
  (
    n768,
    n724,
    n729,
    n736,
    n696
  );


  nand
  g780
  (
    n765,
    n705,
    n738,
    n739,
    n391
  );


  nor
  g781
  (
    n809,
    n735,
    n700,
    n738
  );


  buf
  g782
  (
    n823,
    n745
  );


  not
  g783
  (
    n825,
    n744
  );


  buf
  g784
  (
    n821,
    n751
  );


  buf
  g785
  (
    n822,
    n749
  );


  not
  g786
  (
    n848,
    n746
  );


  not
  g787
  (
    n817,
    n742
  );


  buf
  g788
  (
    n843,
    n743
  );


  buf
  g789
  (
    n831,
    n748
  );


  buf
  g790
  (
    n814,
    n749
  );


  not
  g791
  (
    n840,
    n751
  );


  buf
  g792
  (
    n845,
    n748
  );


  not
  g793
  (
    n828,
    n750
  );


  not
  g794
  (
    n836,
    n749
  );


  buf
  g795
  (
    n844,
    n746
  );


  buf
  g796
  (
    n824,
    n750
  );


  not
  g797
  (
    n832,
    n749
  );


  buf
  g798
  (
    n849,
    n751
  );


  not
  g799
  (
    n842,
    n745
  );


  buf
  g800
  (
    n851,
    n744
  );


  not
  g801
  (
    KeyWire_0_20,
    n742
  );


  not
  g802
  (
    n852,
    n743
  );


  buf
  g803
  (
    n829,
    n750
  );


  not
  g804
  (
    n827,
    n746
  );


  buf
  g805
  (
    n830,
    n750
  );


  buf
  g806
  (
    n847,
    n746
  );


  buf
  g807
  (
    n846,
    n748
  );


  not
  g808
  (
    n850,
    n748
  );


  not
  g809
  (
    n834,
    n744
  );


  not
  g810
  (
    n820,
    n747
  );


  buf
  g811
  (
    n839,
    n747
  );


  buf
  g812
  (
    n837,
    n742
  );


  buf
  g813
  (
    n835,
    n743
  );


  buf
  g814
  (
    n838,
    n751
  );


  buf
  g815
  (
    n841,
    n745
  );


  not
  g816
  (
    KeyWire_0_31,
    n747
  );


  buf
  g817
  (
    n815,
    n742
  );


  not
  g818
  (
    n819,
    n744
  );


  not
  g819
  (
    n826,
    n745
  );


  not
  g820
  (
    n816,
    n747
  );


  not
  g821
  (
    n853,
    n743
  );


  buf
  g822
  (
    n863,
    n814
  );


  not
  g823
  (
    n856,
    n815
  );


  not
  g824
  (
    n859,
    n815
  );


  buf
  g825
  (
    n864,
    n814
  );


  not
  g826
  (
    n855,
    n814
  );


  buf
  g827
  (
    n862,
    n816
  );


  not
  g828
  (
    n860,
    n815
  );


  not
  g829
  (
    n858,
    n816
  );


  not
  g830
  (
    n857,
    n815
  );


  not
  g831
  (
    n861,
    n814
  );


  buf
  g832
  (
    n854,
    n816
  );


  not
  g833
  (
    n882,
    n864
  );


  not
  g834
  (
    n868,
    n651
  );


  buf
  g835
  (
    n879,
    n862
  );


  buf
  g836
  (
    n874,
    n653
  );


  and
  g837
  (
    n865,
    n653,
    n822
  );


  and
  g838
  (
    n883,
    n821,
    n820,
    n655,
    n650
  );


  nor
  g839
  (
    n878,
    n654,
    n818,
    n856
  );


  or
  g840
  (
    n871,
    n394,
    n821,
    n653,
    n652
  );


  and
  g841
  (
    n870,
    n861,
    n651,
    n823,
    n394
  );


  or
  g842
  (
    n881,
    n655,
    n863,
    n817,
    n860
  );


  nor
  g843
  (
    n880,
    n862,
    n819,
    n864
  );


  and
  g844
  (
    n877,
    n823,
    n819,
    n818,
    n654
  );


  or
  g845
  (
    n869,
    n821,
    n820,
    n823,
    n816
  );


  xor
  g846
  (
    n867,
    n855,
    n822,
    n860,
    n652
  );


  nor
  g847
  (
    n875,
    n863,
    n862,
    n394,
    n864
  );


  xor
  g848
  (
    n885,
    n859,
    n655,
    n817,
    n854
  );


  xnor
  g849
  (
    KeyWire_0_27,
    n864,
    n651,
    n817,
    n824
  );


  and
  g850
  (
    n866,
    n654,
    n653,
    n863,
    n857
  );


  and
  g851
  (
    n872,
    n823,
    n858,
    n820,
    n654
  );


  nor
  g852
  (
    n876,
    n818,
    n820,
    n819,
    n652
  );


  xnor
  g853
  (
    n873,
    n863,
    n821,
    n861,
    n822
  );


  and
  g854
  (
    n884,
    n652,
    n817,
    n651,
    n862
  );


  nand
  g855
  (
    n901,
    n886,
    n710,
    n787,
    n794
  );


  or
  g856
  (
    n897,
    n790,
    n777,
    n786,
    n782
  );


  or
  g857
  (
    n952,
    n807,
    n764,
    n795,
    n783
  );


  or
  g858
  (
    n904,
    n865,
    n759,
    n877,
    n778
  );


  nor
  g859
  (
    n958,
    n802,
    n800,
    n791,
    n776
  );


  nor
  g860
  (
    n931,
    n870,
    n799,
    n801,
    n787
  );


  xnor
  g861
  (
    n938,
    n809,
    n789,
    n782,
    n759
  );


  nor
  g862
  (
    n949,
    n764,
    n758,
    n760,
    n762
  );


  nor
  g863
  (
    n922,
    n793,
    n796,
    n885,
    n765
  );


  nand
  g864
  (
    n955,
    n765,
    n791,
    n795,
    n811
  );


  or
  g865
  (
    n917,
    n755,
    n871,
    n795,
    n774
  );


  xor
  g866
  (
    n926,
    n790,
    n880,
    n812,
    n781
  );


  nor
  g867
  (
    n932,
    n868,
    n773,
    n869,
    n800
  );


  and
  g868
  (
    n909,
    n804,
    n867,
    n810,
    n753
  );


  or
  g869
  (
    n950,
    n874,
    n871,
    n868,
    n656
  );


  nand
  g870
  (
    n905,
    n779,
    n870,
    n759,
    n808
  );


  nor
  g871
  (
    n920,
    n785,
    n789,
    n879,
    n781
  );


  xor
  g872
  (
    n896,
    n876,
    n787,
    n777,
    n766
  );


  nor
  g873
  (
    n889,
    n774,
    n776,
    n878,
    n800
  );


  nor
  g874
  (
    n943,
    n656,
    n881,
    n786,
    n805
  );


  nor
  g875
  (
    n954,
    n792,
    n872,
    n754,
    n876
  );


  nand
  g876
  (
    n972,
    n875,
    n869,
    n787,
    n786
  );


  xor
  g877
  (
    n892,
    n709,
    n753,
    n773,
    n757
  );


  nand
  g878
  (
    n970,
    n764,
    n799,
    n708,
    n779
  );


  and
  g879
  (
    n966,
    n871,
    n784,
    n873,
    n879
  );


  or
  g880
  (
    n891,
    n769,
    n813,
    n782,
    n794
  );


  and
  g881
  (
    n934,
    n763,
    n754,
    n772,
    n804
  );


  xor
  g882
  (
    n968,
    n797,
    n753,
    n769,
    n771
  );


  nor
  g883
  (
    n903,
    n797,
    n775,
    n792,
    n794
  );


  xnor
  g884
  (
    n924,
    n803,
    n771,
    n885
  );


  nand
  g885
  (
    KeyWire_0_1,
    n811,
    n760,
    n764,
    n768
  );


  nand
  g886
  (
    n907,
    n765,
    n709,
    n799,
    n763
  );


  nor
  g887
  (
    n914,
    n762,
    n798,
    n753,
    n708
  );


  nor
  g888
  (
    n916,
    n804,
    n755,
    n865,
    n772
  );


  xor
  g889
  (
    n937,
    n754,
    n873,
    n811
  );


  nand
  g890
  (
    n939,
    n875,
    n872,
    n886,
    n808
  );


  xor
  g891
  (
    n963,
    n877,
    n882,
    n796,
    n767
  );


  xnor
  g892
  (
    n967,
    n756,
    n773,
    n870,
    n752
  );


  xor
  g893
  (
    n894,
    n874,
    n789,
    n790,
    n762
  );


  or
  g894
  (
    n887,
    n766,
    n761,
    n802,
    n756
  );


  xor
  g895
  (
    n945,
    n880,
    n783,
    n777,
    n809
  );


  and
  g896
  (
    n890,
    n866,
    n879,
    n776,
    n780
  );


  and
  g897
  (
    n911,
    n792,
    n797,
    n879,
    n802
  );


  nor
  g898
  (
    n971,
    n656,
    n771,
    n783,
    n760
  );


  and
  g899
  (
    n960,
    n884,
    n809,
    n807,
    n878
  );


  nand
  g900
  (
    n918,
    n778,
    n807,
    n873,
    n882
  );


  and
  g901
  (
    n953,
    n756,
    n875,
    n775,
    n793
  );


  xnor
  g902
  (
    n940,
    n874,
    n808,
    n801,
    n878
  );


  nor
  g903
  (
    n973,
    n807,
    n768,
    n754,
    n866
  );


  nor
  g904
  (
    n956,
    n757,
    n804,
    n761,
    n870
  );


  xnor
  g905
  (
    n948,
    n770,
    n775,
    n798,
    n771
  );


  or
  g906
  (
    n936,
    n781,
    n757,
    n785,
    n813
  );


  xnor
  g907
  (
    n965,
    n776,
    n805,
    n772,
    n811
  );


  and
  g908
  (
    n888,
    n875,
    n783,
    n877,
    n767
  );


  nor
  g909
  (
    n908,
    n876,
    n780,
    n777,
    n784
  );


  xnor
  g910
  (
    n951,
    n869,
    n781,
    n883,
    n865
  );


  xor
  g911
  (
    n915,
    n757,
    n762,
    n884,
    n760
  );


  xnor
  g912
  (
    n946,
    n755,
    n770,
    n761,
    n752
  );


  xor
  g913
  (
    n959,
    n883,
    n769,
    n798,
    n778
  );


  or
  g914
  (
    n923,
    n786,
    n881,
    n761
  );


  or
  g915
  (
    n900,
    n793,
    n769,
    n880,
    n708
  );


  xor
  g916
  (
    n929,
    n765,
    n866,
    n795,
    n868
  );


  xnor
  g917
  (
    n942,
    n798,
    n812,
    n791,
    n770
  );


  nor
  g918
  (
    n893,
    n768,
    n867,
    n801,
    n752
  );


  nand
  g919
  (
    n925,
    n809,
    n763,
    n880,
    n758
  );


  nor
  g920
  (
    n919,
    n883,
    n805,
    n806
  );


  nand
  g921
  (
    n930,
    n884,
    n867,
    n773,
    n881
  );


  nand
  g922
  (
    n935,
    n766,
    n788,
    n810,
    n784
  );


  nor
  g923
  (
    n910,
    n800,
    n871,
    n866,
    n882
  );


  xor
  g924
  (
    n961,
    n886,
    n805,
    n756,
    n709
  );


  or
  g925
  (
    n933,
    n812,
    n883,
    n755,
    n806
  );


  or
  g926
  (
    n962,
    n788,
    n708,
    n758,
    n810
  );


  xor
  g927
  (
    n921,
    n759,
    n758,
    n867,
    n788
  );


  and
  g928
  (
    n928,
    n793,
    n785,
    n882,
    n774
  );


  xnor
  g929
  (
    n912,
    n874,
    n655,
    n797,
    n778
  );


  and
  g930
  (
    n906,
    n766,
    n785,
    n876,
    n782
  );


  nand
  g931
  (
    n902,
    n780,
    n813,
    n767,
    n812
  );


  xnor
  g932
  (
    n969,
    n865,
    n801,
    n772,
    n779
  );


  xnor
  g933
  (
    n899,
    n808,
    n763,
    n752,
    n803
  );


  xnor
  g934
  (
    n898,
    n877,
    n792,
    n775,
    n872
  );


  xnor
  g935
  (
    n964,
    n796,
    n885,
    n884,
    n802
  );


  nor
  g936
  (
    n944,
    n770,
    n767,
    n779,
    n780
  );


  xnor
  g937
  (
    n957,
    n878,
    n872,
    n788,
    n810
  );


  xnor
  g938
  (
    n947,
    n789,
    n806,
    n796,
    n709
  );


  xor
  g939
  (
    n927,
    n868,
    n774,
    n869,
    n794
  );


  and
  g940
  (
    n941,
    n791,
    n768,
    n790,
    n799
  );


  nand
  g941
  (
    n895,
    n886,
    n803,
    n784
  );


  or
  g942
  (
    n977,
    n887,
    n893,
    n896,
    n889
  );


  or
  g943
  (
    n975,
    n900,
    n896,
    n895
  );


  and
  g944
  (
    n978,
    n894,
    n897,
    n887,
    n893
  );


  nor
  g945
  (
    n980,
    n895,
    n895,
    n898,
    n900
  );


  nor
  g946
  (
    n985,
    n897,
    n892,
    n900,
    n893
  );


  nand
  g947
  (
    n984,
    n892,
    n894,
    n895,
    n889
  );


  nand
  g948
  (
    n976,
    n889,
    n889,
    n898,
    n887
  );


  xor
  g949
  (
    n981,
    n888,
    n891,
    n899
  );


  xnor
  g950
  (
    n987,
    n898,
    n894,
    n891,
    n888
  );


  nor
  g951
  (
    KeyWire_0_4,
    n887,
    n891,
    n898,
    n888
  );


  nor
  g952
  (
    n986,
    n890,
    n900,
    n897
  );


  xnor
  g953
  (
    n982,
    n888,
    n896,
    n899
  );


  nor
  g954
  (
    n979,
    n893,
    n890
  );


  nand
  g955
  (
    n974,
    n899,
    n894,
    n892
  );


  not
  g956
  (
    n988,
    n986
  );


  buf
  g957
  (
    n990,
    n984
  );


  not
  g958
  (
    n989,
    n985
  );


  buf
  g959
  (
    n991,
    n987
  );


  not
  g960
  (
    n992,
    n658
  );


  not
  g961
  (
    n995,
    n991
  );


  xnor
  g962
  (
    n996,
    n658,
    n657
  );


  and
  g963
  (
    KeyWire_0_2,
    n990,
    n656,
    n657
  );


  xnor
  g964
  (
    n994,
    n989,
    n988,
    n991,
    n658
  );


  xor
  g965
  (
    n1006,
    n906,
    n902,
    n907
  );


  xor
  g966
  (
    n1004,
    n903,
    n994,
    n902
  );


  and
  g967
  (
    n998,
    n902,
    n992,
    n908,
    n903
  );


  nor
  g968
  (
    n1000,
    n993,
    n992,
    n904,
    n901
  );


  or
  g969
  (
    n1005,
    n905,
    n903,
    n993
  );


  xnor
  g970
  (
    n1002,
    n904,
    n906,
    n905
  );


  xnor
  g971
  (
    n999,
    n903,
    n908,
    n992,
    n905
  );


  xor
  g972
  (
    n997,
    n905,
    n901,
    n907
  );


  xnor
  g973
  (
    n1001,
    n992,
    n993,
    n904,
    n907
  );


  nand
  g974
  (
    n1003,
    n907,
    n904,
    n901,
    n906
  );


  not
  g975
  (
    n1014,
    n998
  );


  buf
  g976
  (
    n1025,
    n999
  );


  not
  g977
  (
    n1029,
    n1001
  );


  buf
  g978
  (
    n1026,
    n396
  );


  buf
  g979
  (
    n1012,
    n1000
  );


  buf
  g980
  (
    n1032,
    n1002
  );


  buf
  g981
  (
    n1033,
    n1000
  );


  buf
  g982
  (
    n1024,
    n998
  );


  buf
  g983
  (
    n1008,
    n998
  );


  buf
  g984
  (
    n1018,
    n1001
  );


  not
  g985
  (
    n1023,
    n908
  );


  not
  g986
  (
    n1021,
    n1000
  );


  buf
  g987
  (
    n1007,
    n1000
  );


  buf
  g988
  (
    n1034,
    n1003
  );


  not
  g989
  (
    n1015,
    n911
  );


  buf
  g990
  (
    n1017,
    n997
  );


  not
  g991
  (
    n1028,
    n1003
  );


  buf
  g992
  (
    n1031,
    n908
  );


  buf
  g993
  (
    n1011,
    n910
  );


  xnor
  g994
  (
    n1013,
    n997,
    n998,
    n909
  );


  xnor
  g995
  (
    n1009,
    n909,
    n911,
    n912,
    n1002
  );


  nand
  g996
  (
    n1016,
    n1004,
    n999,
    n909,
    n912
  );


  xor
  g997
  (
    n1020,
    n659,
    n1001,
    n395,
    n396
  );


  nand
  g998
  (
    n1022,
    n911,
    n909,
    n999
  );


  nand
  g999
  (
    n1010,
    n1002,
    n1003,
    n396,
    n910
  );


  xor
  g1000
  (
    n1035,
    n912,
    n997,
    n395,
    n396
  );


  xor
  g1001
  (
    n1027,
    n395,
    n910,
    n1003
  );


  nor
  g1002
  (
    n1019,
    n397,
    n395,
    n659,
    n997
  );


  or
  g1003
  (
    n1030,
    n1002,
    n397,
    n1001,
    n911
  );


  nand
  g1004
  (
    n1052,
    n1013,
    n1027,
    n1031
  );


  nand
  g1005
  (
    n1044,
    n398,
    n400,
    n401
  );


  nor
  g1006
  (
    n1041,
    n1034,
    n1012,
    n1032
  );


  xnor
  g1007
  (
    n1039,
    n1024,
    n399,
    n1031
  );


  or
  g1008
  (
    n1049,
    n1025,
    n1035,
    n1032
  );


  and
  g1009
  (
    n1053,
    n399,
    n398,
    n400
  );


  nand
  g1010
  (
    n1055,
    n1023,
    n401,
    n1010
  );


  and
  g1011
  (
    n1043,
    n401,
    n1031,
    n1029
  );


  xnor
  g1012
  (
    n1054,
    n1034,
    n1030,
    n1033
  );


  xnor
  g1013
  (
    n1040,
    n1034,
    n397,
    n1008
  );


  nand
  g1014
  (
    n1051,
    n1016,
    n1035
  );


  or
  g1015
  (
    n1042,
    n1031,
    n398,
    n1033
  );


  xnor
  g1016
  (
    n1045,
    n401,
    n1007,
    n399
  );


  xnor
  g1017
  (
    n1036,
    n399,
    n1032
  );


  nor
  g1018
  (
    n1038,
    n1011,
    n400
  );


  nand
  g1019
  (
    n1048,
    n1034,
    n1014,
    n398
  );


  and
  g1020
  (
    n1050,
    n1015,
    n1035,
    n1033
  );


  or
  g1021
  (
    n1046,
    n1019,
    n397,
    n1020
  );


  nor
  g1022
  (
    n1037,
    n1018,
    n1033,
    n1017,
    n1021
  );


  xnor
  g1023
  (
    n1047,
    n1009,
    n1026,
    n1022,
    n1028
  );


  nor
  g1024
  (
    n1078,
    n674,
    n671,
    n1039,
    n666
  );


  nor
  g1025
  (
    n1068,
    n678,
    n669,
    n670,
    n664
  );


  xor
  g1026
  (
    n1088,
    n676,
    n1048,
    n667,
    n671
  );


  xnor
  g1027
  (
    n1075,
    n663,
    n676,
    n668
  );


  nand
  g1028
  (
    n1083,
    n1048,
    n1037,
    n677,
    n1039
  );


  or
  g1029
  (
    n1071,
    n675,
    n1047,
    n1040,
    n680
  );


  nand
  g1030
  (
    n1073,
    n668,
    n678,
    n1042,
    n1047
  );


  nand
  g1031
  (
    n1082,
    n680,
    n1046,
    n660,
    n1036
  );


  or
  g1032
  (
    n1077,
    n659,
    n670,
    n1038
  );


  xnor
  g1033
  (
    n1069,
    n1043,
    n669,
    n677,
    n679
  );


  or
  g1034
  (
    n1074,
    n1043,
    n665,
    n663,
    n674
  );


  nor
  g1035
  (
    n1059,
    n669,
    n678,
    n671,
    n676
  );


  and
  g1036
  (
    n1085,
    n1040,
    n660,
    n681,
    n667
  );


  and
  g1037
  (
    n1086,
    n678,
    n1037,
    n673,
    n679
  );


  nand
  g1038
  (
    n1065,
    n665,
    n1045,
    n1041,
    n1042
  );


  xnor
  g1039
  (
    n1062,
    n659,
    n674,
    n673,
    n1038
  );


  nand
  g1040
  (
    n1076,
    n663,
    n675,
    n660,
    n1039
  );


  xor
  g1041
  (
    n1087,
    n661,
    n664,
    n668,
    n1046
  );


  nor
  g1042
  (
    n1072,
    n662,
    n661,
    n1040,
    n664
  );


  nor
  g1043
  (
    n1064,
    n673,
    n662,
    n1036,
    n661
  );


  xnor
  g1044
  (
    n1058,
    n1040,
    n679,
    n663,
    n1036
  );


  and
  g1045
  (
    n1056,
    n674,
    n665,
    n667,
    n662
  );


  or
  g1046
  (
    n1081,
    n1041,
    n670,
    n675,
    n660
  );


  xor
  g1047
  (
    n1066,
    n667,
    n1047,
    n681,
    n669
  );


  xnor
  g1048
  (
    n1090,
    n672,
    n1047,
    n1042,
    n671
  );


  nor
  g1049
  (
    n1084,
    n1045,
    n1036,
    n1037,
    n666
  );


  or
  g1050
  (
    n1079,
    n680,
    n1044,
    n1037,
    n679
  );


  xor
  g1051
  (
    n1061,
    n676,
    n1041,
    n681,
    n677
  );


  nor
  g1052
  (
    n1070,
    n662,
    n1045,
    n1043,
    n1046
  );


  nand
  g1053
  (
    n1057,
    n666,
    n672
  );


  or
  g1054
  (
    n1067,
    n664,
    n670,
    n681,
    n1044
  );


  xnor
  g1055
  (
    n1089,
    n1043,
    n1046,
    n1044,
    n1039
  );


  and
  g1056
  (
    n1060,
    n680,
    n1041,
    n1042,
    n1044
  );


  nand
  g1057
  (
    n1063,
    n675,
    n677,
    n1038,
    n1045
  );


  and
  g1058
  (
    n1080,
    n666,
    n673,
    n661,
    n665
  );


  nor
  g1059
  (
    n1091,
    n1056,
    n682
  );


  buf
  g1060
  (
    n1092,
    n1091
  );


  nor
  g1061
  (
    n1094,
    n1049,
    n1092
  );


  nand
  g1062
  (
    n1093,
    n1049,
    n1048
  );


  not
  g1063
  (
    n1097,
    n1094
  );


  buf
  g1064
  (
    KeyWire_0_8,
    n682
  );


  nand
  g1065
  (
    KeyWire_0_9,
    n1094,
    n1093
  );


  not
  g1066
  (
    n1098,
    n1096
  );


  buf
  g1067
  (
    n1099,
    n1097
  );


  xnor
  g1068
  (
    n1100,
    n1098,
    n1099
  );


  or
  g1069
  (
    n1102,
    n683,
    n1100,
    n912,
    n913
  );


  nand
  g1070
  (
    n1101,
    n1100,
    n683,
    n913
  );


  or
  g1071
  (
    n1103,
    n1101,
    n1102
  );


  not
  g1072
  (
    n1106,
    n1103
  );


  buf
  g1073
  (
    n1105,
    n1103
  );


  xnor
  g1074
  (
    n1104,
    n1099,
    n1103
  );


  xor
  g1075
  (
    n1108,
    n915,
    n915,
    n916,
    n913
  );


  nor
  g1076
  (
    n1107,
    n915,
    n913,
    n1105,
    n1106
  );


  xnor
  g1077
  (
    n1109,
    n914,
    n914,
    n915,
    n1104
  );


  nand
  g1078
  (
    n1110,
    n914,
    n914,
    n1106,
    n916
  );


  xor
  g1079
  (
    n1111,
    n918,
    n917,
    n916
  );


  nand
  g1080
  (
    n1113,
    n917,
    n918,
    n1108
  );


  or
  g1081
  (
    n1114,
    n917,
    n919,
    n916,
    n1107
  );


  and
  g1082
  (
    n1112,
    n918,
    n1109,
    n919,
    n1110
  );


  nor
  g1083
  (
    n1119,
    n1112,
    n1114,
    n919
  );


  xor
  g1084
  (
    n1118,
    n922,
    n1111,
    n1114
  );


  or
  g1085
  (
    n1115,
    n920,
    n920,
    n921,
    n1113
  );


  xnor
  g1086
  (
    n1117,
    n922,
    n920,
    n919
  );


  nor
  g1087
  (
    n1116,
    n922,
    n921
  );


  nand
  g1088
  (
    n1122,
    n830,
    n828,
    n1050,
    n994
  );


  and
  g1089
  (
    n1139,
    n827,
    n825,
    n1116,
    n1050
  );


  nor
  g1090
  (
    n1132,
    n1117,
    n995,
    n1118
  );


  nand
  g1091
  (
    n1137,
    n1116,
    n923,
    n1118,
    n830
  );


  nor
  g1092
  (
    KeyWire_0_23,
    n995,
    n1049,
    n826,
    n830
  );


  xnor
  g1093
  (
    n1124,
    n828,
    n824,
    n1051
  );


  and
  g1094
  (
    n1136,
    n1119,
    n828,
    n996,
    n829
  );


  nand
  g1095
  (
    n1123,
    n1115,
    n996,
    n711,
    n1050
  );


  or
  g1096
  (
    n1127,
    n924,
    n1116,
    n994,
    n710
  );


  xor
  g1097
  (
    n1131,
    n1115,
    n710,
    n1117,
    n826
  );


  nor
  g1098
  (
    n1128,
    n1119,
    n1050,
    n996,
    n825
  );


  xor
  g1099
  (
    n1133,
    n827,
    n923,
    n1116
  );


  xor
  g1100
  (
    n1138,
    n1115,
    n826,
    n829
  );


  and
  g1101
  (
    n1134,
    n923,
    n827,
    n922
  );


  xor
  g1102
  (
    n1130,
    n924,
    n831,
    n825,
    n828
  );


  or
  g1103
  (
    n1129,
    n830,
    n711,
    n1117,
    n1119
  );


  xnor
  g1104
  (
    n1126,
    n1119,
    n924,
    n1117,
    n826
  );


  nor
  g1105
  (
    n1135,
    n1118,
    n829,
    n710,
    n1049
  );


  nor
  g1106
  (
    n1125,
    n825,
    n996,
    n813,
    n824
  );


  xnor
  g1107
  (
    n1120,
    n1115,
    n995,
    n711
  );


  or
  g1108
  (
    n1165,
    n932,
    n1131,
    n1137,
    n1124
  );


  xor
  g1109
  (
    n1148,
    n1136,
    n932,
    n1127,
    n1120
  );


  and
  g1110
  (
    n1167,
    n1132,
    n926,
    n934
  );


  xnor
  g1111
  (
    n1143,
    n932,
    n933,
    n1122,
    n931
  );


  nor
  g1112
  (
    n1169,
    n1128,
    n932,
    n1132,
    n927
  );


  and
  g1113
  (
    n1166,
    n1124,
    n1138,
    n1128,
    n927
  );


  and
  g1114
  (
    n1161,
    n1125,
    n924,
    n1122,
    n1127
  );


  nor
  g1115
  (
    n1145,
    n1137,
    n1125,
    n1138,
    n1129
  );


  nor
  g1116
  (
    n1141,
    n930,
    n1125,
    n1134,
    n1136
  );


  nand
  g1117
  (
    n1144,
    n1126,
    n1123,
    n934,
    n1139
  );


  and
  g1118
  (
    n1168,
    n1121,
    n1132,
    n1124,
    n1135
  );


  nand
  g1119
  (
    n1146,
    n925,
    n1127,
    n1122,
    n929
  );


  nand
  g1120
  (
    n1142,
    n934,
    n1133,
    n930,
    n1128
  );


  nor
  g1121
  (
    n1140,
    n1135,
    n1129,
    n1138,
    n1133
  );


  and
  g1122
  (
    n1164,
    n1120,
    n1127,
    n1134,
    n1138
  );


  and
  g1123
  (
    n1159,
    n1131,
    n1130,
    n925,
    n1128
  );


  xor
  g1124
  (
    n1158,
    n1132,
    n1137,
    n929,
    n1129
  );


  nor
  g1125
  (
    n1155,
    n1124,
    n1139,
    n1121,
    n1135
  );


  nand
  g1126
  (
    n1157,
    n928,
    n1136,
    n931,
    n1125
  );


  xor
  g1127
  (
    n1152,
    n1130,
    n1123,
    n928
  );


  or
  g1128
  (
    n1156,
    n1130,
    n928,
    n1121,
    n925
  );


  xnor
  g1129
  (
    n1151,
    n1139,
    n1120,
    n1123,
    n1126
  );


  xor
  g1130
  (
    n1149,
    n931,
    n1131,
    n1135,
    n1137
  );


  xor
  g1131
  (
    n1150,
    n927,
    n1122,
    n1126,
    n931
  );


  or
  g1132
  (
    n1153,
    n928,
    n934,
    n1133,
    n933
  );


  nand
  g1133
  (
    n1147,
    n933,
    n933,
    n929,
    n1133
  );


  xor
  g1134
  (
    n1160,
    n1121,
    n1131,
    n930,
    n1134
  );


  xor
  g1135
  (
    n1162,
    n930,
    n1120,
    n925,
    n1129
  );


  xor
  g1136
  (
    n1163,
    n1130,
    n926,
    n929
  );


  xnor
  g1137
  (
    n1154,
    n1126,
    n1136,
    n1134,
    n927
  );


  or
  g1138
  (
    n1170,
    n1094,
    n939,
    n937,
    n714
  );


  xnor
  g1139
  (
    n1179,
    n1152,
    n714,
    n938,
    n711
  );


  nand
  g1140
  (
    n1172,
    n683,
    n936,
    n939,
    n935
  );


  nand
  g1141
  (
    n1178,
    n1150,
    n712,
    n938
  );


  xnor
  g1142
  (
    n1171,
    n1149,
    n712,
    n936,
    n935
  );


  nor
  g1143
  (
    n1180,
    n1146,
    n1148,
    n684,
    n1144
  );


  or
  g1144
  (
    n1181,
    n1140,
    n1143,
    n713,
    n939
  );


  nor
  g1145
  (
    n1182,
    n938,
    n1147,
    n684,
    n939
  );


  or
  g1146
  (
    n1174,
    n1145,
    n1142,
    n937,
    n1151
  );


  and
  g1147
  (
    n1177,
    n713,
    n937,
    n936,
    n714
  );


  xor
  g1148
  (
    n1173,
    n937,
    n713,
    n938,
    n684
  );


  or
  g1149
  (
    n1176,
    n1141,
    n1094,
    n712,
    n935
  );


  nor
  g1150
  (
    n1175,
    n684,
    n713,
    n936,
    n935
  );


  not
  g1151
  (
    n1201,
    n1174
  );


  buf
  g1152
  (
    n1191,
    n1180
  );


  buf
  g1153
  (
    n1195,
    n1174
  );


  not
  g1154
  (
    n1219,
    n1173
  );


  not
  g1155
  (
    n1210,
    n941
  );


  buf
  g1156
  (
    n1189,
    n1179
  );


  buf
  g1157
  (
    n1207,
    n1182
  );


  not
  g1158
  (
    n1193,
    n940
  );


  buf
  g1159
  (
    n1213,
    n945
  );


  buf
  g1160
  (
    n1185,
    n1175
  );


  not
  g1161
  (
    n1209,
    n1172
  );


  buf
  g1162
  (
    n1206,
    n942
  );


  not
  g1163
  (
    n1184,
    n944
  );


  not
  g1164
  (
    n1183,
    n943
  );


  buf
  g1165
  (
    n1208,
    n943
  );


  not
  g1166
  (
    n1188,
    n1173
  );


  not
  g1167
  (
    n1196,
    n1170
  );


  not
  g1168
  (
    n1214,
    n1175
  );


  not
  g1169
  (
    n1194,
    n1170
  );


  buf
  g1170
  (
    n1203,
    n1179
  );


  not
  g1171
  (
    n1216,
    n1172
  );


  not
  g1172
  (
    n1218,
    n940
  );


  buf
  g1173
  (
    n1211,
    n1181
  );


  not
  g1174
  (
    n1204,
    n1174
  );


  buf
  g1175
  (
    n1217,
    n941
  );


  xnor
  g1176
  (
    n1190,
    n944,
    n1182,
    n1173
  );


  or
  g1177
  (
    n1215,
    n1176,
    n1177,
    n1175,
    n1178
  );


  or
  g1178
  (
    n1186,
    n1178,
    n945,
    n1171,
    n1176
  );


  nor
  g1179
  (
    n1202,
    n1178,
    n1179,
    n1175
  );


  and
  g1180
  (
    n1197,
    n1170,
    n1170,
    n1181,
    n1176
  );


  xor
  g1181
  (
    n1187,
    n943,
    n944,
    n1178,
    n940
  );


  or
  g1182
  (
    n1220,
    n1171,
    n1181,
    n1182,
    n941
  );


  or
  g1183
  (
    n1198,
    n1176,
    n945,
    n1172,
    n1182
  );


  nand
  g1184
  (
    n1192,
    n945,
    n1171,
    n1173,
    n1177
  );


  xnor
  g1185
  (
    n1200,
    n940,
    n1180,
    n941,
    n1171
  );


  xnor
  g1186
  (
    n1199,
    n943,
    n1181,
    n1177,
    n1180
  );


  xnor
  g1187
  (
    n1212,
    n942,
    n1172,
    n1177,
    n1180
  );


  nor
  g1188
  (
    n1205,
    n1174,
    n944,
    n942
  );


  nor
  g1189
  (
    n1243,
    n1207,
    n1198,
    n971,
    n956
  );


  or
  g1190
  (
    n1233,
    n948,
    n952,
    n946,
    n955
  );


  and
  g1191
  (
    n1248,
    n950,
    n970,
    n958,
    n949
  );


  nand
  g1192
  (
    n1244,
    n957,
    n952,
    n954
  );


  or
  g1193
  (
    n1253,
    n964,
    n1188,
    n1193,
    n962
  );


  nand
  g1194
  (
    n1242,
    n963,
    n967,
    n960,
    n1212
  );


  xnor
  g1195
  (
    n1240,
    n959,
    n964,
    n969,
    n946
  );


  xnor
  g1196
  (
    n1250,
    n972,
    n1195,
    n1200,
    n961
  );


  xnor
  g1197
  (
    n1257,
    n949,
    n972,
    n950,
    n958
  );


  or
  g1198
  (
    n1246,
    n960,
    n1210,
    n953,
    n968
  );


  xor
  g1199
  (
    n1254,
    n968,
    n965,
    n972,
    n1206
  );


  or
  g1200
  (
    n1230,
    n954,
    n1213,
    n969,
    n950
  );


  xnor
  g1201
  (
    n1229,
    n960,
    n1219,
    n947,
    n954
  );


  xnor
  g1202
  (
    n1235,
    n947,
    n969,
    n966,
    n959
  );


  xnor
  g1203
  (
    n1221,
    n1218,
    n953,
    n955,
    n966
  );


  xor
  g1204
  (
    n1255,
    n957,
    n1204,
    n951,
    n1215
  );


  xnor
  g1205
  (
    n1241,
    n970,
    n955,
    n960,
    n1199
  );


  or
  g1206
  (
    n1238,
    n962,
    n1216,
    n968,
    n1187
  );


  xor
  g1207
  (
    n1237,
    n951,
    n965,
    n971,
    n955
  );


  xnor
  g1208
  (
    n1227,
    n1201,
    n956,
    n946,
    n971
  );


  or
  g1209
  (
    n1232,
    n951,
    n1190,
    n966,
    n1197
  );


  xor
  g1210
  (
    n1226,
    n959,
    n950,
    n1194,
    n949
  );


  xor
  g1211
  (
    n1224,
    n1186,
    n1196,
    n1205,
    n968
  );


  nand
  g1212
  (
    n1249,
    n953,
    n948,
    n963,
    n1214
  );


  and
  g1213
  (
    n1251,
    n973,
    n949,
    n958,
    n952
  );


  nor
  g1214
  (
    n1231,
    n956,
    n954,
    n1184,
    n948
  );


  or
  g1215
  (
    n1223,
    n973,
    n961,
    n1189
  );


  xor
  g1216
  (
    n1236,
    n951,
    n947,
    n962,
    n1183
  );


  xnor
  g1217
  (
    n1252,
    n970,
    n1185,
    n963,
    n1209
  );


  nand
  g1218
  (
    n1245,
    n966,
    n965,
    n967,
    n957
  );


  xnor
  g1219
  (
    n1234,
    n967,
    n1211,
    n948,
    n958
  );


  and
  g1220
  (
    n1256,
    n971,
    n969,
    n970,
    n963
  );


  nor
  g1221
  (
    n1228,
    n973,
    n959,
    n1203,
    n946
  );


  nand
  g1222
  (
    n1222,
    n1208,
    n964,
    n957,
    n947
  );


  or
  g1223
  (
    n1225,
    n972,
    n967,
    n964,
    n1192
  );


  xnor
  g1224
  (
    n1247,
    n965,
    n953,
    n1202,
    n1191
  );


  or
  g1225
  (
    n1239,
    n961,
    n956,
    n1217,
    n962
  );


  xor
  g1226
  (
    n1325,
    n1005,
    n1006,
    n1226,
    n1235
  );


  nand
  g1227
  (
    KeyWire_0_10,
    n1244,
    n1221,
    n1225,
    n1254
  );


  xor
  g1228
  (
    n1268,
    n846,
    n1065,
    n1086,
    n1247
  );


  nand
  g1229
  (
    n1320,
    n832,
    n1079,
    n1153,
    n850
  );


  or
  g1230
  (
    n1293,
    n1249,
    n834,
    n1223,
    n1054
  );


  or
  g1231
  (
    n1283,
    n1222,
    n852,
    n1058,
    n1220
  );


  nand
  g1232
  (
    n1313,
    n1233,
    n839,
    n1055,
    n1163
  );


  nor
  g1233
  (
    n1326,
    n838,
    n1237,
    n852,
    n836
  );


  nand
  g1234
  (
    n1305,
    n1253,
    n1247,
    n1088,
    n846
  );


  nand
  g1235
  (
    n1272,
    n1084,
    n841,
    n1256,
    n1165
  );


  nand
  g1236
  (
    n1294,
    n1235,
    n1231,
    n1156,
    n1070
  );


  and
  g1237
  (
    n1316,
    n1230,
    n1005,
    n1160,
    n1237
  );


  or
  g1238
  (
    n1308,
    n1063,
    n848,
    n1168,
    n840
  );


  xnor
  g1239
  (
    n1281,
    n837,
    n1228,
    n842,
    n1237
  );


  or
  g1240
  (
    n1323,
    n848,
    n1060,
    n1080,
    n1053
  );


  xor
  g1241
  (
    n1319,
    n843,
    n1164,
    n1234,
    n853
  );


  xor
  g1242
  (
    n1298,
    n1243,
    n1250,
    n847,
    n1235
  );


  xor
  g1243
  (
    n1330,
    n851,
    n847,
    n1072,
    n1239
  );


  or
  g1244
  (
    n1315,
    n1059,
    n1236,
    n841,
    n838
  );


  nor
  g1245
  (
    n1269,
    n1252,
    n1224,
    n1248,
    n831
  );


  and
  g1246
  (
    n1309,
    n1053,
    n1241,
    n1254,
    n1246
  );


  nand
  g1247
  (
    n1273,
    n1234,
    n1004,
    n852,
    n1157
  );


  and
  g1248
  (
    n1282,
    n1229,
    n1004,
    n1245,
    n1253
  );


  or
  g1249
  (
    n1306,
    n849,
    n1005,
    n852,
    n838
  );


  nand
  g1250
  (
    n1299,
    n1248,
    n1240,
    n1249,
    n1069
  );


  xor
  g1251
  (
    n1317,
    n1251,
    n834,
    n1236,
    n1233
  );


  xor
  g1252
  (
    n1292,
    n1238,
    n1052,
    n1241,
    n1155
  );


  xnor
  g1253
  (
    n1280,
    n1139,
    n1257,
    n1249,
    n1083
  );


  nand
  g1254
  (
    n1286,
    n1161,
    n1243,
    n1251
  );


  xor
  g1255
  (
    n1297,
    n1221,
    n1225,
    n1052
  );


  nand
  g1256
  (
    n1314,
    n1228,
    n840,
    n843,
    n1243
  );


  or
  g1257
  (
    n1275,
    n1071,
    n1226,
    n1246
  );


  or
  g1258
  (
    n1263,
    n1231,
    n1249,
    n1228,
    n1054
  );


  nor
  g1259
  (
    n1324,
    n1075,
    n1240,
    n845,
    n1223
  );


  nor
  g1260
  (
    n1259,
    n1255,
    n1074,
    n1245,
    n1006
  );


  xor
  g1261
  (
    n1276,
    n1236,
    n1052,
    n1159,
    n1055
  );


  nor
  g1262
  (
    n1261,
    n1005,
    n1230,
    n833,
    n1073
  );


  xnor
  g1263
  (
    n1258,
    n843,
    n1247,
    n1234,
    n1228
  );


  nand
  g1264
  (
    n1332,
    n839,
    n1158,
    n844
  );


  nand
  g1265
  (
    n1285,
    n853,
    n833,
    n837,
    n1224
  );


  xnor
  g1266
  (
    n1335,
    n847,
    n832,
    n1238,
    n1256
  );


  nor
  g1267
  (
    n1260,
    n843,
    n1051,
    n1242,
    n842
  );


  and
  g1268
  (
    n1304,
    n831,
    n1162,
    n1242,
    n1232
  );


  and
  g1269
  (
    n1267,
    n844,
    n1006,
    n1224,
    n1238
  );


  nand
  g1270
  (
    n1312,
    n1231,
    n1227,
    n1232
  );


  or
  g1271
  (
    n1302,
    n1244,
    n834,
    n832,
    n846
  );


  and
  g1272
  (
    n1287,
    n846,
    n1246,
    n839,
    n844
  );


  xnor
  g1273
  (
    n1274,
    n851,
    n1062,
    n1082,
    n1222
  );


  xnor
  g1274
  (
    n1295,
    n1081,
    n1233,
    n848,
    n1068
  );


  xor
  g1275
  (
    n1328,
    n1224,
    n1221,
    n1231,
    n1255
  );


  xnor
  g1276
  (
    n1337,
    n1252,
    n1240,
    n1251,
    n1230
  );


  and
  g1277
  (
    n1311,
    n1052,
    n1239,
    n853,
    n1227
  );


  xor
  g1278
  (
    n1333,
    n833,
    n1154,
    n837,
    n1235
  );


  nor
  g1279
  (
    n1307,
    n1232,
    n1250,
    n1006
  );


  and
  g1280
  (
    n1279,
    n1085,
    n1257,
    n1255,
    n839
  );


  xnor
  g1281
  (
    n1329,
    n1223,
    n1244,
    n836,
    n1004
  );


  nor
  g1282
  (
    n1288,
    n836,
    n835,
    n1090,
    n842
  );


  and
  g1283
  (
    n1291,
    n1238,
    n834,
    n836,
    n835
  );


  nor
  g1284
  (
    n1266,
    n1248,
    n1222,
    n1078,
    n1229
  );


  xnor
  g1285
  (
    n1262,
    n833,
    n1066,
    n1239,
    n1244
  );


  xor
  g1286
  (
    n1301,
    n1254,
    n845,
    n1252,
    n1061
  );


  nor
  g1287
  (
    n1296,
    n1254,
    n1253,
    n832,
    n714
  );


  xor
  g1288
  (
    n1336,
    n850,
    n1245,
    n853,
    n831
  );


  nand
  g1289
  (
    n1270,
    n1053,
    n1054,
    n1057,
    n1223
  );


  xnor
  g1290
  (
    n1290,
    n1089,
    n1166,
    n1227,
    n1230
  );


  nand
  g1291
  (
    n1318,
    n1102,
    n851,
    n841,
    n837
  );


  xor
  g1292
  (
    n1303,
    n1256,
    n840,
    n1241
  );


  nor
  g1293
  (
    n1264,
    n1252,
    n1234,
    n847,
    n1053
  );


  and
  g1294
  (
    n1271,
    n1242,
    n1222,
    n1055,
    n1237
  );


  nor
  g1295
  (
    n1278,
    n1054,
    n1255,
    n1229,
    n1242
  );


  xnor
  g1296
  (
    n1327,
    n850,
    n835,
    n849,
    n1169
  );


  xor
  g1297
  (
    n1284,
    n1055,
    n1167,
    n1233,
    n1077
  );


  or
  g1298
  (
    n1322,
    n838,
    n1229,
    n1051,
    n1240
  );


  nand
  g1299
  (
    n1338,
    n1248,
    n1256,
    n1221,
    n1236
  );


  nand
  g1300
  (
    n1321,
    n1225,
    n1226,
    n1241,
    n835
  );


  or
  g1301
  (
    n1310,
    n1239,
    n1067,
    n1253,
    n841
  );


  xor
  g1302
  (
    n1277,
    n849,
    n1064,
    n1257,
    n845
  );


  xor
  g1303
  (
    n1334,
    n1226,
    n1051,
    n1257,
    n1247
  );


  nand
  g1304
  (
    KeyWire_0_13,
    n1245,
    n848,
    n1250,
    n1076
  );


  xor
  g1305
  (
    n1331,
    n842,
    n1087,
    n849,
    n1243
  );


  or
  g1306
  (
    KeyWire_0_18,
    n851,
    n845,
    n1232,
    n850
  );


  nand
  g1307
  (
    n1357,
    n1279,
    n1331,
    n1330,
    n1287
  );


  xnor
  g1308
  (
    n1343,
    n1272,
    n1318,
    n1300,
    n1281
  );


  xnor
  g1309
  (
    n1356,
    n1332,
    n1271,
    n1324,
    n1283
  );


  xnor
  g1310
  (
    n1350,
    n1288,
    n1333,
    n973,
    n1293
  );


  nand
  g1311
  (
    n1342,
    n1332,
    n1276,
    n1330,
    n1336
  );


  nand
  g1312
  (
    n1340,
    n1307,
    n1321,
    n1308,
    n1291
  );


  and
  g1313
  (
    n1353,
    n1335,
    n1336,
    n1327,
    n1305
  );


  nand
  g1314
  (
    n1352,
    n1289,
    n1326,
    n1266,
    n1334
  );


  nor
  g1315
  (
    n1348,
    n1274,
    n1313,
    n1324,
    n1334
  );


  and
  g1316
  (
    n1346,
    n1326,
    n1309,
    n1319,
    n1331
  );


  or
  g1317
  (
    n1359,
    n1320,
    n1336,
    n1310,
    n1333
  );


  xnor
  g1318
  (
    n1363,
    n1337,
    n1295,
    n1330,
    n1306
  );


  and
  g1319
  (
    KeyWire_0_7,
    n1275,
    n1331,
    n1325,
    n1323
  );


  or
  g1320
  (
    n1341,
    n1335,
    n1311,
    n1328,
    n1331
  );


  nand
  g1321
  (
    n1345,
    n1269,
    n1268,
    n1325,
    n1332
  );


  or
  g1322
  (
    n1368,
    n1290,
    n1326,
    n1325,
    n1332
  );


  xor
  g1323
  (
    n1351,
    n1328,
    n1280,
    n1335,
    n1330
  );


  xor
  g1324
  (
    n1344,
    n1336,
    n1337,
    n1282,
    n1278
  );


  or
  g1325
  (
    n1362,
    n1328,
    n1327,
    n1261,
    n1334
  );


  nor
  g1326
  (
    n1347,
    n1323,
    n1329,
    n1286
  );


  or
  g1327
  (
    n1364,
    n1324,
    n1284,
    n1329
  );


  and
  g1328
  (
    n1360,
    n1324,
    n1322,
    n1326,
    n1265
  );


  nand
  g1329
  (
    n1349,
    n1277,
    n1327,
    n1334,
    n1285
  );


  and
  g1330
  (
    n1361,
    n1259,
    n1312,
    n1333,
    n1263
  );


  or
  g1331
  (
    n1365,
    n1267,
    n1292,
    n1317,
    n1298
  );


  xor
  g1332
  (
    n1366,
    n1337,
    n1262,
    n1304,
    n1260
  );


  nand
  g1333
  (
    n1369,
    n1270,
    n1303,
    n1337,
    n1325
  );


  nor
  g1334
  (
    n1355,
    n1314,
    n1302,
    n1315,
    n1297
  );


  xnor
  g1335
  (
    n1367,
    n1333,
    n1273,
    n1316,
    n1328
  );


  xnor
  g1336
  (
    n1358,
    n1301,
    n1264,
    n1296,
    n1258
  );


  nor
  g1337
  (
    n1354,
    n1335,
    n1327,
    n1294,
    n1299
  );


  or
  g1338
  (
    n1371,
    n1354,
    n1345,
    n1361,
    n1363
  );


  and
  g1339
  (
    n1373,
    n1357,
    n1347,
    n1349,
    n1369
  );


  and
  g1340
  (
    n1374,
    n1341,
    n1352,
    n1368,
    n1364
  );


  xor
  g1341
  (
    n1375,
    n1342,
    n1365,
    n1355,
    n1350
  );


  nor
  g1342
  (
    n1376,
    n1367,
    n1358,
    n1359,
    n1339
  );


  xnor
  g1343
  (
    n1372,
    n1353,
    n1340,
    n1366,
    n1344
  );


  nand
  g1344
  (
    n1377,
    n1351,
    n1369,
    n1356,
    n1362
  );


  nand
  g1345
  (
    n1370,
    n1343,
    n1348,
    n1360,
    n1346
  );


  not
  g1346
  (
    n1378,
    n1377
  );


  xnor
  g1347
  (
    n1380,
    n1369,
    n1338,
    n154,
    n1378
  );


  and
  g1348
  (
    n1379,
    n1338,
    n155,
    n1378
  );


  xnor
  g1349
  (
    n1382,
    n1369,
    n1378,
    n155
  );


  xnor
  g1350
  (
    n1381,
    n154,
    n1338,
    n155
  );


  xor
  g1351
  (
    n1383,
    n1379,
    n1382,
    n1380,
    n1381
  );


  xor
  KeyGate_0_0
  (
    n214,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n913,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n993,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n641,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n983,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n251,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n221,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1339,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1096,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1095,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n1289,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n771,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n433,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1265,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n313,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n237,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n211,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n493,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n1300,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n738,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n833,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n162,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n376,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1121,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n294,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n89,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n616,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n886,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n253,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n408,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n724,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n818,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


