

module Stat_1000_202
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n647,
  n629,
  n639,
  n626,
  n622,
  n627,
  n646,
  n640,
  n641,
  n635,
  n633,
  n619,
  n625,
  n644,
  n624,
  n618,
  n631,
  n620,
  n636,
  n638,
  n1017,
  n1026,
  n1027,
  n1028,
  n1020,
  n1021,
  n1022,
  n1024,
  n1023,
  n1019,
  n1025,
  n1032
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n647;output n629;output n639;output n626;output n622;output n627;output n646;output n640;output n641;output n635;output n633;output n619;output n625;output n644;output n624;output n618;output n631;output n620;output n636;output n638;output n1017;output n1026;output n1027;output n1028;output n1020;output n1021;output n1022;output n1024;output n1023;output n1019;output n1025;output n1032;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n621;wire n623;wire n628;wire n630;wire n632;wire n634;wire n637;wire n642;wire n643;wire n645;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1018;wire n1029;wire n1030;wire n1031;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n76,
    n9
  );


  not
  g1
  (
    n59,
    n1
  );


  buf
  g2
  (
    n61,
    n14
  );


  not
  g3
  (
    n41,
    n17
  );


  buf
  g4
  (
    n60,
    n10
  );


  buf
  g5
  (
    n56,
    n2
  );


  not
  g6
  (
    n48,
    n11
  );


  not
  g7
  (
    KeyWire_0_6,
    n6
  );


  not
  g8
  (
    KeyWire_0_5,
    n3
  );


  buf
  g9
  (
    n55,
    n19
  );


  not
  g10
  (
    n72,
    n5
  );


  buf
  g11
  (
    n71,
    n14
  );


  buf
  g12
  (
    n38,
    n15
  );


  buf
  g13
  (
    n39,
    n6
  );


  not
  g14
  (
    n50,
    n4
  );


  not
  g15
  (
    n40,
    n11
  );


  buf
  g16
  (
    n65,
    n14
  );


  buf
  g17
  (
    n73,
    n15
  );


  buf
  g18
  (
    n53,
    n3
  );


  buf
  g19
  (
    n58,
    n8
  );


  not
  g20
  (
    n45,
    n16
  );


  not
  g21
  (
    n63,
    n15
  );


  buf
  g22
  (
    n52,
    n10
  );


  not
  g23
  (
    n33,
    n14
  );


  buf
  g24
  (
    n47,
    n12
  );


  not
  g25
  (
    n54,
    n2
  );


  buf
  g26
  (
    n74,
    n7
  );


  not
  g27
  (
    n35,
    n18
  );


  buf
  g28
  (
    n44,
    n19
  );


  buf
  g29
  (
    n49,
    n9
  );


  buf
  g30
  (
    n66,
    n17
  );


  buf
  g31
  (
    n64,
    n8
  );


  buf
  g32
  (
    n78,
    n5
  );


  buf
  g33
  (
    n37,
    n7
  );


  not
  g34
  (
    n46,
    n16
  );


  not
  g35
  (
    n69,
    n18
  );


  buf
  g36
  (
    n70,
    n16
  );


  buf
  g37
  (
    n62,
    n18
  );


  not
  g38
  (
    n80,
    n13
  );


  not
  g39
  (
    KeyWire_0_15,
    n15
  );


  not
  g40
  (
    n34,
    n1
  );


  not
  g41
  (
    n57,
    n13
  );


  not
  g42
  (
    n36,
    n17
  );


  buf
  g43
  (
    n67,
    n4
  );


  not
  g44
  (
    n75,
    n16
  );


  not
  g45
  (
    n79,
    n12
  );


  not
  g46
  (
    n77,
    n17
  );


  not
  g47
  (
    n68,
    n18
  );


  not
  g48
  (
    n156,
    n74
  );


  not
  g49
  (
    n95,
    n58
  );


  buf
  g50
  (
    n186,
    n38
  );


  not
  g51
  (
    n83,
    n71
  );


  not
  g52
  (
    n263,
    n76
  );


  not
  g53
  (
    n178,
    n57
  );


  buf
  g54
  (
    n141,
    n76
  );


  not
  g55
  (
    n222,
    n52
  );


  not
  g56
  (
    n149,
    n71
  );


  not
  g57
  (
    n210,
    n25
  );


  not
  g58
  (
    n157,
    n48
  );


  buf
  g59
  (
    n246,
    n45
  );


  not
  g60
  (
    n205,
    n74
  );


  not
  g61
  (
    n128,
    n51
  );


  buf
  g62
  (
    n107,
    n73
  );


  not
  g63
  (
    n150,
    n80
  );


  buf
  g64
  (
    n126,
    n71
  );


  not
  g65
  (
    n191,
    n53
  );


  buf
  g66
  (
    n147,
    n80
  );


  buf
  g67
  (
    n249,
    n44
  );


  not
  g68
  (
    n198,
    n44
  );


  not
  g69
  (
    n132,
    n66
  );


  not
  g70
  (
    n239,
    n44
  );


  not
  g71
  (
    n102,
    n56
  );


  not
  g72
  (
    n154,
    n41
  );


  not
  g73
  (
    n99,
    n65
  );


  buf
  g74
  (
    n214,
    n24
  );


  buf
  g75
  (
    n100,
    n47
  );


  buf
  g76
  (
    n93,
    n62
  );


  buf
  g77
  (
    n167,
    n78
  );


  not
  g78
  (
    n169,
    n67
  );


  buf
  g79
  (
    n195,
    n55
  );


  not
  g80
  (
    n170,
    n24
  );


  not
  g81
  (
    n230,
    n47
  );


  buf
  g82
  (
    n243,
    n33
  );


  not
  g83
  (
    n136,
    n43
  );


  not
  g84
  (
    n152,
    n43
  );


  buf
  g85
  (
    n112,
    n23
  );


  not
  g86
  (
    n87,
    n51
  );


  buf
  g87
  (
    n188,
    n65
  );


  not
  g88
  (
    KeyWire_0_13,
    n76
  );


  not
  g89
  (
    n137,
    n70
  );


  not
  g90
  (
    n176,
    n42
  );


  buf
  g91
  (
    n245,
    n72
  );


  buf
  g92
  (
    n119,
    n59
  );


  buf
  g93
  (
    n106,
    n50
  );


  not
  g94
  (
    n221,
    n45
  );


  not
  g95
  (
    n262,
    n62
  );


  buf
  g96
  (
    n180,
    n21
  );


  not
  g97
  (
    n108,
    n22
  );


  not
  g98
  (
    n181,
    n69
  );


  buf
  g99
  (
    n81,
    n39
  );


  buf
  g100
  (
    n86,
    n45
  );


  buf
  g101
  (
    n201,
    n47
  );


  buf
  g102
  (
    n145,
    n38
  );


  not
  g103
  (
    n165,
    n41
  );


  buf
  g104
  (
    n98,
    n72
  );


  not
  g105
  (
    n173,
    n48
  );


  not
  g106
  (
    n192,
    n77
  );


  buf
  g107
  (
    n225,
    n34
  );


  not
  g108
  (
    n94,
    n22
  );


  buf
  g109
  (
    n127,
    n77
  );


  buf
  g110
  (
    n104,
    n46
  );


  not
  g111
  (
    n190,
    n20
  );


  not
  g112
  (
    n143,
    n25
  );


  not
  g113
  (
    n259,
    n46
  );


  not
  g114
  (
    n237,
    n79
  );


  not
  g115
  (
    n233,
    n69
  );


  not
  g116
  (
    n135,
    n61
  );


  buf
  g117
  (
    n117,
    n37
  );


  not
  g118
  (
    n82,
    n58
  );


  not
  g119
  (
    n200,
    n70
  );


  not
  g120
  (
    n241,
    n25
  );


  not
  g121
  (
    n163,
    n71
  );


  buf
  g122
  (
    n164,
    n61
  );


  not
  g123
  (
    n203,
    n77
  );


  not
  g124
  (
    n260,
    n66
  );


  not
  g125
  (
    n116,
    n68
  );


  not
  g126
  (
    n84,
    n40
  );


  not
  g127
  (
    n121,
    n79
  );


  buf
  g128
  (
    n264,
    n63
  );


  not
  g129
  (
    n251,
    n67
  );


  buf
  g130
  (
    n90,
    n66
  );


  not
  g131
  (
    n197,
    n59
  );


  buf
  g132
  (
    n124,
    n54
  );


  buf
  g133
  (
    n118,
    n54
  );


  not
  g134
  (
    n158,
    n78
  );


  not
  g135
  (
    n92,
    n40
  );


  not
  g136
  (
    n134,
    n36
  );


  not
  g137
  (
    n168,
    n36
  );


  not
  g138
  (
    n184,
    n69
  );


  not
  g139
  (
    n105,
    n56
  );


  not
  g140
  (
    n258,
    n42
  );


  buf
  g141
  (
    n254,
    n23
  );


  buf
  g142
  (
    n226,
    n61
  );


  not
  g143
  (
    n266,
    n60
  );


  not
  g144
  (
    n196,
    n60
  );


  buf
  g145
  (
    n224,
    n37
  );


  not
  g146
  (
    n125,
    n74
  );


  buf
  g147
  (
    n256,
    n24
  );


  buf
  g148
  (
    n270,
    n20
  );


  not
  g149
  (
    n130,
    n75
  );


  buf
  g150
  (
    n159,
    n73
  );


  buf
  g151
  (
    n122,
    n79
  );


  not
  g152
  (
    n151,
    n56
  );


  not
  g153
  (
    n223,
    n59
  );


  buf
  g154
  (
    n185,
    n65
  );


  not
  g155
  (
    n161,
    n49
  );


  not
  g156
  (
    n255,
    n57
  );


  buf
  g157
  (
    n183,
    n54
  );


  not
  g158
  (
    n171,
    n79
  );


  not
  g159
  (
    n240,
    n40
  );


  buf
  g160
  (
    KeyWire_0_2,
    n72
  );


  buf
  g161
  (
    n189,
    n38
  );


  not
  g162
  (
    n229,
    n22
  );


  buf
  g163
  (
    n236,
    n20
  );


  buf
  g164
  (
    n216,
    n39
  );


  buf
  g165
  (
    n267,
    n56
  );


  buf
  g166
  (
    n232,
    n25
  );


  not
  g167
  (
    KeyWire_0_1,
    n19
  );


  not
  g168
  (
    n209,
    n34
  );


  buf
  g169
  (
    n269,
    n52
  );


  not
  g170
  (
    n231,
    n70
  );


  buf
  g171
  (
    n172,
    n34
  );


  buf
  g172
  (
    n187,
    n60
  );


  buf
  g173
  (
    n215,
    n37
  );


  not
  g174
  (
    n109,
    n76
  );


  buf
  g175
  (
    n177,
    n69
  );


  not
  g176
  (
    n166,
    n21
  );


  not
  g177
  (
    n175,
    n50
  );


  buf
  g178
  (
    n265,
    n42
  );


  not
  g179
  (
    n242,
    n61
  );


  buf
  g180
  (
    KeyWire_0_20,
    n64
  );


  not
  g181
  (
    n140,
    n19
  );


  buf
  g182
  (
    n144,
    n64
  );


  buf
  g183
  (
    n208,
    n24
  );


  not
  g184
  (
    n217,
    n47
  );


  buf
  g185
  (
    n115,
    n78
  );


  not
  g186
  (
    n227,
    n33
  );


  not
  g187
  (
    n133,
    n66
  );


  not
  g188
  (
    n247,
    n73
  );


  not
  g189
  (
    n212,
    n26
  );


  not
  g190
  (
    n234,
    n35
  );


  not
  g191
  (
    n162,
    n37
  );


  not
  g192
  (
    n146,
    n26
  );


  not
  g193
  (
    n179,
    n52
  );


  buf
  g194
  (
    n110,
    n45
  );


  buf
  g195
  (
    n85,
    n33
  );


  buf
  g196
  (
    n204,
    n64
  );


  buf
  g197
  (
    n155,
    n39
  );


  buf
  g198
  (
    n97,
    n57
  );


  buf
  g199
  (
    n218,
    n58
  );


  buf
  g200
  (
    n182,
    n35
  );


  buf
  g201
  (
    n199,
    n55
  );


  buf
  g202
  (
    n228,
    n60
  );


  buf
  g203
  (
    n250,
    n43
  );


  not
  g204
  (
    n202,
    n54
  );


  not
  g205
  (
    n238,
    n77
  );


  not
  g206
  (
    n194,
    n65
  );


  not
  g207
  (
    n96,
    n63
  );


  not
  g208
  (
    n88,
    n68
  );


  buf
  g209
  (
    n207,
    n42
  );


  not
  g210
  (
    n129,
    n35
  );


  not
  g211
  (
    n114,
    n53
  );


  not
  g212
  (
    n193,
    n59
  );


  buf
  g213
  (
    n244,
    n49
  );


  buf
  g214
  (
    n142,
    n55
  );


  not
  g215
  (
    n219,
    n35
  );


  buf
  g216
  (
    n138,
    n62
  );


  buf
  g217
  (
    n206,
    n38
  );


  buf
  g218
  (
    n220,
    n34
  );


  not
  g219
  (
    n153,
    n62
  );


  buf
  g220
  (
    n91,
    n36
  );


  not
  g221
  (
    n252,
    n58
  );


  buf
  g222
  (
    n211,
    n70
  );


  not
  g223
  (
    n111,
    n75
  );


  not
  g224
  (
    n89,
    n67
  );


  buf
  g225
  (
    n103,
    n23
  );


  not
  g226
  (
    n160,
    n68
  );


  not
  g227
  (
    n253,
    n75
  );


  not
  g228
  (
    n261,
    n36
  );


  buf
  g229
  (
    n174,
    n67
  );


  nand
  g230
  (
    n113,
    n22,
    n41
  );


  nand
  g231
  (
    n123,
    n73,
    n48,
    n75,
    n68
  );


  and
  g232
  (
    n268,
    n53,
    n63,
    n46,
    n40
  );


  xor
  g233
  (
    n257,
    n20,
    n33,
    n51,
    n52
  );


  or
  g234
  (
    n148,
    n23,
    n49,
    n44,
    n50
  );


  nor
  g235
  (
    n213,
    n80,
    n80,
    n39,
    n63
  );


  xnor
  g236
  (
    n131,
    n78,
    n53,
    n43,
    n46
  );


  nor
  g237
  (
    n139,
    n48,
    n50,
    n57,
    n55
  );


  and
  g238
  (
    n271,
    n21,
    n41,
    n72,
    n74
  );


  nor
  g239
  (
    n248,
    n21,
    n51,
    n49,
    n64
  );


  or
  g240
  (
    n455,
    n247,
    n174,
    n196,
    n145
  );


  nor
  g241
  (
    n376,
    n209,
    n251,
    n169,
    n249
  );


  xnor
  g242
  (
    n287,
    n103,
    n172,
    n211,
    n213
  );


  or
  g243
  (
    n400,
    n244,
    n173,
    n226,
    n209
  );


  and
  g244
  (
    n425,
    n171,
    n231,
    n106,
    n125
  );


  nor
  g245
  (
    n385,
    n135,
    n242,
    n243,
    n191
  );


  nor
  g246
  (
    n382,
    n220,
    n146,
    n213,
    n231
  );


  nand
  g247
  (
    n295,
    n268,
    n149,
    n238,
    n258
  );


  xnor
  g248
  (
    n446,
    n253,
    n163,
    n239,
    n226
  );


  and
  g249
  (
    n405,
    n108,
    n220,
    n226,
    n173
  );


  and
  g250
  (
    n423,
    n246,
    n219,
    n85,
    n89
  );


  xnor
  g251
  (
    n329,
    n103,
    n134,
    n148,
    n157
  );


  xnor
  g252
  (
    n313,
    n82,
    n218,
    n242,
    n158
  );


  xnor
  g253
  (
    n448,
    n171,
    n86,
    n110,
    n199
  );


  and
  g254
  (
    n442,
    n166,
    n247,
    n186,
    n199
  );


  or
  g255
  (
    n374,
    n238,
    n219,
    n170,
    n161
  );


  nand
  g256
  (
    n424,
    n189,
    n258,
    n217,
    n95
  );


  and
  g257
  (
    n351,
    n154,
    n82,
    n245,
    n128
  );


  and
  g258
  (
    n370,
    n90,
    n113,
    n258,
    n213
  );


  nand
  g259
  (
    n378,
    n159,
    n120,
    n197,
    n255
  );


  nand
  g260
  (
    n434,
    n110,
    n265,
    n96,
    n266
  );


  xnor
  g261
  (
    n431,
    n219,
    n198,
    n154,
    n114
  );


  and
  g262
  (
    n430,
    n259,
    n112,
    n248,
    n126
  );


  nor
  g263
  (
    n393,
    n111,
    n230,
    n84,
    n198
  );


  and
  g264
  (
    n310,
    n239,
    n263,
    n105,
    n98
  );


  xnor
  g265
  (
    n443,
    n98,
    n244,
    n157,
    n208
  );


  xnor
  g266
  (
    n353,
    n215,
    n167,
    n137,
    n143
  );


  nor
  g267
  (
    n418,
    n168,
    n201,
    n212,
    n102
  );


  or
  g268
  (
    n403,
    n185,
    n95,
    n243,
    n181
  );


  or
  g269
  (
    n459,
    n127,
    n262,
    n142,
    n175
  );


  nand
  g270
  (
    n362,
    n198,
    n97,
    n254,
    n100
  );


  or
  g271
  (
    n314,
    n267,
    n205,
    n264,
    n212
  );


  nor
  g272
  (
    n460,
    n240,
    n166,
    n227,
    n93
  );


  nor
  g273
  (
    n392,
    n133,
    n81,
    n82,
    n92
  );


  and
  g274
  (
    n309,
    n242,
    n127,
    n136,
    n103
  );


  and
  g275
  (
    n342,
    n109,
    n108,
    n182,
    n138
  );


  xnor
  g276
  (
    n320,
    n207,
    n261,
    n162,
    n120
  );


  and
  g277
  (
    n368,
    n152,
    n186,
    n100,
    n156
  );


  xor
  g278
  (
    n419,
    n252,
    n116,
    n246,
    n263
  );


  or
  g279
  (
    n274,
    n228,
    n129,
    n144,
    n225
  );


  xnor
  g280
  (
    n328,
    n256,
    n137,
    n253,
    n99
  );


  xor
  g281
  (
    n277,
    n174,
    n252,
    n208,
    n225
  );


  or
  g282
  (
    n447,
    n267,
    n145,
    n130,
    n212
  );


  xnor
  g283
  (
    n359,
    n155,
    n122,
    n99,
    n210
  );


  xnor
  g284
  (
    n438,
    n111,
    n156,
    n240,
    n127
  );


  xnor
  g285
  (
    n413,
    n161,
    n159,
    n123,
    n151
  );


  xnor
  g286
  (
    n389,
    n149,
    n233,
    n115,
    n195
  );


  xor
  g287
  (
    n441,
    n258,
    n196,
    n168,
    n209
  );


  nor
  g288
  (
    n308,
    n163,
    n230,
    n229,
    n100
  );


  or
  g289
  (
    n322,
    n182,
    n216,
    n155,
    n109
  );


  or
  g290
  (
    n439,
    n153,
    n241,
    n164,
    n229
  );


  and
  g291
  (
    n428,
    n125,
    n220,
    n120,
    n87
  );


  or
  g292
  (
    n420,
    n252,
    n217,
    n157,
    n133
  );


  or
  g293
  (
    n394,
    n257,
    n157,
    n254,
    n164
  );


  xnor
  g294
  (
    n347,
    n188,
    n260,
    n116,
    n122
  );


  nand
  g295
  (
    n432,
    n191,
    n88,
    n216,
    n104
  );


  nor
  g296
  (
    n332,
    n108,
    n172,
    n264,
    n86
  );


  nand
  g297
  (
    n409,
    n199,
    n150,
    n222,
    n94
  );


  or
  g298
  (
    n421,
    n174,
    n150,
    n87,
    n171
  );


  xnor
  g299
  (
    n412,
    n202,
    n190,
    n233,
    n255
  );


  nor
  g300
  (
    n346,
    n206,
    n138,
    n124,
    n109
  );


  nor
  g301
  (
    n361,
    n172,
    n112,
    n87,
    n148
  );


  nor
  g302
  (
    n334,
    n223,
    n238,
    n191,
    n101
  );


  nand
  g303
  (
    n316,
    n202,
    n221,
    n247,
    n235
  );


  xor
  g304
  (
    n371,
    n163,
    n93,
    n181,
    n146
  );


  xnor
  g305
  (
    n285,
    n231,
    n187,
    n121,
    n118
  );


  nor
  g306
  (
    KeyWire_0_11,
    n204,
    n248,
    n211,
    n194
  );


  nor
  g307
  (
    KeyWire_0_4,
    n261,
    n196,
    n254,
    n175
  );


  nor
  g308
  (
    n324,
    n131,
    n263,
    n203,
    n184
  );


  or
  g309
  (
    n396,
    n116,
    n128,
    n226,
    n156
  );


  and
  g310
  (
    KeyWire_0_27,
    n181,
    n184,
    n165,
    n250
  );


  or
  g311
  (
    n433,
    n169,
    n165,
    n104,
    n237
  );


  nand
  g312
  (
    n354,
    n192,
    n155,
    n236,
    n224
  );


  nand
  g313
  (
    n283,
    n155,
    n228,
    n81,
    n99
  );


  xnor
  g314
  (
    n407,
    n147,
    n154,
    n119,
    n117
  );


  xor
  g315
  (
    n436,
    n143,
    n261,
    n185,
    n107
  );


  and
  g316
  (
    n402,
    n225,
    n220,
    n235,
    n173
  );


  nor
  g317
  (
    n302,
    n180,
    n205,
    n250,
    n141
  );


  nor
  g318
  (
    n390,
    n109,
    n202,
    n97,
    n187
  );


  xor
  g319
  (
    n321,
    n218,
    n88,
    n189
  );


  xor
  g320
  (
    n326,
    n119,
    n135,
    n256,
    n233
  );


  and
  g321
  (
    n364,
    n243,
    n144,
    n150,
    n265
  );


  and
  g322
  (
    n417,
    n123,
    n127,
    n179,
    n252
  );


  or
  g323
  (
    n404,
    n254,
    n107,
    n189,
    n102
  );


  or
  g324
  (
    n276,
    n165,
    n113,
    n118,
    n106
  );


  and
  g325
  (
    n349,
    n264,
    n84,
    n190,
    n246
  );


  and
  g326
  (
    n427,
    n102,
    n247,
    n152,
    n215
  );


  and
  g327
  (
    n444,
    n268,
    n162,
    n84,
    n105
  );


  xor
  g328
  (
    n344,
    n193,
    n242,
    n149,
    n201
  );


  nand
  g329
  (
    n435,
    n123,
    n173,
    n167
  );


  and
  g330
  (
    n311,
    n200,
    n179,
    n140,
    n170
  );


  nand
  g331
  (
    n414,
    n119,
    n141,
    n147,
    n168
  );


  xor
  g332
  (
    n299,
    n122,
    n117,
    n142,
    n134
  );


  nor
  g333
  (
    n301,
    n85,
    n164,
    n91,
    n179
  );


  and
  g334
  (
    n398,
    n105,
    n204,
    n208,
    n135
  );


  nor
  g335
  (
    KeyWire_0_28,
    n131,
    n251,
    n209,
    n228
  );


  xnor
  g336
  (
    n360,
    n194,
    n126,
    n140,
    n89
  );


  nor
  g337
  (
    KeyWire_0_3,
    n141,
    n153,
    n182,
    n217
  );


  nand
  g338
  (
    n381,
    n171,
    n153,
    n132,
    n94
  );


  and
  g339
  (
    KeyWire_0_21,
    n203,
    n169,
    n227,
    n175
  );


  or
  g340
  (
    n350,
    n86,
    n215,
    n223,
    n263
  );


  xnor
  g341
  (
    n294,
    n98,
    n234,
    n116,
    n93
  );


  or
  g342
  (
    n356,
    n200,
    n249,
    n90,
    n158
  );


  or
  g343
  (
    n325,
    n126,
    n138,
    n240,
    n105
  );


  nor
  g344
  (
    n293,
    n146,
    n94,
    n135,
    n192
  );


  and
  g345
  (
    n387,
    n83,
    n210,
    n152,
    n131
  );


  xnor
  g346
  (
    n339,
    n219,
    n260,
    n176,
    n229
  );


  nor
  g347
  (
    n386,
    n122,
    n160,
    n86,
    n174
  );


  nor
  g348
  (
    n373,
    n266,
    n257,
    n112,
    n186
  );


  nand
  g349
  (
    n307,
    n115,
    n172,
    n144,
    n197
  );


  nor
  g350
  (
    n429,
    n218,
    n178,
    n191,
    n84
  );


  nand
  g351
  (
    n337,
    n130,
    n90,
    n110,
    n202
  );


  or
  g352
  (
    n290,
    n239,
    n96,
    n83,
    n108
  );


  xor
  g353
  (
    n336,
    n245,
    n262,
    n91,
    n136
  );


  nand
  g354
  (
    n297,
    n137,
    n195,
    n266,
    n156
  );


  nand
  g355
  (
    n345,
    n183,
    n161,
    n196,
    n176
  );


  nor
  g356
  (
    n395,
    n249,
    n183,
    n241,
    n99
  );


  xor
  g357
  (
    n292,
    n162,
    n180,
    n239,
    n248
  );


  xor
  g358
  (
    n366,
    n175,
    n260,
    n139,
    n217
  );


  or
  g359
  (
    n319,
    n218,
    n221,
    n214,
    n222
  );


  or
  g360
  (
    n312,
    n259,
    n82,
    n170,
    n210
  );


  or
  g361
  (
    n401,
    n139,
    n257,
    n200,
    n148
  );


  xnor
  g362
  (
    n379,
    n129,
    n201,
    n153,
    n125
  );


  xnor
  g363
  (
    n315,
    n101,
    n229,
    n95,
    n102
  );


  xnor
  g364
  (
    n289,
    n152,
    n245,
    n197,
    n142
  );


  and
  g365
  (
    n304,
    n193,
    n83,
    n251,
    n145
  );


  nor
  g366
  (
    n458,
    n193,
    n130,
    n106,
    n176
  );


  xnor
  g367
  (
    n365,
    n114,
    n151,
    n241,
    n250
  );


  nand
  g368
  (
    n451,
    n199,
    n158,
    n206,
    n267
  );


  xnor
  g369
  (
    n279,
    n159,
    n221,
    n81,
    n224
  );


  xor
  g370
  (
    n340,
    n138,
    n148,
    n262,
    n170
  );


  nor
  g371
  (
    n281,
    n214,
    n133,
    n134,
    n184
  );


  nor
  g372
  (
    n291,
    n111,
    n169,
    n188,
    n89
  );


  nand
  g373
  (
    KeyWire_0_30,
    n203,
    n160,
    n228,
    n237
  );


  and
  g374
  (
    n452,
    n129,
    n151,
    n134,
    n164
  );


  nand
  g375
  (
    n449,
    n246,
    n238,
    n100,
    n190
  );


  or
  g376
  (
    n416,
    n154,
    n114,
    n92,
    n106
  );


  xor
  g377
  (
    n372,
    n92,
    n257,
    n188,
    n151
  );


  xnor
  g378
  (
    n357,
    n194,
    n256,
    n178,
    n222
  );


  xnor
  g379
  (
    n288,
    n266,
    n96,
    n198,
    n110
  );


  xor
  g380
  (
    n284,
    n97,
    n160,
    n136,
    n121
  );


  xnor
  g381
  (
    n330,
    n214,
    n167,
    n126,
    n166
  );


  xnor
  g382
  (
    n282,
    n215,
    n234,
    n85,
    n177
  );


  xor
  g383
  (
    n275,
    n140,
    n139,
    n187,
    n103
  );


  nor
  g384
  (
    n305,
    n124,
    n143,
    n214,
    n211
  );


  or
  g385
  (
    n355,
    n165,
    n201,
    n237,
    n224
  );


  or
  g386
  (
    n377,
    n128,
    n150,
    n183,
    n115
  );


  and
  g387
  (
    n384,
    n183,
    n177,
    n158,
    n205
  );


  xnor
  g388
  (
    n338,
    n231,
    n235,
    n249,
    n230
  );


  xor
  g389
  (
    n318,
    n85,
    n176,
    n195,
    n177
  );


  xor
  g390
  (
    n273,
    n268,
    n139,
    n120,
    n124
  );


  xor
  g391
  (
    n406,
    n253,
    n104,
    n186,
    n131
  );


  or
  g392
  (
    n333,
    n112,
    n136,
    n91
  );


  nand
  g393
  (
    n411,
    n178,
    n166,
    n204,
    n187
  );


  nor
  g394
  (
    n453,
    n212,
    n117,
    n180,
    n210
  );


  nor
  g395
  (
    n454,
    n95,
    n189,
    n132,
    n207
  );


  or
  g396
  (
    n415,
    n92,
    n236,
    n204,
    n216
  );


  xor
  g397
  (
    n363,
    n168,
    n94,
    n244,
    n236
  );


  nand
  g398
  (
    n410,
    n124,
    n188,
    n251,
    n137
  );


  or
  g399
  (
    n450,
    n207,
    n223,
    n255,
    n140
  );


  nand
  g400
  (
    n397,
    n118,
    n259,
    n162,
    n193
  );


  xnor
  g401
  (
    n399,
    n118,
    n111,
    n232,
    n248
  );


  and
  g402
  (
    n303,
    n213,
    n206,
    n240,
    n234
  );


  xor
  g403
  (
    n278,
    n145,
    n253,
    n190,
    n250
  );


  or
  g404
  (
    n367,
    n83,
    n121,
    n260,
    n227
  );


  and
  g405
  (
    n380,
    n264,
    n87,
    n113,
    n259
  );


  xnor
  g406
  (
    n358,
    n255,
    n128,
    n129,
    n256
  );


  xor
  g407
  (
    n348,
    n241,
    n107,
    n130,
    n159
  );


  nor
  g408
  (
    n286,
    n182,
    n185,
    n216,
    n101
  );


  xor
  g409
  (
    n306,
    n223,
    n207,
    n208,
    n104
  );


  and
  g410
  (
    n327,
    n90,
    n230,
    n181,
    n265
  );


  nor
  g411
  (
    n341,
    n146,
    n261,
    n194,
    n117
  );


  xor
  g412
  (
    n445,
    n132,
    n144,
    n180,
    n88
  );


  nand
  g413
  (
    n388,
    n107,
    n232,
    n197,
    n114
  );


  nand
  g414
  (
    n375,
    n101,
    n211,
    n224,
    n235
  );


  or
  g415
  (
    n369,
    n185,
    n113,
    n125,
    n96
  );


  or
  g416
  (
    n437,
    n195,
    n222,
    n121,
    n160
  );


  and
  g417
  (
    n456,
    n143,
    n119,
    n93,
    n184
  );


  or
  g418
  (
    n352,
    n232,
    n225,
    n245,
    n234
  );


  nor
  g419
  (
    n383,
    n267,
    n200,
    n163,
    n142
  );


  xor
  g420
  (
    n408,
    n268,
    n149,
    n192,
    n237
  );


  and
  g421
  (
    KeyWire_0_19,
    n192,
    n203,
    n97,
    n262
  );


  and
  g422
  (
    n343,
    n147,
    n265,
    n179,
    n233
  );


  xor
  g423
  (
    n317,
    n178,
    n177,
    n161,
    n133
  );


  xnor
  g424
  (
    n422,
    n89,
    n227,
    n123,
    n141
  );


  nand
  g425
  (
    n296,
    n244,
    n147,
    n236,
    n221
  );


  xnor
  g426
  (
    n391,
    n243,
    n232,
    n206,
    n115
  );


  and
  g427
  (
    n440,
    n81,
    n205,
    n132,
    n98
  );


  nand
  g428
  (
    n555,
    n298,
    n401
  );


  nand
  g429
  (
    n515,
    n278,
    n420
  );


  xnor
  g430
  (
    n540,
    n390,
    n403
  );


  and
  g431
  (
    n569,
    n334,
    n410
  );


  and
  g432
  (
    n499,
    n275,
    n406
  );


  xor
  g433
  (
    n470,
    n432,
    n439
  );


  or
  g434
  (
    n564,
    n368,
    n382
  );


  nand
  g435
  (
    n496,
    n396,
    n366
  );


  nor
  g436
  (
    n541,
    n323,
    n450
  );


  xor
  g437
  (
    n543,
    n311,
    n377
  );


  xor
  g438
  (
    n495,
    n408,
    n328
  );


  xnor
  g439
  (
    n554,
    n376,
    n289
  );


  xor
  g440
  (
    n597,
    n406,
    n421
  );


  xor
  g441
  (
    n530,
    n276,
    n417
  );


  and
  g442
  (
    n508,
    n444,
    n379
  );


  xor
  g443
  (
    n471,
    n352,
    n351
  );


  xor
  g444
  (
    n586,
    n358,
    n361
  );


  xor
  g445
  (
    n480,
    n367,
    n373
  );


  nand
  g446
  (
    n521,
    n330,
    n293
  );


  nor
  g447
  (
    n548,
    n385,
    n325
  );


  nor
  g448
  (
    n588,
    n333,
    n407
  );


  nor
  g449
  (
    n552,
    n415,
    n381
  );


  nand
  g450
  (
    n498,
    n290,
    n434
  );


  xor
  g451
  (
    n463,
    n435,
    n455
  );


  nand
  g452
  (
    n523,
    n285,
    n360
  );


  and
  g453
  (
    n587,
    n445,
    n354
  );


  xor
  g454
  (
    n553,
    n430,
    n297
  );


  or
  g455
  (
    KeyWire_0_22,
    n446,
    n381
  );


  nor
  g456
  (
    n502,
    n378,
    n424
  );


  nand
  g457
  (
    n488,
    n418,
    n305
  );


  and
  g458
  (
    n565,
    n337,
    n318
  );


  xor
  g459
  (
    n501,
    n320,
    n279
  );


  nand
  g460
  (
    n614,
    n446,
    n342
  );


  and
  g461
  (
    n500,
    n277,
    n374
  );


  or
  g462
  (
    n504,
    n452,
    n445
  );


  nand
  g463
  (
    n612,
    n356,
    n336
  );


  nand
  g464
  (
    n577,
    n306,
    n370
  );


  and
  g465
  (
    n531,
    n379,
    n442
  );


  and
  g466
  (
    n582,
    n431,
    n380
  );


  nand
  g467
  (
    n556,
    n399,
    n393
  );


  and
  g468
  (
    n469,
    n353,
    n412
  );


  and
  g469
  (
    n466,
    n443,
    n418
  );


  nand
  g470
  (
    n465,
    n302,
    n427
  );


  xor
  g471
  (
    KeyWire_0_8,
    n353,
    n389
  );


  and
  g472
  (
    n494,
    n357,
    n359
  );


  nand
  g473
  (
    n561,
    n331,
    n389
  );


  xnor
  g474
  (
    n461,
    n420,
    n329
  );


  or
  g475
  (
    n615,
    n369,
    n448
  );


  nor
  g476
  (
    n482,
    n448,
    n366
  );


  nor
  g477
  (
    n545,
    n427,
    n384
  );


  and
  g478
  (
    n598,
    n296,
    n447
  );


  nand
  g479
  (
    n572,
    n443,
    n421
  );


  xnor
  g480
  (
    n481,
    n307,
    n382
  );


  xor
  g481
  (
    n528,
    n372,
    n440
  );


  xnor
  g482
  (
    n516,
    n317,
    n294
  );


  xnor
  g483
  (
    n576,
    n404,
    n438
  );


  xor
  g484
  (
    n478,
    n303,
    n436
  );


  xor
  g485
  (
    n510,
    n343,
    n363
  );


  nor
  g486
  (
    n583,
    n332,
    n451
  );


  xor
  g487
  (
    n574,
    n325,
    n332
  );


  and
  g488
  (
    n533,
    n310,
    n453
  );


  or
  g489
  (
    n479,
    n347,
    n401
  );


  or
  g490
  (
    n490,
    n328,
    n334
  );


  xor
  g491
  (
    n497,
    n383,
    n385
  );


  and
  g492
  (
    n613,
    n335,
    n322
  );


  nor
  g493
  (
    n567,
    n361,
    n308
  );


  and
  g494
  (
    n603,
    n286,
    n304
  );


  and
  g495
  (
    n529,
    n430,
    n340
  );


  nor
  g496
  (
    n562,
    n383,
    n402
  );


  xnor
  g497
  (
    n525,
    n419,
    n404
  );


  nand
  g498
  (
    n493,
    n454,
    n429
  );


  xor
  g499
  (
    n536,
    n437,
    n354
  );


  and
  g500
  (
    n522,
    n422,
    n363
  );


  or
  g501
  (
    n585,
    n437,
    n343
  );


  nand
  g502
  (
    n537,
    n288,
    n292
  );


  nand
  g503
  (
    KeyWire_0_26,
    n428,
    n358
  );


  nor
  g504
  (
    n484,
    n399,
    n315
  );


  nand
  g505
  (
    n589,
    n364,
    n384
  );


  xor
  g506
  (
    n491,
    n396,
    n394
  );


  xnor
  g507
  (
    n584,
    n392,
    n326
  );


  nand
  g508
  (
    n563,
    n449,
    n336
  );


  and
  g509
  (
    n573,
    n349,
    n274
  );


  xor
  g510
  (
    n532,
    n330,
    n321
  );


  nor
  g511
  (
    n596,
    n360,
    n367
  );


  xnor
  g512
  (
    n611,
    n419,
    n326
  );


  and
  g513
  (
    n578,
    n309,
    n402
  );


  xor
  g514
  (
    n507,
    n408,
    n451
  );


  nand
  g515
  (
    n602,
    n350,
    n447
  );


  or
  g516
  (
    n594,
    n284,
    n338
  );


  nor
  g517
  (
    KeyWire_0_0,
    n413,
    n392
  );


  xnor
  g518
  (
    n503,
    n416,
    n388
  );


  or
  g519
  (
    n610,
    n327,
    n452
  );


  nor
  g520
  (
    n566,
    n281,
    n394
  );


  xnor
  g521
  (
    n617,
    n411,
    n287
  );


  xnor
  g522
  (
    n616,
    n314,
    n301
  );


  xnor
  g523
  (
    n506,
    n423,
    n414
  );


  nand
  g524
  (
    n505,
    n386,
    n337
  );


  nand
  g525
  (
    n467,
    n426,
    n417
  );


  xnor
  g526
  (
    n542,
    n411,
    n391
  );


  or
  g527
  (
    n549,
    n395,
    n378
  );


  and
  g528
  (
    n534,
    n346,
    n397
  );


  nand
  g529
  (
    n591,
    n412,
    n424
  );


  nand
  g530
  (
    KeyWire_0_9,
    n346,
    n291
  );


  and
  g531
  (
    n517,
    n347,
    n344
  );


  nand
  g532
  (
    n512,
    n441,
    n316
  );


  xor
  g533
  (
    n539,
    n362,
    n282
  );


  nor
  g534
  (
    n593,
    n295,
    n352
  );


  xor
  g535
  (
    n607,
    n371,
    n407
  );


  xor
  g536
  (
    n568,
    n342,
    n313
  );


  or
  g537
  (
    KeyWire_0_12,
    n338,
    n432
  );


  and
  g538
  (
    n605,
    n344,
    n395
  );


  nor
  g539
  (
    n476,
    n454,
    n390
  );


  nand
  g540
  (
    n608,
    n327,
    n438
  );


  and
  g541
  (
    n520,
    n387,
    n441
  );


  xor
  g542
  (
    n601,
    n433,
    n405
  );


  nor
  g543
  (
    n609,
    n387,
    n324
  );


  or
  g544
  (
    n524,
    n431,
    n365
  );


  xor
  g545
  (
    n526,
    n339,
    n312
  );


  or
  g546
  (
    n477,
    n350,
    n413
  );


  xor
  g547
  (
    n475,
    n369,
    n348
  );


  and
  g548
  (
    n513,
    n273,
    n416
  );


  and
  g549
  (
    n590,
    n351,
    n393
  );


  nor
  g550
  (
    n560,
    n398,
    n409
  );


  nor
  g551
  (
    n468,
    n377,
    n339
  );


  and
  g552
  (
    n519,
    n436,
    n442
  );


  xnor
  g553
  (
    n551,
    n372,
    n375
  );


  nand
  g554
  (
    n606,
    n329,
    n425
  );


  xnor
  g555
  (
    n559,
    n405,
    n375
  );


  nor
  g556
  (
    n570,
    n283,
    n299
  );


  nand
  g557
  (
    n581,
    n386,
    n423
  );


  xnor
  g558
  (
    n485,
    n449,
    n435
  );


  and
  g559
  (
    n600,
    n280,
    n341
  );


  nand
  g560
  (
    n464,
    n300,
    n355
  );


  and
  g561
  (
    n580,
    n453,
    n373
  );


  xnor
  g562
  (
    n599,
    n398,
    n434
  );


  nor
  g563
  (
    n538,
    n340,
    n450
  );


  xnor
  g564
  (
    n592,
    n345,
    n374
  );


  nor
  g565
  (
    n472,
    n409,
    n357
  );


  or
  g566
  (
    n571,
    n439,
    n391
  );


  nor
  g567
  (
    n558,
    n428,
    n426
  );


  xnor
  g568
  (
    KeyWire_0_18,
    n440,
    n433
  );


  nand
  g569
  (
    n595,
    n370,
    n333
  );


  xor
  g570
  (
    n535,
    n415,
    n400
  );


  nand
  g571
  (
    n489,
    n410,
    n368
  );


  and
  g572
  (
    n462,
    n364,
    n425
  );


  or
  g573
  (
    n547,
    n397,
    n345
  );


  nand
  g574
  (
    n518,
    n356,
    n348
  );


  nand
  g575
  (
    n474,
    n403,
    n362
  );


  nor
  g576
  (
    n527,
    n371,
    n380
  );


  nor
  g577
  (
    n492,
    n355,
    n324
  );


  or
  g578
  (
    n487,
    n400,
    n388
  );


  and
  g579
  (
    n575,
    n414,
    n444
  );


  xor
  g580
  (
    n550,
    n319,
    n359
  );


  nand
  g581
  (
    n486,
    n376,
    n331
  );


  and
  g582
  (
    n546,
    n341,
    n365
  );


  xnor
  g583
  (
    n579,
    n349,
    n335
  );


  nand
  g584
  (
    n514,
    n429,
    n422
  );


  nand
  g585
  (
    n634,
    n544,
    n556,
    n513,
    n485
  );


  and
  g586
  (
    n622,
    n525,
    n463,
    n553,
    n527
  );


  or
  g587
  (
    n621,
    n572,
    n573,
    n517,
    n557
  );


  nand
  g588
  (
    n639,
    n523,
    n563,
    n497,
    n474
  );


  xor
  g589
  (
    n629,
    n467,
    n535,
    n516,
    n464
  );


  nand
  g590
  (
    n636,
    n462,
    n502,
    n548,
    n461
  );


  or
  g591
  (
    n624,
    n560,
    n514,
    n511,
    n489
  );


  and
  g592
  (
    n633,
    n490,
    n532,
    n540,
    n515
  );


  or
  g593
  (
    n640,
    n479,
    n475,
    n480,
    n472
  );


  nand
  g594
  (
    n627,
    n471,
    n547,
    n530,
    n566
  );


  or
  g595
  (
    n620,
    n512,
    n550,
    n486,
    n508
  );


  xnor
  g596
  (
    n643,
    n487,
    n478,
    n470,
    n529
  );


  or
  g597
  (
    n632,
    n526,
    n507,
    n466,
    n509
  );


  xnor
  g598
  (
    n626,
    n518,
    n546,
    n542,
    n500
  );


  or
  g599
  (
    n635,
    n558,
    n476,
    n537,
    n571
  );


  xor
  g600
  (
    n619,
    n545,
    n481,
    n567,
    n522
  );


  nor
  g601
  (
    n630,
    n504,
    n573,
    n571,
    n565
  );


  or
  g602
  (
    n631,
    n506,
    n482,
    n503,
    n465
  );


  nor
  g603
  (
    n623,
    n496,
    n568,
    n572,
    n488
  );


  xnor
  g604
  (
    n641,
    n483,
    n536,
    n562,
    n569
  );


  xnor
  g605
  (
    n628,
    n477,
    n469,
    n494,
    n538
  );


  xor
  g606
  (
    n646,
    n499,
    n541,
    n524,
    n552
  );


  xor
  g607
  (
    n625,
    n520,
    n539,
    n492,
    n498
  );


  nor
  g608
  (
    n642,
    n510,
    n569,
    n519,
    n551
  );


  or
  g609
  (
    n647,
    n534,
    n495,
    n570,
    n501
  );


  nand
  g610
  (
    n644,
    n554,
    n555,
    n568,
    n491
  );


  xor
  g611
  (
    n618,
    n561,
    n549,
    n559,
    n570
  );


  or
  g612
  (
    n637,
    n564,
    n533,
    n543,
    n521
  );


  nor
  g613
  (
    n638,
    n473,
    n505,
    n484,
    n493
  );


  and
  g614
  (
    n645,
    n468,
    n531,
    n567,
    n528
  );


  buf
  g615
  (
    n657,
    n639
  );


  buf
  g616
  (
    n656,
    n642
  );


  not
  g617
  (
    n650,
    n644
  );


  not
  g618
  (
    n652,
    n640
  );


  buf
  g619
  (
    n655,
    n643
  );


  not
  g620
  (
    n648,
    n641
  );


  not
  g621
  (
    n653,
    n645
  );


  not
  g622
  (
    n651,
    n638
  );


  not
  g623
  (
    n649,
    n646
  );


  not
  g624
  (
    n654,
    n647
  );


  buf
  g625
  (
    n658,
    n270
  );


  buf
  g626
  (
    n661,
    n270
  );


  buf
  g627
  (
    n685,
    n457
  );


  not
  g628
  (
    n664,
    n653
  );


  buf
  g629
  (
    n686,
    n574
  );


  buf
  g630
  (
    n677,
    n656
  );


  not
  g631
  (
    n666,
    n656
  );


  not
  g632
  (
    n689,
    n651
  );


  buf
  g633
  (
    n672,
    n654
  );


  not
  g634
  (
    n695,
    n271
  );


  buf
  g635
  (
    n684,
    n27
  );


  not
  g636
  (
    n674,
    n458
  );


  buf
  g637
  (
    n669,
    n26
  );


  not
  g638
  (
    n668,
    n652
  );


  buf
  g639
  (
    n667,
    n649
  );


  not
  g640
  (
    n671,
    n654
  );


  not
  g641
  (
    n681,
    n456
  );


  buf
  g642
  (
    n690,
    n648
  );


  buf
  g643
  (
    n679,
    n651
  );


  not
  g644
  (
    n678,
    n654
  );


  not
  g645
  (
    n660,
    n29
  );


  not
  g646
  (
    n694,
    n459
  );


  not
  g647
  (
    n670,
    n648
  );


  buf
  g648
  (
    n662,
    n457
  );


  buf
  g649
  (
    n659,
    n657
  );


  buf
  g650
  (
    n687,
    n269
  );


  nand
  g651
  (
    n673,
    n27,
    n648,
    n657,
    n650
  );


  xnor
  g652
  (
    n665,
    n650,
    n27,
    n455,
    n456
  );


  xnor
  g653
  (
    n693,
    n656,
    n655,
    n648,
    n652
  );


  and
  g654
  (
    n676,
    n649,
    n269,
    n651,
    n655
  );


  and
  g655
  (
    n675,
    n657,
    n26,
    n28,
    n649
  );


  or
  g656
  (
    n683,
    n652,
    n271,
    n270,
    n653
  );


  xor
  g657
  (
    n680,
    n649,
    n650,
    n28
  );


  xor
  g658
  (
    n682,
    n459,
    n27,
    n654,
    n655
  );


  nor
  g659
  (
    n691,
    n653,
    n652,
    n269,
    n574
  );


  and
  g660
  (
    n663,
    n270,
    n653,
    n28
  );


  or
  g661
  (
    n692,
    n656,
    n269,
    n651,
    n29
  );


  xor
  g662
  (
    n688,
    n657,
    n655,
    n458,
    n29
  );


  not
  g663
  (
    n699,
    n662
  );


  not
  g664
  (
    n713,
    n669
  );


  buf
  g665
  (
    n712,
    n671
  );


  not
  g666
  (
    n714,
    n665
  );


  buf
  g667
  (
    n708,
    n667
  );


  buf
  g668
  (
    n700,
    n668
  );


  buf
  g669
  (
    n710,
    n658
  );


  buf
  g670
  (
    n696,
    n668
  );


  buf
  g671
  (
    n704,
    n663
  );


  not
  g672
  (
    n709,
    n659
  );


  or
  g673
  (
    n697,
    n658,
    n670,
    n661,
    n664
  );


  or
  g674
  (
    n706,
    n659,
    n659,
    n663,
    n668
  );


  xor
  g675
  (
    n715,
    n658,
    n661,
    n664,
    n666
  );


  or
  g676
  (
    n705,
    n659,
    n671,
    n662,
    n661
  );


  xnor
  g677
  (
    n703,
    n665,
    n660,
    n661
  );


  or
  g678
  (
    n716,
    n662,
    n663,
    n658,
    n665
  );


  nand
  g679
  (
    n707,
    n665,
    n666,
    n668,
    n667
  );


  xor
  g680
  (
    n702,
    n667,
    n669,
    n664
  );


  xnor
  g681
  (
    n711,
    n664,
    n662,
    n670
  );


  or
  g682
  (
    n701,
    n660,
    n663,
    n667,
    n670
  );


  xnor
  g683
  (
    n698,
    n669,
    n660,
    n666
  );


  xnor
  g684
  (
    n735,
    n695,
    n704
  );


  nor
  g685
  (
    n728,
    n674,
    n711,
    n675,
    n692
  );


  nor
  g686
  (
    n752,
    n686,
    n689,
    n692,
    n685
  );


  nand
  g687
  (
    KeyWire_0_14,
    n675,
    n704,
    n701,
    n714
  );


  and
  g688
  (
    KeyWire_0_10,
    n690,
    n681,
    n712,
    n676
  );


  nor
  g689
  (
    n730,
    n680,
    n682,
    n706
  );


  or
  g690
  (
    n732,
    n713,
    n677,
    n680,
    n705
  );


  and
  g691
  (
    n734,
    n684,
    n707,
    n688,
    n691
  );


  nand
  g692
  (
    n747,
    n672,
    n703,
    n691,
    n687
  );


  nand
  g693
  (
    n717,
    n577,
    n697,
    n685,
    n699
  );


  xnor
  g694
  (
    n736,
    n688,
    n685,
    n682,
    n672
  );


  or
  g695
  (
    n733,
    n682,
    n683,
    n674,
    n678
  );


  nor
  g696
  (
    n748,
    n681,
    n693,
    n683,
    n684
  );


  xor
  g697
  (
    n723,
    n673,
    n694,
    n671,
    n708
  );


  or
  g698
  (
    n744,
    n693,
    n698,
    n711,
    n678
  );


  nor
  g699
  (
    n718,
    n716,
    n688,
    n677,
    n675
  );


  nand
  g700
  (
    n746,
    n712,
    n690,
    n695,
    n700
  );


  or
  g701
  (
    n725,
    n695,
    n693,
    n674,
    n689
  );


  nand
  g702
  (
    n740,
    n689,
    n707,
    n680,
    n577
  );


  xnor
  g703
  (
    n751,
    n702,
    n708,
    n679,
    n684
  );


  and
  g704
  (
    n727,
    n715,
    n688,
    n676,
    n694
  );


  or
  g705
  (
    n738,
    n713,
    n714,
    n710,
    n696
  );


  or
  g706
  (
    n739,
    n673,
    n686,
    n678,
    n676
  );


  nand
  g707
  (
    n753,
    n705,
    n675,
    n706,
    n681
  );


  nand
  g708
  (
    n749,
    n680,
    n689,
    n673,
    n575
  );


  nand
  g709
  (
    n722,
    n691,
    n686,
    n677,
    n672
  );


  nor
  g710
  (
    n719,
    n692,
    n679,
    n715
  );


  nand
  g711
  (
    n731,
    n677,
    n695,
    n671,
    n687
  );


  xnor
  g712
  (
    n726,
    n686,
    n678,
    n683,
    n681
  );


  and
  g713
  (
    n741,
    n710,
    n672,
    n679,
    n709
  );


  nor
  g714
  (
    n745,
    n702,
    n694,
    n701,
    n691
  );


  nor
  g715
  (
    n729,
    n690,
    n575,
    n687
  );


  and
  g716
  (
    n737,
    n673,
    n683,
    n685,
    n576
  );


  or
  g717
  (
    n742,
    n684,
    n676,
    n709,
    n698
  );


  or
  g718
  (
    n724,
    n696,
    n703,
    n692,
    n694
  );


  or
  g719
  (
    n721,
    n716,
    n693,
    n576,
    n690
  );


  xor
  g720
  (
    n743,
    n674,
    n700,
    n697,
    n699
  );


  nand
  g721
  (
    n771,
    n580,
    n726,
    n584,
    n728
  );


  or
  g722
  (
    n765,
    n723,
    n581,
    n731
  );


  xnor
  g723
  (
    n770,
    n720,
    n583,
    n719,
    n727
  );


  xnor
  g724
  (
    n762,
    n718,
    n721,
    n725,
    n726
  );


  nor
  g725
  (
    n763,
    n717,
    n720,
    n579,
    n722
  );


  xnor
  g726
  (
    n761,
    n719,
    n722,
    n723,
    n579
  );


  xnor
  g727
  (
    n769,
    n725,
    n717,
    n724,
    n731
  );


  and
  g728
  (
    n755,
    n718,
    n727,
    n729
  );


  xnor
  g729
  (
    n754,
    n719,
    n584,
    n578,
    n717
  );


  xnor
  g730
  (
    n756,
    n582,
    n730,
    n723,
    n731
  );


  xor
  g731
  (
    n760,
    n728,
    n728,
    n720,
    n578
  );


  xor
  g732
  (
    n768,
    n726,
    n723,
    n725,
    n730
  );


  nor
  g733
  (
    n758,
    n727,
    n717,
    n585,
    n724
  );


  xnor
  g734
  (
    n757,
    n730,
    n726,
    n719,
    n718
  );


  nor
  g735
  (
    n772,
    n724,
    n583,
    n718,
    n729
  );


  nor
  g736
  (
    n767,
    n722,
    n728,
    n729,
    n582
  );


  nand
  g737
  (
    n766,
    n585,
    n725,
    n721
  );


  and
  g738
  (
    n764,
    n730,
    n731,
    n722,
    n721
  );


  and
  g739
  (
    n759,
    n724,
    n720,
    n729,
    n580
  );


  xnor
  g740
  (
    n784,
    n772,
    n755,
    n737,
    n752
  );


  xnor
  g741
  (
    n776,
    n740,
    n732,
    n766
  );


  xor
  g742
  (
    n800,
    n753,
    n741,
    n769,
    n770
  );


  nor
  g743
  (
    n783,
    n737,
    n749,
    n746,
    n753
  );


  or
  g744
  (
    n792,
    n758,
    n737,
    n748,
    n772
  );


  xnor
  g745
  (
    n804,
    n765,
    n770,
    n734,
    n742
  );


  xnor
  g746
  (
    n790,
    n754,
    n741,
    n733,
    n763
  );


  nor
  g747
  (
    n793,
    n742,
    n746,
    n743,
    n764
  );


  xor
  g748
  (
    n774,
    n747,
    n762,
    n771,
    n743
  );


  and
  g749
  (
    n803,
    n770,
    n733,
    n754
  );


  xor
  g750
  (
    n791,
    n734,
    n760,
    n736,
    n750
  );


  nand
  g751
  (
    n789,
    n768,
    n764,
    n755
  );


  or
  g752
  (
    KeyWire_0_23,
    n756,
    n742,
    n748,
    n768
  );


  xnor
  g753
  (
    n788,
    n740,
    n767,
    n738,
    n751
  );


  nand
  g754
  (
    n805,
    n745,
    n748,
    n769,
    n747
  );


  nor
  g755
  (
    n809,
    n753,
    n744,
    n758,
    n735
  );


  nand
  g756
  (
    n778,
    n760,
    n769,
    n765,
    n764
  );


  or
  g757
  (
    n806,
    n768,
    n739,
    n735,
    n736
  );


  nor
  g758
  (
    n798,
    n737,
    n738,
    n750,
    n762
  );


  and
  g759
  (
    n808,
    n762,
    n740,
    n771,
    n751
  );


  nor
  g760
  (
    n781,
    n765,
    n767,
    n752,
    n746
  );


  xor
  g761
  (
    n775,
    n767,
    n765,
    n743,
    n771
  );


  or
  g762
  (
    n797,
    n739,
    n739,
    n743,
    n750
  );


  xor
  g763
  (
    n807,
    n749,
    n763,
    n744,
    n752
  );


  and
  g764
  (
    n780,
    n732,
    n757,
    n761,
    n763
  );


  and
  g765
  (
    n795,
    n744,
    n738,
    n732,
    n733
  );


  xnor
  g766
  (
    n782,
    n738,
    n749,
    n741,
    n750
  );


  or
  g767
  (
    n785,
    n766,
    n768,
    n742,
    n746
  );


  xor
  g768
  (
    n779,
    n751,
    n772,
    n763,
    n745
  );


  nor
  g769
  (
    n802,
    n757,
    n741,
    n747,
    n740
  );


  and
  g770
  (
    n786,
    n756,
    n735,
    n770,
    n749
  );


  xnor
  g771
  (
    n787,
    n762,
    n752,
    n759,
    n745
  );


  and
  g772
  (
    n801,
    n748,
    n734,
    n766,
    n751
  );


  nor
  g773
  (
    n773,
    n772,
    n747,
    n767,
    n744
  );


  xnor
  g774
  (
    n799,
    n745,
    n736,
    n769,
    n759
  );


  xnor
  g775
  (
    n777,
    n761,
    n753,
    n739,
    n736
  );


  nand
  g776
  (
    n796,
    n732,
    n771,
    n735,
    n734
  );


  buf
  g777
  (
    n817,
    n803
  );


  buf
  g778
  (
    n819,
    n801
  );


  buf
  g779
  (
    KeyWire_0_17,
    n800
  );


  buf
  g780
  (
    n836,
    n773
  );


  buf
  g781
  (
    n828,
    n803
  );


  buf
  g782
  (
    n815,
    n586
  );


  buf
  g783
  (
    n830,
    n779
  );


  buf
  g784
  (
    n839,
    n781
  );


  buf
  g785
  (
    n813,
    n776
  );


  not
  g786
  (
    n831,
    n589
  );


  not
  g787
  (
    n846,
    n776
  );


  not
  g788
  (
    n833,
    n586
  );


  not
  g789
  (
    n822,
    n797
  );


  not
  g790
  (
    n818,
    n802
  );


  not
  g791
  (
    n844,
    n782
  );


  not
  g792
  (
    n814,
    n779
  );


  buf
  g793
  (
    n826,
    n790
  );


  xnor
  g794
  (
    n820,
    n806,
    n804,
    n793
  );


  nor
  g795
  (
    n823,
    n799,
    n798,
    n786,
    n587
  );


  xnor
  g796
  (
    n812,
    n807,
    n802,
    n787,
    n588
  );


  xnor
  g797
  (
    KeyWire_0_25,
    n805,
    n798,
    n807,
    n784
  );


  and
  g798
  (
    n811,
    n804,
    n780,
    n590,
    n782
  );


  and
  g799
  (
    n840,
    n777,
    n775,
    n781,
    n780
  );


  nor
  g800
  (
    n810,
    n788,
    n791,
    n799,
    n805
  );


  and
  g801
  (
    KeyWire_0_16,
    n796,
    n796,
    n775,
    n807
  );


  xnor
  g802
  (
    n835,
    n800,
    n808,
    n784,
    n786
  );


  and
  g803
  (
    n825,
    n806,
    n777,
    n802,
    n808
  );


  and
  g804
  (
    n821,
    n589,
    n783,
    n591,
    n778
  );


  xor
  g805
  (
    n837,
    n800,
    n803,
    n806,
    n591
  );


  xnor
  g806
  (
    n838,
    n783,
    n799,
    n806,
    n789
  );


  nor
  g807
  (
    n845,
    n791,
    n789,
    n799,
    n801
  );


  or
  g808
  (
    n841,
    n788,
    n590,
    n796,
    n798
  );


  xnor
  g809
  (
    n848,
    n795,
    n774,
    n792,
    n803
  );


  nand
  g810
  (
    n816,
    n793,
    n792,
    n801,
    n800
  );


  and
  g811
  (
    n829,
    n801,
    n785,
    n794,
    n802
  );


  and
  g812
  (
    n847,
    n807,
    n790,
    n804,
    n798
  );


  nor
  g813
  (
    n849,
    n787,
    n797,
    n805
  );


  nand
  g814
  (
    n834,
    n588,
    n805,
    n804,
    n794
  );


  or
  g815
  (
    n824,
    n774,
    n797,
    n795,
    n773
  );


  and
  g816
  (
    n842,
    n587,
    n778,
    n785,
    n796
  );


  and
  g817
  (
    n864,
    n820,
    n821,
    n822,
    n819
  );


  nor
  g818
  (
    n868,
    n822,
    n811,
    n828,
    n809
  );


  nor
  g819
  (
    n854,
    n825,
    n809,
    n821,
    n811
  );


  xnor
  g820
  (
    n857,
    n824,
    n811,
    n813,
    n829
  );


  xor
  g821
  (
    n850,
    n822,
    n825,
    n814,
    n810
  );


  nand
  g822
  (
    n852,
    n823,
    n595,
    n815,
    n594
  );


  nor
  g823
  (
    n872,
    n592,
    n817,
    n816,
    n825
  );


  or
  g824
  (
    n861,
    n594,
    n817,
    n823,
    n827
  );


  or
  g825
  (
    n862,
    n821,
    n824,
    n823,
    n809
  );


  or
  g826
  (
    n859,
    n810,
    n820,
    n826,
    n595
  );


  nor
  g827
  (
    n866,
    n815,
    n829,
    n827,
    n828
  );


  xnor
  g828
  (
    n863,
    n810,
    n815,
    n814,
    n593
  );


  xor
  g829
  (
    n871,
    n830,
    n820,
    n818,
    n829
  );


  and
  g830
  (
    n855,
    n812,
    n826,
    n813,
    n830
  );


  xor
  g831
  (
    n860,
    n828,
    n818,
    n808,
    n593
  );


  or
  g832
  (
    n873,
    n814,
    n814,
    n819,
    n817
  );


  or
  g833
  (
    n856,
    n815,
    n809,
    n813,
    n824
  );


  nor
  g834
  (
    n867,
    n824,
    n812,
    n810,
    n811
  );


  xnor
  g835
  (
    n869,
    n827,
    n818,
    n821,
    n812
  );


  xnor
  g836
  (
    n853,
    n826,
    n828,
    n816,
    n829
  );


  or
  g837
  (
    n858,
    n813,
    n816,
    n823,
    n817
  );


  xor
  g838
  (
    n851,
    n812,
    n819,
    n825,
    n808
  );


  xnor
  g839
  (
    n865,
    n827,
    n592,
    n816,
    n820
  );


  xor
  g840
  (
    n870,
    n826,
    n822,
    n819,
    n818
  );


  not
  g841
  (
    n879,
    n831
  );


  buf
  g842
  (
    n904,
    n848
  );


  buf
  g843
  (
    n889,
    n846
  );


  buf
  g844
  (
    n890,
    n839
  );


  buf
  g845
  (
    n932,
    n851
  );


  buf
  g846
  (
    n876,
    n833
  );


  buf
  g847
  (
    n919,
    n873
  );


  not
  g848
  (
    n880,
    n873
  );


  not
  g849
  (
    n896,
    n854
  );


  not
  g850
  (
    n924,
    n865
  );


  not
  g851
  (
    n888,
    n860
  );


  not
  g852
  (
    n900,
    n861
  );


  not
  g853
  (
    n914,
    n834
  );


  buf
  g854
  (
    n884,
    n856
  );


  not
  g855
  (
    n905,
    n834
  );


  not
  g856
  (
    n917,
    n835
  );


  buf
  g857
  (
    n931,
    n862
  );


  not
  g858
  (
    n911,
    n861
  );


  buf
  g859
  (
    n927,
    n841
  );


  buf
  g860
  (
    n925,
    n859
  );


  buf
  g861
  (
    n883,
    n844
  );


  not
  g862
  (
    n908,
    n841
  );


  not
  g863
  (
    n899,
    n845
  );


  buf
  g864
  (
    n874,
    n841
  );


  not
  g865
  (
    n922,
    n872
  );


  not
  g866
  (
    n921,
    n842
  );


  buf
  g867
  (
    n886,
    n832
  );


  not
  g868
  (
    n923,
    n847
  );


  buf
  g869
  (
    n934,
    n851
  );


  buf
  g870
  (
    n891,
    n849
  );


  buf
  g871
  (
    n895,
    n858
  );


  nand
  g872
  (
    n875,
    n872,
    n838
  );


  nand
  g873
  (
    n907,
    n853,
    n839,
    n870,
    n835
  );


  xor
  g874
  (
    n916,
    n832,
    n859,
    n858,
    n873
  );


  and
  g875
  (
    n881,
    n870,
    n872,
    n849,
    n843
  );


  nor
  g876
  (
    n933,
    n831,
    n871,
    n599,
    n834
  );


  nor
  g877
  (
    n893,
    n836,
    n844,
    n871,
    n846
  );


  xnor
  g878
  (
    n928,
    n845,
    n842,
    n841,
    n850
  );


  or
  g879
  (
    n892,
    n846,
    n597,
    n856,
    n852
  );


  nor
  g880
  (
    n885,
    n864,
    n867,
    n849,
    n866
  );


  xnor
  g881
  (
    n887,
    n831,
    n837,
    n860,
    n868
  );


  xnor
  g882
  (
    n918,
    n869,
    n867,
    n833,
    n871
  );


  nor
  g883
  (
    n920,
    n852,
    n848,
    n870,
    n863
  );


  and
  g884
  (
    n906,
    n836,
    n843,
    n30
  );


  xor
  g885
  (
    n878,
    n840,
    n833,
    n838,
    n839
  );


  xnor
  g886
  (
    n903,
    n831,
    n845,
    n598
  );


  nor
  g887
  (
    n894,
    n857,
    n848,
    n869,
    n864
  );


  and
  g888
  (
    n930,
    n29,
    n847,
    n846,
    n868
  );


  xor
  g889
  (
    n902,
    n863,
    n835,
    n832
  );


  or
  g890
  (
    n901,
    n867,
    n862,
    n599,
    n847
  );


  nor
  g891
  (
    n912,
    n833,
    n596,
    n849,
    n30
  );


  xnor
  g892
  (
    n926,
    n30,
    n853,
    n837,
    n865
  );


  or
  g893
  (
    n929,
    n873,
    n834,
    n597,
    n872
  );


  nand
  g894
  (
    n897,
    n871,
    n868,
    n855
  );


  xor
  g895
  (
    n910,
    n847,
    n836,
    n840,
    n845
  );


  and
  g896
  (
    n935,
    n842,
    n842,
    n837,
    n844
  );


  xor
  g897
  (
    n915,
    n832,
    n30,
    n850,
    n596
  );


  or
  g898
  (
    n882,
    n868,
    n839,
    n31,
    n843
  );


  nand
  g899
  (
    n898,
    n848,
    n844,
    n830,
    n837
  );


  xor
  g900
  (
    n913,
    n857,
    n869,
    n840
  );


  xnor
  g901
  (
    n909,
    n866,
    n830,
    n867,
    n838
  );


  xor
  g902
  (
    n877,
    n854,
    n840,
    n870,
    n836
  );


  nand
  g903
  (
    n977,
    n933,
    n935,
    n906,
    n887
  );


  nor
  g904
  (
    n971,
    n901,
    n934,
    n883,
    n903
  );


  xor
  g905
  (
    KeyWire_0_31,
    n272,
    n883,
    n913,
    n879
  );


  xnor
  g906
  (
    n996,
    n888,
    n921,
    n879,
    n935
  );


  nor
  g907
  (
    n958,
    n907,
    n917,
    n932
  );


  and
  g908
  (
    n975,
    n887,
    n915,
    n905,
    n889
  );


  or
  g909
  (
    n990,
    n883,
    n889,
    n888,
    n901
  );


  xnor
  g910
  (
    n951,
    n910,
    n889,
    n924,
    n922
  );


  or
  g911
  (
    n955,
    n882,
    n897,
    n920,
    n925
  );


  xnor
  g912
  (
    n945,
    n935,
    n930,
    n921,
    n908
  );


  and
  g913
  (
    n952,
    n897,
    n272,
    n880,
    n924
  );


  and
  g914
  (
    n939,
    n875,
    n890,
    n914,
    n899
  );


  or
  g915
  (
    n944,
    n882,
    n911,
    n933,
    n891
  );


  xor
  g916
  (
    n961,
    n884,
    n920,
    n878,
    n885
  );


  nand
  g917
  (
    n938,
    n932,
    n879,
    n883,
    n875
  );


  xnor
  g918
  (
    n962,
    n877,
    n888,
    n923,
    n896
  );


  xor
  g919
  (
    n981,
    n893,
    n878,
    n884,
    n935
  );


  and
  g920
  (
    n963,
    n884,
    n910,
    n907,
    n903
  );


  and
  g921
  (
    n974,
    n920,
    n905,
    n909,
    n911
  );


  nor
  g922
  (
    n967,
    n919,
    n915,
    n921,
    n911
  );


  xnor
  g923
  (
    n986,
    n903,
    n934,
    n892,
    n930
  );


  xor
  g924
  (
    n946,
    n915,
    n895,
    n875,
    n902
  );


  and
  g925
  (
    n992,
    n912,
    n891,
    n928,
    n901
  );


  xor
  g926
  (
    n983,
    n908,
    n894,
    n895,
    n902
  );


  or
  g927
  (
    n940,
    n913,
    n929,
    n918,
    n878
  );


  and
  g928
  (
    n997,
    n925,
    n894,
    n930,
    n931
  );


  xnor
  g929
  (
    n956,
    n926,
    n882,
    n885,
    n894
  );


  nor
  g930
  (
    n993,
    n890,
    n874,
    n891,
    n924
  );


  nor
  g931
  (
    n950,
    n907,
    n894,
    n895,
    n876
  );


  or
  g932
  (
    n979,
    n899,
    n921,
    n916,
    n881
  );


  and
  g933
  (
    n973,
    n886,
    n891,
    n898,
    n932
  );


  and
  g934
  (
    n969,
    n927,
    n895,
    n881,
    n918
  );


  and
  g935
  (
    n948,
    n931,
    n899,
    n902,
    n917
  );


  or
  g936
  (
    n957,
    n916,
    n880,
    n908,
    n917
  );


  nor
  g937
  (
    n941,
    n900,
    n879,
    n909,
    n924
  );


  xor
  g938
  (
    n972,
    n876,
    n884,
    n901,
    n914
  );


  xnor
  g939
  (
    n968,
    n934,
    n926,
    n915,
    n877
  );


  or
  g940
  (
    n984,
    n874,
    n911,
    n922,
    n930
  );


  or
  g941
  (
    n947,
    n885,
    n900,
    n905,
    n896
  );


  and
  g942
  (
    n980,
    n928,
    n913,
    n919
  );


  xor
  g943
  (
    n978,
    n887,
    n923,
    n922,
    n876
  );


  nand
  g944
  (
    n985,
    n874,
    n898,
    n886,
    n928
  );


  xnor
  g945
  (
    n942,
    n271,
    n900,
    n902,
    n923
  );


  or
  g946
  (
    n991,
    n880,
    n916,
    n933,
    n918
  );


  nor
  g947
  (
    n982,
    n932,
    n887,
    n904,
    n892
  );


  or
  g948
  (
    n995,
    n897,
    n882,
    n934,
    n920
  );


  nor
  g949
  (
    n937,
    n885,
    n931,
    n914,
    n910
  );


  xor
  g950
  (
    n994,
    n900,
    n904,
    n877,
    n908
  );


  nor
  g951
  (
    n988,
    n907,
    n892,
    n874,
    n886
  );


  and
  g952
  (
    n949,
    n923,
    n913,
    n929,
    n890
  );


  nand
  g953
  (
    n954,
    n912,
    n905,
    n928,
    n914
  );


  nor
  g954
  (
    n970,
    n878,
    n922,
    n909,
    n912
  );


  nor
  g955
  (
    n989,
    n927,
    n906,
    n897
  );


  xnor
  g956
  (
    n936,
    n893,
    n929,
    n888,
    n892
  );


  or
  g957
  (
    n964,
    n881,
    n925,
    n904,
    n893
  );


  nand
  g958
  (
    n965,
    n877,
    n881,
    n925,
    n903
  );


  nand
  g959
  (
    n959,
    n926,
    n933,
    n889,
    n876
  );


  nor
  g960
  (
    n966,
    n880,
    n931,
    n918,
    n886
  );


  or
  g961
  (
    n953,
    n912,
    n896,
    n898,
    n899
  );


  xnor
  g962
  (
    n987,
    n909,
    n926,
    n896,
    n893
  );


  and
  g963
  (
    n976,
    n904,
    n927,
    n898,
    n271
  );


  nor
  g964
  (
    n998,
    n890,
    n927,
    n916,
    n906
  );


  and
  g965
  (
    n960,
    n919,
    n910,
    n929,
    n875
  );


  nor
  g966
  (
    n1001,
    n978,
    n959,
    n985,
    n960
  );


  and
  g967
  (
    n1006,
    n957,
    n31,
    n956,
    n966
  );


  or
  g968
  (
    n1003,
    n973,
    n970,
    n971,
    n950
  );


  or
  g969
  (
    n1000,
    n979,
    n990,
    n998,
    n944
  );


  xor
  g970
  (
    n1007,
    n989,
    n974,
    n992,
    n32
  );


  xor
  g971
  (
    n1009,
    n948,
    n938,
    n994,
    n962
  );


  nand
  g972
  (
    n1016,
    n997,
    n961,
    n968,
    n998
  );


  xnor
  g973
  (
    n999,
    n964,
    n995,
    n958,
    n996
  );


  xnor
  g974
  (
    KeyWire_0_7,
    n936,
    n31,
    n946,
    n997
  );


  or
  g975
  (
    n1005,
    n947,
    n983,
    n975,
    n980
  );


  or
  g976
  (
    n1015,
    n949,
    n993,
    n996,
    n952
  );


  nand
  g977
  (
    n1011,
    n943,
    n986,
    n941,
    n982
  );


  and
  g978
  (
    KeyWire_0_29,
    n955,
    n981,
    n965,
    n32
  );


  xor
  g979
  (
    n1014,
    n977,
    n32,
    n972,
    n937
  );


  nor
  g980
  (
    n1010,
    n945,
    n939,
    n984,
    n991
  );


  xor
  g981
  (
    n1004,
    n976,
    n969,
    n953,
    n963
  );


  nand
  g982
  (
    n1008,
    n942,
    n954,
    n967,
    n988
  );


  nand
  g983
  (
    n1002,
    n951,
    n940,
    n31,
    n987
  );


  nand
  g984
  (
    n1026,
    n613,
    n1004,
    n1006,
    n1016
  );


  or
  g985
  (
    n1022,
    n1008,
    n612,
    n1014,
    n604
  );


  xor
  g986
  (
    KeyWire_0_24,
    n1003,
    n612,
    n614,
    n605
  );


  nand
  g987
  (
    n1020,
    n999,
    n1002,
    n1012,
    n601
  );


  or
  g988
  (
    n1027,
    n1015,
    n1009,
    n600,
    n1007
  );


  xnor
  g989
  (
    n1019,
    n607,
    n605,
    n1000,
    n602
  );


  and
  g990
  (
    n1028,
    n1001,
    n603,
    n610,
    n614
  );


  nand
  g991
  (
    n1018,
    n611,
    n608,
    n603,
    n1013
  );


  or
  g992
  (
    n1023,
    n1005,
    n611,
    n1011,
    n1010
  );


  xor
  g993
  (
    n1017,
    n609,
    n606,
    n602
  );


  or
  g994
  (
    n1024,
    n600,
    n604,
    n610,
    n613
  );


  nand
  g995
  (
    n1025,
    n609,
    n607,
    n601,
    n608
  );


  xor
  g996
  (
    n1029,
    n616,
    n1028,
    n615
  );


  nor
  g997
  (
    n1030,
    n1029,
    n32,
    n272,
    n616
  );


  and
  g998
  (
    n1031,
    n272,
    n460,
    n1029
  );


  xor
  g999
  (
    n1032,
    n1030,
    n617,
    n1031
  );


  xor
  KeyGate_0_0
  (
    n483,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n272,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n101,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n280,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n457,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n51,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n42,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1013,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n604,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n473,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n720,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n298,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n544,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n235,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n750,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n43,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n843,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n827,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n557,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n323,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n120,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n335,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n509,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n794,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1021,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n832,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n511,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n300,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n426,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1012,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n331,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n943,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


