// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_301 written by SynthGen on 2021/04/05 11:24:04
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_301 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n836, n835, n2834, n2856, n2809, n2830, n2911, n2926,
 n2945, n2767, n2819, n2917, n2792, n2894, n2838, n2751,
 n2884, n2861, n2824, n3023, n3022, n3021, n3026, n3030,
 n3031, n3028, n3027, n3025, n3029, n3020, n3032, n3024);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n836, n835, n2834, n2856, n2809, n2830, n2911, n2926,
 n2945, n2767, n2819, n2917, n2792, n2894, n2838, n2751,
 n2884, n2861, n2824, n3023, n3022, n3021, n3026, n3030,
 n3031, n3028, n3027, n3025, n3029, n3020, n3032, n3024;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
 n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
 n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
 n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
 n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
 n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
 n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
 n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
 n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
 n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
 n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
 n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
 n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
 n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
 n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
 n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
 n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
 n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
 n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
 n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
 n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
 n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
 n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
 n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
 n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
 n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
 n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
 n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
 n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
 n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
 n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
 n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
 n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
 n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
 n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
 n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
 n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
 n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
 n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
 n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
 n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
 n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
 n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
 n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
 n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
 n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
 n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
 n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
 n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
 n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
 n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
 n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
 n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
 n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
 n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
 n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
 n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
 n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
 n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
 n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
 n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
 n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
 n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
 n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
 n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
 n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
 n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
 n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
 n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
 n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
 n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
 n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
 n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
 n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
 n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
 n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
 n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
 n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
 n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
 n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
 n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
 n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
 n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
 n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
 n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
 n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
 n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
 n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
 n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
 n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
 n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
 n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
 n2747, n2748, n2749, n2750, n2752, n2753, n2754, n2755,
 n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
 n2764, n2765, n2766, n2768, n2769, n2770, n2771, n2772,
 n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
 n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
 n2789, n2790, n2791, n2793, n2794, n2795, n2796, n2797,
 n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
 n2806, n2807, n2808, n2810, n2811, n2812, n2813, n2814,
 n2815, n2816, n2817, n2818, n2820, n2821, n2822, n2823,
 n2825, n2826, n2827, n2828, n2829, n2831, n2832, n2833,
 n2835, n2836, n2837, n2839, n2840, n2841, n2842, n2843,
 n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
 n2852, n2853, n2854, n2855, n2857, n2858, n2859, n2860,
 n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
 n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
 n2878, n2879, n2880, n2881, n2882, n2883, n2885, n2886,
 n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2895,
 n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
 n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2912,
 n2913, n2914, n2915, n2916, n2918, n2919, n2920, n2921,
 n2922, n2923, n2924, n2925, n2927, n2928, n2929, n2930,
 n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
 n2939, n2940, n2941, n2942, n2943, n2944, n2946, n2947,
 n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
 n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
 n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
 n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
 n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
 n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
 n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
 n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
 n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019;

not  g0 (n35, n2);
not  g1 (n33, n1);
buf  g2 (n45, n3);
buf  g3 (n43, n2);
buf  g4 (n44, n4);
buf  g5 (n36, n4);
buf  g6 (n46, n1);
not  g7 (n40, n2);
buf  g8 (n34, n2);
not  g9 (n41, n1);
not  g10 (n38, n1);
buf  g11 (n37, n3);
not  g12 (n42, n3);
not  g13 (n39, n3);
not  g14 (n90, n33);
buf  g15 (n79, n39);
buf  g16 (n59, n40);
not  g17 (n101, n41);
buf  g18 (n84, n39);
not  g19 (n82, n44);
buf  g20 (n53, n44);
buf  g21 (n75, n42);
not  g22 (n74, n39);
not  g23 (n63, n39);
not  g24 (n47, n41);
not  g25 (n97, n33);
buf  g26 (n61, n34);
buf  g27 (n68, n38);
buf  g28 (n78, n43);
not  g29 (n87, n41);
buf  g30 (n98, n46);
not  g31 (n50, n45);
not  g32 (n95, n35);
buf  g33 (n66, n38);
not  g34 (n65, n44);
buf  g35 (n62, n34);
not  g36 (n77, n46);
not  g37 (n76, n38);
buf  g38 (n58, n36);
buf  g39 (n80, n44);
buf  g40 (n51, n35);
buf  g41 (n91, n36);
not  g42 (n83, n43);
not  g43 (n96, n40);
buf  g44 (n86, n42);
buf  g45 (n72, n41);
not  g46 (n92, n35);
buf  g47 (n94, n45);
not  g48 (n102, n34);
not  g49 (n64, n37);
buf  g50 (n99, n37);
buf  g51 (n67, n43);
buf  g52 (n69, n43);
not  g53 (n71, n42);
buf  g54 (n88, n34);
not  g55 (n93, n40);
not  g56 (n48, n42);
not  g57 (n100, n33);
not  g58 (n60, n45);
buf  g59 (n85, n36);
buf  g60 (n55, n37);
buf  g61 (n81, n33);
buf  g62 (n57, n45);
buf  g63 (n52, n38);
not  g64 (n70, n46);
not  g65 (n56, n36);
buf  g66 (n54, n40);
buf  g67 (n73, n46);
not  g68 (n89, n37);
buf  g69 (n49, n35);
not  g70 (n131, n69);
buf  g71 (n136, n11);
buf  g72 (n321, n79);
buf  g73 (n195, n49);
not  g74 (n188, n14);
not  g75 (n175, n28);
not  g76 (n242, n62);
not  g77 (n125, n48);
not  g78 (n116, n56);
buf  g79 (n164, n51);
buf  g80 (n315, n99);
not  g81 (n268, n72);
buf  g82 (n294, n102);
not  g83 (n161, n26);
buf  g84 (n218, n48);
buf  g85 (n222, n88);
buf  g86 (n243, n73);
not  g87 (n182, n82);
not  g88 (n160, n21);
not  g89 (n290, n68);
buf  g90 (n120, n78);
not  g91 (n274, n75);
buf  g92 (n248, n18);
not  g93 (n192, n23);
not  g94 (n185, n72);
buf  g95 (n260, n94);
not  g96 (n305, n66);
not  g97 (n326, n11);
buf  g98 (n264, n9);
not  g99 (n210, n54);
buf  g100 (n133, n49);
buf  g101 (n158, n80);
buf  g102 (n289, n64);
buf  g103 (n267, n25);
not  g104 (n173, n13);
buf  g105 (n270, n78);
buf  g106 (n244, n55);
not  g107 (n127, n20);
not  g108 (n319, n13);
not  g109 (n146, n51);
not  g110 (n278, n31);
not  g111 (n181, n17);
buf  g112 (n186, n23);
buf  g113 (n292, n20);
not  g114 (n130, n65);
buf  g115 (n230, n58);
buf  g116 (n323, n60);
buf  g117 (n107, n72);
buf  g118 (n108, n53);
buf  g119 (n303, n91);
buf  g120 (n214, n6);
not  g121 (n159, n22);
buf  g122 (n145, n50);
not  g123 (n128, n61);
not  g124 (n265, n16);
not  g125 (n257, n10);
not  g126 (n124, n89);
buf  g127 (n311, n68);
buf  g128 (n154, n27);
buf  g129 (n252, n10);
buf  g130 (n203, n68);
buf  g131 (n259, n79);
not  g132 (n201, n98);
not  g133 (n149, n94);
not  g134 (n307, n66);
not  g135 (n152, n70);
not  g136 (n304, n71);
buf  g137 (n122, n7);
not  g138 (n117, n30);
buf  g139 (n314, n4);
not  g140 (n166, n31);
buf  g141 (n282, n19);
not  g142 (n198, n54);
buf  g143 (n151, n84);
not  g144 (n235, n11);
not  g145 (n121, n93);
not  g146 (n273, n87);
not  g147 (n172, n91);
not  g148 (n148, n20);
not  g149 (n299, n76);
buf  g150 (n165, n85);
not  g151 (n232, n72);
not  g152 (n224, n101);
not  g153 (n247, n89);
buf  g154 (n286, n70);
not  g155 (n221, n11);
buf  g156 (n256, n15);
not  g157 (n219, n21);
buf  g158 (n228, n9);
buf  g159 (n212, n81);
buf  g160 (n104, n24);
buf  g161 (n170, n57);
not  g162 (n280, n16);
not  g163 (n324, n79);
not  g164 (n255, n93);
buf  g165 (n313, n70);
buf  g166 (n277, n27);
buf  g167 (n111, n53);
buf  g168 (n291, n93);
buf  g169 (n225, n65);
buf  g170 (n258, n54);
not  g171 (n129, n60);
not  g172 (n246, n75);
buf  g173 (n168, n100);
not  g174 (n254, n77);
not  g175 (n302, n56);
buf  g176 (n295, n100);
not  g177 (n110, n28);
buf  g178 (n223, n18);
buf  g179 (n191, n78);
not  g180 (n276, n77);
buf  g181 (n287, n93);
buf  g182 (n275, n83);
buf  g183 (n113, n92);
not  g184 (n140, n7);
not  g185 (n137, n57);
not  g186 (n251, n10);
buf  g187 (n147, n97);
not  g188 (n157, n25);
buf  g189 (n178, n61);
buf  g190 (n301, n57);
buf  g191 (n320, n92);
buf  g192 (n112, n12);
buf  g193 (n293, n62);
buf  g194 (n153, n86);
buf  g195 (n187, n65);
buf  g196 (n249, n8);
buf  g197 (n213, n102);
not  g198 (n205, n26);
not  g199 (n238, n82);
not  g200 (n163, n101);
buf  g201 (n132, n80);
buf  g202 (n318, n50);
buf  g203 (n123, n98);
buf  g204 (n208, n12);
not  g205 (n176, n82);
buf  g206 (n202, n18);
buf  g207 (n272, n32);
not  g208 (n279, n47);
not  g209 (n240, n7);
buf  g210 (n231, n62);
buf  g211 (n306, n100);
not  g212 (n239, n28);
buf  g213 (n271, n22);
buf  g214 (n150, n79);
buf  g215 (n183, n90);
buf  g216 (n288, n17);
buf  g217 (n262, n83);
not  g218 (n103, n66);
not  g219 (n250, n90);
not  g220 (n322, n95);
not  g221 (n194, n98);
buf  g222 (n215, n12);
buf  g223 (n245, n84);
buf  g224 (n236, n58);
not  g225 (n237, n26);
not  g226 (n162, n50);
buf  g227 (n227, n49);
not  g228 (n126, n64);
buf  g229 (n284, n86);
buf  g230 (n184, n16);
buf  g231 (n144, n86);
not  g232 (n234, n5);
buf  g233 (n109, n18);
not  g234 (n114, n75);
not  g235 (n189, n71);
buf  g236 (n190, n47);
buf  g237 (n216, n59);
buf  g238 (n199, n75);
not  g239 (n312, n71);
not  g240 (n206, n81);
not  g241 (n200, n91);
buf  g242 (n134, n74);
not  g243 (n263, n5);
not  g244 (n142, n96);
buf  g245 (n119, n6);
not  g246 (n143, n76);
buf  g247 (n138, n27);
not  g248 (n309, n69);
not  g249 (n139, n52);
buf  g250 (n217, n53);
buf  g251 (n118, n64);
not  g252 (n297, n76);
buf  g253 (n266, n16);
buf  g254 (n105, n92);
buf  g255 (n296, n83);
or   g256 (n298, n13, n60, n91, n90);
xor  g257 (n141, n31, n101, n17, n73);
nand g258 (n285, n29, n52, n25, n4);
xnor g259 (n226, n13, n25, n73, n88);
and  g260 (n177, n22, n55, n86, n87);
nor  g261 (n229, n21, n67, n97, n64);
or   g262 (n179, n63, n12, n27, n24);
nand g263 (n196, n55, n8, n63, n81);
or   g264 (n204, n70, n47, n95, n8);
nand g265 (n281, n19, n89, n77, n101);
nand g266 (n253, n21, n30, n59, n97);
nand g267 (n241, n23, n62, n78, n5);
xor  g268 (n211, n87, n19, n59, n53);
and  g269 (n233, n99, n99, n10, n63);
xnor g270 (n106, n17, n67, n23, n15);
xor  g271 (n283, n65, n31, n54, n52);
nor  g272 (n174, n22, n63, n9, n29);
xnor g273 (n325, n32, n95, n87, n74);
or   g274 (n310, n14, n76, n49, n102);
nor  g275 (n115, n74, n95, n29, n97);
or   g276 (n220, n15, n32, n50, n88);
xnor g277 (n135, n66, n14, n55, n73);
and  g278 (n269, n20, n51, n26, n57);
and  g279 (n180, n96, n102, n85, n69);
nand g280 (n171, n24, n96, n15, n56);
nor  g281 (n300, n88, n51, n7, n80);
xor  g282 (n197, n61, n6, n59, n80);
nand g283 (n316, n24, n48, n90, n100);
xnor g284 (n317, n84, n96, n5, n32);
or   g285 (n167, n77, n48, n67, n58);
xor  g286 (n209, n82, n81, n61, n28);
xor  g287 (n308, n85, n47, n6, n71);
or   g288 (n261, n58, n99, n8, n98);
nor  g289 (n156, n30, n84, n74, n9);
and  g290 (n155, n56, n19, n30, n52);
nor  g291 (n169, n92, n83, n69, n94);
and  g292 (n207, n67, n14, n94, n85);
xnor g293 (n193, n29, n68, n89, n60);
not  g294 (n659, n243);
not  g295 (n485, n160);
buf  g296 (n540, n231);
buf  g297 (n523, n121);
buf  g298 (n574, n305);
not  g299 (n661, n133);
not  g300 (n682, n120);
not  g301 (n596, n241);
not  g302 (n364, n262);
not  g303 (n627, n176);
not  g304 (n347, n117);
not  g305 (n403, n275);
buf  g306 (n438, n302);
not  g307 (n569, n247);
buf  g308 (n373, n184);
not  g309 (n463, n229);
buf  g310 (n366, n135);
not  g311 (n621, n133);
not  g312 (n631, n135);
not  g313 (n550, n164);
buf  g314 (n418, n195);
buf  g315 (n465, n185);
buf  g316 (n649, n125);
buf  g317 (n422, n265);
not  g318 (n359, n166);
not  g319 (n539, n117);
not  g320 (n332, n162);
not  g321 (n484, n222);
not  g322 (n394, n269);
buf  g323 (n614, n211);
buf  g324 (n608, n159);
buf  g325 (n691, n278);
not  g326 (n491, n157);
not  g327 (n507, n212);
not  g328 (n522, n117);
buf  g329 (n663, n225);
buf  g330 (n449, n263);
buf  g331 (n556, n299);
not  g332 (n527, n109);
not  g333 (n592, n142);
buf  g334 (n428, n124);
buf  g335 (n365, n142);
not  g336 (n693, n291);
not  g337 (n666, n260);
buf  g338 (n562, n310);
buf  g339 (n407, n175);
not  g340 (n679, n238);
buf  g341 (n481, n289);
not  g342 (n599, n258);
not  g343 (n353, n275);
buf  g344 (n391, n244);
not  g345 (n429, n309);
buf  g346 (n678, n148);
buf  g347 (n456, n159);
buf  g348 (n575, n111);
not  g349 (n656, n134);
buf  g350 (n335, n288);
buf  g351 (n541, n119);
buf  g352 (n392, n314);
buf  g353 (n652, n129);
buf  g354 (n681, n169);
not  g355 (n553, n227);
buf  g356 (n367, n115);
buf  g357 (n567, n162);
buf  g358 (n607, n214);
buf  g359 (n483, n183);
buf  g360 (n546, n114);
not  g361 (n447, n151);
buf  g362 (n441, n292);
buf  g363 (n588, n129);
not  g364 (n396, n265);
buf  g365 (n609, n218);
not  g366 (n532, n173);
not  g367 (n606, n196);
buf  g368 (n421, n188);
buf  g369 (n511, n207);
not  g370 (n426, n183);
buf  g371 (n440, n177);
buf  g372 (n338, n134);
not  g373 (n515, n269);
buf  g374 (n343, n164);
buf  g375 (n412, n119);
buf  g376 (n685, n103);
buf  g377 (n328, n298);
not  g378 (n387, n190);
buf  g379 (n439, n157);
not  g380 (n500, n149);
not  g381 (n499, n122);
not  g382 (n459, n251);
not  g383 (n637, n218);
not  g384 (n629, n205);
not  g385 (n572, n136);
buf  g386 (n482, n276);
buf  g387 (n543, n216);
not  g388 (n529, n111);
not  g389 (n424, n215);
not  g390 (n472, n269);
buf  g391 (n657, n202);
not  g392 (n398, n242);
not  g393 (n436, n237);
not  g394 (n686, n198);
not  g395 (n565, n283);
buf  g396 (n602, n254);
buf  g397 (n630, n169);
not  g398 (n535, n203);
buf  g399 (n524, n130);
not  g400 (n677, n242);
not  g401 (n570, n147);
not  g402 (n384, n149);
not  g403 (n698, n264);
buf  g404 (n377, n167);
buf  g405 (n597, n315);
buf  g406 (n390, n283);
buf  g407 (n411, n308);
buf  g408 (n568, n272);
not  g409 (n452, n231);
not  g410 (n494, n110);
buf  g411 (n445, n180);
not  g412 (n497, n124);
buf  g413 (n478, n181);
buf  g414 (n531, n207);
not  g415 (n383, n250);
not  g416 (n382, n120);
not  g417 (n525, n136);
buf  g418 (n549, n145);
buf  g419 (n635, n303);
not  g420 (n669, n107);
not  g421 (n676, n192);
buf  g422 (n405, n244);
buf  g423 (n537, n253);
not  g424 (n351, n217);
not  g425 (n650, n277);
not  g426 (n559, n261);
not  g427 (n598, n131);
xnor g428 (n651, n278, n226, n208);
and  g429 (n643, n205, n236, n156);
nand g430 (n689, n239, n267, n243);
or   g431 (n696, n228, n299, n171);
xnor g432 (n336, n126, n291, n300);
nand g433 (n545, n230, n278, n191);
xor  g434 (n520, n170, n224, n163);
nand g435 (n466, n103, n163, n304);
nor  g436 (n622, n209, n221, n133);
and  g437 (n521, n274, n188, n277);
xor  g438 (n395, n205, n233, n139);
or   g439 (n605, n180, n254, n251);
nand g440 (n516, n110, n200, n220);
nor  g441 (n610, n174, n214, n175);
nor  g442 (n389, n142, n180, n139);
or   g443 (n397, n138, n259, n262);
xnor g444 (n352, n271, n121, n293);
xor  g445 (n446, n260, n272, n200);
and  g446 (n408, n166, n114, n178);
xor  g447 (n542, n248, n231, n191);
or   g448 (n538, n189, n262, n283);
or   g449 (n416, n172, n147, n105);
nor  g450 (n579, n277, n298, n227);
nor  g451 (n348, n192, n158, n216);
xnor g452 (n654, n145, n259, n296);
nor  g453 (n502, n295, n220, n144);
and  g454 (n697, n173, n124, n165);
nor  g455 (n628, n245, n306, n228);
or   g456 (n474, n309, n310, n132);
nand g457 (n356, n315, n128, n224);
and  g458 (n618, n297, n195);
nor  g459 (n477, n214, n312, n213);
xnor g460 (n683, n161, n274, n136);
nand g461 (n340, n110, n288, n240);
nand g462 (n358, n314, n174, n284);
nand g463 (n554, n108, n238, n198);
or   g464 (n379, n201, n251, n268);
and  g465 (n647, n267, n105, n279);
xor  g466 (n415, n248, n282, n226);
nand g467 (n334, n304, n293, n187);
xor  g468 (n638, n191, n301, n125);
or   g469 (n586, n285, n273, n187);
nand g470 (n639, n308, n278, n217);
and  g471 (n413, n280, n313, n270);
nor  g472 (n557, n207, n135, n294);
xor  g473 (n400, n176, n123, n287);
nand g474 (n688, n305, n239, n224);
or   g475 (n528, n106, n300, n230);
nor  g476 (n563, n265, n252, n228);
xor  g477 (n604, n155, n304, n286);
or   g478 (n458, n196, n206, n235);
and  g479 (n694, n184, n112, n160);
nor  g480 (n496, n173, n310, n276);
nor  g481 (n468, n189, n151, n134);
xnor g482 (n615, n297, n286, n153);
xnor g483 (n517, n178, n270, n146);
xor  g484 (n664, n266, n298, n153);
nand g485 (n623, n307, n226, n273);
xnor g486 (n504, n307, n281, n141);
xor  g487 (n514, n270, n196, n234);
nand g488 (n508, n292, n153, n256);
and  g489 (n354, n161, n241, n281);
or   g490 (n393, n178, n131, n300);
nand g491 (n624, n307, n166, n140);
xnor g492 (n626, n160, n208, n211);
or   g493 (n362, n118, n288, n249);
and  g494 (n680, n236, n247, n293);
or   g495 (n658, n227, n208, n139);
and  g496 (n388, n156, n138, n127);
xor  g497 (n488, n260, n120, n121);
and  g498 (n427, n314, n199, n264);
and  g499 (n577, n271, n103, n194);
xor  g500 (n648, n165, n279, n284);
nor  g501 (n330, n289, n194, n186);
nand g502 (n641, n145, n197, n260);
or   g503 (n632, n233, n219, n301);
nand g504 (n699, n313, n273, n289);
nor  g505 (n600, n182, n179, n250);
and  g506 (n595, n105, n219, n108);
or   g507 (n473, n178, n134, n156);
xnor g508 (n489, n168, n113, n157);
or   g509 (n672, n311, n123, n186);
xnor g510 (n479, n209, n244, n272);
or   g511 (n437, n306, n210, n184);
and  g512 (n402, n201, n119, n150);
nand g513 (n547, n191, n243, n255);
xnor g514 (n645, n162, n310, n139);
or   g515 (n555, n112, n198, n164);
xnor g516 (n480, n158, n131, n295);
nor  g517 (n687, n198, n200, n169);
and  g518 (n552, n206, n252, n302);
and  g519 (n566, n240, n206, n160);
or   g520 (n337, n263, n225, n183);
and  g521 (n460, n225, n290, n193);
or   g522 (n594, n248, n235, n150);
or   g523 (n423, n206, n127, n285);
xnor g524 (n616, n275, n120, n233);
xnor g525 (n611, n203, n213, n253);
or   g526 (n573, n118, n303, n159);
and  g527 (n576, n140, n157, n146);
nor  g528 (n692, n199, n112, n171);
and  g529 (n551, n182, n235, n220);
xor  g530 (n518, n186, n108, n179);
xnor g531 (n584, n128, n118, n246);
and  g532 (n432, n230, n294, n177);
xnor g533 (n603, n274, n104, n257);
nand g534 (n385, n304, n106, n264);
nor  g535 (n339, n262, n156, n189);
xor  g536 (n327, n177, n114, n194);
nand g537 (n469, n195, n229, n313);
or   g538 (n589, n155, n121, n131);
xnor g539 (n512, n106, n155, n210);
xor  g540 (n667, n239, n253, n163);
nor  g541 (n329, n167, n216, n112);
nor  g542 (n526, n171, n297, n109);
nand g543 (n560, n282, n308, n242);
nor  g544 (n430, n171, n172, n274);
or   g545 (n417, n213, n108, n140);
xnor g546 (n487, n231, n292, n249);
nor  g547 (n619, n290, n168, n282);
or   g548 (n674, n149, n240, n221);
nor  g549 (n419, n309, n234, n308);
nand g550 (n585, n122, n132, n234);
xnor g551 (n640, n148, n255, n238);
and  g552 (n344, n161, n151, n116);
xnor g553 (n561, n190, n268, n301);
xor  g554 (n675, n137, n254, n187);
or   g555 (n544, n152, n275, n297);
nand g556 (n498, n130, n140, n219);
or   g557 (n475, n261, n271, n245);
xnor g558 (n476, n110, n261, n115);
nand g559 (n444, n265, n215, n246);
xor  g560 (n633, n124, n216, n306);
and  g561 (n457, n223, n232, n237);
xnor g562 (n425, n286, n109, n111);
xor  g563 (n363, n280, n311, n256);
or   g564 (n355, n145, n123, n107);
nor  g565 (n493, n126, n279, n149);
or   g566 (n533, n170, n192, n209);
nand g567 (n453, n172, n220, n138);
nor  g568 (n587, n144, n193, n219);
xor  g569 (n503, n203, n150, n237);
or   g570 (n401, n148, n215, n299);
xnor g571 (n662, n284, n141, n276);
nor  g572 (n369, n199, n184, n256);
or   g573 (n591, n153, n176, n115);
xnor g574 (n349, n221, n212, n239);
or   g575 (n451, n263, n109, n212);
xor  g576 (n668, n127, n122, n141);
and  g577 (n519, n158, n229, n280);
xnor g578 (n653, n181, n243, n246);
and  g579 (n690, n232, n180, n291);
and  g580 (n536, n221, n210, n197);
and  g581 (n461, n225, n287, n252);
xnor g582 (n590, n143, n222, n104);
nand g583 (n660, n263, n175, n289);
nor  g584 (n374, n185, n276, n312);
xor  g585 (n492, n204, n207, n236);
xor  g586 (n464, n127, n128, n267);
xor  g587 (n486, n193, n217, n266);
xor  g588 (n462, n129, n201, n272);
nor  g589 (n448, n144, n204, n197);
xnor g590 (n581, n266, n215, n190);
xor  g591 (n442, n305, n256, n130);
nand g592 (n345, n183, n181, n258);
nand g593 (n564, n204, n117, n294);
or   g594 (n357, n152, n227, n235);
or   g595 (n350, n273, n151, n172);
and  g596 (n582, n213, n129, n179);
or   g597 (n455, n177, n251, n189);
and  g598 (n386, n232, n282, n201);
xnor g599 (n467, n224, n200, n287);
nor  g600 (n578, n285, n202, n271);
and  g601 (n375, n204, n230, n190);
xor  g602 (n414, n113, n208, n255);
nand g603 (n505, n252, n296, n202);
nor  g604 (n371, n266, n106, n254);
xor  g605 (n495, n305, n126, n311);
xor  g606 (n513, n313, n253, n185);
nor  g607 (n454, n107, n174);
or   g608 (n580, n115, n315, n226);
xnor g609 (n410, n154, n138, n264);
xnor g610 (n342, n279, n233, n181);
xnor g611 (n613, n290, n286, n223);
or   g612 (n646, n187, n107, n182);
and  g613 (n636, n259, n249, n133);
xor  g614 (n333, n165, n268, n141);
and  g615 (n625, n188, n250, n291);
nand g616 (n665, n281, n167, n162);
and  g617 (n509, n104, n158, n113);
xnor g618 (n433, n209, n222, n306);
nand g619 (n471, n159, n196, n300);
nand g620 (n404, n296, n152, n132);
or   g621 (n378, n175, n197, n150);
or   g622 (n593, n176, n288, n218);
xor  g623 (n435, n132, n296, n116);
and  g624 (n490, n270, n188, n105);
nor  g625 (n548, n277, n247, n250);
nand g626 (n376, n155, n169, n126);
xnor g627 (n671, n234, n114, n285);
nand g628 (n380, n142, n103, n212);
nand g629 (n510, n229, n295, n280);
xor  g630 (n530, n259, n202, n152);
and  g631 (n368, n248, n214, n194);
or   g632 (n571, n223, n294, n301);
nand g633 (n695, n154, n268, n179);
nand g634 (n341, n163, n257, n143);
nor  g635 (n331, n173, n154, n232);
or   g636 (n506, n284, n203, n168);
and  g637 (n617, n170, n144, n299);
xnor g638 (n634, n257, n143, n193);
xnor g639 (n655, n261, n182, n137);
xor  g640 (n620, n217, n211, n125);
nand g641 (n381, n290, n135, n302);
nor  g642 (n501, n303, n245, n147);
nor  g643 (n360, n258, n116, n211);
nor  g644 (n409, n245, n298, n247);
nand g645 (n443, n186, n292, n244);
and  g646 (n583, n119, n143, n148);
or   g647 (n431, n154, n166, n258);
and  g648 (n406, n287, n303, n113);
xor  g649 (n470, n311, n123, n236);
xor  g650 (n450, n295, n185, n283);
and  g651 (n642, n192, n223, n146);
xnor g652 (n601, n210, n168, n130);
nand g653 (n612, n161, n249, n104);
xor  g654 (n434, n137, n222, n136);
and  g655 (n361, n293, n165, n137);
xnor g656 (n346, n205, n170, n199);
nand g657 (n420, n238, n302, n128);
nor  g658 (n673, n147, n309, n241);
and  g659 (n558, n242, n111, n307);
xnor g660 (n684, n164, n281, n257);
nand g661 (n372, n255, n146, n246);
nor  g662 (n644, n237, n118, n241);
xor  g663 (n534, n267, n122, n125);
nor  g664 (n399, n218, n269, n228);
nand g665 (n370, n312, n314, n240);
and  g666 (n670, n167, n312, n116);
not  g667 (n700, n327);
buf  g668 (n701, n328);
xor  g669 (n709, n317, n317, n316, n315);
and  g670 (n704, n317, n701, n320, n700);
xnor g671 (n703, n320, n321, n319);
xnor g672 (n706, n701, n317, n316, n318);
xor  g673 (n705, n316, n321, n319, n701);
xnor g674 (n707, n318, n701, n700, n319);
xor  g675 (n708, n700, n316, n318, n320);
and  g676 (n702, n319, n318, n700, n320);
buf  g677 (n713, n702);
buf  g678 (n720, n707);
not  g679 (n726, n703);
not  g680 (n710, n702);
not  g681 (n714, n708);
not  g682 (n718, n707);
not  g683 (n716, n704);
buf  g684 (n719, n708);
not  g685 (n712, n705);
not  g686 (n711, n705);
not  g687 (n722, n706);
not  g688 (n724, n709);
buf  g689 (n723, n709);
not  g690 (n721, n707);
buf  g691 (n725, n703);
buf  g692 (n717, n707);
buf  g693 (n729, n706);
buf  g694 (n715, n708);
buf  g695 (n728, n708);
not  g696 (n727, n704);
and  g697 (n745, n551, n371, n722, n715);
xnor g698 (n804, n410, n723, n339, n386);
xnor g699 (n790, n537, n561, n516, n497);
or   g700 (n789, n729, n361, n509, n723);
or   g701 (n791, n407, n425, n409, n524);
or   g702 (n792, n547, n417, n532, n507);
nor  g703 (n750, n391, n345, n719, n430);
or   g704 (n775, n413, n534, n467, n481);
and  g705 (n788, n720, n470, n455, n403);
xor  g706 (n762, n432, n422, n562, n510);
xor  g707 (n739, n718, n727, n544, n471);
nor  g708 (n785, n727, n442, n487, n402);
xnor g709 (n749, n336, n712, n349, n494);
nand g710 (n807, n431, n445, n722, n388);
nand g711 (n767, n500, n394, n726, n486);
and  g712 (n755, n433, n722, n550, n711);
nor  g713 (n748, n530, n367, n513, n727);
nor  g714 (n769, n549, n380, n724, n483);
and  g715 (n760, n458, n463, n563, n716);
or   g716 (n747, n557, n713, n440, n548);
xnor g717 (n780, n713, n415, n715, n517);
and  g718 (n768, n399, n728, n385, n358);
xor  g719 (n798, n721, n480, n560, n717);
nand g720 (n777, n514, n333, n521, n565);
xor  g721 (n752, n721, n533, n419, n460);
nand g722 (n802, n504, n710, n351);
or   g723 (n776, n710, n484, n546, n712);
xnor g724 (n754, n446, n474, n451, n482);
xnor g725 (n786, n365, n395, n334, n447);
nor  g726 (n771, n724, n329, n717, n441);
nor  g727 (n809, n359, n438, n712, n342);
nor  g728 (n746, n376, n729, n356, n363);
nor  g729 (n763, n427, n383, n728, n337);
and  g730 (n806, n392, n475, n508, n536);
xor  g731 (n797, n357, n520, n396, n478);
or   g732 (n736, n477, n722, n526, n725);
or   g733 (n744, n476, n429, n715, n436);
nand g734 (n770, n456, n490, n343, n717);
xor  g735 (n765, n381, n457, n378, n437);
or   g736 (n751, n718, n461, n364, n558);
and  g737 (n774, n728, n439, n531, n713);
xor  g738 (n730, n428, n512, n491, n559);
nor  g739 (n741, n372, n464, n479, n462);
xnor g740 (n773, n408, n714, n720, n347);
xor  g741 (n757, n726, n424, n382, n426);
nand g742 (n766, n450, n555, n404, n718);
nand g743 (n793, n724, n720, n414, n465);
and  g744 (n801, n728, n726, n375, n453);
and  g745 (n759, n389, n459, n353, n539);
xnor g746 (n737, n355, n398, n535, n466);
nand g747 (n734, n529, n331, n449, n711);
or   g748 (n731, n418, n543, n711, n400);
and  g749 (n787, n368, n454, n713, n488);
and  g750 (n732, n352, n452, n554, n729);
nor  g751 (n758, n444, n553, n373, n725);
xor  g752 (n761, n468, n489, n729, n377);
xnor g753 (n782, n726, n370, n350, n397);
xor  g754 (n738, n719, n401, n714, n716);
xor  g755 (n803, n515, n330, n362, n519);
xor  g756 (n756, n719, n721, n435, n725);
and  g757 (n742, n511, n525, n496, n527);
xnor g758 (n783, n335, n716, n538, n469);
nand g759 (n799, n354, n564, n523, n406);
xnor g760 (n778, n721, n411, n340, n540);
nor  g761 (n796, n503, n420, n495, n716);
and  g762 (n808, n360, n393, n718, n542);
xnor g763 (n764, n405, n473, n556, n723);
xnor g764 (n743, n379, n715, n712, n492);
or   g765 (n733, n725, n710, n443, n714);
or   g766 (n740, n714, n568, n341, n720);
nand g767 (n784, n723, n387, n724, n369);
and  g768 (n800, n541, n522, n506, n566);
nand g769 (n772, n412, n421, n552, n346);
xor  g770 (n753, n545, n499, n366, n727);
xnor g771 (n779, n505, n717, n448, n498);
xor  g772 (n795, n332, n416, n501, n423);
xor  g773 (n805, n384, n485, n344, n338);
xnor g774 (n781, n493, n719, n528, n502);
or   g775 (n794, n711, n374, n518, n567);
nor  g776 (n735, n390, n348, n472, n434);
not  g777 (n818, n747);
buf  g778 (n827, n740);
buf  g779 (n824, n736);
not  g780 (n830, n734);
not  g781 (n811, n749);
buf  g782 (n819, n751);
not  g783 (n816, n739);
buf  g784 (n828, n730);
buf  g785 (n825, n742);
not  g786 (n833, n737);
not  g787 (n832, n741);
buf  g788 (n826, n753);
buf  g789 (n814, n735);
buf  g790 (n829, n738);
not  g791 (n815, n748);
buf  g792 (n817, n744);
not  g793 (n812, n731);
buf  g794 (n823, n750);
not  g795 (n821, n745);
not  g796 (n822, n746);
buf  g797 (n813, n743);
buf  g798 (n820, n752);
buf  g799 (n810, n733);
not  g800 (n831, n732);
nor  g801 (n836, n757, n763, n810, n755);
xnor g802 (n834, n759, n754, n811, n758);
or   g803 (n837, n760, n764, n761, n756);
nand g804 (n835, n811, n810, n765, n762);
xor  g805 (n839, n769, n836, n770, n767);
and  g806 (n838, n766, n837, n768, n771);
xnor g807 (n847, n817, n818, n813);
and  g808 (n842, n814, n815, n838);
xor  g809 (n845, n839, n817, n816, n812);
xnor g810 (n841, n816, n816, n813, n815);
nor  g811 (n844, n817, n839, n815, n814);
or   g812 (n840, n839, n814, n816, n817);
xnor g813 (n846, n815, n812, n838, n814);
or   g814 (n843, n839, n818, n838);
not  g815 (n856, n843);
buf  g816 (n867, n846);
not  g817 (n868, n776);
not  g818 (n877, n843);
buf  g819 (n850, n845);
buf  g820 (n879, n843);
not  g821 (n849, n847);
not  g822 (n866, n772);
not  g823 (n852, n846);
not  g824 (n864, n840);
not  g825 (n851, n845);
buf  g826 (n862, n847);
buf  g827 (n863, n774);
buf  g828 (n869, n842);
buf  g829 (n859, n773);
buf  g830 (n858, n840);
buf  g831 (n854, n846);
not  g832 (n848, n841);
buf  g833 (n860, n774);
not  g834 (n874, n842);
not  g835 (n872, n775);
not  g836 (n871, n842);
buf  g837 (n853, n841);
not  g838 (n855, n840);
not  g839 (n857, n843);
not  g840 (n876, n773);
not  g841 (n865, n841);
buf  g842 (n861, n844);
or   g843 (n878, n844, n841, n845);
nand g844 (n873, n846, n847, n775);
and  g845 (n875, n845, n847, n844);
or   g846 (n870, n844, n842, n840);
nand g847 (n911, n855, n848, n780);
xnor g848 (n887, n831, n820, n832);
or   g849 (n893, n779, n830, n851, n848);
or   g850 (n894, n828, n854, n849);
xor  g851 (n895, n571, n821, n858, n573);
or   g852 (n899, n823, n830, n850, n853);
xnor g853 (n886, n861, n855, n821, n824);
or   g854 (n904, n822, n860, n777);
or   g855 (n897, n778, n829, n827, n831);
and  g856 (n900, n823, n863, n853, n857);
xnor g857 (n892, n862, n850, n849);
xnor g858 (n908, n832, n862, n780, n829);
or   g859 (n910, n857, n861, n820, n859);
xor  g860 (n891, n826, n860, n854, n827);
xor  g861 (n882, n857, n832, n824);
xnor g862 (n914, n855, n851, n859, n569);
nand g863 (n884, n856, n822, n862, n826);
or   g864 (n898, n820, n852, n819, n781);
or   g865 (n880, n819, n861, n825, n851);
or   g866 (n888, n854, n827, n862, n831);
nand g867 (n902, n848, n823, n828, n859);
or   g868 (n901, n854, n853, n828, n852);
xnor g869 (n890, n858, n825, n856, n829);
nor  g870 (n913, n859, n819, n820, n858);
and  g871 (n903, n831, n779, n827, n829);
and  g872 (n896, n833, n822, n860, n821);
nand g873 (n906, n778, n782, n852, n819);
nand g874 (n885, n821, n822, n576, n782);
or   g875 (n905, n858, n825, n852, n824);
xnor g876 (n909, n860, n830, n848, n851);
and  g877 (n912, n850, n849, n823, n856);
nor  g878 (n883, n574, n857, n828, n781);
xor  g879 (n889, n861, n856, n572, n776);
and  g880 (n881, n825, n826, n830, n855);
or   g881 (n907, n570, n575, n826, n853);
nor  g882 (n935, n890, n614, n881, n601);
nand g883 (n915, n615, n625, n616, n608);
and  g884 (n932, n612, n786, n577, n603);
xor  g885 (n929, n600, n622, n883, n597);
nand g886 (n918, n783, n885, n611, n889);
nand g887 (n919, n605, n899, n880, n594);
nand g888 (n921, n587, n784, n602, n599);
nor  g889 (n927, n590, n579, n897, n584);
nor  g890 (n924, n610, n618, n595, n896);
nor  g891 (n930, n626, n788, n786, n606);
nand g892 (n931, n892, n624, n789, n581);
xnor g893 (n928, n607, n788, n598, n787);
and  g894 (n922, n585, n785, n783, n893);
xnor g895 (n920, n580, n609, n623, n785);
and  g896 (n926, n891, n888, n882, n886);
nand g897 (n923, n583, n621, n596, n784);
xor  g898 (n917, n895, n578, n887, n588);
nand g899 (n916, n604, n589, n617, n593);
xnor g900 (n934, n592, n894, n582, n898);
and  g901 (n933, n900, n884, n591, n619);
xor  g902 (n925, n586, n787, n613, n620);
not  g903 (n939, n915);
buf  g904 (n943, n916);
not  g905 (n936, n915);
buf  g906 (n938, n916);
buf  g907 (n941, n915);
buf  g908 (n940, n916);
not  g909 (n937, n915);
buf  g910 (n942, n916);
not  g911 (n945, n863);
xor  g912 (n948, n867, n790, n789, n911);
or   g913 (n963, n873, n870, n798, n876);
nand g914 (n950, n865, n875, n874);
or   g915 (n967, n872, n864, n939, n791);
and  g916 (n972, n943, n908, n796, n938);
xor  g917 (n961, n914, n864, n794, n877);
nor  g918 (n954, n875, n937, n792, n941);
xor  g919 (n959, n910, n797, n790, n871);
xnor g920 (n973, n936, n865, n866, n941);
nor  g921 (n958, n877, n941, n876, n936);
xor  g922 (n955, n905, n909, n943, n941);
or   g923 (n947, n870, n871, n867);
or   g924 (n957, n936, n792, n873, n943);
or   g925 (n949, n940, n936, n799, n797);
nor  g926 (n975, n869, n868, n794, n942);
and  g927 (n953, n866, n942, n940, n791);
and  g928 (n956, n865, n901, n864, n869);
or   g929 (n965, n875, n912, n939, n940);
or   g930 (n964, n864, n876, n865, n793);
and  g931 (n960, n798, n868, n937, n871);
nand g932 (n968, n938, n903, n868, n795);
xor  g933 (n971, n873, n869, n866);
and  g934 (n944, n874, n873, n938, n868);
xnor g935 (n970, n871, n796, n904, n869);
nand g936 (n969, n940, n939, n874);
xnor g937 (n966, n870, n902, n875, n872);
xnor g938 (n946, n877, n937, n913, n906);
and  g939 (n974, n872, n872, n876, n942);
xor  g940 (n951, n937, n795, n943, n877);
xnor g941 (n952, n867, n907, n870, n863);
nand g942 (n962, n938, n863, n942, n793);
nand g943 (n977, n918, n919);
xnor g944 (n984, n919, n917);
nand g945 (n979, n945, n919, n922, n918);
or   g946 (n983, n921, n923, n917, n920);
nor  g947 (n985, n948, n918, n945, n917);
xnor g948 (n982, n948, n946, n919, n917);
nor  g949 (n980, n923, n922, n944);
and  g950 (n976, n920, n922);
nor  g951 (n978, n946, n947, n920, n921);
nand g952 (n981, n918, n921, n947);
and  g953 (n989, n800, n803, n977, n804);
nor  g954 (n986, n803, n976, n805, n800);
or   g955 (n987, n977, n799, n804, n801);
or   g956 (n988, n801, n802, n978);
xor  g957 (n992, n951, n989, n950, n949);
xnor g958 (n990, n952, n629, n953, n988);
nand g959 (n991, n989, n952, n987, n953);
and  g960 (n993, n950, n954, n628, n951);
and  g961 (n994, n954, n949, n986, n627);
xor  g962 (n1002, n983, n990, n636, n992);
xnor g963 (n1005, n633, n992, n962, n982);
nand g964 (n1006, n964, n960, n630, n968);
and  g965 (n1009, n965, n958, n979, n983);
xnor g966 (n1012, n964, n982, n993, n985);
xor  g967 (n996, n994, n991, n993, n992);
nor  g968 (n1013, n833, n981, n980);
nor  g969 (n995, n994, n967, n957, n961);
nor  g970 (n1010, n634, n992, n993, n972);
xnor g971 (n1004, n993, n984, n959, n961);
xnor g972 (n1003, n971, n981, n966, n635);
nor  g973 (n999, n963, n631, n985, n632);
nor  g974 (n998, n994, n994, n991, n979);
nand g975 (n997, n967, n991, n978, n990);
and  g976 (n1014, n956, n990, n965, n962);
xnor g977 (n1001, n957, n968, n970, n971);
nand g978 (n1007, n833, n991, n958, n637);
xor  g979 (n1000, n960, n956, n955);
nor  g980 (n1011, n984, n959, n966, n969);
xnor g981 (n1008, n969, n970, n963, n990);
not  g982 (n1027, n923);
not  g983 (n1024, n1000);
not  g984 (n1019, n999);
buf  g985 (n1022, n924);
not  g986 (n1026, n923);
not  g987 (n1023, n1000);
not  g988 (n1021, n998);
not  g989 (n1015, n996);
buf  g990 (n1020, n995);
buf  g991 (n1018, n997);
not  g992 (n1025, n999);
buf  g993 (n1017, n995);
nand g994 (n1016, n1001, n996, n997, n998);
not  g995 (n1040, n1024);
not  g996 (n1028, n653);
not  g997 (n1034, n640);
not  g998 (n1042, n1026);
buf  g999 (n1044, n1025);
not  g1000 (n1037, n639);
and  g1001 (n1039, n1022, n641, n1023);
or   g1002 (n1032, n323, n324, n1027, n1020);
nor  g1003 (n1038, n1025, n324, n642, n646);
xnor g1004 (n1035, n647, n324, n322, n1024);
nand g1005 (n1030, n650, n323, n321, n648);
and  g1006 (n1029, n652, n638, n651, n644);
nand g1007 (n1033, n1021, n323, n645, n1016);
and  g1008 (n1031, n1019, n1017, n805, n1026);
xor  g1009 (n1041, n323, n654, n1015, n322);
nand g1010 (n1043, n324, n649, n1027, n643);
xnor g1011 (n1036, n1018, n325, n322);
buf  g1012 (n1071, n1037);
buf  g1013 (n1059, n1032);
not  g1014 (n1067, n1028);
not  g1015 (n1056, n1031);
buf  g1016 (n1049, n1029);
not  g1017 (n1070, n1036);
not  g1018 (n1051, n1034);
not  g1019 (n1063, n1035);
not  g1020 (n1047, n1032);
buf  g1021 (n1073, n1030);
not  g1022 (n1054, n1037);
not  g1023 (n1068, n1031);
not  g1024 (n1065, n1029);
buf  g1025 (n1057, n1032);
buf  g1026 (n1081, n1033);
not  g1027 (n1080, n1035);
buf  g1028 (n1069, n1029);
buf  g1029 (n1062, n1033);
buf  g1030 (n1077, n1036);
not  g1031 (n1060, n1030);
buf  g1032 (n1075, n1029);
buf  g1033 (n1058, n1031);
not  g1034 (n1079, n1030);
not  g1035 (n1064, n1032);
not  g1036 (n1046, n1036);
buf  g1037 (n1078, n1035);
not  g1038 (n1055, n1030);
buf  g1039 (n1052, n1035);
buf  g1040 (n1053, n1033);
buf  g1041 (n1082, n1036);
not  g1042 (n1076, n1031);
not  g1043 (n1050, n1034);
buf  g1044 (n1066, n1033);
not  g1045 (n1074, n1034);
buf  g1046 (n1061, n1028);
buf  g1047 (n1072, n1028);
not  g1048 (n1048, n1034);
not  g1049 (n1045, n1028);
buf  g1050 (n1160, n1064);
buf  g1051 (n1191, n1060);
buf  g1052 (n1148, n660);
not  g1053 (n1208, n1003);
buf  g1054 (n1103, n1055);
not  g1055 (n1099, n833);
buf  g1056 (n1223, n1051);
buf  g1057 (n1220, n1059);
not  g1058 (n1226, n1073);
buf  g1059 (n1086, n1066);
not  g1060 (n1140, n878);
buf  g1061 (n1200, n1008);
not  g1062 (n1206, n1063);
not  g1063 (n1182, n1008);
not  g1064 (n1158, n1049);
not  g1065 (n1130, n1075);
buf  g1066 (n1137, n665);
buf  g1067 (n1089, n659);
buf  g1068 (n1088, n1066);
buf  g1069 (n1084, n1068);
buf  g1070 (n1104, n1061);
buf  g1071 (n1203, n1065);
not  g1072 (n1231, n1054);
not  g1073 (n1216, n1076);
not  g1074 (n1233, n1062);
buf  g1075 (n1218, n975);
not  g1076 (n1168, n1080);
buf  g1077 (n1107, n1069);
buf  g1078 (n1128, n1067);
buf  g1079 (n1146, n1009);
buf  g1080 (n1147, n1014);
buf  g1081 (n1134, n1081);
not  g1082 (n1087, n1066);
buf  g1083 (n1222, n1053);
not  g1084 (n1194, n1014);
buf  g1085 (n1142, n1055);
not  g1086 (n1085, n1012);
not  g1087 (n1116, n1049);
buf  g1088 (n1141, n1013);
buf  g1089 (n1110, n1078);
buf  g1090 (n1170, n1045);
not  g1091 (n1169, n973);
not  g1092 (n1090, n1077);
not  g1093 (n1114, n1067);
buf  g1094 (n1151, n1003);
buf  g1095 (n1209, n668);
not  g1096 (n1163, n666);
buf  g1097 (n1213, n1058);
not  g1098 (n1180, n1056);
not  g1099 (n1214, n1074);
buf  g1100 (n1139, n1067);
not  g1101 (n1164, n1007);
not  g1102 (n1228, n1053);
buf  g1103 (n1129, n1047);
not  g1104 (n1111, n1061);
not  g1105 (n1205, n1073);
not  g1106 (n1196, n1051);
not  g1107 (n1192, n1072);
buf  g1108 (n1133, n1077);
buf  g1109 (n1189, n1013);
not  g1110 (n1119, n1080);
buf  g1111 (n1136, n1050);
buf  g1112 (n1113, n1079);
not  g1113 (n1156, n1004);
buf  g1114 (n1095, n1064);
not  g1115 (n1125, n1007);
buf  g1116 (n1166, n1064);
buf  g1117 (n1221, n1080);
not  g1118 (n1234, n1008);
buf  g1119 (n1121, n1068);
buf  g1120 (n1132, n1048);
not  g1121 (n1175, n1065);
buf  g1122 (n1190, n1006);
not  g1123 (n1162, n1001);
not  g1124 (n1108, n879);
buf  g1125 (n1092, n664);
not  g1126 (n1091, n1081);
not  g1127 (n1201, n1045);
buf  g1128 (n1131, n1011);
not  g1129 (n1219, n655);
not  g1130 (n1210, n1055);
buf  g1131 (n1172, n1004);
buf  g1132 (n1135, n1047);
not  g1133 (n1215, n1011);
buf  g1134 (n1159, n1068);
buf  g1135 (n1177, n1057);
not  g1136 (n1188, n1008);
buf  g1137 (n1183, n669);
buf  g1138 (n1217, n1075);
buf  g1139 (n1143, n1053);
not  g1140 (n1098, n1052);
buf  g1141 (n1186, n1081);
not  g1142 (n1152, n1076);
buf  g1143 (n1187, n1069);
buf  g1144 (n1176, n661);
not  g1145 (n1093, n1002);
not  g1146 (n1149, n879);
buf  g1147 (n1124, n1005);
buf  g1148 (n1126, n1072);
buf  g1149 (n1211, n1047);
buf  g1150 (n1145, n1045);
buf  g1151 (n1227, n1060);
buf  g1152 (n1100, n1050);
buf  g1153 (n1232, n1074);
buf  g1154 (n1154, n1058);
not  g1155 (n1153, n1078);
buf  g1156 (n1198, n1072);
not  g1157 (n1185, n1013);
not  g1158 (n1096, n1079);
not  g1159 (n1199, n1046);
buf  g1160 (n1171, n1059);
nor  g1161 (n1184, n1002, n878, n1003);
xnor g1162 (n1174, n1046, n1058, n1011);
xor  g1163 (n1083, n1050, n1010, n1074);
nor  g1164 (n1165, n657, n974, n1079);
nand g1165 (n1202, n1005, n1003, n1063);
and  g1166 (n1181, n1082, n1045, n879);
xor  g1167 (n1138, n1059, n1063, n1014);
nand g1168 (n1109, n1077, n1076, n1070);
xnor g1169 (n1150, n1078, n1068, n1066);
or   g1170 (n1117, n1046, n1057, n972);
nor  g1171 (n1122, n1049, n1079, n656);
nand g1172 (n1155, n1076, n1007, n1052);
nor  g1173 (n1112, n1049, n1059, n667);
nand g1174 (n1230, n1075, n878, n1065);
and  g1175 (n1193, n1071, n1077, n1012);
and  g1176 (n1127, n878, n663, n1010);
nand g1177 (n1115, n1064, n1070, n1057);
xor  g1178 (n1094, n1056, n662, n1073);
xnor g1179 (n1097, n973, n1062);
nor  g1180 (n1178, n1052, n1011, n1069);
or   g1181 (n1123, n1071, n1007, n1013);
nand g1182 (n1229, n1060, n1063, n1053);
nor  g1183 (n1144, n1071, n1006, n1058);
xor  g1184 (n1106, n879, n1012, n1071);
nand g1185 (n1207, n1056, n1004, n1009);
or   g1186 (n1102, n1081, n1078, n1054);
xnor g1187 (n1120, n1006, n1061, n1010);
and  g1188 (n1197, n1052, n1055, n1065);
nand g1189 (n1105, n1046, n1070, n1009);
nand g1190 (n1173, n1056, n974, n1009);
xnor g1191 (n1224, n975, n658, n1051);
nand g1192 (n1161, n670, n1006, n1054);
xnor g1193 (n1204, n1050, n1054, n1082);
nand g1194 (n1195, n1010, n1005);
xor  g1195 (n1212, n1004, n1062, n1061);
or   g1196 (n1179, n1012, n1082, n1051);
nand g1197 (n1101, n1082, n1057, n1080);
nor  g1198 (n1167, n1073, n1048);
nor  g1199 (n1118, n1075, n1067, n1060);
or   g1200 (n1225, n1072, n1048, n1047);
nor  g1201 (n1157, n1070, n1074, n1069);
not  g1202 (n1503, n1213);
buf  g1203 (n1618, n1178);
buf  g1204 (n1406, n1173);
not  g1205 (n1356, n1143);
not  g1206 (n1782, n1123);
buf  g1207 (n1532, n1117);
buf  g1208 (n1714, n1124);
not  g1209 (n1315, n933);
buf  g1210 (n1757, n1146);
not  g1211 (n1778, n1194);
buf  g1212 (n1664, n1228);
buf  g1213 (n1403, n1219);
buf  g1214 (n1601, n1201);
not  g1215 (n1421, n1098);
not  g1216 (n1373, n934);
not  g1217 (n1385, n1179);
buf  g1218 (n1268, n935);
not  g1219 (n1819, n1139);
not  g1220 (n1581, n1128);
buf  g1221 (n1394, n673);
buf  g1222 (n1296, n709);
buf  g1223 (n1368, n1041);
buf  g1224 (n1247, n1204);
buf  g1225 (n1418, n676);
not  g1226 (n1352, n1180);
not  g1227 (n1483, n1186);
buf  g1228 (n1486, n1154);
buf  g1229 (n1338, n1156);
not  g1230 (n1316, n1123);
not  g1231 (n1446, n1230);
buf  g1232 (n1716, n685);
buf  g1233 (n1604, n1101);
buf  g1234 (n1454, n1160);
buf  g1235 (n1517, n1181);
not  g1236 (n1362, n1099);
not  g1237 (n1340, n1143);
not  g1238 (n1476, n1199);
not  g1239 (n1659, n1093);
buf  g1240 (n1330, n934);
not  g1241 (n1564, n928);
not  g1242 (n1263, n1229);
not  g1243 (n1497, n1159);
buf  g1244 (n1829, n1209);
not  g1245 (n1802, n1090);
buf  g1246 (n1646, n1208);
not  g1247 (n1603, n1209);
buf  g1248 (n1720, n1183);
not  g1249 (n1390, n1164);
not  g1250 (n1482, n1111);
not  g1251 (n1347, n1089);
buf  g1252 (n1520, n1165);
not  g1253 (n1702, n1042);
buf  g1254 (n1360, n1132);
not  g1255 (n1401, n1113);
not  g1256 (n1681, n1180);
not  g1257 (n1253, n1112);
buf  g1258 (n1332, n1107);
not  g1259 (n1558, n1093);
buf  g1260 (n1777, n1219);
not  g1261 (n1323, n1142);
buf  g1262 (n1422, n1113);
buf  g1263 (n1796, n1220);
buf  g1264 (n1764, n1198);
not  g1265 (n1313, n1198);
buf  g1266 (n1522, n1117);
buf  g1267 (n1699, n1221);
not  g1268 (n1440, n1159);
not  g1269 (n1776, n1041);
not  g1270 (n1426, n1144);
not  g1271 (n1585, n1128);
buf  g1272 (n1578, n1123);
buf  g1273 (n1249, n1169);
buf  g1274 (n1358, n1231);
not  g1275 (n1238, n1131);
not  g1276 (n1607, n1104);
not  g1277 (n1396, n1175);
buf  g1278 (n1734, n1148);
buf  g1279 (n1631, n1121);
buf  g1280 (n1653, n1234);
not  g1281 (n1754, n1109);
not  g1282 (n1402, n1163);
buf  g1283 (n1798, n1126);
not  g1284 (n1553, n1230);
buf  g1285 (n1665, n1103);
buf  g1286 (n1719, n1172);
buf  g1287 (n1586, n1121);
buf  g1288 (n1837, n1217);
buf  g1289 (n1420, n1193);
buf  g1290 (n1668, n1108);
not  g1291 (n1371, n1084);
not  g1292 (n1821, n1095);
buf  g1293 (n1807, n1088);
not  g1294 (n1800, n1139);
not  g1295 (n1339, n1206);
not  g1296 (n1513, n1218);
not  g1297 (n1689, n1171);
buf  g1298 (n1695, n709);
buf  g1299 (n1608, n1134);
not  g1300 (n1364, n1202);
buf  g1301 (n1820, n1183);
buf  g1302 (n1515, n1185);
buf  g1303 (n1295, n1168);
not  g1304 (n1438, n1163);
buf  g1305 (n1671, n1218);
not  g1306 (n1495, n1166);
buf  g1307 (n1629, n932);
not  g1308 (n1376, n1099);
not  g1309 (n1471, n1146);
not  g1310 (n1828, n1040);
not  g1311 (n1737, n1119);
buf  g1312 (n1544, n1042);
not  g1313 (n1441, n1136);
not  g1314 (n1708, n1148);
buf  g1315 (n1272, n1094);
not  g1316 (n1254, n1200);
not  g1317 (n1657, n1115);
not  g1318 (n1538, n690);
not  g1319 (n1599, n1214);
buf  g1320 (n1416, n1152);
buf  g1321 (n1459, n1230);
buf  g1322 (n1572, n1192);
buf  g1323 (n1815, n1113);
not  g1324 (n1597, n1209);
not  g1325 (n1816, n932);
not  g1326 (n1799, n1085);
buf  g1327 (n1269, n688);
buf  g1328 (n1662, n1178);
buf  g1329 (n1589, n924);
not  g1330 (n1381, n1201);
buf  g1331 (n1431, n927);
not  g1332 (n1826, n1228);
buf  g1333 (n1616, n1174);
not  g1334 (n1488, n1141);
not  g1335 (n1701, n1135);
buf  g1336 (n1678, n1228);
buf  g1337 (n1617, n1148);
buf  g1338 (n1327, n1137);
buf  g1339 (n1453, n1089);
not  g1340 (n1504, n1039);
buf  g1341 (n1600, n807);
not  g1342 (n1491, n1234);
not  g1343 (n1451, n1170);
not  g1344 (n1633, n1226);
not  g1345 (n1640, n1231);
buf  g1346 (n1817, n680);
not  g1347 (n1615, n1162);
buf  g1348 (n1781, n1177);
buf  g1349 (n1670, n1104);
not  g1350 (n1801, n1153);
buf  g1351 (n1317, n1210);
buf  g1352 (n1243, n1206);
buf  g1353 (n1655, n1207);
buf  g1354 (n1256, n1183);
not  g1355 (n1466, n1214);
buf  g1356 (n1548, n1171);
not  g1357 (n1355, n1171);
buf  g1358 (n1606, n1120);
buf  g1359 (n1525, n1099);
not  g1360 (n1709, n1202);
buf  g1361 (n1264, n1190);
buf  g1362 (n1569, n932);
buf  g1363 (n1583, n1144);
not  g1364 (n1713, n1166);
buf  g1365 (n1444, n1098);
buf  g1366 (n1588, n1103);
not  g1367 (n1291, n1226);
buf  g1368 (n1625, n1122);
not  g1369 (n1759, n807);
not  g1370 (n1388, n931);
buf  g1371 (n1561, n1165);
not  g1372 (n1259, n1227);
not  g1373 (n1345, n1039);
not  g1374 (n1326, n1038);
not  g1375 (n1750, n1091);
not  g1376 (n1370, n930);
not  g1377 (n1484, n1232);
buf  g1378 (n1706, n1105);
not  g1379 (n1407, n1134);
not  g1380 (n1301, n1194);
buf  g1381 (n1363, n1167);
not  g1382 (n1822, n1041);
not  g1383 (n1310, n1125);
buf  g1384 (n1686, n926);
buf  g1385 (n1287, n672);
not  g1386 (n1580, n1167);
not  g1387 (n1721, n1092);
not  g1388 (n1470, n1182);
not  g1389 (n1728, n1184);
not  g1390 (n1305, n929);
buf  g1391 (n1809, n1149);
not  g1392 (n1622, n806);
buf  g1393 (n1511, n926);
buf  g1394 (n1423, n1200);
buf  g1395 (n1410, n1125);
not  g1396 (n1274, n1147);
not  g1397 (n1519, n1085);
not  g1398 (n1814, n1098);
not  g1399 (n1751, n926);
buf  g1400 (n1457, n1188);
buf  g1401 (n1582, n1115);
buf  g1402 (n1354, n1177);
buf  g1403 (n1343, n1181);
not  g1404 (n1242, n1129);
buf  g1405 (n1775, n1207);
not  g1406 (n1369, n1118);
not  g1407 (n1712, n1125);
buf  g1408 (n1649, n1043);
not  g1409 (n1490, n1222);
not  g1410 (n1424, n1172);
not  g1411 (n1680, n682);
buf  g1412 (n1705, n1232);
not  g1413 (n1683, n1229);
not  g1414 (n1790, n1083);
buf  g1415 (n1530, n678);
buf  g1416 (n1425, n1137);
buf  g1417 (n1630, n1214);
not  g1418 (n1285, n1207);
not  g1419 (n1435, n1095);
buf  g1420 (n1736, n1131);
not  g1421 (n1284, n681);
buf  g1422 (n1346, n1170);
buf  g1423 (n1248, n1182);
buf  g1424 (n1672, n1157);
not  g1425 (n1591, n1136);
not  g1426 (n1745, n1130);
buf  g1427 (n1437, n671);
buf  g1428 (n1833, n1170);
not  g1429 (n1500, n1140);
buf  g1430 (n1767, n1185);
not  g1431 (n1567, n1145);
not  g1432 (n1378, n1164);
buf  g1433 (n1730, n1122);
not  g1434 (n1614, n1182);
buf  g1435 (n1570, n1129);
buf  g1436 (n1258, n930);
not  g1437 (n1468, n1096);
buf  g1438 (n1690, n1190);
not  g1439 (n1474, n933);
buf  g1440 (n1475, n1138);
not  g1441 (n1723, n1178);
not  g1442 (n1357, n1161);
not  g1443 (n1328, n1202);
buf  g1444 (n1344, n927);
buf  g1445 (n1696, n1195);
buf  g1446 (n1465, n1217);
buf  g1447 (n1350, n1100);
not  g1448 (n1729, n1193);
not  g1449 (n1290, n1127);
not  g1450 (n1641, n1038);
buf  g1451 (n1842, n1224);
not  g1452 (n1688, n1095);
not  g1453 (n1240, n1044);
not  g1454 (n1840, n1133);
buf  g1455 (n1417, n1106);
buf  g1456 (n1623, n1119);
buf  g1457 (n1462, n1088);
not  g1458 (n1666, n1117);
not  g1459 (n1594, n1205);
buf  g1460 (n1294, n1176);
not  g1461 (n1747, n1226);
not  g1462 (n1322, n1116);
buf  g1463 (n1439, n1143);
buf  g1464 (n1555, n1152);
buf  g1465 (n1733, n1084);
buf  g1466 (n1400, n809);
buf  g1467 (n1707, n1201);
not  g1468 (n1693, n1092);
not  g1469 (n1537, n1205);
buf  g1470 (n1523, n1197);
not  g1471 (n1415, n1102);
not  g1472 (n1261, n1096);
not  g1473 (n1501, n1207);
not  g1474 (n1460, n1184);
not  g1475 (n1489, n1157);
buf  g1476 (n1741, n1044);
not  g1477 (n1375, n1218);
buf  g1478 (n1732, n1103);
not  g1479 (n1677, n1090);
buf  g1480 (n1717, n1122);
buf  g1481 (n1703, n1227);
not  g1482 (n1514, n1190);
not  g1483 (n1300, n1128);
not  g1484 (n1550, n1138);
not  g1485 (n1832, n1203);
buf  g1486 (n1433, n1225);
not  g1487 (n1783, n1178);
buf  g1488 (n1241, n1213);
buf  g1489 (n1769, n1184);
buf  g1490 (n1792, n1118);
not  g1491 (n1469, n1201);
buf  g1492 (n1236, n927);
buf  g1493 (n1383, n1187);
buf  g1494 (n1823, n1175);
buf  g1495 (n1838, n1227);
buf  g1496 (n1559, n935);
not  g1497 (n1250, n674);
not  g1498 (n1804, n1096);
not  g1499 (n1795, n929);
not  g1500 (n1627, n1196);
not  g1501 (n1565, n1206);
not  g1502 (n1306, n934);
buf  g1503 (n1244, n1222);
buf  g1504 (n1361, n1126);
buf  g1505 (n1726, n1110);
buf  g1506 (n1687, n679);
buf  g1507 (n1557, n1119);
buf  g1508 (n1549, n1141);
not  g1509 (n1637, n1135);
buf  g1510 (n1320, n1225);
not  g1511 (n1539, n1089);
not  g1512 (n1456, n1223);
buf  g1513 (n1333, n1090);
buf  g1514 (n1508, n1149);
buf  g1515 (n1788, n1116);
buf  g1516 (n1443, n1097);
not  g1517 (n1309, n1151);
not  g1518 (n1529, n1217);
not  g1519 (n1644, n1145);
not  g1520 (n1598, n1093);
not  g1521 (n1542, n928);
not  g1522 (n1379, n1088);
not  g1523 (n1735, n1087);
not  g1524 (n1450, n1154);
not  g1525 (n1293, n1037);
not  g1526 (n1762, n687);
not  g1527 (n1808, n1182);
buf  g1528 (n1793, n1192);
buf  g1529 (n1643, n1137);
buf  g1530 (n1506, n1111);
buf  g1531 (n1786, n1148);
not  g1532 (n1679, n1223);
buf  g1533 (n1251, n1188);
buf  g1534 (n1560, n1155);
buf  g1535 (n1731, n1141);
not  g1536 (n1611, n1232);
buf  g1537 (n1391, n931);
not  g1538 (n1276, n1138);
not  g1539 (n1335, n689);
not  g1540 (n1658, n1206);
not  g1541 (n1645, n1221);
not  g1542 (n1647, n1190);
buf  g1543 (n1442, n1133);
buf  g1544 (n1758, n1134);
not  g1545 (n1694, n1133);
buf  g1546 (n1556, n1154);
not  g1547 (n1413, n1118);
buf  g1548 (n1289, n1147);
not  g1549 (n1307, n1175);
not  g1550 (n1571, n1117);
not  g1551 (n1587, n1215);
buf  g1552 (n1235, n1100);
buf  g1553 (n1429, n1086);
not  g1554 (n1551, n1160);
not  g1555 (n1770, n1119);
not  g1556 (n1304, n1173);
buf  g1557 (n1535, n1110);
not  g1558 (n1768, n1167);
buf  g1559 (n1408, n1168);
not  g1560 (n1761, n1177);
not  g1561 (n1281, n1212);
buf  g1562 (n1448, n1212);
not  g1563 (n1395, n1039);
not  g1564 (n1784, n1106);
buf  g1565 (n1697, n1014);
not  g1566 (n1266, n1153);
not  g1567 (n1563, n1146);
not  g1568 (n1834, n1210);
buf  g1569 (n1684, n1111);
buf  g1570 (n1257, n924);
not  g1571 (n1738, n1090);
not  g1572 (n1610, n1150);
buf  g1573 (n1367, n1114);
not  g1574 (n1652, n1122);
buf  g1575 (n1752, n1180);
buf  g1576 (n1359, n1121);
not  g1577 (n1780, n1040);
not  g1578 (n1656, n1153);
not  g1579 (n1593, n1233);
not  g1580 (n1545, n1151);
not  g1581 (n1541, n1042);
not  g1582 (n1624, n1038);
not  g1583 (n1318, n1180);
not  g1584 (n1463, n1147);
not  g1585 (n1324, n1192);
not  g1586 (n1831, n1151);
buf  g1587 (n1521, n1194);
not  g1588 (n1676, n1126);
buf  g1589 (n1458, n1211);
not  g1590 (n1419, n1043);
not  g1591 (n1494, n1137);
not  g1592 (n1279, n1231);
buf  g1593 (n1634, n1223);
buf  g1594 (n1766, n1191);
not  g1595 (n1547, n1129);
buf  g1596 (n1436, n1216);
not  g1597 (n1428, n1166);
not  g1598 (n1432, n1114);
not  g1599 (n1704, n1109);
not  g1600 (n1461, n1197);
buf  g1601 (n1638, n683);
not  g1602 (n1239, n1234);
buf  g1603 (n1812, n1108);
buf  g1604 (n1669, n1086);
buf  g1605 (n1811, n1222);
not  g1606 (n1533, n1216);
buf  g1607 (n1540, n1142);
not  g1608 (n1312, n1135);
buf  g1609 (n1493, n1176);
buf  g1610 (n1813, n1105);
buf  g1611 (n1464, n1133);
buf  g1612 (n1478, n1174);
buf  g1613 (n1824, n1094);
buf  g1614 (n1568, n1224);
buf  g1615 (n1331, n1147);
not  g1616 (n1510, n1110);
not  g1617 (n1382, n1150);
buf  g1618 (n1692, n1086);
buf  g1619 (n1612, n1219);
not  g1620 (n1673, n1085);
not  g1621 (n1505, n1228);
buf  g1622 (n1642, n1164);
not  g1623 (n1252, n1146);
buf  g1624 (n1739, n809);
buf  g1625 (n1772, n1096);
not  g1626 (n1595, n1172);
buf  g1627 (n1445, n1230);
buf  g1628 (n1434, n1233);
not  g1629 (n1405, n1089);
not  g1630 (n1841, n1219);
buf  g1631 (n1660, n1041);
buf  g1632 (n1377, n1152);
not  g1633 (n1384, n1083);
buf  g1634 (n1502, n1162);
not  g1635 (n1492, n1130);
not  g1636 (n1746, n925);
buf  g1637 (n1280, n1105);
not  g1638 (n1543, n1212);
not  g1639 (n1654, n1169);
buf  g1640 (n1397, n1114);
buf  g1641 (n1648, n931);
not  g1642 (n1427, n1088);
not  g1643 (n1743, n1225);
buf  g1644 (n1265, n1213);
buf  g1645 (n1771, n1220);
not  g1646 (n1255, n1084);
not  g1647 (n1325, n1231);
not  g1648 (n1651, n1107);
buf  g1649 (n1636, n1100);
not  g1650 (n1353, n1108);
not  g1651 (n1742, n1093);
buf  g1652 (n1753, n1186);
buf  g1653 (n1314, n1135);
buf  g1654 (n1479, n1142);
not  g1655 (n1626, n677);
buf  g1656 (n1584, n927);
buf  g1657 (n1602, n1114);
buf  g1658 (n1789, n1159);
buf  g1659 (n1632, n1197);
buf  g1660 (n1319, n1136);
not  g1661 (n1380, n1158);
buf  g1662 (n1534, n1150);
buf  g1663 (n1298, n1218);
not  g1664 (n1685, n1094);
not  g1665 (n1398, n1040);
buf  g1666 (n1605, n1044);
not  g1667 (n1485, n933);
not  g1668 (n1774, n1128);
not  g1669 (n1740, n1232);
not  g1670 (n1827, n1234);
not  g1671 (n1260, n1094);
buf  g1672 (n1609, n1140);
buf  g1673 (n1496, n1039);
not  g1674 (n1785, n1210);
buf  g1675 (n1365, n1087);
not  g1676 (n1682, n1086);
not  g1677 (n1283, n1112);
not  g1678 (n1577, n1220);
buf  g1679 (n1246, n1183);
buf  g1680 (n1321, n1042);
buf  g1681 (n1765, n1125);
not  g1682 (n1722, n1197);
buf  g1683 (n1341, n1129);
not  g1684 (n1393, n1162);
not  g1685 (n1499, n1097);
not  g1686 (n1297, n1199);
buf  g1687 (n1661, n1176);
buf  g1688 (n1805, n1213);
buf  g1689 (n1399, n1127);
buf  g1690 (n1273, n1155);
buf  g1691 (n1710, n1120);
not  g1692 (n1270, n1136);
buf  g1693 (n1498, n1157);
not  g1694 (n1412, n1199);
not  g1695 (n1336, n1173);
not  g1696 (n1552, n1186);
buf  g1697 (n1487, n1208);
not  g1698 (n1756, n1095);
buf  g1699 (n1275, n808);
not  g1700 (n1667, n1205);
buf  g1701 (n1619, n1108);
buf  g1702 (n1299, n1104);
buf  g1703 (n1524, n1165);
buf  g1704 (n1725, n1103);
not  g1705 (n1760, n1156);
not  g1706 (n1386, n1132);
buf  g1707 (n1674, n1187);
not  g1708 (n1286, n1185);
buf  g1709 (n1639, n1155);
buf  g1710 (n1303, n1184);
not  g1711 (n1698, n1224);
not  g1712 (n1480, n1164);
not  g1713 (n1271, n1043);
buf  g1714 (n1835, n1179);
not  g1715 (n1282, n1216);
not  g1716 (n1797, n684);
not  g1717 (n1366, n1085);
not  g1718 (n1447, n1211);
buf  g1719 (n1806, n1099);
buf  g1720 (n1839, n932);
not  g1721 (n1635, n1198);
buf  g1722 (n1803, n1158);
buf  g1723 (n1554, n934);
buf  g1724 (n1262, n1115);
not  g1725 (n1414, n1043);
buf  g1726 (n1278, n1144);
buf  g1727 (n1715, n1102);
buf  g1728 (n1791, n1134);
not  g1729 (n1245, n1194);
not  g1730 (n1650, n1109);
not  g1731 (n1536, n1151);
not  g1732 (n1748, n1162);
not  g1733 (n1836, n1152);
buf  g1734 (n1579, n1127);
buf  g1735 (n1628, n1106);
buf  g1736 (n1575, n1233);
not  g1737 (n1302, n1092);
buf  g1738 (n1592, n1109);
buf  g1739 (n1467, n1092);
not  g1740 (n1576, n1211);
buf  g1741 (n1573, n1132);
not  g1742 (n1596, n1204);
not  g1743 (n1337, n1208);
buf  g1744 (n1620, n1163);
buf  g1745 (n1744, n1110);
buf  g1746 (n1348, n1113);
not  g1747 (n1810, n1188);
buf  g1748 (n1389, n1203);
not  g1749 (n1342, n1223);
buf  g1750 (n1613, n1037);
buf  g1751 (n1267, n1161);
buf  g1752 (n1311, n1118);
not  g1753 (n1449, n1121);
buf  g1754 (n1509, n1187);
not  g1755 (n1526, n1107);
and  g1756 (n1372, n1138, n1166, n1155);
nand g1757 (n1292, n929, n808, n1123);
nor  g1758 (n1566, n1204, n1149, n1210);
and  g1759 (n1718, n1212, n1102, n686);
xnor g1760 (n1727, n1227, n1222, n1163);
and  g1761 (n1825, n1204, n675, n1106);
nand g1762 (n1452, n1208, n1112, n1168);
xor  g1763 (n1724, n1215, n1124, n1130);
or   g1764 (n1411, n1132, n1115, n1215);
nand g1765 (n1351, n1168, n1214, n1102);
nand g1766 (n1562, n1160, n1186, n1161);
or   g1767 (n1387, n1145, n1097, n1217);
nand g1768 (n1334, n1221, n1084, n1196);
xor  g1769 (n1277, n1191, n1189, n1193);
and  g1770 (n1329, n1196, n1167, n1097);
xnor g1771 (n1818, n1116, n1130, n1175);
nor  g1772 (n1763, n1189, n1141, n1104);
xor  g1773 (n1574, n1200, n926, n1173);
or   g1774 (n1308, n1202, n1038, n1225);
xor  g1775 (n1516, n1189, n1091, n1157);
nor  g1776 (n1409, n1143, n1105, n1116);
nor  g1777 (n1481, n1149, n1196, n1159);
and  g1778 (n1773, n1112, n930);
xor  g1779 (n1237, n1198, n1120, n1153);
or   g1780 (n1473, n1156, n931, n1139);
nor  g1781 (n1477, n1189, n925, n1209);
nand g1782 (n1546, n1160, n1127, n1107);
xnor g1783 (n1288, n1229, n1203, n1124);
xor  g1784 (n1711, n1124, n1195, n1120);
xnor g1785 (n1472, n928, n1179, n1101);
or   g1786 (n1779, n1211, n1224, n1215);
xor  g1787 (n1749, n1220, n925, n1187);
xnor g1788 (n1830, n1091, n1098, n1174);
xnor g1789 (n1700, n1221, n1195, n1176);
nor  g1790 (n1531, n1101, n1087, n1181);
xnor g1791 (n1675, n1200, n1203, n1126);
xor  g1792 (n1392, n1040, n1091, n933);
xor  g1793 (n1349, n1174, n1181, n1229);
and  g1794 (n1518, n1199, n1192, n1158);
or   g1795 (n1430, n1111, n1140, n935);
xnor g1796 (n1787, n1101, n1191, n1142);
xor  g1797 (n1512, n1188, n1144, n1087);
nand g1798 (n1691, n1083, n929, n1131);
xnor g1799 (n1527, n1044, n1233, n925);
or   g1800 (n1590, n1156, n924, n1170);
nor  g1801 (n1404, n1140, n1161, n1145);
xnor g1802 (n1755, n1185, n1193, n1158);
and  g1803 (n1663, n1179, n1191, n1169);
or   g1804 (n1794, n1205, n1177, n1171);
xnor g1805 (n1528, n1195, n1169, n1172);
or   g1806 (n1507, n1100, n1131, n928);
and  g1807 (n1455, n1216, n806, n1083);
and  g1808 (n1621, n1165, n1150, n1154);
or   g1809 (n1374, n1139, n1226, n935);
buf  g1810 (n2629, n1708);
not  g1811 (n2543, n1241);
not  g1812 (n1903, n1332);
not  g1813 (n2306, n1596);
buf  g1814 (n2628, n1740);
not  g1815 (n2279, n1365);
not  g1816 (n2396, n1721);
buf  g1817 (n2024, n1516);
not  g1818 (n2058, n1690);
buf  g1819 (n1858, n1767);
not  g1820 (n2046, n1510);
not  g1821 (n2555, n1252);
buf  g1822 (n2726, n1410);
not  g1823 (n2666, n1766);
not  g1824 (n2007, n1311);
buf  g1825 (n2157, n1663);
not  g1826 (n2452, n1452);
not  g1827 (n1959, n1376);
not  g1828 (n2594, n1514);
not  g1829 (n2415, n1505);
not  g1830 (n2340, n1822);
not  g1831 (n2683, n1765);
not  g1832 (n2489, n1668);
not  g1833 (n1998, n1276);
not  g1834 (n2626, n1284);
buf  g1835 (n2606, n1419);
buf  g1836 (n2152, n1822);
buf  g1837 (n2656, n1527);
not  g1838 (n2394, n1681);
not  g1839 (n2663, n1465);
not  g1840 (n2307, n1769);
buf  g1841 (n1999, n1823);
buf  g1842 (n2295, n1298);
not  g1843 (n2060, n1271);
buf  g1844 (n2168, n1813);
buf  g1845 (n2159, n1746);
not  g1846 (n2069, n1581);
buf  g1847 (n1883, n1408);
buf  g1848 (n2181, n1532);
buf  g1849 (n1851, n1411);
buf  g1850 (n2232, n1297);
not  g1851 (n2611, n1338);
buf  g1852 (n2638, n1572);
buf  g1853 (n2634, n1794);
buf  g1854 (n2383, n1302);
not  g1855 (n2380, n1248);
buf  g1856 (n2689, n1348);
not  g1857 (n2425, n1770);
buf  g1858 (n2403, n1409);
buf  g1859 (n2175, n1571);
buf  g1860 (n2353, n1734);
buf  g1861 (n1844, n1583);
not  g1862 (n2038, n1640);
buf  g1863 (n1940, n1246);
buf  g1864 (n2068, n1594);
not  g1865 (n2511, n1248);
not  g1866 (n2222, n1337);
buf  g1867 (n2164, n1373);
not  g1868 (n2223, n1584);
not  g1869 (n2410, n1737);
buf  g1870 (n2449, n1622);
not  g1871 (n1977, n1668);
not  g1872 (n2070, n1730);
not  g1873 (n2576, n1319);
not  g1874 (n2532, n1524);
buf  g1875 (n2318, n1324);
not  g1876 (n1860, n1292);
not  g1877 (n2109, n1573);
buf  g1878 (n2121, n1488);
not  g1879 (n2720, n1577);
buf  g1880 (n2022, n1293);
not  g1881 (n2325, n1749);
buf  g1882 (n2578, n1398);
buf  g1883 (n2389, n1588);
not  g1884 (n2268, n1341);
not  g1885 (n2304, n1609);
not  g1886 (n2215, n1683);
buf  g1887 (n2561, n1239);
buf  g1888 (n2125, n1513);
not  g1889 (n2635, n1587);
not  g1890 (n2676, n1818);
not  g1891 (n2385, n1352);
not  g1892 (n2319, n1364);
buf  g1893 (n2133, n1656);
not  g1894 (n2148, n1347);
not  g1895 (n2252, n1604);
buf  g1896 (n2542, n1523);
buf  g1897 (n2377, n1328);
not  g1898 (n2324, n1327);
buf  g1899 (n2495, n1610);
buf  g1900 (n1951, n1626);
buf  g1901 (n2326, n1663);
not  g1902 (n2146, n1720);
buf  g1903 (n2539, n1291);
buf  g1904 (n2242, n1837);
not  g1905 (n2723, n1821);
buf  g1906 (n2355, n1747);
buf  g1907 (n2469, n1244);
not  g1908 (n2248, n1590);
not  g1909 (n2020, n1756);
buf  g1910 (n2023, n1625);
buf  g1911 (n2103, n1667);
not  g1912 (n2030, n1505);
buf  g1913 (n2059, n1556);
buf  g1914 (n2475, n1705);
buf  g1915 (n2518, n1319);
buf  g1916 (n2501, n1719);
not  g1917 (n1929, n1413);
not  g1918 (n1941, n1776);
buf  g1919 (n2513, n1463);
not  g1920 (n2566, n1309);
buf  g1921 (n2291, n1633);
buf  g1922 (n2616, n1513);
not  g1923 (n1969, n1484);
not  g1924 (n1921, n1463);
buf  g1925 (n2470, n1799);
not  g1926 (n1985, n1307);
not  g1927 (n2311, n1505);
not  g1928 (n1948, n1455);
not  g1929 (n2280, n1447);
not  g1930 (n2116, n1462);
not  g1931 (n2687, n1632);
not  g1932 (n2560, n1448);
buf  g1933 (n2296, n1602);
buf  g1934 (n2399, n1500);
not  g1935 (n2436, n1526);
buf  g1936 (n1902, n1264);
not  g1937 (n1995, n1396);
buf  g1938 (n2715, n1490);
buf  g1939 (n2350, n1726);
not  g1940 (n2259, n1628);
not  g1941 (n2710, n1693);
buf  g1942 (n1952, n1449);
buf  g1943 (n2457, n1250);
buf  g1944 (n2659, n1344);
not  g1945 (n2364, n1455);
buf  g1946 (n2285, n1277);
not  g1947 (n2272, n1529);
not  g1948 (n2716, n1330);
buf  g1949 (n1886, n1406);
not  g1950 (n1911, n1716);
buf  g1951 (n2450, n1520);
buf  g1952 (n2547, n1409);
buf  g1953 (n2000, n1595);
buf  g1954 (n2056, n1370);
buf  g1955 (n2655, n1320);
not  g1956 (n2680, n1392);
not  g1957 (n2199, n1532);
buf  g1958 (n2603, n1475);
buf  g1959 (n1912, n1395);
buf  g1960 (n2612, n1650);
buf  g1961 (n2714, n1682);
buf  g1962 (n1955, n1333);
buf  g1963 (n2081, n1309);
buf  g1964 (n2333, n1299);
not  g1965 (n2675, n1689);
buf  g1966 (n2093, n1757);
not  g1967 (n1984, n1280);
not  g1968 (n2685, n1486);
buf  g1969 (n2115, n1424);
buf  g1970 (n2390, n1755);
buf  g1971 (n2526, n1315);
not  g1972 (n2163, n1710);
buf  g1973 (n2132, n1445);
buf  g1974 (n2682, n1646);
buf  g1975 (n2329, n1335);
not  g1976 (n2673, n1553);
buf  g1977 (n1932, n1514);
not  g1978 (n1987, n1364);
buf  g1979 (n2700, n1709);
buf  g1980 (n1847, n1474);
not  g1981 (n2235, n1356);
buf  g1982 (n1978, n1765);
buf  g1983 (n2359, n1738);
buf  g1984 (n2497, n1568);
buf  g1985 (n2719, n1666);
buf  g1986 (n2423, n1387);
buf  g1987 (n2491, n1482);
buf  g1988 (n2379, n1673);
buf  g1989 (n2386, n1827);
buf  g1990 (n1931, n1288);
not  g1991 (n2602, n1479);
buf  g1992 (n2257, n1499);
buf  g1993 (n2391, n1493);
not  g1994 (n2493, n1432);
buf  g1995 (n2357, n1381);
not  g1996 (n1910, n692);
buf  g1997 (n1970, n1647);
buf  g1998 (n2564, n1269);
not  g1999 (n2104, n1729);
not  g2000 (n2535, n1734);
buf  g2001 (n2482, n1527);
buf  g2002 (n1947, n1390);
not  g2003 (n2702, n1326);
buf  g2004 (n2674, n1437);
buf  g2005 (n2447, n1592);
not  g2006 (n1857, n1523);
not  g2007 (n2127, n1751);
buf  g2008 (n1906, n1758);
not  g2009 (n1963, n1454);
not  g2010 (n2332, n1764);
not  g2011 (n2553, n1462);
not  g2012 (n2647, n1793);
buf  g2013 (n2147, n1634);
buf  g2014 (n2586, n1357);
buf  g2015 (n2565, n1267);
buf  g2016 (n1865, n1308);
buf  g2017 (n2284, n1260);
buf  g2018 (n1992, n1443);
not  g2019 (n2530, n1746);
not  g2020 (n2588, n1325);
not  g2021 (n2417, n1594);
buf  g2022 (n2098, n1542);
buf  g2023 (n2176, n1605);
buf  g2024 (n2365, n1310);
not  g2025 (n2260, n1481);
buf  g2026 (n1997, n1543);
buf  g2027 (n2211, n1399);
buf  g2028 (n2229, n1806);
not  g2029 (n2621, n1240);
not  g2030 (n2584, n1262);
buf  g2031 (n2510, n1384);
buf  g2032 (n2312, n1372);
buf  g2033 (n2155, n1470);
buf  g2034 (n1950, n1357);
buf  g2035 (n2221, n1691);
buf  g2036 (n2108, n1763);
buf  g2037 (n2266, n1402);
buf  g2038 (n1949, n1235);
buf  g2039 (n2562, n1745);
not  g2040 (n2551, n1397);
not  g2041 (n2618, n1489);
buf  g2042 (n2521, n1467);
buf  g2043 (n2426, n1294);
not  g2044 (n2652, n1476);
not  g2045 (n1942, n1720);
buf  g2046 (n2462, n1243);
not  g2047 (n2598, n1587);
buf  g2048 (n2393, n1580);
not  g2049 (n2028, n1533);
not  g2050 (n2574, n1395);
buf  g2051 (n2485, n1412);
not  g2052 (n2192, n1346);
buf  g2053 (n2338, n1418);
buf  g2054 (n2301, n1258);
buf  g2055 (n2254, n1589);
not  g2056 (n2004, n1727);
not  g2057 (n1960, n1597);
not  g2058 (n2467, n1793);
buf  g2059 (n1908, n1378);
buf  g2060 (n2299, n1362);
not  g2061 (n2191, n1289);
not  g2062 (n1894, n1604);
buf  g2063 (n1891, n1319);
not  g2064 (n1868, n1834);
not  g2065 (n2165, n1478);
not  g2066 (n1887, n1702);
not  g2067 (n2520, n1300);
not  g2068 (n1899, n1772);
buf  g2069 (n2473, n1667);
buf  g2070 (n1982, n1330);
not  g2071 (n2455, n1691);
not  g2072 (n2119, n1631);
buf  g2073 (n1928, n1251);
not  g2074 (n1943, n1486);
buf  g2075 (n1938, n1603);
buf  g2076 (n2045, n1251);
not  g2077 (n2206, n1741);
buf  g2078 (n2270, n1629);
not  g2079 (n2435, n1678);
buf  g2080 (n1979, n1355);
not  g2081 (n2585, n1798);
not  g2082 (n2694, n1484);
not  g2083 (n2697, n1311);
buf  g2084 (n2110, n1497);
not  g2085 (n2481, n1545);
not  g2086 (n2079, n1731);
buf  g2087 (n1976, n1712);
not  g2088 (n2593, n1574);
not  g2089 (n2131, n1580);
not  g2090 (n1901, n1258);
buf  g2091 (n2292, n1703);
buf  g2092 (n2233, n1729);
buf  g2093 (n2416, n1629);
buf  g2094 (n2264, n1478);
buf  g2095 (n2218, n1779);
not  g2096 (n2278, n1238);
buf  g2097 (n2552, n1832);
not  g2098 (n2166, n1535);
not  g2099 (n2609, n1379);
buf  g2100 (n2113, n1275);
buf  g2101 (n2508, n1269);
not  g2102 (n2063, n1695);
not  g2103 (n2571, n1615);
not  g2104 (n2140, n1379);
not  g2105 (n2135, n1397);
not  g2106 (n2371, n1386);
buf  g2107 (n1919, n1599);
not  g2108 (n2048, n1534);
buf  g2109 (n2153, n1680);
buf  g2110 (n2706, n1719);
not  g2111 (n2424, n1612);
buf  g2112 (n2533, n1618);
buf  g2113 (n2499, n1452);
buf  g2114 (n2506, n1735);
not  g2115 (n2114, n1725);
buf  g2116 (n1850, n1771);
buf  g2117 (n2712, n1797);
not  g2118 (n2367, n1800);
not  g2119 (n2352, n1352);
not  g2120 (n1882, n1400);
not  g2121 (n2692, n1696);
buf  g2122 (n2498, n1503);
buf  g2123 (n1926, n1271);
buf  g2124 (n1877, n1279);
buf  g2125 (n1974, n1614);
buf  g2126 (n2182, n1378);
not  g2127 (n2136, n1511);
buf  g2128 (n2039, n1627);
buf  g2129 (n2019, n1350);
not  g2130 (n2607, n1785);
not  g2131 (n2736, n1425);
not  g2132 (n1934, n1398);
buf  g2133 (n2536, n1366);
not  g2134 (n2650, n1778);
buf  g2135 (n1864, n1376);
buf  g2136 (n2504, n1564);
not  g2137 (n2351, n1471);
buf  g2138 (n2043, n1548);
buf  g2139 (n2360, n1246);
not  g2140 (n2213, n1373);
not  g2141 (n2143, n1273);
buf  g2142 (n2073, n1404);
not  g2143 (n2373, n1695);
buf  g2144 (n2062, n1381);
not  g2145 (n2094, n1398);
not  g2146 (n2003, n1624);
buf  g2147 (n1915, n1689);
buf  g2148 (n2476, n1353);
buf  g2149 (n2014, n1555);
buf  g2150 (n1871, n1437);
buf  g2151 (n2179, n1371);
buf  g2152 (n2186, n1442);
buf  g2153 (n2323, n1781);
buf  g2154 (n1863, n1822);
buf  g2155 (n2649, n1438);
not  g2156 (n2640, n1769);
not  g2157 (n2434, n1724);
buf  g2158 (n2074, n1651);
buf  g2159 (n2225, n1256);
buf  g2160 (n2220, n1424);
not  g2161 (n2583, n1760);
buf  g2162 (n2412, n1811);
not  g2163 (n2183, n1280);
buf  g2164 (n2321, n1293);
not  g2165 (n2134, n1732);
not  g2166 (n2505, n1787);
buf  g2167 (n2619, n1542);
not  g2168 (n2741, n1347);
buf  g2169 (n1973, n1283);
not  g2170 (n2657, n1377);
not  g2171 (n1856, n1271);
not  g2172 (n2636, n1375);
buf  g2173 (n1975, n1817);
not  g2174 (n2029, n1393);
not  g2175 (n2298, n1236);
not  g2176 (n2654, n1464);
not  g2177 (n2642, n1632);
not  g2178 (n1994, n1785);
buf  g2179 (n2128, n1328);
not  g2180 (n2732, n1480);
not  g2181 (n1956, n1589);
not  g2182 (n2397, n1765);
buf  g2183 (n2465, n1533);
buf  g2184 (n2310, n1612);
not  g2185 (n1944, n1643);
buf  g2186 (n2651, n1782);
buf  g2187 (n2721, n696);
buf  g2188 (n2243, n1620);
not  g2189 (n2053, n1339);
not  g2190 (n2558, n1801);
not  g2191 (n2514, n1354);
buf  g2192 (n2707, n1766);
buf  g2193 (n2239, n1635);
nand g2194 (n2228, n1616, n1334, n1606, n1358);
xnor g2195 (n2545, n1668, n1288, n1739, n1353);
nor  g2196 (n2083, n1360, n1273, n1334, n1319);
nand g2197 (n1946, n697, n1269, n1558, n1335);
xnor g2198 (n2293, n1365, n1609, n1466, n1623);
nand g2199 (n2021, n1500, n1747, n1830, n1491);
or   g2200 (n2055, n1336, n1407, n1344, n1705);
xnor g2201 (n2503, n1683, n1484, n1363, n1461);
xor  g2202 (n2086, n1384, n1761, n1402, n1338);
xnor g2203 (n2013, n1720, n1752, n1321, n1423);
xor  g2204 (n2077, n1692, n1323, n1828, n1776);
and  g2205 (n2017, n1802, n1268, n1528, n1777);
xor  g2206 (n2249, n1499, n1470, n1641, n1763);
and  g2207 (n2231, n1654, n1744, n1443, n1493);
or   g2208 (n1888, n1333, n1574, n1416, n1439);
or   g2209 (n2251, n1576, n1594, n1842, n1482);
nand g2210 (n1900, n1404, n1454, n1332, n1448);
or   g2211 (n2639, n1274, n1435, n1356, n1536);
or   g2212 (n2361, n1701, n1673, n1470, n1607);
nor  g2213 (n1914, n1648, n1450, n1762, n1301);
and  g2214 (n2448, n1592, n1433, n1389, n1544);
nand g2215 (n2690, n1323, n1316, n1331, n1533);
nand g2216 (n2372, n1774, n1273, n1431, n1722);
xor  g2217 (n2509, n1413, n1652, n1670, n1828);
or   g2218 (n2724, n1717, n1473, n1522, n1405);
or   g2219 (n1905, n1774, n1368, n1832, n1276);
xor  g2220 (n2557, n1759, n1376, n1541, n1498);
xor  g2221 (n2262, n1556, n1298, n1638, n1747);
xnor g2222 (n1993, n1353, n1247, n1784, n1701);
and  g2223 (n2015, n1720, n1244, n1452, n1815);
xor  g2224 (n1962, n1530, n1446, n1743, n1351);
xnor g2225 (n1872, n1367, n1662, n1770, n1237);
or   g2226 (n2538, n1440, n1775, n1384, n1422);
nor  g2227 (n2366, n1507, n1268, n1357, n1350);
xnor g2228 (n2573, n1407, n1509, n1583, n1464);
xor  g2229 (n2065, n1486, n1295, n1543, n1691);
and  g2230 (n2207, n1557, n1274, n1800, n1470);
or   g2231 (n2572, n1241, n1423, n1339, n1535);
xor  g2232 (n1924, n1485, n1575, n1508, n1483);
and  g2233 (n2336, n1305, n1587, n1786, n1332);
xnor g2234 (n2054, n1463, n1396, n1306);
xor  g2235 (n2144, n1570, n1278, n1347, n1477);
xnor g2236 (n2463, n1718, n1824, n1731, n1659);
xor  g2237 (n2120, n1468, n1279, n1536, n1550);
nand g2238 (n2265, n1261, n1265, n1650, n1451);
or   g2239 (n2196, n1831, n1345, n1690, n1323);
and  g2240 (n2568, n1730, n1657, n1834, n1628);
nand g2241 (n2283, n1267, n1301, n1251, n1264);
nor  g2242 (n2172, n1472, n1644, n1830, n1480);
and  g2243 (n2502, n1366, n1784, n1321, n1539);
xnor g2244 (n2614, n1306, n1549, n1465, n1672);
or   g2245 (n2544, n1808, n1528, n1243, n1315);
xor  g2246 (n2203, n1582, n326, n1389, n1441);
nor  g2247 (n2420, n1456, n1379, n1741, n1302);
xnor g2248 (n2646, n1255, n1337, n1582, n1286);
or   g2249 (n2316, n1600, n1476, n1282, n1578);
or   g2250 (n2263, n1641, n1617, n1840, n1759);
nand g2251 (n1861, n1744, n1611, n1364, n1702);
xor  g2252 (n2531, n1302, n1394, n1343, n1386);
xor  g2253 (n2582, n1508, n1541, n1602, n1816);
and  g2254 (n2672, n1636, n1666, n1285, n1312);
or   g2255 (n2224, n1648, n1771, n1773, n1322);
and  g2256 (n2488, n1521, n1549, n1410, n1670);
xnor g2257 (n2313, n1563, n1487, n1726, n1395);
xor  g2258 (n2688, n1530, n1406, n1839, n1818);
nand g2259 (n1898, n1620, n1411, n1405, n1634);
nor  g2260 (n2212, n1454, n1655, n1418, n1314);
nand g2261 (n2234, n1550, n1752, n1262, n1780);
xnor g2262 (n2742, n1658, n325, n1427, n1747);
or   g2263 (n2031, n1709, n1621, n1278, n1750);
or   g2264 (n2731, n1444, n1666, n1322, n1830);
and  g2265 (n2075, n1809, n1436, n1303, n1356);
nand g2266 (n2430, n1734, n1677, n1650, n1759);
xor  g2267 (n2184, n1655, n1340, n1542, n1366);
or   g2268 (n1889, n1681, n1694, n1579, n1460);
nand g2269 (n2101, n1649, n1451, n1287, n1755);
or   g2270 (n2197, n1785, n1418, n1799, n1729);
and  g2271 (n2126, n1688, n1476, n1358, n1509);
xnor g2272 (n2549, n1617, n1774, n1437, n1285);
or   g2273 (n1867, n1238, n1321, n1270, n1669);
or   g2274 (n2276, n1235, n1643, n1361, n1275);
or   g2275 (n2471, n1564, n1715, n1425, n1246);
nor  g2276 (n2294, n1257, n1775, n1314, n1363);
nor  g2277 (n2458, n1242, n1304, n1548, n1537);
xnor g2278 (n2484, n1323, n1296, n1788, n1354);
xnor g2279 (n2718, n1326, n1688, n1479, n1782);
xnor g2280 (n2516, n1745, n1696, n1811, n1388);
or   g2281 (n1869, n1253, n1381, n1280, n1476);
and  g2282 (n2138, n1757, n1239, n1695, n1634);
and  g2283 (n2123, n1788, n1724, n1512, n1645);
xor  g2284 (n2089, n1469, n1535, n1421, n1565);
xor  g2285 (n2730, n1665, n1497, n1499, n1477);
or   g2286 (n2117, n1262, n1367, n1781, n1321);
nor  g2287 (n1923, n1673, n1394, n1261, n1503);
or   g2288 (n2216, n1276, n1758, n1435, n1409);
xor  g2289 (n2151, n1346, n1586, n1559, n1728);
and  g2290 (n2250, n1762, n1604, n1493, n1549);
and  g2291 (n2198, n1259, n1560, n1318, n1365);
xor  g2292 (n2559, n1780, n1816, n1590, n1266);
nand g2293 (n2615, n1307, n1579, n1540, n1803);
or   g2294 (n2042, n1812, n1593, n1517, n1721);
xor  g2295 (n1971, n1364, n1652, n1477, n1412);
nor  g2296 (n1893, n1635, n1343, n1515, n1805);
and  g2297 (n2178, n1400, n1533, n1676, n1713);
or   g2298 (n2644, n1556, n1781, n1525, n1687);
xnor g2299 (n1917, n1536, n1638, n1821, n1820);
or   g2300 (n2738, n1461, n1837, n1524, n1571);
xor  g2301 (n2490, n1414, n1340, n1303, n1661);
xor  g2302 (n2040, n1670, n1694, n1305, n1562);
or   g2303 (n1904, n1273, n1735, n1580, n1528);
nand g2304 (n2414, n1658, n1448, n1277, n1317);
xnor g2305 (n2725, n1415, n1802, n1763, n1450);
nor  g2306 (n2209, n1299, n1664, n1442, n1836);
xor  g2307 (n1862, n1236, n1473, n1615, n1504);
or   g2308 (n2107, n1552, n1360, n1835, n1312);
nor  g2309 (n2431, n1403, n1329, n1648, n1754);
or   g2310 (n2454, n1518, n1320, n1675, n1760);
xor  g2311 (n2267, n1789, n1718, n1795, n1424);
xor  g2312 (n1878, n1591, n1282, n1812, n1275);
nor  g2313 (n1852, n1667, n1727, n1354, n1462);
and  g2314 (n1983, n1416, n1363, n1353, n1812);
xnor g2315 (n1996, n1733, n326, n1728, n1662);
xor  g2316 (n2139, n1623, n1509, n1829, n1419);
nor  g2317 (n2515, n1808, n1620, n1438, n1387);
nor  g2318 (n2044, n1385, n1397, n1570, n1663);
nand g2319 (n2388, n1366, n1547, n1248, n1801);
and  g2320 (n2289, n1581, n1308, n1575, n1685);
nor  g2321 (n2335, n1702, n1350, n1529, n1781);
or   g2322 (n2026, n1833, n1444, n1410, n1672);
xnor g2323 (n2601, n1680, n1440, n1644, n1684);
and  g2324 (n1972, n1791, n1495, n1415, n1738);
xnor g2325 (n2344, n1445, n1767, n1698, n1372);
nor  g2326 (n1875, n1453, n1306, n1621, n1296);
and  g2327 (n1907, n1442, n1360, n1611, n1625);
nor  g2328 (n1897, n1664, n1608, n1527, n1714);
xnor g2329 (n2354, n1704, n1727, n1324, n1657);
nor  g2330 (n2701, n1292, n1614, n1314, n1731);
nor  g2331 (n2102, n1806, n1753, n1469, n1688);
or   g2332 (n2546, n1598, n1295, n1573, n1668);
xor  g2333 (n2214, n1761, n1560, n1799, n1345);
xnor g2334 (n2064, n1552, n1431, n1402, n1710);
xor  g2335 (n1988, n1467, n1725, n1383, n1342);
xnor g2336 (n2327, n1351, n1333, n1808, n1603);
nand g2337 (n2085, n1796, n1240, n1409, n1711);
xnor g2338 (n2382, n1336, n1427, n1352, n1438);
or   g2339 (n1909, n1335, n1840, n1599, n1429);
or   g2340 (n2667, n1610, n1525, n1408, n1708);
or   g2341 (n1954, n1685, n1382, n1671, n1732);
nand g2342 (n2241, n1310, n1776, n1613, n1543);
xnor g2343 (n2012, n1810, n1567, n1250, n1502);
nand g2344 (n2018, n1602, n1479, n1388, n1258);
and  g2345 (n2671, n1740, n1826, n1535, n1480);
or   g2346 (n2577, n1679, n1355, n1581, n1729);
or   g2347 (n2150, n1813, n1638, n1567, n1414);
xnor g2348 (n2438, n1544, n1325, n1797, n1820);
xnor g2349 (n2717, n1419, n1263, n1301, n1534);
xor  g2350 (n2534, n1672, n698, n1798);
xor  g2351 (n2623, n1806, n1827, n1836, n1332);
nor  g2352 (n2400, n1562, n1517, n1523, n1595);
xnor g2353 (n2087, n1562, n1508, n1775, n1598);
xnor g2354 (n2401, n1344, n1700, n1383, n1349);
xnor g2355 (n2145, n1466, n1636, n1401, n1342);
and  g2356 (n2275, n1562, n1801, n1613, n1772);
or   g2357 (n2236, n1778, n1814, n1621, n1565);
and  g2358 (n2187, n1297, n1390, n1504, n1428);
and  g2359 (n1935, n1833, n1241, n1827, n1778);
nor  g2360 (n2432, n1359, n1823, n1773, n1686);
nor  g2361 (n2238, n1369, n1623, n1300, n1365);
nand g2362 (n2091, n1384, n1239, n1359, n1768);
nand g2363 (n2303, n1827, n1740, n1626, n1337);
xor  g2364 (n2405, n1678, n1474, n1257, n1619);
xnor g2365 (n2591, n1270, n1265, n1719, n1272);
xor  g2366 (n2729, n1600, n1661, n1839, n1564);
nand g2367 (n1884, n1500, n1647, n1458, n1507);
nor  g2368 (n1986, n1838, n1259, n1542, n1695);
xor  g2369 (n2477, n1763, n1610, n1488, n1368);
nor  g2370 (n2660, n1385, n1764, n1490, n1547);
xor  g2371 (n2204, n1413, n1748, n1572, n1375);
xnor g2372 (n2678, n1706, n1401, n1479, n1295);
and  g2373 (n2076, n1433, n1245, n1250, n1423);
and  g2374 (n2711, n1304, n1616, n1583, n1316);
nor  g2375 (n2297, n1496, n1468, n1267, n1576);
or   g2376 (n2658, n1682, n1594, n1826, n1328);
and  g2377 (n2219, n1588, n1769, n1715, n1478);
xor  g2378 (n2337, n1281, n1552, n1498, n1642);
nor  g2379 (n2739, n1835, n1481, n1503, n1449);
or   g2380 (n2662, n1396, n1676, n1504, n1456);
nor  g2381 (n2130, n1835, n1821, n1631, n1327);
nand g2382 (n2072, n1700, n1471, n1733, n1412);
nand g2383 (n1855, n1696, n1829, n1558, n1680);
or   g2384 (n2699, n1398, n1737, n1401, n1472);
or   g2385 (n1961, n1672, n1725, n1496, n1617);
xor  g2386 (n2255, n1660, n1422, n1471, n1736);
or   g2387 (n1913, n1711, n1289, n1361, n1639);
xor  g2388 (n2630, n1426, n1717, n1819, n1522);
or   g2389 (n2100, n1768, n1660, n1619, n1266);
and  g2390 (n2409, n1712, n1261, n1792, n1671);
nand g2391 (n2519, n1606, n1299, n1235, n1399);
nor  g2392 (n2478, n1597, n1768, n1565, n1773);
and  g2393 (n2088, n1711, n1546, n1797, n1482);
xor  g2394 (n2129, n1288, n1338, n1659, n1586);
xnor g2395 (n2387, n1811, n1513, n1817, n1245);
or   g2396 (n2613, n1656, n1753, n1294, n1348);
nor  g2397 (n2362, n1724, n1694, n1684, n1698);
xnor g2398 (n2681, n1410, n1497, n1420, n1430);
xnor g2399 (n1967, n1700, n1566, n1567, n1381);
xor  g2400 (n2610, n1838, n1380, n1741, n1373);
xor  g2401 (n2443, n1590, n1659, n1447, n1416);
xor  g2402 (n2686, n1510, n1254, n1758, n1334);
nand g2403 (n2099, n1532, n1709, n1429, n1841);
and  g2404 (n2277, n326, n325, n1268, n1301);
and  g2405 (n2439, n1400, n1489, n1531, n1597);
and  g2406 (n2037, n1530, n1521, n1427, n1713);
and  g2407 (n2705, n1391, n1631, n1502, n1388);
nor  g2408 (n2090, n1256, n1391, n1348, n1280);
or   g2409 (n2548, n1282, n1417, n1343, n1837);
or   g2410 (n1965, n1735, n1434, n1436, n1564);
xnor g2411 (n1991, n1810, n1497, n1425, n1293);
nand g2412 (n2078, n1421, n1281, n1249, n1389);
nand g2413 (n2653, n1487, n1786, n1422, n1624);
nor  g2414 (n2317, n1450, n1739, n1254, n1674);
nor  g2415 (n2253, n1805, n1600, n1284, n1584);
or   g2416 (n2445, n1515, n1453, n1270, n1550);
xor  g2417 (n2608, n1290, n1468, n1553, n1828);
or   g2418 (n2288, n1699, n1713, n1504, n1786);
xor  g2419 (n1873, n1428, n1639, n1484, n1820);
xnor g2420 (n2625, n1665, n1663, n1807, n1445);
xor  g2421 (n2177, n1283, n1488, n1439, n1512);
xnor g2422 (n1958, n1632, n1461, n1627, n1746);
nand g2423 (n2507, n1683, n1371, n1238, n1608);
xor  g2424 (n2668, n1374, n1483, n1704, n1481);
or   g2425 (n2734, n1469, n1331, n1377, n1573);
nor  g2426 (n2061, n1804, n1615, n1817, n1792);
nand g2427 (n1879, n1581, n1767, n1387, n1259);
or   g2428 (n2210, n1591, n1498, n1537, n1688);
nand g2429 (n2322, n1784, n1730, n1835, n1489);
nand g2430 (n2595, n1599, n1573, n1507, n1755);
nor  g2431 (n1927, n1519, n1303, n1788, n1512);
and  g2432 (n2727, n1304, n1473, n1671, n1255);
or   g2433 (n2273, n1578, n1465, n1440, n1242);
or   g2434 (n2036, n1293, n1550, n1519, n1784);
xnor g2435 (n2358, n1704, n1320, n1577, n1445);
and  g2436 (n2105, n1514, n1292, n1769, n1789);
or   g2437 (n2460, n1513, n1282, n1436, n1679);
and  g2438 (n1953, n1657, n1692, n1443, n1495);
nor  g2439 (n2691, n1756, n1630, n1538);
nor  g2440 (n2487, n1612, n1809, n1516, n1422);
xor  g2441 (n2541, n1669, n1400, n1457, n1635);
and  g2442 (n2468, n1752, n1348, n1657, n1644);
xnor g2443 (n2095, n1429, n1703, n1559, n1378);
xnor g2444 (n2314, n1281, n1423, n1406, n1508);
nand g2445 (n2528, n1789, n1645, n1611, n1515);
and  g2446 (n1968, n1731, n1815, n1655, n1739);
nor  g2447 (n2227, n1481, n1783, n1455, n1754);
xor  g2448 (n2032, n1383, n1254, n1235, n1468);
xor  g2449 (n2346, n1453, n1838, n1266, n1616);
xor  g2450 (n1843, n1394, n1339, n1841, n1665);
xor  g2451 (n2348, n1315, n1247, n1675, n1537);
and  g2452 (n2446, n1300, n1665, n1649, n1269);
xnor g2453 (n2406, n1815, n1793, n1444, n1502);
or   g2454 (n2245, n326, n1804, n1362, n1702);
xor  g2455 (n2696, n1477, n1589, n1723, n1629);
nand g2456 (n2112, n1587, n1801, n1463, n1575);
and  g2457 (n2500, n1305, n1339, n1252, n1732);
nor  g2458 (n2392, n1432, n1618, n1510, n1534);
xnor g2459 (n2174, n1674, n1816, n1494, n1289);
xor  g2460 (n2669, n1245, n1637, n1519, n1825);
and  g2461 (n2185, n1382, n1640, n1617, n1697);
xor  g2462 (n2740, n1553, n1329, n1302, n1336);
nand g2463 (n2522, n1642, n1320, n1585, n1290);
or   g2464 (n2258, n1355, n1592, n1715, n1743);
nor  g2465 (n2496, n1825, n1524, n1706, n1286);
nand g2466 (n2735, n1698, n1489, n1643, n1511);
xnor g2467 (n2708, n1706, n1257, n1786, n1344);
or   g2468 (n2025, n1285, n1386, n1464, n1611);
nor  g2469 (n1964, n1748, n1646, n1606, n1333);
xor  g2470 (n2590, n1814, n1705, n1640, n1324);
nor  g2471 (n2453, n1837, n1392, n1558, n1263);
xnor g2472 (n2661, n1526, n1544, n1646, n1679);
xnor g2473 (n2300, n1298, n1713, n1809, n1627);
xor  g2474 (n2356, n1485, n1692, n1787, n1426);
xnor g2475 (n1896, n1305, n1714, n1258, n1674);
xor  g2476 (n1866, n1247, n1420, n1577, n1579);
nor  g2477 (n2050, n1664, n1286, n1744, n1506);
xnor g2478 (n2527, n1698, n1310, n1689, n1491);
nand g2479 (n2537, n1238, n1561, n1375, n1473);
and  g2480 (n2418, n1328, n1716, n1487, n1415);
nand g2481 (n2092, n1256, n1403, n1670, n1257);
xnor g2482 (n2208, n1441, n1592, n1494, n1491);
nor  g2483 (n1880, n1813, n1414, n1566, n1681);
xor  g2484 (n2142, n1447, n1246, n1785, n1449);
or   g2485 (n2474, n1244, n1388, n1511, n1601);
nand g2486 (n2051, n1369, n1684, n1735, n1765);
xor  g2487 (n2641, n1466, n1710, n1653, n1350);
nor  g2488 (n2244, n1420, n1770, n1279, n1297);
or   g2489 (n2563, n1703, n1753, n1638, n1778);
nand g2490 (n2341, n1554, n1327, n1498, n1287);
xor  g2491 (n1939, n1304, n1626, n1669, n1789);
xor  g2492 (n2554, n1425, n1561, n1387, n1842);
or   g2493 (n2451, n1684, n1336, n1599, n1622);
xnor g2494 (n2643, n1826, n1414, n1248, n1514);
and  g2495 (n2540, n1649, n1619, n1716, n1490);
nand g2496 (n2124, n1291, n1236, n1548, n1549);
and  g2497 (n2605, n1749, n1658, n1338, n1318);
xnor g2498 (n2246, n1814, n1316, n1506, n1755);
xnor g2499 (n2320, n1417, n1803, n1596, n1788);
and  g2500 (n2343, n1825, n1618, n1312, n1404);
nand g2501 (n2084, n1243, n1417, n1296, n1428);
xnor g2502 (n2339, n1840, n1545, n1707, n1728);
and  g2503 (n2071, n1692, n1352, n1475, n1391);
nor  g2504 (n1980, n1355, n1432, n1733, n1419);
nand g2505 (n2427, n1630, n1519, n1459, n1241);
or   g2506 (n1937, n1322, n1436, n1435, n1582);
or   g2507 (n2180, n1433, n1538, n1669, n1717);
or   g2508 (n2282, n1567, n1812, n1739, n1588);
and  g2509 (n2111, n691, n1495, n1821, n1389);
and  g2510 (n2411, n1598, n1313, n1362, n1803);
or   g2511 (n2141, n1525, n1466, n1839, n1613);
and  g2512 (n2398, n1403, n1263, n1600, n1782);
nor  g2513 (n2413, n1561, n1374, n1686, n1251);
and  g2514 (n2737, n1290, n1287, n693, n1803);
nand g2515 (n2575, n1367, n1736, n1359, n1699);
or   g2516 (n2492, n1253, n1360, n1547, n1546);
xor  g2517 (n2011, n1628, n1624, n1776, n695);
xor  g2518 (n2589, n1496, n1349, n1242, n1809);
and  g2519 (n2395, n1240, n1568, n1278, n1724);
xnor g2520 (n2149, n1794, n1395, n1738, n1530);
xor  g2521 (n1874, n1823, n1701, n1370, n1450);
xnor g2522 (n2052, n1405, n1272, n1745, n1242);
xor  g2523 (n1881, n1834, n1651, n1515, n1676);
or   g2524 (n2378, n1413, n1391, n1770, n1687);
and  g2525 (n2698, n1449, n1693, n1607, n1377);
or   g2526 (n2631, n1430, n1370, n1509, n1518);
and  g2527 (n2315, n1760, n1299, n1718, n1308);
xnor g2528 (n2347, n1585, n1283, n1829, n1654);
and  g2529 (n2648, n1621, n1411, n1472, n1325);
and  g2530 (n2433, n1792, n1454, n1751, n1761);
nor  g2531 (n2041, n1679, n1307, n1704, n1406);
or   g2532 (n2345, n1772, n1780, n1538, n1625);
or   g2533 (n2308, n1261, n1495, n1511, n1240);
xnor g2534 (n1895, n1654, n1578, n1619, n1361);
nor  g2535 (n2016, n1329, n1501, n1491, n1376);
nand g2536 (n2158, n1543, n1831, n1359, n1677);
nand g2537 (n1849, n1804, n1696, n1572, n1534);
nor  g2538 (n2137, n1317, n1347, n1520, n1439);
nand g2539 (n2189, n1833, n1746, n1492, n1361);
xor  g2540 (n2006, n1728, n1707, n1811, n1331);
nor  g2541 (n2437, n1705, n1767, n1756, n1546);
or   g2542 (n2637, n1591, n1294, n1661, n1255);
and  g2543 (n2684, n1448, n1279, n1560, n1456);
xnor g2544 (n2670, n1814, n1815, n1771, n1833);
nor  g2545 (n2034, n1417, n1522, n1494, n1707);
xnor g2546 (n2422, n1678, n1629, n1386, n1633);
or   g2547 (n1845, n1510, n1583, n1750, n1744);
or   g2548 (n2617, n1741, n1578, n1800, n1551);
nor  g2549 (n2057, n1501, n1577, n1690, n1609);
xor  g2550 (n2587, n1662, n1380, n1816, n1478);
xnor g2551 (n2170, n1602, n1651, n1748, n1451);
or   g2552 (n2033, n1807, n1545, n1593, n1540);
or   g2553 (n2363, n1385, n1645, n1690, n1499);
or   g2554 (n1918, n1447, n1714, n1431, n1795);
or   g2555 (n1876, n1298, n1576, n1469, n1675);
or   g2556 (n2429, n1237, n1326, n1290, n1405);
xnor g2557 (n2160, n1345, n1819, n1777, n1774);
nand g2558 (n2230, n1329, n1260, n1289, n1442);
nand g2559 (n2665, n1752, n1474, n1439, n1750);
xor  g2560 (n2287, n1779, n1838, n1595, n1610);
nand g2561 (n1859, n1307, n1807, n1588, n1551);
xor  g2562 (n1981, n1520, n1764, n1593, n1396);
xnor g2563 (n2305, n1346, n1637, n1256, n1708);
xor  g2564 (n2604, n1557, n1351, n1596, n1407);
xor  g2565 (n1930, n1358, n1428, n1590, n1608);
and  g2566 (n2201, n1603, n1291, n1324, n1749);
xnor g2567 (n2570, n1673, n1397, n1697, n1311);
nand g2568 (n2466, n1642, n1277, n1807, n1719);
nor  g2569 (n1848, n1393, n1609, n1582, n1272);
nand g2570 (n2369, n1658, n1780, n1452, n1327);
and  g2571 (n2728, n1394, n1363, n1633, n1272);
or   g2572 (n2097, n1671, n1440, n1745, n1685);
xor  g2573 (n2704, n1244, n1624, n1601, n1368);
xor  g2574 (n2567, n1512, n1310, n1766, n1631);
or   g2575 (n2035, n1699, n1559, n1370, n1642);
xor  g2576 (n2402, n1309, n1628, n1369, n1736);
or   g2577 (n2290, n1378, n1694, n1622, n1330);
nor  g2578 (n2200, n1796, n1677, n1775, n1712);
nand g2579 (n2596, n1292, n1790, n1603, n1570);
xor  g2580 (n1846, n1792, n1379, n1832, n1762);
xnor g2581 (n2407, n1501, n1805, n1790, n1325);
nor  g2582 (n1925, n1797, n1818, n1506, n1521);
nand g2583 (n2556, n1686, n1726, n1496, n1714);
xnor g2584 (n2375, n1297, n1438, n1791, n1766);
or   g2585 (n2444, n1652, n1596, n1601, n1557);
nor  g2586 (n2122, n1399, n1601, n1791, n1401);
nor  g2587 (n2190, n1635, n1554, n1317, n1451);
xnor g2588 (n1933, n1783, n1754, n1616, n1415);
nor  g2589 (n2627, n699, n1551, n1721, n1653);
or   g2590 (n2483, n1287, n1418, n1431, n1693);
nand g2591 (n2274, n1485, n1503, n1373, n1277);
and  g2592 (n2695, n1828, n1595, n1486, n1529);
nor  g2593 (n2261, n1412, n1826, n1313, n1475);
and  g2594 (n2066, n1711, n1383, n1799, n1810);
nor  g2595 (n2376, n1529, n1480, n1340, n1569);
nor  g2596 (n2428, n1236, n1718, n1335, n1501);
and  g2597 (n2580, n1434, n1264, n1822, n1683);
nand g2598 (n2286, n1461, n1517, n1524, n1633);
xnor g2599 (n2456, n1566, n1345, n1678, n1547);
or   g2600 (n2106, n1408, n1630, n1607, n1758);
nor  g2601 (n2193, n1531, n1483, n1441, n1804);
xor  g2602 (n2525, n1507, n1522, n1557, n1723);
or   g2603 (n2217, n1751, n1790, n1262, n1732);
or   g2604 (n2067, n1726, n1372, n1385, n1526);
xor  g2605 (n1854, n1403, n1579, n1460, n1286);
nand g2606 (n2010, n1620, n1824, n1485, n1575);
xor  g2607 (n2154, n1456, n1730, n1315, n1536);
and  g2608 (n2173, n325, n1598, n1585, n1318);
xor  g2609 (n2368, n1250, n1824, n1723, n1580);
xor  g2610 (n2517, n1607, n1604, n1798, n1829);
xnor g2611 (n2349, n1357, n1680, n1740, n1525);
and  g2612 (n1892, n1459, n1467, n1613, n1458);
and  g2613 (n2188, n1834, n1341, n1314, n1253);
xor  g2614 (n2195, n1808, n1483, n1337, n1446);
nand g2615 (n2009, n1349, n1553, n1830, n1626);
or   g2616 (n2421, n1420, n1699, n1559, n1836);
xor  g2617 (n2082, n1805, n1831, n1540, n1825);
or   g2618 (n2302, n1608, n1539, n1382, n1605);
nor  g2619 (n2713, n1748, n1555, n1721, n1404);
xnor g2620 (n2550, n1540, n1490, n1569, n1648);
nand g2621 (n2461, n1743, n1493, n1462, n1313);
xor  g2622 (n2384, n1725, n1586, n1528, n1382);
or   g2623 (n2664, n1716, n1734, n1527, n1283);
xnor g2624 (n1990, n1563, n1457, n1538, n1460);
xnor g2625 (n2027, n1782, n1813, n1275, n1773);
nor  g2626 (n2118, n1374, n1643, n1722, n1710);
nor  g2627 (n2479, n1492, n1255, n1796, n1639);
nand g2628 (n2599, n1313, n1407, n1342, n1831);
nor  g2629 (n2381, n1756, n1736, n1372, n1761);
or   g2630 (n2247, n1842, n1664, n1288, n1641);
and  g2631 (n2049, n1800, n1544, n1691, n1737);
xnor g2632 (n2342, n1421, n1817, n1660, n1646);
xor  g2633 (n2002, n1651, n1284, n1453, n1546);
nand g2634 (n2709, n1520, n1270, n1787, n1568);
nand g2635 (n2370, n1457, n1399, n1686, n1676);
xor  g2636 (n2001, n1265, n1475, n1625, n1249);
nor  g2637 (n2256, n1703, n1584, n1342, n1518);
xnor g2638 (n2620, n1245, n1341, n1380, n1585);
xor  g2639 (n2486, n1754, n1267, n1330, n1260);
and  g2640 (n2162, n1655, n1790, n1606, n1806);
or   g2641 (n2419, n1685, n1518, n1733, n1618);
nor  g2642 (n2597, n1839, n1840, n1505, n1659);
xnor g2643 (n2600, n1563, n1492, n1517);
nor  g2644 (n2464, n1455, n1375, n1777, n1623);
or   g2645 (n2442, n1441, n1722, n1243, n1371);
nor  g2646 (n2331, n1750, n1777, n1446, n1565);
or   g2647 (n2404, n694, n1552, n1424, n1458);
xor  g2648 (n1916, n1369, n1742, n1751, n1569);
xor  g2649 (n2226, n1742, n1708, n1795, n1239);
and  g2650 (n2161, n1523, n1701, n1426, n1465);
or   g2651 (n2632, n1371, n1749, n1738, n1416);
nor  g2652 (n1853, n1555, n1667, n1662, n1802);
nor  g2653 (n2494, n1539, n1576, n1584, n1253);
xnor g2654 (n2733, n1675, n1464, n1687, n1586);
xnor g2655 (n2330, n1753, n1331, n1561, n1697);
xnor g2656 (n1920, n1322, n1392, n1558, n1563);
nand g2657 (n2309, n1650, n1615, n1358, n1836);
xor  g2658 (n2693, n1637, n1841, n1532, n1393);
xor  g2659 (n2205, n1285, n1252, n1303, n1757);
and  g2660 (n2328, n1660, n1794, n1640, n1783);
xnor g2661 (n1870, n1237, n1263, n1349, n1649);
xor  g2662 (n2269, n1260, n1351, n1819, n1712);
nand g2663 (n2096, n1802, n1521, n1760, n1254);
and  g2664 (n2171, n1727, n1368, n1652, n1356);
xor  g2665 (n2047, n1706, n1605, n1661, n1444);
and  g2666 (n2459, n1697, n1795, n1354, n1471);
nor  g2667 (n1936, n1259, n1715, n1764, n1656);
nand g2668 (n2008, n1709, n1589, n1274, n1309);
xnor g2669 (n2645, n1639, n1343, n1656, n1783);
xnor g2670 (n2703, n1430, n1737, n1408, n1793);
xnor g2671 (n1885, n1637, n1571, n1446, n1636);
nand g2672 (n2080, n1653, n1541, n1487, n1654);
xnor g2673 (n2169, n1393, n1402, n1666, n1612);
xor  g2674 (n2579, n1252, n1614, n1674, n1653);
and  g2675 (n2633, n1842, n1377, n1334, n1593);
nand g2676 (n1957, n1437, n1295, n1551, n1516);
or   g2677 (n2441, n1411, n1312, n1597, n1707);
nor  g2678 (n2529, n1432, n1341, n1488, n1500);
nand g2679 (n2480, n1265, n1682, n1531, n1284);
nand g2680 (n1989, n1467, n1380, n1474, n1458);
and  g2681 (n2156, n1723, n1268, n1291, n1311);
xor  g2682 (n2622, n1266, n1819, n1820, n1318);
nor  g2683 (n2408, n1281, n1554, n1346, n1482);
and  g2684 (n2334, n1832, n1237, n1627, n1647);
xnor g2685 (n2440, n1278, n1433, n1681, n1271);
nor  g2686 (n2512, n1571, n1687, n1614, n1340);
and  g2687 (n2202, n1308, n1434, n1390, n1459);
and  g2688 (n2569, n1824, n1300, n1772, n1794);
or   g2689 (n2240, n1768, n1247, n1516, n1574);
xnor g2690 (n2005, n1435, n1541, n1636, n1548);
xor  g2691 (n1890, n1494, n1791, n1796, n1555);
xnor g2692 (n2167, n1294, n1274, n1460, n1457);
xor  g2693 (n2524, n1743, n1554, n1742, n1566);
nor  g2694 (n2281, n1693, n1574, n1264, n1742);
or   g2695 (n2677, n1632, n1502, n1622, n1390);
nor  g2696 (n2523, n1841, n1316, n1296, n1591);
nand g2697 (n2271, n1644, n1434, n1570, n1374);
nand g2698 (n2472, n1677, n1572, n1443, n1605);
nand g2699 (n1945, n1556, n1689, n1568, n1526);
xor  g2700 (n2679, n1823, n1429, n1362, n1392);
nand g2701 (n2194, n1757, n1569, n1722, n1317);
nor  g2702 (n1966, n1367, n1472, n1700, n1810);
or   g2703 (n1922, n1427, n1717, n1634, n1537);
and  g2704 (n2722, n1539, n1682, n1249);
xor  g2705 (n2581, n1779, n1426, n1545, n1818);
xor  g2706 (n2592, n1771, n1531, n1459, n1762);
nand g2707 (n2624, n1647, n1779, n1641, n1506);
or   g2708 (n2374, n1759, n1430, n1787, n1645);
xnor g2709 (n2237, n1421, n1276, n1326, n1560);
xor  g2710 (n2759, n2583, n2649, n2240, n2472);
xnor g2711 (n2843, n2328, n1938, n2007, n2391);
nor  g2712 (n2877, n2461, n1883, n2224, n2248);
and  g2713 (n2948, n1921, n2553, n2283, n1999);
nand g2714 (n2938, n1848, n1893, n1924, n2421);
nor  g2715 (n2859, n2424, n2161, n2302, n2419);
xnor g2716 (n2762, n2278, n1869, n2318, n2418);
xnor g2717 (n2826, n2093, n2732, n2355, n2662);
nand g2718 (n2802, n2217, n2001, n2625, n2674);
nand g2719 (n2896, n2104, n2544, n1992, n2048);
xor  g2720 (n2797, n2180, n2020, n1941, n2075);
xor  g2721 (n2815, n2229, n2575, n2271, n2399);
or   g2722 (n2747, n2463, n2037, n2734, n2322);
nor  g2723 (n2867, n2353, n2651, n2617, n2367);
xnor g2724 (n2920, n2289, n2022, n2584, n2525);
xor  g2725 (n2894, n2492, n2469, n2491, n2496);
xor  g2726 (n2927, n2394, n2687, n1975, n2276);
nor  g2727 (n2880, n2202, n2608, n1881, n2524);
and  g2728 (n2871, n2571, n2639, n2646, n2573);
nand g2729 (n2842, n2210, n2142, n2017, n2696);
xnor g2730 (n2918, n2168, n2249, n2281, n1948);
xnor g2731 (n2804, n2432, n2666, n2585, n2434);
and  g2732 (n2813, n2582, n2170, n2008, n2404);
and  g2733 (n2828, n2659, n2056, n2678, n2543);
nor  g2734 (n2866, n2262, n2728, n2580, n2264);
xor  g2735 (n2757, n2645, n1991, n2416, n2272);
nor  g2736 (n2962, n2489, n1933, n2122, n2237);
or   g2737 (n2822, n2299, n2174, n2140, n2233);
xor  g2738 (n2890, n2077, n2657, n2596, n2603);
nand g2739 (n2929, n2516, n2201, n2088, n2471);
xor  g2740 (n2964, n2736, n1942, n2671, n2589);
xor  g2741 (n2936, n2092, n2107, n2166, n2258);
or   g2742 (n2963, n2673, n2396, n1854, n2356);
xnor g2743 (n2892, n2268, n2214, n2740, n2400);
or   g2744 (n2772, n2035, n2119, n1979, n2117);
nand g2745 (n2833, n1954, n2371, n1982, n2440);
nand g2746 (n2899, n2043, n2655, n2733, n2708);
xnor g2747 (n2841, n2096, n2621, n2228, n1958);
nand g2748 (n2916, n2537, n2338, n2449, n2000);
or   g2749 (n2887, n2422, n1960, n2635, n2173);
and  g2750 (n2906, n2405, n2231, n2197, n1949);
nor  g2751 (n2873, n2724, n1931, n2482, n2612);
nand g2752 (n2967, n2343, n2390, n2392, n2504);
nor  g2753 (n2799, n2716, n2118, n2175, n2176);
nor  g2754 (n2809, n2604, n2131, n2642, n1962);
and  g2755 (n2817, n2535, n2501, n2026, n2212);
xor  g2756 (n2749, n2196, n1852, n1936, n2398);
nand g2757 (n2898, n2622, n2607, n1914, n2374);
nand g2758 (n2746, n2663, n2742, n1873, n2234);
xnor g2759 (n2954, n2139, n2133, n2610, n2187);
xnor g2760 (n2825, n1973, n2699, n2366, n2206);
and  g2761 (n2788, n2102, n1970, n2448, n2559);
nor  g2762 (n2770, n2536, n2569, n2063, n2619);
or   g2763 (n2876, n2379, n2047, n2316, n1887);
and  g2764 (n2888, n2285, n2567, n2339, n2042);
nand g2765 (n2748, n2305, n2055, n2557, n2221);
xnor g2766 (n2956, n2114, n1910, n2383, n2279);
nand g2767 (n2824, n1985, n2222, n2467, n2576);
xnor g2768 (n2782, n2451, n2199, n2251, n2123);
nor  g2769 (n2926, n1909, n1906, n2508, n2522);
or   g2770 (n2919, n2713, n2479, n2311, n1971);
or   g2771 (n2756, n1986, n2453, n2541, n2255);
nand g2772 (n2844, n2287, n2074, n2406, n2694);
xor  g2773 (n2901, n2637, n2465, n1972, n2125);
xor  g2774 (n2860, n2679, n2417, n2433, n2376);
xor  g2775 (n2847, n2677, n2510, n2534, n2286);
nand g2776 (n2765, n2352, n2223, n1871, n2160);
and  g2777 (n2811, n2384, n2599, n2359, n2475);
xor  g2778 (n2784, n2632, n2638, n2079, n2239);
nand g2779 (n2839, n2113, n2130, n2216, n2413);
xnor g2780 (n2837, n2314, n1969, n2200, n2532);
or   g2781 (n2800, n2184, n1859, n2073, n2336);
nor  g2782 (n2853, n2132, n2207, n2193, n2623);
nand g2783 (n2775, n2739, n2257, n2238, n2360);
and  g2784 (n2777, n2064, n2148, n2235, n2085);
and  g2785 (n2925, n2128, n2049, n2014, n2312);
nor  g2786 (n2870, n2277, n2083, n2034, n2372);
or   g2787 (n2801, n1862, n2024, n1880, n2362);
nor  g2788 (n2760, n1901, n2426, n2293, n2052);
xor  g2789 (n2763, n2566, n2253, n1884, n2420);
or   g2790 (n2908, n2065, n2704, n2163, n2613);
nand g2791 (n2862, n1951, n2317, n2511, n2038);
or   g2792 (n2803, n2296, n2149, n2298, n2552);
xor  g2793 (n2856, n2533, n2466, n2388, n2514);
nand g2794 (n2814, n2560, n2507, n2668, n2661);
xor  g2795 (n2780, n2630, n2361, n2436, n2072);
xnor g2796 (n2829, n2615, n2150, n2660, n2445);
xor  g2797 (n2924, n2647, n2454, n2058, n1998);
nand g2798 (n2818, n2016, n2636, n2194, n2124);
xor  g2799 (n2806, n2529, n2040, n2045, n1963);
xor  g2800 (n2827, n2246, n2452, n2313, n1965);
nand g2801 (n2965, n2368, n2597, n1851, n1959);
nor  g2802 (n2744, n2209, n2681, n1858, n2334);
nor  g2803 (n2850, n2342, n2204, n2171, n1930);
nor  g2804 (n2861, n2387, n2067, n2493, n2377);
and  g2805 (n2937, n2628, n2078, n2331, n2477);
and  g2806 (n2830, n1964, n2731, n2593, n1892);
nand g2807 (n2957, n1866, n1987, n2301, n2151);
xor  g2808 (n2789, n1879, n2005, n1856, n2137);
nand g2809 (n2879, n2698, n2664, n2087, n2550);
nand g2810 (n2947, n1950, n2715, n2185, n2198);
nand g2811 (n2851, n1870, n2592, n2155, n2270);
and  g2812 (n2914, n2680, n2021, n2308, n2157);
xnor g2813 (n2928, n2478, n2203, n2676, n2578);
xnor g2814 (n2889, n2494, n2480, n1983, n1947);
or   g2815 (n2904, n2503, n2505, n1894, n2211);
and  g2816 (n2755, n2069, n2627, n1853, n2685);
nand g2817 (n2753, n2460, n2428, n1882, n2588);
nand g2818 (n2805, n2332, n1925, n2030, n2675);
and  g2819 (n2907, n2714, n2488, n2425, n2284);
nand g2820 (n2774, n2054, n1943, n2089, n2523);
and  g2821 (n2840, n2564, n2294, n2225, n2656);
nor  g2822 (n2790, n2561, n2385, n2178, n2126);
xor  g2823 (n2934, n2654, n2689, n2036, n1913);
xor  g2824 (n2786, n2023, n2003, n2141, n1995);
xnor g2825 (n2821, n1927, n2407, n2230, n1976);
nand g2826 (n2878, n2373, n2241, n2586, n2183);
and  g2827 (n2791, n2315, n2252, n2723, n1996);
and  g2828 (n2798, n2147, n2401, n2061, n1946);
and  g2829 (n2783, n2098, n1896, n2236, n2068);
nor  g2830 (n2951, n2509, n2046, n2669, n2062);
and  g2831 (n2778, n2520, n1867, n2389, n2134);
and  g2832 (n2958, n1863, n2004, n2429, n2354);
or   g2833 (n2903, n2295, n2340, n2190, n2050);
nand g2834 (n2751, n2365, n2327, n2375, n2730);
nand g2835 (n2750, n2690, n2410, n1874, n2718);
xnor g2836 (n2881, n2084, n2347, n2563, n2414);
or   g2837 (n2885, n1865, n2542, n2324, n1868);
and  g2838 (n2776, n2476, n2691, n2227, n1897);
nor  g2839 (n2913, n2634, n2136, n2297, n2033);
and  g2840 (n2931, n2409, n2403, n2572, n2412);
or   g2841 (n2909, n2152, n2427, n1916, n1945);
nand g2842 (n2942, n2738, n1989, n2261, n2737);
or   g2843 (n2820, n2620, n2039, n2288, n2456);
nand g2844 (n2882, n2146, n2013, n1915, n1847);
xnor g2845 (n2868, n1952, n2591, n1926, n2344);
nand g2846 (n2810, n2051, n1978, n2162, n2540);
and  g2847 (n2943, n1935, n1898, n2473, n2602);
nor  g2848 (n2854, n1994, n2325, n2310, n2722);
nor  g2849 (n2796, n2244, n1939, n2626, n2629);
nor  g2850 (n2812, n2565, n2435, n2497, n2682);
xnor g2851 (n2874, n2512, n2127, n2499, n2330);
nor  g2852 (n2966, n2652, n2266, n2701, n2551);
and  g2853 (n2917, n2382, n2111, n2164, n2380);
nand g2854 (n2766, n2727, n1929, n2010, n1911);
or   g2855 (n2864, n2018, n2665, n1877, n2468);
xor  g2856 (n2941, n2019, n2725, n2219, n2070);
nor  g2857 (n2767, n1981, n2095, n2444, n2282);
nand g2858 (n2743, n1932, n1993, n2697, n1928);
xnor g2859 (n2836, n1956, n2695, n2658, n2370);
or   g2860 (n2831, n2208, n2129, n2643, n2326);
or   g2861 (n2764, n2280, n2254, n2115, n2579);
and  g2862 (n2745, n1849, n2693, n2378, n1977);
or   g2863 (n2961, n2459, n2439, n2430, n1953);
or   g2864 (n2832, n2528, n2464, n1878, n2577);
nor  g2865 (n2950, n2397, n1922, n2100, n2594);
nand g2866 (n2807, n2082, n2306, n1968, n2172);
and  g2867 (n2923, n2348, n2135, n2321, n2481);
xor  g2868 (n2823, n2487, n2337, n2053, n2495);
nor  g2869 (n2779, n2386, n2470, n2349, n2028);
or   g2870 (n2792, n2275, n2177, n2547, n2291);
nor  g2871 (n2835, n2179, n2556, n2393, n1917);
nand g2872 (n2944, n2012, n2688, n2631, n2143);
and  g2873 (n2891, n2539, n2066, n2519, n2729);
or   g2874 (n2838, n1974, n2099, n2605, n2364);
nand g2875 (n2769, n2555, n1988, n2320, n2545);
nand g2876 (n2794, n2717, n2598, n2554, n2726);
nor  g2877 (n2911, n2335, n2188, n1957, n2618);
xnor g2878 (n2915, n2243, n2329, n1844, n1890);
xnor g2879 (n2946, n2721, n2735, n2027, n1919);
xnor g2880 (n2932, n1980, n2345, n2041, n2226);
xnor g2881 (n2905, n2002, n2260, n2106, n2521);
nand g2882 (n2858, n2103, n2006, n2080, n2581);
nand g2883 (n2752, n2269, n2256, n2307, n2015);
nor  g2884 (n2857, n2548, n1864, n2502, n1944);
or   g2885 (n2852, n2112, n1872, n1966, n1918);
and  g2886 (n2886, n2097, n2319, n2358, n2458);
nand g2887 (n2921, n2076, n2159, n1907, n2144);
or   g2888 (n2930, n1861, n2186, n2446, n2672);
and  g2889 (n2960, n2741, n2250, n2498, n2438);
and  g2890 (n2863, n2683, n2562, n2044, n1888);
nor  g2891 (n2754, n1889, n2108, n1961, n2259);
nor  g2892 (n2939, n2232, n2091, n1857, n2057);
nor  g2893 (n2959, n2587, n2490, n2350, n2641);
xor  g2894 (n2869, n2181, n2700, n2457, n2402);
or   g2895 (n2773, n2702, n1843, n2484, n2110);
and  g2896 (n2771, n1908, n1899, n1934, n2154);
xnor g2897 (n2910, n2483, n2703, n1885, n2121);
nor  g2898 (n2902, n2712, n2408, n2709, n2292);
nand g2899 (n2795, n2094, n2167, n2624, n1967);
nor  g2900 (n2872, n2303, n2300, n2443, n2450);
xnor g2901 (n2883, n2441, n2032, n1940, n2411);
nor  g2902 (n2935, n1990, n1900, n2357, n2462);
or   g2903 (n2819, n2169, n2506, n1904, n2570);
and  g2904 (n2808, n2025, n2156, n2595, n2531);
nand g2905 (n2955, n2218, n2684, n2601, n1903);
nor  g2906 (n2893, n2546, n2447, n2538, n1875);
nor  g2907 (n2897, n2609, n1997, n1891, n2060);
and  g2908 (n2895, n2059, n2145, n2670, n2109);
nand g2909 (n2846, n2719, n2720, n2530, n2195);
xnor g2910 (n2953, n2431, n2346, n1937, n2395);
or   g2911 (n2849, n2423, n2158, n2500, n2247);
xor  g2912 (n2884, n1886, n2616, n1984, n1860);
nand g2913 (n2834, n1850, n2633, n2515, n2614);
nor  g2914 (n2793, n2692, n2031, n2706, n2574);
nand g2915 (n2865, n1855, n2437, n2263, n2265);
and  g2916 (n2785, n2274, n2242, n2153, n2526);
nor  g2917 (n2787, n2309, n2381, n2191, n2486);
xor  g2918 (n2949, n2455, n2105, n1876, n2369);
xnor g2919 (n2945, n2165, n2590, n2333, n2513);
and  g2920 (n2781, n2290, n1912, n2653, n2558);
xnor g2921 (n2922, n2415, n2474, n2485, n2205);
and  g2922 (n2761, n2648, n2182, n2341, n2517);
nor  g2923 (n2940, n2215, n2220, n2273, n2650);
xnor g2924 (n2855, n2009, n1905, n1846, n2363);
nor  g2925 (n2875, n2568, n1920, n2323, n2245);
nand g2926 (n2933, n2189, n2116, n2640, n2011);
or   g2927 (n2900, n1955, n1923, n2081, n2304);
xor  g2928 (n2952, n2667, n2686, n2442, n2611);
and  g2929 (n2848, n1895, n1902, n2120, n2518);
xnor g2930 (n2758, n2086, n2071, n2710, n2600);
xnor g2931 (n2768, n2192, n2527, n1845, n2101);
xor  g2932 (n2845, n2644, n2707, n2705, n2138);
and  g2933 (n2912, n2267, n2711, n2213, n2090);
and  g2934 (n2816, n2549, n2351, n2029, n2606);
xnor g2935 (n3001, n2926, n2783, n2906, n2878);
xnor g2936 (n2987, n2854, n2956, n2841, n2951);
or   g2937 (n3003, n2916, n2831, n2860, n2792);
nand g2938 (n2972, n2902, n2830, n2789, n2829);
nand g2939 (n2974, n2781, n2923, n2832, n2953);
and  g2940 (n2977, n2877, n2957, n2779, n2936);
and  g2941 (n2993, n2839, n2768, n2798, n2778);
or   g2942 (n2991, n2895, n2822, n2924, n2771);
nand g2943 (n2976, n2797, n2824, n2919, n2856);
nand g2944 (n2985, n2809, n2804, n2944, n2932);
and  g2945 (n3010, n2875, n2950, n2811, n2800);
or   g2946 (n3007, n2894, n2796, n2935, n2888);
or   g2947 (n2978, n2846, n2937, n2799, n2867);
and  g2948 (n3006, n2886, n2784, n2772, n2823);
nand g2949 (n2995, n2967, n2853, n2871, n2929);
xor  g2950 (n3000, n2764, n2920, n2807, n2949);
nand g2951 (n2968, n2941, n2850, n2838, n2948);
nor  g2952 (n2986, n2819, n2833, n2794, n2909);
nand g2953 (n3016, n2880, n2777, n2868, n2842);
xor  g2954 (n2998, n2965, n2766, n2896, n2887);
nor  g2955 (n3019, n2814, n2911, n2770, n2802);
nor  g2956 (n2989, n2862, n2858, n2905, n2866);
and  g2957 (n2999, n2918, n2925, n2820, n2912);
and  g2958 (n3011, n2775, n2891, n2913, n2910);
xor  g2959 (n3004, n2892, n2843, n2961, n2761);
and  g2960 (n2984, n2782, n2879, n2834, n2801);
and  g2961 (n3009, n2847, n2921, n2855, n2952);
nor  g2962 (n2971, n2857, n2861, n2931, n2803);
nor  g2963 (n2981, n2908, n2940, n2845, n2884);
xnor g2964 (n3002, n2828, n2760, n2863, n2859);
or   g2965 (n2969, n2881, n2785, n2795, n2899);
nand g2966 (n2996, n2767, n2942, n2765, n2939);
or   g2967 (n2988, n2898, n2762, n2897, n2901);
xnor g2968 (n2992, n2790, n2934, n2851, n2933);
and  g2969 (n2994, n2883, n2874, n2773, n2930);
nand g2970 (n2982, n2849, n2818, n2914, n2805);
nor  g2971 (n3005, n2864, n2915, n2787, n2840);
or   g2972 (n3017, n2844, n2904, n2872, n2959);
nor  g2973 (n2973, n2869, n2963, n2870, n2808);
xnor g2974 (n2983, n2873, n2769, n2837, n2958);
and  g2975 (n3015, n2806, n2810, n2821, n2890);
nor  g2976 (n2975, n2900, n2786, n2812, n2907);
and  g2977 (n2990, n2928, n2763, n2865, n2774);
xor  g2978 (n2979, n2964, n2954, n2825, n2966);
or   g2979 (n3018, n2889, n2793, n2903, n2885);
or   g2980 (n3012, n2815, n2791, n2780, n2946);
or   g2981 (n3014, n2826, n2813, n2917, n2960);
nand g2982 (n3008, n2852, n2827, n2962, n2816);
or   g2983 (n2997, n2882, n2836, n2943, n2922);
xor  g2984 (n2980, n2927, n2848, n2938, n2817);
or   g2985 (n3013, n2893, n2835, n2788, n2955);
nand g2986 (n2970, n2947, n2876, n2776, n2945);
nand g2987 (n3031, n2980, n2989, n3019, n2996);
nand g2988 (n3024, n2997, n3006, n3016, n2978);
xnor g2989 (n3023, n3009, n2998, n3005, n2975);
nor  g2990 (n3021, n2969, n2976, n3017, n2988);
xnor g2991 (n3020, n3001, n2972, n2985, n3015);
and  g2992 (n3028, n2992, n3012, n2971, n2984);
and  g2993 (n3022, n2999, n2970, n3004, n2983);
xnor g2994 (n3027, n2987, n2977, n2973, n2994);
xor  g2995 (n3029, n2982, n2991, n3008, n3010);
xnor g2996 (n3025, n3018, n3011, n2981, n2974);
and  g2997 (n3030, n3000, n2990, n2968, n3013);
xnor g2998 (n3032, n2995, n2979, n2986, n3003);
or   g2999 (n3026, n2993, n3014, n3007, n3002);
endmodule
