

module Stat_1670_321
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n45,
  n46,
  n47,
  n48,
  n49,
  n50,
  n51,
  n52,
  n53,
  n54,
  n55,
  n56,
  n57,
  n58,
  n59,
  n1399,
  n1404,
  n1389,
  n1409,
  n1396,
  n1393,
  n1387,
  n1388,
  n1410,
  n1386,
  n1412,
  n1406,
  n1398,
  n1395,
  n1402,
  n1401,
  n1413,
  n1405,
  n1421,
  n1420,
  n1419,
  n1415,
  n1455,
  n1463,
  n1448,
  n1460,
  n1451,
  n1464,
  n1687,
  n1686,
  n1690,
  n1691,
  n1689,
  n1697,
  n1694,
  n1692,
  n1698,
  n1695,
  n1688,
  n1693,
  n1729,
  n1720,
  n1722,
  n1727,
  n1724,
  n1728,
  n1725,
  n1726,
  n1723,
  n1721
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input n40;input n41;input n42;input n43;input n44;input n45;input n46;input n47;input n48;input n49;input n50;input n51;input n52;input n53;input n54;input n55;input n56;input n57;input n58;input n59;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1399;output n1404;output n1389;output n1409;output n1396;output n1393;output n1387;output n1388;output n1410;output n1386;output n1412;output n1406;output n1398;output n1395;output n1402;output n1401;output n1413;output n1405;output n1421;output n1420;output n1419;output n1415;output n1455;output n1463;output n1448;output n1460;output n1451;output n1464;output n1687;output n1686;output n1690;output n1691;output n1689;output n1697;output n1694;output n1692;output n1698;output n1695;output n1688;output n1693;output n1729;output n1720;output n1722;output n1727;output n1724;output n1728;output n1725;output n1726;output n1723;output n1721;
  wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1390;wire n1391;wire n1392;wire n1394;wire n1397;wire n1400;wire n1403;wire n1407;wire n1408;wire n1411;wire n1414;wire n1416;wire n1417;wire n1418;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1449;wire n1450;wire n1452;wire n1453;wire n1454;wire n1456;wire n1457;wire n1458;wire n1459;wire n1461;wire n1462;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1696;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;

  buf
  g0
  (
    n95,
    n16
  );


  buf
  g1
  (
    n238,
    n40
  );


  not
  g2
  (
    n68,
    n24
  );


  buf
  g3
  (
    n65,
    n37
  );


  buf
  g4
  (
    n105,
    n6
  );


  buf
  g5
  (
    n150,
    n23
  );


  not
  g6
  (
    n97,
    n1
  );


  buf
  g7
  (
    n140,
    n5
  );


  buf
  g8
  (
    n183,
    n47
  );


  not
  g9
  (
    n133,
    n17
  );


  buf
  g10
  (
    n162,
    n32
  );


  not
  g11
  (
    n126,
    n10
  );


  buf
  g12
  (
    n146,
    n29
  );


  buf
  g13
  (
    n158,
    n19
  );


  not
  g14
  (
    n74,
    n20
  );


  not
  g15
  (
    n159,
    n35
  );


  not
  g16
  (
    n96,
    n41
  );


  buf
  g17
  (
    n231,
    n4
  );


  buf
  g18
  (
    n134,
    n27
  );


  not
  g19
  (
    n157,
    n31
  );


  not
  g20
  (
    n243,
    n34
  );


  not
  g21
  (
    n176,
    n48
  );


  buf
  g22
  (
    n115,
    n44
  );


  not
  g23
  (
    n108,
    n32
  );


  not
  g24
  (
    n237,
    n36
  );


  not
  g25
  (
    n191,
    n26
  );


  buf
  g26
  (
    n227,
    n17
  );


  not
  g27
  (
    n79,
    n25
  );


  buf
  g28
  (
    n236,
    n25
  );


  buf
  g29
  (
    n161,
    n11
  );


  not
  g30
  (
    n145,
    n10
  );


  buf
  g31
  (
    n230,
    n46
  );


  buf
  g32
  (
    n201,
    n44
  );


  buf
  g33
  (
    KeyWire_0_11,
    n40
  );


  not
  g34
  (
    KeyWire_0_19,
    n29
  );


  not
  g35
  (
    n148,
    n20
  );


  buf
  g36
  (
    n112,
    n28
  );


  buf
  g37
  (
    n91,
    n8
  );


  not
  g38
  (
    n246,
    n28
  );


  buf
  g39
  (
    n141,
    n34
  );


  not
  g40
  (
    n207,
    n19
  );


  not
  g41
  (
    n211,
    n24
  );


  buf
  g42
  (
    n216,
    n11
  );


  buf
  g43
  (
    n113,
    n18
  );


  not
  g44
  (
    n168,
    n38
  );


  not
  g45
  (
    n88,
    n31
  );


  buf
  g46
  (
    KeyWire_0_43,
    n9
  );


  buf
  g47
  (
    n117,
    n3
  );


  buf
  g48
  (
    n217,
    n37
  );


  not
  g49
  (
    n64,
    n35
  );


  buf
  g50
  (
    n110,
    n30
  );


  not
  g51
  (
    n189,
    n27
  );


  not
  g52
  (
    n125,
    n44
  );


  buf
  g53
  (
    KeyWire_0_48,
    n46
  );


  buf
  g54
  (
    n80,
    n2
  );


  buf
  g55
  (
    n239,
    n15
  );


  not
  g56
  (
    n206,
    n47
  );


  not
  g57
  (
    n225,
    n46
  );


  buf
  g58
  (
    n234,
    n29
  );


  not
  g59
  (
    KeyWire_0_16,
    n2
  );


  not
  g60
  (
    n147,
    n43
  );


  buf
  g61
  (
    n198,
    n33
  );


  buf
  g62
  (
    n61,
    n39
  );


  buf
  g63
  (
    n190,
    n1
  );


  not
  g64
  (
    n247,
    n40
  );


  buf
  g65
  (
    n196,
    n21
  );


  buf
  g66
  (
    KeyWire_0_32,
    n42
  );


  buf
  g67
  (
    n182,
    n45
  );


  buf
  g68
  (
    n193,
    n2
  );


  not
  g69
  (
    n99,
    n21
  );


  not
  g70
  (
    n185,
    n15
  );


  not
  g71
  (
    n241,
    n30
  );


  buf
  g72
  (
    n62,
    n39
  );


  not
  g73
  (
    n130,
    n7
  );


  not
  g74
  (
    n200,
    n8
  );


  buf
  g75
  (
    n155,
    n37
  );


  buf
  g76
  (
    n177,
    n42
  );


  buf
  g77
  (
    n173,
    n6
  );


  not
  g78
  (
    n233,
    n9
  );


  buf
  g79
  (
    n175,
    n12
  );


  buf
  g80
  (
    n154,
    n3
  );


  not
  g81
  (
    n204,
    n20
  );


  buf
  g82
  (
    n249,
    n30
  );


  not
  g83
  (
    n192,
    n46
  );


  buf
  g84
  (
    n214,
    n16
  );


  buf
  g85
  (
    n184,
    n45
  );


  buf
  g86
  (
    n86,
    n14
  );


  not
  g87
  (
    n208,
    n32
  );


  buf
  g88
  (
    n81,
    n2
  );


  buf
  g89
  (
    n226,
    n35
  );


  buf
  g90
  (
    n222,
    n14
  );


  buf
  g91
  (
    n122,
    n28
  );


  buf
  g92
  (
    n245,
    n47
  );


  buf
  g93
  (
    n136,
    n9
  );


  buf
  g94
  (
    n218,
    n23
  );


  not
  g95
  (
    n235,
    n41
  );


  not
  g96
  (
    n151,
    n43
  );


  buf
  g97
  (
    KeyWire_0_54,
    n47
  );


  not
  g98
  (
    n228,
    n32
  );


  buf
  g99
  (
    n197,
    n1
  );


  buf
  g100
  (
    n94,
    n10
  );


  buf
  g101
  (
    n165,
    n7
  );


  buf
  g102
  (
    n195,
    n30
  );


  not
  g103
  (
    n220,
    n12
  );


  buf
  g104
  (
    n128,
    n9
  );


  not
  g105
  (
    n84,
    n48
  );


  buf
  g106
  (
    n72,
    n41
  );


  buf
  g107
  (
    n129,
    n3
  );


  buf
  g108
  (
    n172,
    n13
  );


  buf
  g109
  (
    n209,
    n18
  );


  not
  g110
  (
    n106,
    n19
  );


  buf
  g111
  (
    n109,
    n8
  );


  not
  g112
  (
    n123,
    n27
  );


  buf
  g113
  (
    n102,
    n38
  );


  buf
  g114
  (
    KeyWire_0_9,
    n19
  );


  buf
  g115
  (
    n166,
    n42
  );


  not
  g116
  (
    n242,
    n44
  );


  buf
  g117
  (
    n85,
    n22
  );


  buf
  g118
  (
    n100,
    n36
  );


  not
  g119
  (
    n181,
    n24
  );


  buf
  g120
  (
    n127,
    n17
  );


  not
  g121
  (
    n63,
    n6
  );


  not
  g122
  (
    n250,
    n48
  );


  buf
  g123
  (
    n90,
    n33
  );


  buf
  g124
  (
    n170,
    n4
  );


  not
  g125
  (
    n121,
    n8
  );


  buf
  g126
  (
    n164,
    n5
  );


  buf
  g127
  (
    n69,
    n21
  );


  not
  g128
  (
    n76,
    n38
  );


  not
  g129
  (
    n114,
    n12
  );


  not
  g130
  (
    n248,
    n14
  );


  buf
  g131
  (
    n167,
    n21
  );


  not
  g132
  (
    n124,
    n11
  );


  not
  g133
  (
    n139,
    n43
  );


  not
  g134
  (
    n116,
    n38
  );


  not
  g135
  (
    n93,
    n40
  );


  not
  g136
  (
    n187,
    n7
  );


  not
  g137
  (
    n131,
    n29
  );


  buf
  g138
  (
    n156,
    n27
  );


  buf
  g139
  (
    n169,
    n16
  );


  buf
  g140
  (
    n149,
    n10
  );


  buf
  g141
  (
    n240,
    n26
  );


  not
  g142
  (
    n142,
    n41
  );


  buf
  g143
  (
    n98,
    n24
  );


  buf
  g144
  (
    n87,
    n14
  );


  not
  g145
  (
    n77,
    n35
  );


  buf
  g146
  (
    n163,
    n33
  );


  not
  g147
  (
    n82,
    n36
  );


  not
  g148
  (
    n103,
    n18
  );


  not
  g149
  (
    n104,
    n11
  );


  not
  g150
  (
    KeyWire_0_57,
    n42
  );


  not
  g151
  (
    n160,
    n36
  );


  buf
  g152
  (
    n171,
    n5
  );


  buf
  g153
  (
    n180,
    n4
  );


  buf
  g154
  (
    n138,
    n13
  );


  not
  g155
  (
    n143,
    n15
  );


  not
  g156
  (
    n152,
    n1
  );


  buf
  g157
  (
    n179,
    n34
  );


  buf
  g158
  (
    n219,
    n23
  );


  buf
  g159
  (
    n101,
    n26
  );


  buf
  g160
  (
    n202,
    n18
  );


  buf
  g161
  (
    n135,
    n45
  );


  buf
  g162
  (
    n132,
    n37
  );


  not
  g163
  (
    n71,
    n5
  );


  not
  g164
  (
    n174,
    n4
  );


  buf
  g165
  (
    n205,
    n45
  );


  buf
  g166
  (
    n144,
    n22
  );


  not
  g167
  (
    n229,
    n28
  );


  not
  g168
  (
    n199,
    n16
  );


  not
  g169
  (
    n153,
    n26
  );


  buf
  g170
  (
    n66,
    n7
  );


  buf
  g171
  (
    n212,
    n43
  );


  not
  g172
  (
    n210,
    n15
  );


  not
  g173
  (
    n194,
    n20
  );


  not
  g174
  (
    n186,
    n3
  );


  not
  g175
  (
    n203,
    n23
  );


  buf
  g176
  (
    n224,
    n13
  );


  buf
  g177
  (
    n107,
    n13
  );


  not
  g178
  (
    n244,
    n22
  );


  not
  g179
  (
    n111,
    n22
  );


  not
  g180
  (
    n118,
    n39
  );


  not
  g181
  (
    n178,
    n33
  );


  not
  g182
  (
    n83,
    n31
  );


  buf
  g183
  (
    n213,
    n25
  );


  buf
  g184
  (
    n137,
    n12
  );


  buf
  g185
  (
    n221,
    n6
  );


  not
  g186
  (
    n215,
    n17
  );


  not
  g187
  (
    n232,
    n25
  );


  not
  g188
  (
    n223,
    n39
  );


  buf
  g189
  (
    n73,
    n34
  );


  not
  g190
  (
    n70,
    n31
  );


  buf
  g191
  (
    n594,
    n228
  );


  not
  g192
  (
    n252,
    n115
  );


  not
  g193
  (
    n409,
    n178
  );


  buf
  g194
  (
    n602,
    n64
  );


  buf
  g195
  (
    n503,
    n182
  );


  not
  g196
  (
    n628,
    n86
  );


  not
  g197
  (
    n874,
    n200
  );


  buf
  g198
  (
    n831,
    n89
  );


  buf
  g199
  (
    n856,
    n122
  );


  buf
  g200
  (
    n528,
    n184
  );


  not
  g201
  (
    n819,
    n246
  );


  buf
  g202
  (
    n416,
    n207
  );


  buf
  g203
  (
    n852,
    n215
  );


  not
  g204
  (
    n943,
    n162
  );


  not
  g205
  (
    n458,
    n162
  );


  not
  g206
  (
    n728,
    n136
  );


  buf
  g207
  (
    n540,
    n138
  );


  not
  g208
  (
    n312,
    n155
  );


  not
  g209
  (
    n273,
    n226
  );


  not
  g210
  (
    n837,
    n216
  );


  not
  g211
  (
    n700,
    n83
  );


  buf
  g212
  (
    n502,
    n129
  );


  buf
  g213
  (
    n938,
    n159
  );


  not
  g214
  (
    n604,
    n173
  );


  buf
  g215
  (
    n414,
    n127
  );


  not
  g216
  (
    n842,
    n118
  );


  buf
  g217
  (
    n769,
    n216
  );


  buf
  g218
  (
    n906,
    n144
  );


  not
  g219
  (
    n671,
    n124
  );


  buf
  g220
  (
    n721,
    n184
  );


  not
  g221
  (
    n459,
    n63
  );


  not
  g222
  (
    n849,
    n175
  );


  buf
  g223
  (
    n821,
    n247
  );


  buf
  g224
  (
    n761,
    n215
  );


  not
  g225
  (
    n888,
    n94
  );


  not
  g226
  (
    n467,
    n147
  );


  not
  g227
  (
    n687,
    n117
  );


  buf
  g228
  (
    n488,
    n122
  );


  not
  g229
  (
    n832,
    n151
  );


  not
  g230
  (
    n393,
    n198
  );


  buf
  g231
  (
    n506,
    n200
  );


  not
  g232
  (
    n263,
    n204
  );


  not
  g233
  (
    n715,
    n220
  );


  buf
  g234
  (
    n392,
    n65
  );


  not
  g235
  (
    n863,
    n80
  );


  buf
  g236
  (
    n569,
    n139
  );


  not
  g237
  (
    n316,
    n60
  );


  buf
  g238
  (
    n447,
    n199
  );


  not
  g239
  (
    n265,
    n173
  );


  not
  g240
  (
    n878,
    n144
  );


  buf
  g241
  (
    n281,
    n148
  );


  not
  g242
  (
    n702,
    n228
  );


  buf
  g243
  (
    n696,
    n76
  );


  buf
  g244
  (
    n944,
    n174
  );


  not
  g245
  (
    n693,
    n132
  );


  not
  g246
  (
    n601,
    n189
  );


  not
  g247
  (
    n428,
    n202
  );


  not
  g248
  (
    n526,
    n122
  );


  buf
  g249
  (
    n306,
    n217
  );


  not
  g250
  (
    n855,
    n146
  );


  not
  g251
  (
    n551,
    n81
  );


  not
  g252
  (
    n897,
    n119
  );


  not
  g253
  (
    n286,
    n249
  );


  buf
  g254
  (
    n909,
    n70
  );


  buf
  g255
  (
    n725,
    n95
  );


  not
  g256
  (
    n554,
    n69
  );


  buf
  g257
  (
    n560,
    n113
  );


  not
  g258
  (
    n453,
    n221
  );


  buf
  g259
  (
    n775,
    n142
  );


  not
  g260
  (
    n864,
    n174
  );


  not
  g261
  (
    n866,
    n79
  );


  not
  g262
  (
    n319,
    n67
  );


  buf
  g263
  (
    n507,
    n180
  );


  not
  g264
  (
    n672,
    n236
  );


  not
  g265
  (
    n344,
    n204
  );


  buf
  g266
  (
    KeyWire_0_1,
    n72
  );


  not
  g267
  (
    n361,
    n176
  );


  not
  g268
  (
    n950,
    n116
  );


  not
  g269
  (
    n352,
    n131
  );


  buf
  g270
  (
    n271,
    n148
  );


  not
  g271
  (
    n420,
    n178
  );


  not
  g272
  (
    n916,
    n128
  );


  buf
  g273
  (
    n620,
    n155
  );


  not
  g274
  (
    n653,
    n129
  );


  not
  g275
  (
    KeyWire_0_42,
    n145
  );


  not
  g276
  (
    n773,
    n203
  );


  not
  g277
  (
    n270,
    n227
  );


  buf
  g278
  (
    n913,
    n166
  );


  buf
  g279
  (
    n487,
    n241
  );


  buf
  g280
  (
    n741,
    n145
  );


  buf
  g281
  (
    n353,
    n146
  );


  not
  g282
  (
    n946,
    n96
  );


  buf
  g283
  (
    n455,
    n180
  );


  buf
  g284
  (
    n814,
    n236
  );


  not
  g285
  (
    n749,
    n187
  );


  buf
  g286
  (
    n905,
    n153
  );


  buf
  g287
  (
    n766,
    n179
  );


  buf
  g288
  (
    n522,
    n143
  );


  not
  g289
  (
    n266,
    n192
  );


  not
  g290
  (
    n678,
    n248
  );


  not
  g291
  (
    n808,
    n223
  );


  not
  g292
  (
    n435,
    n190
  );


  not
  g293
  (
    n391,
    n98
  );


  not
  g294
  (
    n436,
    n225
  );


  not
  g295
  (
    KeyWire_0_4,
    n101
  );


  buf
  g296
  (
    n389,
    n238
  );


  buf
  g297
  (
    n763,
    n196
  );


  not
  g298
  (
    n685,
    n163
  );


  buf
  g299
  (
    KeyWire_0_62,
    n216
  );


  not
  g300
  (
    n876,
    n98
  );


  buf
  g301
  (
    n631,
    n201
  );


  not
  g302
  (
    n291,
    n70
  );


  buf
  g303
  (
    n709,
    n112
  );


  buf
  g304
  (
    n807,
    n152
  );


  not
  g305
  (
    n304,
    n154
  );


  not
  g306
  (
    n401,
    n182
  );


  buf
  g307
  (
    n844,
    n206
  );


  not
  g308
  (
    n327,
    n106
  );


  buf
  g309
  (
    n408,
    n59
  );


  buf
  g310
  (
    n272,
    n162
  );


  buf
  g311
  (
    n918,
    n98
  );


  buf
  g312
  (
    n673,
    n101
  );


  not
  g313
  (
    n630,
    n142
  );


  not
  g314
  (
    n744,
    n198
  );


  buf
  g315
  (
    n865,
    n183
  );


  not
  g316
  (
    n752,
    n240
  );


  buf
  g317
  (
    n830,
    n118
  );


  not
  g318
  (
    n886,
    n229
  );


  not
  g319
  (
    n377,
    n163
  );


  not
  g320
  (
    KeyWire_0_28,
    n157
  );


  buf
  g321
  (
    n434,
    n165
  );


  not
  g322
  (
    n629,
    n220
  );


  buf
  g323
  (
    n278,
    n164
  );


  buf
  g324
  (
    n606,
    n215
  );


  buf
  g325
  (
    KeyWire_0_3,
    n58
  );


  buf
  g326
  (
    n268,
    n88
  );


  not
  g327
  (
    n952,
    n111
  );


  not
  g328
  (
    n829,
    n143
  );


  buf
  g329
  (
    n903,
    n73
  );


  buf
  g330
  (
    n937,
    n165
  );


  buf
  g331
  (
    n565,
    n109
  );


  not
  g332
  (
    n921,
    n186
  );


  buf
  g333
  (
    n663,
    n172
  );


  buf
  g334
  (
    n386,
    n107
  );


  buf
  g335
  (
    n746,
    n125
  );


  not
  g336
  (
    n394,
    n240
  );


  buf
  g337
  (
    n654,
    n127
  );


  buf
  g338
  (
    n465,
    n154
  );


  not
  g339
  (
    n890,
    n142
  );


  buf
  g340
  (
    n380,
    n112
  );


  buf
  g341
  (
    n647,
    n143
  );


  buf
  g342
  (
    n798,
    n205
  );


  buf
  g343
  (
    n529,
    n171
  );


  buf
  g344
  (
    n315,
    n190
  );


  not
  g345
  (
    n412,
    n144
  );


  buf
  g346
  (
    n833,
    n130
  );


  buf
  g347
  (
    n759,
    n201
  );


  buf
  g348
  (
    KeyWire_0_30,
    n147
  );


  buf
  g349
  (
    n823,
    n128
  );


  buf
  g350
  (
    n485,
    n187
  );


  not
  g351
  (
    n931,
    n138
  );


  not
  g352
  (
    n584,
    n67
  );


  buf
  g353
  (
    n469,
    n183
  );


  not
  g354
  (
    n718,
    n107
  );


  buf
  g355
  (
    n332,
    n209
  );


  buf
  g356
  (
    n768,
    n95
  );


  not
  g357
  (
    n556,
    n81
  );


  buf
  g358
  (
    n638,
    n192
  );


  not
  g359
  (
    n813,
    n141
  );


  not
  g360
  (
    n433,
    n173
  );


  buf
  g361
  (
    n688,
    n243
  );


  buf
  g362
  (
    n517,
    n141
  );


  buf
  g363
  (
    n816,
    n212
  );


  buf
  g364
  (
    n357,
    n90
  );


  buf
  g365
  (
    n484,
    n233
  );


  buf
  g366
  (
    n719,
    n181
  );


  buf
  g367
  (
    n939,
    n75
  );


  not
  g368
  (
    n738,
    n49
  );


  not
  g369
  (
    n340,
    n134
  );


  buf
  g370
  (
    n843,
    n115
  );


  not
  g371
  (
    n841,
    n91
  );


  buf
  g372
  (
    n658,
    n193
  );


  not
  g373
  (
    n577,
    n113
  );


  buf
  g374
  (
    n379,
    n170
  );


  buf
  g375
  (
    n796,
    n247
  );


  buf
  g376
  (
    n904,
    n134
  );


  buf
  g377
  (
    n660,
    n97
  );


  not
  g378
  (
    n583,
    n117
  );


  not
  g379
  (
    n720,
    n208
  );


  not
  g380
  (
    n568,
    n123
  );


  not
  g381
  (
    n486,
    n117
  );


  buf
  g382
  (
    n600,
    n82
  );


  buf
  g383
  (
    n321,
    n71
  );


  not
  g384
  (
    n729,
    n99
  );


  buf
  g385
  (
    n809,
    n89
  );


  not
  g386
  (
    n282,
    n232
  );


  buf
  g387
  (
    n885,
    n237
  );


  buf
  g388
  (
    n614,
    n206
  );


  not
  g389
  (
    n413,
    n177
  );


  not
  g390
  (
    n680,
    n211
  );


  not
  g391
  (
    n839,
    n66
  );


  buf
  g392
  (
    n346,
    n75
  );


  not
  g393
  (
    n457,
    n241
  );


  buf
  g394
  (
    n451,
    n160
  );


  buf
  g395
  (
    n564,
    n197
  );


  not
  g396
  (
    n562,
    n89
  );


  buf
  g397
  (
    n732,
    n73
  );


  buf
  g398
  (
    n771,
    n67
  );


  buf
  g399
  (
    n812,
    n250
  );


  buf
  g400
  (
    n802,
    n100
  );


  not
  g401
  (
    n264,
    n210
  );


  buf
  g402
  (
    n284,
    n209
  );


  buf
  g403
  (
    n355,
    n51
  );


  buf
  g404
  (
    n861,
    n103
  );


  buf
  g405
  (
    n645,
    n191
  );


  not
  g406
  (
    KeyWire_0_49,
    n140
  );


  not
  g407
  (
    n786,
    n219
  );


  buf
  g408
  (
    KeyWire_0_26,
    n120
  );


  not
  g409
  (
    n847,
    n224
  );


  not
  g410
  (
    n704,
    n140
  );


  not
  g411
  (
    n835,
    n227
  );


  not
  g412
  (
    n884,
    n146
  );


  not
  g413
  (
    n280,
    n90
  );


  not
  g414
  (
    n499,
    n126
  );


  not
  g415
  (
    n877,
    n89
  );


  not
  g416
  (
    n500,
    n207
  );


  buf
  g417
  (
    n634,
    n133
  );


  not
  g418
  (
    n307,
    n128
  );


  not
  g419
  (
    n850,
    n105
  );


  buf
  g420
  (
    n607,
    n202
  );


  buf
  g421
  (
    n427,
    n56
  );


  not
  g422
  (
    n575,
    n220
  );


  buf
  g423
  (
    n561,
    n133
  );


  buf
  g424
  (
    n454,
    n115
  );


  buf
  g425
  (
    n623,
    n118
  );


  not
  g426
  (
    n374,
    n73
  );


  buf
  g427
  (
    n716,
    n175
  );


  buf
  g428
  (
    n533,
    n91
  );


  buf
  g429
  (
    n549,
    n209
  );


  buf
  g430
  (
    n682,
    n152
  );


  not
  g431
  (
    n633,
    n51
  );


  not
  g432
  (
    n818,
    n218
  );


  not
  g433
  (
    n776,
    n49
  );


  not
  g434
  (
    n883,
    n212
  );


  buf
  g435
  (
    n547,
    n218
  );


  not
  g436
  (
    n603,
    n156
  );


  buf
  g437
  (
    n448,
    n79
  );


  buf
  g438
  (
    n846,
    n236
  );


  not
  g439
  (
    n748,
    n246
  );


  buf
  g440
  (
    n932,
    n231
  );


  not
  g441
  (
    n872,
    n161
  );


  not
  g442
  (
    n400,
    n107
  );


  not
  g443
  (
    n713,
    n185
  );


  not
  g444
  (
    n490,
    n203
  );


  buf
  g445
  (
    n388,
    n211
  );


  not
  g446
  (
    n461,
    n223
  );


  not
  g447
  (
    n417,
    n78
  );


  buf
  g448
  (
    n815,
    n185
  );


  buf
  g449
  (
    n643,
    n246
  );


  not
  g450
  (
    n300,
    n151
  );


  not
  g451
  (
    n871,
    n63
  );


  not
  g452
  (
    n418,
    n92
  );


  not
  g453
  (
    n853,
    n86
  );


  not
  g454
  (
    n423,
    n82
  );


  not
  g455
  (
    n530,
    n104
  );


  not
  g456
  (
    n919,
    n81
  );


  not
  g457
  (
    n305,
    n53
  );


  not
  g458
  (
    n641,
    n55
  );


  not
  g459
  (
    n825,
    n62
  );


  not
  g460
  (
    n664,
    n149
  );


  not
  g461
  (
    n322,
    n69
  );


  not
  g462
  (
    n364,
    n121
  );


  buf
  g463
  (
    n898,
    n121
  );


  not
  g464
  (
    n758,
    n120
  );


  not
  g465
  (
    n302,
    n105
  );


  not
  g466
  (
    n296,
    n217
  );


  not
  g467
  (
    n899,
    n155
  );


  not
  g468
  (
    n681,
    n123
  );


  not
  g469
  (
    n902,
    n110
  );


  not
  g470
  (
    n621,
    n118
  );


  not
  g471
  (
    n525,
    n60
  );


  buf
  g472
  (
    n376,
    n55
  );


  not
  g473
  (
    n303,
    n249
  );


  not
  g474
  (
    n475,
    n50
  );


  not
  g475
  (
    n735,
    n153
  );


  not
  g476
  (
    n430,
    n150
  );


  buf
  g477
  (
    n552,
    n175
  );


  not
  g478
  (
    n705,
    n109
  );


  not
  g479
  (
    n314,
    n51
  );


  buf
  g480
  (
    n924,
    n92
  );


  not
  g481
  (
    n385,
    n79
  );


  not
  g482
  (
    n698,
    n86
  );


  not
  g483
  (
    n879,
    n88
  );


  not
  g484
  (
    n820,
    n239
  );


  buf
  g485
  (
    n949,
    n178
  );


  not
  g486
  (
    n449,
    n53
  );


  buf
  g487
  (
    n891,
    n190
  );


  not
  g488
  (
    n287,
    n241
  );


  not
  g489
  (
    n318,
    n154
  );


  not
  g490
  (
    n369,
    n126
  );


  not
  g491
  (
    KeyWire_0_36,
    n104
  );


  not
  g492
  (
    n537,
    n139
  );


  not
  g493
  (
    n471,
    n174
  );


  buf
  g494
  (
    n787,
    n156
  );


  buf
  g495
  (
    n293,
    n58
  );


  buf
  g496
  (
    n857,
    n99
  );


  not
  g497
  (
    n799,
    n119
  );


  buf
  g498
  (
    n396,
    n157
  );


  buf
  g499
  (
    n745,
    n82
  );


  not
  g500
  (
    n512,
    n189
  );


  buf
  g501
  (
    n767,
    n209
  );


  not
  g502
  (
    n928,
    n123
  );


  not
  g503
  (
    n593,
    n83
  );


  not
  g504
  (
    n498,
    n222
  );


  buf
  g505
  (
    n740,
    n80
  );


  not
  g506
  (
    n324,
    n171
  );


  not
  g507
  (
    n652,
    n111
  );


  not
  g508
  (
    n708,
    n132
  );


  not
  g509
  (
    n407,
    n148
  );


  buf
  g510
  (
    n636,
    n232
  );


  not
  g511
  (
    n801,
    n62
  );


  buf
  g512
  (
    n858,
    n165
  );


  buf
  g513
  (
    n848,
    n244
  );


  not
  g514
  (
    KeyWire_0_17,
    n167
  );


  buf
  g515
  (
    n800,
    n85
  );


  buf
  g516
  (
    KeyWire_0_41,
    n90
  );


  not
  g517
  (
    n262,
    n138
  );


  buf
  g518
  (
    n954,
    n243
  );


  buf
  g519
  (
    n609,
    n217
  );


  not
  g520
  (
    n881,
    n53
  );


  buf
  g521
  (
    n942,
    n235
  );


  not
  g522
  (
    n689,
    n171
  );


  buf
  g523
  (
    n387,
    n186
  );


  not
  g524
  (
    n497,
    n236
  );


  not
  g525
  (
    n515,
    n239
  );


  buf
  g526
  (
    n941,
    n177
  );


  not
  g527
  (
    n650,
    n157
  );


  buf
  g528
  (
    n365,
    n116
  );


  buf
  g529
  (
    n882,
    n158
  );


  buf
  g530
  (
    n780,
    n87
  );


  not
  g531
  (
    KeyWire_0_40,
    n176
  );


  not
  g532
  (
    n625,
    n163
  );


  buf
  g533
  (
    n723,
    n194
  );


  not
  g534
  (
    n253,
    n129
  );


  buf
  g535
  (
    n701,
    n194
  );


  buf
  g536
  (
    n462,
    n55
  );


  not
  g537
  (
    n274,
    n94
  );


  not
  g538
  (
    n743,
    n78
  );


  not
  g539
  (
    n350,
    n230
  );


  not
  g540
  (
    n466,
    n105
  );


  buf
  g541
  (
    n495,
    n222
  );


  buf
  g542
  (
    n695,
    n161
  );


  buf
  g543
  (
    n790,
    n206
  );


  buf
  g544
  (
    n589,
    n238
  );


  not
  g545
  (
    KeyWire_0_39,
    n54
  );


  buf
  g546
  (
    n411,
    n181
  );


  buf
  g547
  (
    n956,
    n225
  );


  not
  g548
  (
    n578,
    n249
  );


  not
  g549
  (
    n784,
    n185
  );


  buf
  g550
  (
    n256,
    n188
  );


  not
  g551
  (
    n862,
    n165
  );


  not
  g552
  (
    n599,
    n84
  );


  buf
  g553
  (
    n331,
    n164
  );


  not
  g554
  (
    n452,
    n96
  );


  not
  g555
  (
    n267,
    n213
  );


  not
  g556
  (
    n781,
    n224
  );


  not
  g557
  (
    n867,
    n126
  );


  buf
  g558
  (
    n940,
    n110
  );


  not
  g559
  (
    n510,
    n250
  );


  not
  g560
  (
    n622,
    n82
  );


  not
  g561
  (
    n782,
    n231
  );


  not
  g562
  (
    n269,
    n124
  );


  not
  g563
  (
    n777,
    n108
  );


  buf
  g564
  (
    n677,
    n126
  );


  not
  g565
  (
    n734,
    n147
  );


  buf
  g566
  (
    n580,
    n213
  );


  buf
  g567
  (
    n509,
    n110
  );


  buf
  g568
  (
    n757,
    n131
  );


  not
  g569
  (
    n429,
    n227
  );


  buf
  g570
  (
    n785,
    n235
  );


  not
  g571
  (
    n432,
    n184
  );


  buf
  g572
  (
    n581,
    n125
  );


  buf
  g573
  (
    n887,
    n55
  );


  not
  g574
  (
    n405,
    n186
  );


  not
  g575
  (
    n328,
    n167
  );


  not
  g576
  (
    n923,
    n150
  );


  not
  g577
  (
    n557,
    n54
  );


  buf
  g578
  (
    n826,
    n78
  );


  not
  g579
  (
    n840,
    n127
  );


  not
  g580
  (
    n667,
    n215
  );


  buf
  g581
  (
    n597,
    n94
  );


  buf
  g582
  (
    n733,
    n235
  );


  buf
  g583
  (
    n662,
    n57
  );


  not
  g584
  (
    n440,
    n221
  );


  buf
  g585
  (
    n424,
    n157
  );


  not
  g586
  (
    n679,
    n61
  );


  not
  g587
  (
    n559,
    n201
  );


  not
  g588
  (
    n463,
    n212
  );


  not
  g589
  (
    n824,
    n247
  );


  buf
  g590
  (
    n421,
    n186
  );


  not
  g591
  (
    n290,
    n76
  );


  not
  g592
  (
    n922,
    n50
  );


  not
  g593
  (
    n615,
    n91
  );


  buf
  g594
  (
    n501,
    n155
  );


  not
  g595
  (
    n550,
    n116
  );


  not
  g596
  (
    n348,
    n153
  );


  buf
  g597
  (
    n325,
    n64
  );


  buf
  g598
  (
    n838,
    n63
  );


  buf
  g599
  (
    n669,
    n172
  );


  not
  g600
  (
    n257,
    n147
  );


  not
  g601
  (
    n338,
    n152
  );


  buf
  g602
  (
    n496,
    n56
  );


  buf
  g603
  (
    KeyWire_0_53,
    n133
  );


  not
  g604
  (
    n691,
    n210
  );


  not
  g605
  (
    n783,
    n144
  );


  buf
  g606
  (
    n367,
    n137
  );


  not
  g607
  (
    n665,
    n242
  );


  buf
  g608
  (
    n920,
    n49
  );


  buf
  g609
  (
    n446,
    n192
  );


  buf
  g610
  (
    n566,
    n93
  );


  buf
  g611
  (
    n613,
    n130
  );


  not
  g612
  (
    n298,
    n192
  );


  not
  g613
  (
    n901,
    n97
  );


  not
  g614
  (
    n406,
    n166
  );


  not
  g615
  (
    n817,
    n187
  );


  buf
  g616
  (
    n894,
    n60
  );


  not
  g617
  (
    n299,
    n171
  );


  buf
  g618
  (
    n859,
    n231
  );


  not
  g619
  (
    n684,
    n242
  );


  buf
  g620
  (
    n404,
    n235
  );


  buf
  g621
  (
    n774,
    n61
  );


  not
  g622
  (
    n955,
    n96
  );


  not
  g623
  (
    n828,
    n179
  );


  not
  g624
  (
    n292,
    n64
  );


  buf
  g625
  (
    n611,
    n177
  );


  not
  g626
  (
    n753,
    n83
  );


  buf
  g627
  (
    n450,
    n197
  );


  buf
  g628
  (
    KeyWire_0_60,
    n63
  );


  not
  g629
  (
    n572,
    n92
  );


  not
  g630
  (
    n772,
    n97
  );


  not
  g631
  (
    n311,
    n232
  );


  buf
  g632
  (
    n373,
    n191
  );


  buf
  g633
  (
    n548,
    n100
  );


  not
  g634
  (
    n754,
    n216
  );


  not
  g635
  (
    n489,
    n149
  );


  buf
  g636
  (
    n410,
    n66
  );


  buf
  g637
  (
    n854,
    n158
  );


  buf
  g638
  (
    n362,
    n59
  );


  not
  g639
  (
    n339,
    n232
  );


  not
  g640
  (
    n345,
    n67
  );


  not
  g641
  (
    n553,
    n161
  );


  not
  g642
  (
    n624,
    n129
  );


  not
  g643
  (
    n366,
    n205
  );


  buf
  g644
  (
    n351,
    n93
  );


  buf
  g645
  (
    n492,
    n156
  );


  not
  g646
  (
    n582,
    n188
  );


  not
  g647
  (
    n779,
    n214
  );


  buf
  g648
  (
    n531,
    n234
  );


  not
  g649
  (
    n301,
    n204
  );


  buf
  g650
  (
    n792,
    n69
  );


  not
  g651
  (
    n592,
    n200
  );


  not
  g652
  (
    KeyWire_0_23,
    n211
  );


  not
  g653
  (
    n523,
    n88
  );


  buf
  g654
  (
    n326,
    n208
  );


  buf
  g655
  (
    n917,
    n248
  );


  buf
  g656
  (
    n644,
    n85
  );


  not
  g657
  (
    n930,
    n58
  );


  not
  g658
  (
    n686,
    n226
  );


  buf
  g659
  (
    n683,
    n172
  );


  buf
  g660
  (
    n822,
    n64
  );


  buf
  g661
  (
    n726,
    n49
  );


  not
  g662
  (
    n608,
    n120
  );


  buf
  g663
  (
    n539,
    n80
  );


  not
  g664
  (
    n532,
    n54
  );


  buf
  g665
  (
    n690,
    n62
  );


  buf
  g666
  (
    n659,
    n60
  );


  not
  g667
  (
    n827,
    n75
  );


  not
  g668
  (
    n508,
    n242
  );


  not
  g669
  (
    n474,
    n170
  );


  not
  g670
  (
    n288,
    n206
  );


  not
  g671
  (
    n347,
    n62
  );


  buf
  g672
  (
    n699,
    n136
  );


  buf
  g673
  (
    n524,
    n140
  );


  not
  g674
  (
    n933,
    n106
  );


  not
  g675
  (
    n586,
    n196
  );


  not
  g676
  (
    KeyWire_0_56,
    n104
  );


  not
  g677
  (
    n415,
    n57
  );


  buf
  g678
  (
    n869,
    n229
  );


  buf
  g679
  (
    n310,
    n222
  );


  buf
  g680
  (
    n851,
    n200
  );


  not
  g681
  (
    n889,
    n114
  );


  buf
  g682
  (
    n341,
    n221
  );


  buf
  g683
  (
    KeyWire_0_38,
    n48
  );


  buf
  g684
  (
    n648,
    n210
  );


  not
  g685
  (
    n543,
    n168
  );


  not
  g686
  (
    n910,
    n183
  );


  buf
  g687
  (
    n398,
    n168
  );


  buf
  g688
  (
    n646,
    n112
  );


  not
  g689
  (
    n520,
    n100
  );


  not
  g690
  (
    n674,
    n102
  );


  not
  g691
  (
    n632,
    n180
  );


  not
  g692
  (
    n627,
    n202
  );


  buf
  g693
  (
    n491,
    n71
  );


  buf
  g694
  (
    KeyWire_0_63,
    n88
  );


  buf
  g695
  (
    n494,
    n160
  );


  buf
  g696
  (
    n395,
    n114
  );


  not
  g697
  (
    n742,
    n226
  );


  not
  g698
  (
    n383,
    n234
  );


  buf
  g699
  (
    n595,
    n98
  );


  not
  g700
  (
    n258,
    n194
  );


  buf
  g701
  (
    n555,
    n103
  );


  buf
  g702
  (
    n516,
    n237
  );


  not
  g703
  (
    n399,
    n114
  );


  buf
  g704
  (
    n576,
    n68
  );


  buf
  g705
  (
    n254,
    n172
  );


  buf
  g706
  (
    n541,
    n121
  );


  buf
  g707
  (
    n482,
    n93
  );


  buf
  g708
  (
    n707,
    n218
  );


  buf
  g709
  (
    n538,
    n95
  );


  not
  g710
  (
    n596,
    n194
  );


  buf
  g711
  (
    KeyWire_0_50,
    n148
  );


  buf
  g712
  (
    n505,
    n159
  );


  buf
  g713
  (
    n478,
    n244
  );


  buf
  g714
  (
    n651,
    n58
  );


  not
  g715
  (
    n285,
    n90
  );


  not
  g716
  (
    KeyWire_0_15,
    n177
  );


  not
  g717
  (
    n895,
    n73
  );


  not
  g718
  (
    n639,
    n170
  );


  buf
  g719
  (
    n333,
    n207
  );


  not
  g720
  (
    n927,
    n199
  );


  not
  g721
  (
    n731,
    n78
  );


  buf
  g722
  (
    n860,
    n214
  );


  buf
  g723
  (
    n911,
    n160
  );


  not
  g724
  (
    n567,
    n208
  );


  buf
  g725
  (
    n793,
    n108
  );


  not
  g726
  (
    n751,
    n245
  );


  buf
  g727
  (
    n579,
    n191
  );


  not
  g728
  (
    n706,
    n77
  );


  buf
  g729
  (
    n703,
    n195
  );


  not
  g730
  (
    n384,
    n214
  );


  buf
  g731
  (
    n438,
    n210
  );


  buf
  g732
  (
    n546,
    n85
  );


  not
  g733
  (
    n612,
    n159
  );


  not
  g734
  (
    n958,
    n230
  );


  buf
  g735
  (
    n598,
    n135
  );


  buf
  g736
  (
    n764,
    n226
  );


  not
  g737
  (
    n873,
    n135
  );


  buf
  g738
  (
    n585,
    n149
  );


  not
  g739
  (
    n363,
    n191
  );


  buf
  g740
  (
    n390,
    n146
  );


  not
  g741
  (
    n655,
    n154
  );


  buf
  g742
  (
    n349,
    n240
  );


  buf
  g743
  (
    n381,
    n86
  );


  not
  g744
  (
    n275,
    n130
  );


  not
  g745
  (
    n358,
    n225
  );


  not
  g746
  (
    n953,
    n113
  );


  buf
  g747
  (
    n590,
    n102
  );


  not
  g748
  (
    n750,
    n128
  );


  not
  g749
  (
    n893,
    n229
  );


  buf
  g750
  (
    n694,
    n77
  );


  buf
  g751
  (
    n619,
    n218
  );


  buf
  g752
  (
    n479,
    n65
  );


  not
  g753
  (
    n276,
    n228
  );


  buf
  g754
  (
    n914,
    n57
  );


  buf
  g755
  (
    n359,
    n193
  );


  buf
  g756
  (
    n260,
    n114
  );


  not
  g757
  (
    n868,
    n87
  );


  buf
  g758
  (
    n736,
    n132
  );


  not
  g759
  (
    n402,
    n166
  );


  buf
  g760
  (
    n762,
    n61
  );


  buf
  g761
  (
    n445,
    n198
  );


  not
  g762
  (
    n343,
    n150
  );


  not
  g763
  (
    n334,
    n103
  );


  not
  g764
  (
    n472,
    n166
  );


  buf
  g765
  (
    n804,
    n124
  );


  not
  g766
  (
    n710,
    n139
  );


  buf
  g767
  (
    n765,
    n162
  );


  not
  g768
  (
    n342,
    n237
  );


  not
  g769
  (
    n329,
    n245
  );


  not
  g770
  (
    n473,
    n119
  );


  buf
  g771
  (
    n915,
    n71
  );


  not
  g772
  (
    n929,
    n109
  );


  buf
  g773
  (
    n570,
    n213
  );


  not
  g774
  (
    n797,
    n181
  );


  not
  g775
  (
    n661,
    n132
  );


  not
  g776
  (
    n717,
    n122
  );


  not
  g777
  (
    n336,
    n183
  );


  buf
  g778
  (
    n375,
    n52
  );


  buf
  g779
  (
    n431,
    n195
  );


  buf
  g780
  (
    n957,
    n189
  );


  buf
  g781
  (
    n419,
    n202
  );


  buf
  g782
  (
    n514,
    n65
  );


  buf
  g783
  (
    n563,
    n93
  );


  not
  g784
  (
    n947,
    n184
  );


  not
  g785
  (
    n900,
    n110
  );


  not
  g786
  (
    n656,
    n50
  );


  buf
  g787
  (
    n692,
    n61
  );


  not
  g788
  (
    n483,
    n117
  );


  buf
  g789
  (
    n760,
    n74
  );


  not
  g790
  (
    n527,
    n57
  );


  buf
  g791
  (
    n712,
    n85
  );


  buf
  g792
  (
    n545,
    n116
  );


  buf
  g793
  (
    n536,
    n74
  );


  buf
  g794
  (
    n437,
    n238
  );


  buf
  g795
  (
    n397,
    n169
  );


  not
  g796
  (
    n588,
    n131
  );


  not
  g797
  (
    n378,
    n105
  );


  not
  g798
  (
    n521,
    n125
  );


  buf
  g799
  (
    n255,
    n103
  );


  buf
  g800
  (
    n335,
    n87
  );


  not
  g801
  (
    n739,
    n52
  );


  not
  g802
  (
    n788,
    n199
  );


  not
  g803
  (
    n468,
    n77
  );


  buf
  g804
  (
    n323,
    n54
  );


  not
  g805
  (
    n605,
    n59
  );


  not
  g806
  (
    n542,
    n180
  );


  not
  g807
  (
    n313,
    n167
  );


  buf
  g808
  (
    n297,
    n234
  );


  not
  g809
  (
    KeyWire_0_18,
    n59
  );


  not
  g810
  (
    n666,
    n168
  );


  not
  g811
  (
    n422,
    n113
  );


  not
  g812
  (
    n317,
    n136
  );


  buf
  g813
  (
    n443,
    n97
  );


  not
  g814
  (
    n936,
    n225
  );


  not
  g815
  (
    n806,
    n160
  );


  not
  g816
  (
    n756,
    n87
  );


  not
  g817
  (
    n535,
    n56
  );


  buf
  g818
  (
    n945,
    n239
  );


  buf
  g819
  (
    n657,
    n50
  );


  buf
  g820
  (
    n778,
    n196
  );


  not
  g821
  (
    n794,
    n249
  );


  buf
  g822
  (
    n513,
    n137
  );


  not
  g823
  (
    n320,
    n115
  );


  buf
  g824
  (
    n934,
    n240
  );


  buf
  g825
  (
    n810,
    n106
  );


  buf
  g826
  (
    n360,
    n108
  );


  buf
  g827
  (
    n714,
    n169
  );


  not
  g828
  (
    n737,
    n133
  );


  not
  g829
  (
    n571,
    n167
  );


  not
  g830
  (
    n724,
    n72
  );


  buf
  g831
  (
    n261,
    n68
  );


  buf
  g832
  (
    n309,
    n185
  );


  not
  g833
  (
    n481,
    n74
  );


  not
  g834
  (
    n403,
    n120
  );


  buf
  g835
  (
    n697,
    n124
  );


  not
  g836
  (
    n948,
    n234
  );


  not
  g837
  (
    n730,
    n241
  );


  buf
  g838
  (
    KeyWire_0_44,
    n245
  );


  not
  g839
  (
    n591,
    n72
  );


  buf
  g840
  (
    n834,
    n79
  );


  buf
  g841
  (
    n511,
    n211
  );


  not
  g842
  (
    n892,
    n213
  );


  buf
  g843
  (
    n573,
    n219
  );


  buf
  g844
  (
    n805,
    n108
  );


  not
  g845
  (
    n371,
    n219
  );


  not
  g846
  (
    n444,
    n99
  );


  not
  g847
  (
    n670,
    n224
  );


  buf
  g848
  (
    n789,
    n139
  );


  not
  g849
  (
    n558,
    n214
  );


  not
  g850
  (
    n295,
    n243
  );


  not
  g851
  (
    n791,
    n203
  );


  buf
  g852
  (
    n896,
    n178
  );


  buf
  g853
  (
    n382,
    n228
  );


  buf
  g854
  (
    n456,
    n69
  );


  not
  g855
  (
    n441,
    n143
  );


  buf
  g856
  (
    n279,
    n207
  );


  buf
  g857
  (
    n464,
    n136
  );


  not
  g858
  (
    n845,
    n159
  );


  buf
  g859
  (
    n626,
    n107
  );


  not
  g860
  (
    n642,
    n68
  );


  not
  g861
  (
    KeyWire_0_31,
    n197
  );


  buf
  g862
  (
    n587,
    n169
  );


  not
  g863
  (
    n668,
    n187
  );


  buf
  g864
  (
    n493,
    n138
  );


  not
  g865
  (
    n337,
    n193
  );


  buf
  g866
  (
    n283,
    n135
  );


  xnor
  g867
  (
    n649,
    n101,
    n75,
    n121,
    n188
  );


  and
  g868
  (
    n534,
    n109,
    n244,
    n212
  );


  nor
  g869
  (
    n439,
    n152,
    n201,
    n164,
    n242
  );


  xor
  g870
  (
    n574,
    n175,
    n151,
    n222,
    n176
  );


  or
  g871
  (
    n676,
    n248,
    n112,
    n84,
    n205
  );


  nor
  g872
  (
    n356,
    n205,
    n70,
    n243,
    n174
  );


  xnor
  g873
  (
    n251,
    n158,
    n193,
    n96,
    n217
  );


  nor
  g874
  (
    n544,
    n91,
    n208,
    n145,
    n51
  );


  and
  g875
  (
    n426,
    n84,
    n248,
    n95,
    n123
  );


  xnor
  g876
  (
    KeyWire_0_55,
    n189,
    n142,
    n233,
    n52
  );


  nor
  g877
  (
    n368,
    n145,
    n221,
    n179,
    n163
  );


  and
  g878
  (
    n951,
    n131,
    n141,
    n68,
    n111
  );


  nand
  g879
  (
    n880,
    n190,
    n140,
    n182,
    n125
  );


  or
  g880
  (
    n675,
    n70,
    n203,
    n111,
    n135
  );


  nor
  g881
  (
    n836,
    n229,
    n227,
    n179,
    n99
  );


  or
  g882
  (
    n747,
    n150,
    n223,
    n100,
    n247
  );


  or
  g883
  (
    n926,
    n65,
    n164,
    n196,
    n149
  );


  and
  g884
  (
    n277,
    n72,
    n134,
    n168,
    n250
  );


  xnor
  g885
  (
    n722,
    n119,
    n80,
    n237,
    n102
  );


  or
  g886
  (
    n875,
    n153,
    n127,
    n223,
    n53
  );


  xnor
  g887
  (
    n518,
    n231,
    n246,
    n76,
    n197
  );


  xnor
  g888
  (
    n755,
    n181,
    n101,
    n233,
    n56
  );


  nor
  g889
  (
    n640,
    n220,
    n158,
    n92,
    n77
  );


  xor
  g890
  (
    n477,
    n230,
    n182,
    n130,
    n195
  );


  nand
  g891
  (
    n870,
    n188,
    n137,
    n106
  );


  nor
  g892
  (
    n617,
    n94,
    n104,
    n66,
    n151
  );


  or
  g893
  (
    n770,
    n219,
    n224,
    n83,
    n233
  );


  nand
  g894
  (
    n289,
    n84,
    n245,
    n239,
    n156
  );


  xnor
  g895
  (
    n711,
    n238,
    n199,
    n74,
    n204
  );


  xor
  g896
  (
    n460,
    n176,
    n195,
    n198,
    n76
  );


  nor
  g897
  (
    n425,
    n71,
    n102,
    n141,
    n161
  );


  nor
  g898
  (
    n616,
    n230,
    n134,
    n52,
    n66
  );


  nand
  g899
  (
    n908,
    n173,
    n170,
    n81,
    n169
  );


  buf
  g900
  (
    n1052,
    n258
  );


  not
  g901
  (
    n1024,
    n336
  );


  not
  g902
  (
    n1077,
    n327
  );


  buf
  g903
  (
    n985,
    n349
  );


  buf
  g904
  (
    n960,
    n334
  );


  not
  g905
  (
    n1012,
    n310
  );


  buf
  g906
  (
    n989,
    n357
  );


  buf
  g907
  (
    n981,
    n293
  );


  buf
  g908
  (
    n1026,
    n265
  );


  not
  g909
  (
    n978,
    n303
  );


  buf
  g910
  (
    n961,
    n262
  );


  buf
  g911
  (
    n1008,
    n259
  );


  not
  g912
  (
    n1023,
    n278
  );


  buf
  g913
  (
    n1064,
    n317
  );


  not
  g914
  (
    n1075,
    n368
  );


  buf
  g915
  (
    n992,
    n318
  );


  not
  g916
  (
    n991,
    n364
  );


  buf
  g917
  (
    n1065,
    n320
  );


  buf
  g918
  (
    n1063,
    n252
  );


  not
  g919
  (
    n1037,
    n305
  );


  buf
  g920
  (
    n1035,
    n281
  );


  buf
  g921
  (
    n982,
    n298
  );


  buf
  g922
  (
    n1034,
    n362
  );


  buf
  g923
  (
    n1047,
    n356
  );


  not
  g924
  (
    n1003,
    n329
  );


  buf
  g925
  (
    n996,
    n276
  );


  buf
  g926
  (
    n1053,
    n299
  );


  buf
  g927
  (
    n969,
    n354
  );


  buf
  g928
  (
    n1018,
    n351
  );


  not
  g929
  (
    n1071,
    n269
  );


  not
  g930
  (
    n1066,
    n330
  );


  buf
  g931
  (
    n1060,
    n315
  );


  not
  g932
  (
    n1030,
    n280
  );


  buf
  g933
  (
    n993,
    n251
  );


  buf
  g934
  (
    n976,
    n308
  );


  not
  g935
  (
    n1062,
    n339
  );


  buf
  g936
  (
    n1015,
    n307
  );


  buf
  g937
  (
    n997,
    n360
  );


  buf
  g938
  (
    n983,
    n286
  );


  not
  g939
  (
    KeyWire_0_13,
    n343
  );


  buf
  g940
  (
    n1036,
    n254
  );


  not
  g941
  (
    n1004,
    n345
  );


  buf
  g942
  (
    n1021,
    n367
  );


  buf
  g943
  (
    n999,
    n260
  );


  not
  g944
  (
    n1049,
    n355
  );


  not
  g945
  (
    n972,
    n287
  );


  buf
  g946
  (
    n1050,
    n319
  );


  not
  g947
  (
    KeyWire_0_27,
    n359
  );


  not
  g948
  (
    n965,
    n328
  );


  not
  g949
  (
    n1076,
    n285
  );


  not
  g950
  (
    n984,
    n361
  );


  not
  g951
  (
    KeyWire_0_10,
    n272
  );


  not
  g952
  (
    n988,
    n335
  );


  buf
  g953
  (
    n994,
    n353
  );


  not
  g954
  (
    n1009,
    n277
  );


  buf
  g955
  (
    n1006,
    n289
  );


  buf
  g956
  (
    n1038,
    n270
  );


  buf
  g957
  (
    n970,
    n342
  );


  buf
  g958
  (
    n1016,
    n314
  );


  not
  g959
  (
    n1054,
    n267
  );


  buf
  g960
  (
    n1042,
    n350
  );


  buf
  g961
  (
    n995,
    n256
  );


  buf
  g962
  (
    n1029,
    n302
  );


  not
  g963
  (
    n973,
    n284
  );


  not
  g964
  (
    n1068,
    n264
  );


  buf
  g965
  (
    n974,
    n322
  );


  not
  g966
  (
    n975,
    n283
  );


  buf
  g967
  (
    KeyWire_0_24,
    n358
  );


  buf
  g968
  (
    n987,
    n268
  );


  not
  g969
  (
    n1040,
    n290
  );


  not
  g970
  (
    n1057,
    n338
  );


  buf
  g971
  (
    n1025,
    n295
  );


  buf
  g972
  (
    n1014,
    n292
  );


  buf
  g973
  (
    n1069,
    n275
  );


  buf
  g974
  (
    n986,
    n347
  );


  buf
  g975
  (
    n1043,
    n309
  );


  not
  g976
  (
    n1059,
    n332
  );


  buf
  g977
  (
    n1044,
    n291
  );


  not
  g978
  (
    n966,
    n296
  );


  not
  g979
  (
    n1002,
    n294
  );


  buf
  g980
  (
    n1072,
    n348
  );


  buf
  g981
  (
    n1061,
    n311
  );


  not
  g982
  (
    n1019,
    n271
  );


  not
  g983
  (
    n1041,
    n255
  );


  buf
  g984
  (
    n1067,
    n253
  );


  not
  g985
  (
    n1020,
    n346
  );


  not
  g986
  (
    n1074,
    n344
  );


  buf
  g987
  (
    n1046,
    n331
  );


  buf
  g988
  (
    n1027,
    n301
  );


  buf
  g989
  (
    n998,
    n279
  );


  not
  g990
  (
    n977,
    n363
  );


  buf
  g991
  (
    n968,
    n352
  );


  buf
  g992
  (
    n1005,
    n288
  );


  buf
  g993
  (
    n980,
    n325
  );


  not
  g994
  (
    n962,
    n323
  );


  not
  g995
  (
    n990,
    n340
  );


  not
  g996
  (
    n1039,
    n366
  );


  not
  g997
  (
    n971,
    n297
  );


  not
  g998
  (
    n1022,
    n274
  );


  not
  g999
  (
    n1070,
    n326
  );


  not
  g1000
  (
    n1073,
    n300
  );


  buf
  g1001
  (
    n1028,
    n306
  );


  buf
  g1002
  (
    n1048,
    n324
  );


  not
  g1003
  (
    n1032,
    n273
  );


  buf
  g1004
  (
    n1056,
    n341
  );


  not
  g1005
  (
    n1017,
    n312
  );


  buf
  g1006
  (
    n1001,
    n263
  );


  buf
  g1007
  (
    n1055,
    n304
  );


  buf
  g1008
  (
    n964,
    n316
  );


  buf
  g1009
  (
    n1033,
    n333
  );


  buf
  g1010
  (
    n979,
    n257
  );


  not
  g1011
  (
    n967,
    n313
  );


  not
  g1012
  (
    n1013,
    n365
  );


  not
  g1013
  (
    n1051,
    n266
  );


  not
  g1014
  (
    n1045,
    n321
  );


  not
  g1015
  (
    n1007,
    n282
  );


  not
  g1016
  (
    n1058,
    n261
  );


  not
  g1017
  (
    n1010,
    n337
  );


  or
  g1018
  (
    n1081,
    n413,
    n375,
    n969,
    n383
  );


  nor
  g1019
  (
    n1082,
    n393,
    n414,
    n401,
    n396
  );


  nand
  g1020
  (
    n1090,
    n372,
    n972,
    n974,
    n964
  );


  and
  g1021
  (
    n1092,
    n961,
    n975,
    n384,
    n411
  );


  xor
  g1022
  (
    n1086,
    n371,
    n391,
    n387,
    n405
  );


  and
  g1023
  (
    n1088,
    n399,
    n407,
    n386,
    n380
  );


  nand
  g1024
  (
    n1079,
    n398,
    n970,
    n963,
    n965
  );


  nand
  g1025
  (
    n1089,
    n379,
    n388,
    n416,
    n392
  );


  xnor
  g1026
  (
    n1083,
    n390,
    n408,
    n377,
    n395
  );


  and
  g1027
  (
    n1078,
    n376,
    n373,
    n397,
    n370
  );


  nand
  g1028
  (
    n1080,
    n966,
    n385,
    n971,
    n960
  );


  nand
  g1029
  (
    n1093,
    n403,
    n374,
    n410,
    n382
  );


  xnor
  g1030
  (
    n1084,
    n973,
    n968,
    n409,
    n394
  );


  xnor
  g1031
  (
    n1087,
    n406,
    n369,
    n404,
    n402
  );


  xnor
  g1032
  (
    n1085,
    n381,
    n378,
    n400,
    n967
  );


  nor
  g1033
  (
    n1091,
    n412,
    n962,
    n389,
    n415
  );


  nand
  g1034
  (
    n1122,
    n981,
    n1044,
    n1088,
    n1041
  );


  xnor
  g1035
  (
    KeyWire_0_6,
    n1045,
    n993,
    n1027,
    n1043
  );


  nand
  g1036
  (
    n1103,
    n1083,
    n1033,
    n1046,
    n987
  );


  and
  g1037
  (
    n1104,
    n1038,
    n1006,
    n1089,
    n1022
  );


  nor
  g1038
  (
    n1108,
    n1009,
    n1026,
    n994,
    n1088
  );


  and
  g1039
  (
    n1095,
    n1039,
    n1045,
    n1011,
    n1023
  );


  xor
  g1040
  (
    n1101,
    n1037,
    n1014,
    n1005,
    n1078
  );


  nand
  g1041
  (
    n1119,
    n1029,
    n1091,
    n1044,
    n1036
  );


  nor
  g1042
  (
    n1111,
    n977,
    n999,
    n1084,
    n1028
  );


  and
  g1043
  (
    n1120,
    n1080,
    n1019,
    n1007,
    n1003
  );


  xor
  g1044
  (
    n1097,
    n1045,
    n1016,
    n1024,
    n986
  );


  nor
  g1045
  (
    n1102,
    n1032,
    n1087,
    n1089,
    n1090
  );


  nor
  g1046
  (
    n1115,
    n998,
    n1020,
    n991,
    n1041
  );


  nor
  g1047
  (
    n1116,
    n1079,
    n980,
    n1087,
    n1085
  );


  nor
  g1048
  (
    n1118,
    n979,
    n1015,
    n1002,
    n1042
  );


  and
  g1049
  (
    n1096,
    n1041,
    n992,
    n1012,
    n982
  );


  nand
  g1050
  (
    n1121,
    n1087,
    n1090,
    n988,
    n1004
  );


  xnor
  g1051
  (
    n1113,
    n996,
    n1017,
    n1088,
    n1086
  );


  xor
  g1052
  (
    n1100,
    n976,
    n1081,
    n1043,
    n1000
  );


  nand
  g1053
  (
    n1107,
    n1087,
    n1086,
    n1042,
    n1010
  );


  nand
  g1054
  (
    n1094,
    n990,
    n1090,
    n1089,
    n1034
  );


  nor
  g1055
  (
    n1117,
    n1082,
    n1018,
    n1043,
    n1042
  );


  nand
  g1056
  (
    n1112,
    n1044,
    n1089,
    n1042,
    n1088
  );


  and
  g1057
  (
    n1105,
    n978,
    n1041,
    n1013,
    n984
  );


  or
  g1058
  (
    n1099,
    n1035,
    n989,
    n1008,
    n997
  );


  nand
  g1059
  (
    n1098,
    n1046,
    n1001,
    n995,
    n1090
  );


  or
  g1060
  (
    n1106,
    n1025,
    n1085,
    n1043,
    n1021
  );


  xnor
  g1061
  (
    n1114,
    n1040,
    n1030,
    n1091,
    n983
  );


  nand
  g1062
  (
    n1109,
    n1044,
    n1031,
    n1045,
    n985
  );


  buf
  g1063
  (
    n1129,
    n1048
  );


  buf
  g1064
  (
    n1126,
    n1091
  );


  buf
  g1065
  (
    n1136,
    n1109
  );


  buf
  g1066
  (
    n1133,
    n1105
  );


  buf
  g1067
  (
    n1134,
    n1098
  );


  not
  g1068
  (
    n1123,
    n1107
  );


  not
  g1069
  (
    n1137,
    n1106
  );


  buf
  g1070
  (
    n1127,
    n1100
  );


  not
  g1071
  (
    n1131,
    n1047
  );


  buf
  g1072
  (
    n1130,
    n1096
  );


  and
  g1073
  (
    n1124,
    n1108,
    n1047
  );


  xnor
  g1074
  (
    n1138,
    n1048,
    n1099,
    n1097,
    n1049
  );


  or
  g1075
  (
    n1135,
    n1049,
    n1049,
    n1103,
    n1048
  );


  and
  g1076
  (
    n1128,
    n1049,
    n1104,
    n1046
  );


  nor
  g1077
  (
    n1125,
    n1101,
    n1048,
    n1102,
    n1094
  );


  xnor
  g1078
  (
    KeyWire_0_25,
    n1047,
    n1047,
    n1091,
    n1095
  );


  nand
  g1079
  (
    n1164,
    n526,
    n433,
    n442,
    n1126
  );


  xnor
  g1080
  (
    n1170,
    n1133,
    n1120,
    n490,
    n499
  );


  and
  g1081
  (
    n1162,
    n528,
    n523,
    n509,
    n1138
  );


  or
  g1082
  (
    n1151,
    n455,
    n431,
    n519,
    n498
  );


  xor
  g1083
  (
    n1180,
    n1136,
    n452,
    n454,
    n1134
  );


  xor
  g1084
  (
    n1152,
    n423,
    n437,
    n1131,
    n480
  );


  xnor
  g1085
  (
    KeyWire_0_7,
    n473,
    n478,
    n504,
    n427
  );


  nand
  g1086
  (
    n1145,
    n1111,
    n483,
    n463,
    n445
  );


  nor
  g1087
  (
    n1155,
    n489,
    n482,
    n448,
    n1130
  );


  and
  g1088
  (
    n1179,
    n1132,
    n1110,
    n527,
    n1131
  );


  or
  g1089
  (
    n1148,
    n522,
    n1138,
    n520,
    n1129
  );


  xnor
  g1090
  (
    n1177,
    n496,
    n1128,
    n525,
    n497
  );


  nor
  g1091
  (
    KeyWire_0_2,
    n1137,
    n517,
    n502,
    n429
  );


  nand
  g1092
  (
    n1142,
    n447,
    n1137,
    n1133
  );


  xor
  g1093
  (
    n1158,
    n1136,
    n1133,
    n451,
    n1112
  );


  and
  g1094
  (
    n1175,
    n417,
    n1129,
    n459,
    n1127
  );


  and
  g1095
  (
    n1167,
    n1138,
    n485,
    n479,
    n471
  );


  xnor
  g1096
  (
    n1143,
    n1136,
    n464,
    n470,
    n515
  );


  xnor
  g1097
  (
    n1140,
    n432,
    n446,
    n1118,
    n516
  );


  xnor
  g1098
  (
    n1159,
    n1132,
    n1136,
    n458,
    n1135
  );


  or
  g1099
  (
    n1144,
    n450,
    n512,
    n1134,
    n1128
  );


  nand
  g1100
  (
    n1165,
    n1115,
    n422,
    n1125,
    n476
  );


  xor
  g1101
  (
    n1141,
    n441,
    n1135,
    n494,
    n1125
  );


  xnor
  g1102
  (
    n1157,
    n420,
    n467,
    n484,
    n508
  );


  and
  g1103
  (
    n1147,
    n434,
    n492,
    n1117,
    n449
  );


  xnor
  g1104
  (
    n1163,
    n477,
    n440,
    n475,
    n465
  );


  xnor
  g1105
  (
    n1174,
    n1119,
    n518,
    n530,
    n424
  );


  or
  g1106
  (
    n1169,
    n425,
    n461,
    n507,
    n481
  );


  xor
  g1107
  (
    n1171,
    n495,
    n468,
    n436,
    n430
  );


  nor
  g1108
  (
    n1150,
    n1127,
    n1135,
    n531
  );


  or
  g1109
  (
    n1149,
    n419,
    n510,
    n435,
    n503
  );


  xor
  g1110
  (
    n1161,
    n500,
    n460,
    n438,
    n426
  );


  and
  g1111
  (
    n1154,
    n486,
    n453,
    n472,
    n1138
  );


  xnor
  g1112
  (
    n1156,
    n462,
    n1133,
    n506,
    n1130
  );


  xor
  g1113
  (
    n1146,
    n1123,
    n511,
    n466,
    n505
  );


  or
  g1114
  (
    n1173,
    n491,
    n514,
    n1126,
    n457
  );


  nand
  g1115
  (
    n1176,
    n1134,
    n487,
    n444,
    n1113
  );


  xnor
  g1116
  (
    n1168,
    n1114,
    n439,
    n474,
    n1124
  );


  or
  g1117
  (
    KeyWire_0_52,
    n469,
    n521,
    n1134,
    n488
  );


  and
  g1118
  (
    n1139,
    n529,
    n421,
    n418,
    n513
  );


  nor
  g1119
  (
    n1178,
    n493,
    n501,
    n1116,
    n443
  );


  xor
  g1120
  (
    n1153,
    n428,
    n1137,
    n456,
    n524
  );


  not
  g1121
  (
    n1208,
    n1140
  );


  not
  g1122
  (
    n1192,
    n1144
  );


  buf
  g1123
  (
    n1197,
    n1149
  );


  not
  g1124
  (
    n1201,
    n1142
  );


  buf
  g1125
  (
    n1199,
    n1154
  );


  buf
  g1126
  (
    n1185,
    n1150
  );


  buf
  g1127
  (
    n1211,
    n1146
  );


  buf
  g1128
  (
    n1212,
    n1051
  );


  buf
  g1129
  (
    n1189,
    n1150
  );


  not
  g1130
  (
    n1220,
    n1142
  );


  buf
  g1131
  (
    n1196,
    n1147
  );


  not
  g1132
  (
    n1200,
    n1147
  );


  not
  g1133
  (
    n1190,
    n1153
  );


  buf
  g1134
  (
    n1216,
    n1140
  );


  not
  g1135
  (
    n1181,
    n1149
  );


  buf
  g1136
  (
    n1202,
    n1155
  );


  buf
  g1137
  (
    n1186,
    n1155
  );


  buf
  g1138
  (
    n1182,
    n1148
  );


  buf
  g1139
  (
    n1194,
    n1152
  );


  buf
  g1140
  (
    n1184,
    n1147
  );


  buf
  g1141
  (
    n1206,
    n1140
  );


  buf
  g1142
  (
    n1183,
    n1141
  );


  buf
  g1143
  (
    n1215,
    n1152
  );


  not
  g1144
  (
    n1195,
    n1145
  );


  not
  g1145
  (
    n1193,
    n1145
  );


  buf
  g1146
  (
    n1217,
    n1149
  );


  buf
  g1147
  (
    n1203,
    n1050
  );


  and
  g1148
  (
    n1204,
    n1140,
    n1139,
    n1154,
    n1145
  );


  xor
  g1149
  (
    n1187,
    n1144,
    n1151,
    n532
  );


  and
  g1150
  (
    n1219,
    n1142,
    n1148,
    n1149,
    n1154
  );


  and
  g1151
  (
    n1191,
    n1156,
    n1150,
    n1050,
    n1147
  );


  or
  g1152
  (
    n1213,
    n1153,
    n1146,
    n1152
  );


  nand
  g1153
  (
    n1207,
    n1155,
    n1151
  );


  xor
  g1154
  (
    n1188,
    n1148,
    n1153,
    n1150,
    n1139
  );


  nand
  g1155
  (
    n1209,
    n1145,
    n1156,
    n1146
  );


  xnor
  g1156
  (
    n1198,
    n1148,
    n1143,
    n1142,
    n1141
  );


  xnor
  g1157
  (
    n1214,
    n1143,
    n1143,
    n1139,
    n1051
  );


  xnor
  g1158
  (
    n1205,
    n1143,
    n1139,
    n1141,
    n1154
  );


  xor
  g1159
  (
    n1210,
    n1157,
    n1144,
    n1146
  );


  and
  g1160
  (
    n1218,
    n1153,
    n1156,
    n1141,
    n1050
  );


  nand
  g1161
  (
    n1232,
    n1161,
    n1162,
    n1197,
    n1170
  );


  nor
  g1162
  (
    n1238,
    n1175,
    n1161,
    n1169,
    n1190
  );


  or
  g1163
  (
    n1222,
    n1193,
    n1174,
    n1167,
    n1160
  );


  nand
  g1164
  (
    n1236,
    n1205,
    n1186,
    n1191,
    n1160
  );


  nor
  g1165
  (
    n1223,
    n1159,
    n1204,
    n1173,
    n1166
  );


  nor
  g1166
  (
    n1234,
    n1158,
    n1165,
    n1169,
    n1173
  );


  xnor
  g1167
  (
    n1225,
    n1158,
    n1161,
    n1203,
    n1166
  );


  nor
  g1168
  (
    n1226,
    n1202,
    n1158,
    n1172,
    n1163
  );


  nor
  g1169
  (
    n1239,
    n1167,
    n1172,
    n1169,
    n1198
  );


  and
  g1170
  (
    n1241,
    n1195,
    n1160,
    n1159,
    n1164
  );


  xor
  g1171
  (
    n1231,
    n1160,
    n1194,
    n1169,
    n1162
  );


  nor
  g1172
  (
    n1228,
    n1172,
    n1159,
    n1173,
    n1168
  );


  or
  g1173
  (
    n1227,
    n1187,
    n1166,
    n1172,
    n1159
  );


  xor
  g1174
  (
    n1243,
    n1196,
    n1158,
    n1164,
    n1171
  );


  nor
  g1175
  (
    n1240,
    n1174,
    n1175,
    n1181,
    n1185
  );


  xor
  g1176
  (
    n1235,
    n1161,
    n1174,
    n1164,
    n1199
  );


  xnor
  g1177
  (
    n1233,
    n1168,
    n1188,
    n1184,
    n1175
  );


  xor
  g1178
  (
    n1242,
    n1167,
    n1171,
    n1165,
    n1157
  );


  and
  g1179
  (
    n1245,
    n1164,
    n1163,
    n1200,
    n1165
  );


  or
  g1180
  (
    n1229,
    n1173,
    n1192,
    n1157,
    n1168
  );


  xnor
  g1181
  (
    n1221,
    n1163,
    n1189,
    n1182,
    n1162
  );


  and
  g1182
  (
    n1224,
    n1165,
    n1183,
    n1170
  );


  or
  g1183
  (
    n1244,
    n1162,
    n1171,
    n1170,
    n1157
  );


  or
  g1184
  (
    n1230,
    n1167,
    n1175,
    n1174,
    n1201
  );


  xor
  g1185
  (
    n1237,
    n1171,
    n1166,
    n1168,
    n1163
  );


  buf
  g1186
  (
    n1266,
    n1234
  );


  buf
  g1187
  (
    n1263,
    n1227
  );


  not
  g1188
  (
    n1256,
    n1235
  );


  not
  g1189
  (
    n1251,
    n1236
  );


  not
  g1190
  (
    n1252,
    n1229
  );


  not
  g1191
  (
    n1267,
    n1228
  );


  not
  g1192
  (
    n1260,
    n1242
  );


  buf
  g1193
  (
    n1265,
    n1243
  );


  not
  g1194
  (
    n1250,
    n1241
  );


  not
  g1195
  (
    n1255,
    n1240
  );


  not
  g1196
  (
    n1248,
    n1230
  );


  buf
  g1197
  (
    n1259,
    n1222
  );


  not
  g1198
  (
    n1247,
    n1226
  );


  buf
  g1199
  (
    n1258,
    n1237
  );


  buf
  g1200
  (
    n1246,
    n1223
  );


  not
  g1201
  (
    n1264,
    n1233
  );


  not
  g1202
  (
    n1269,
    n1238
  );


  buf
  g1203
  (
    KeyWire_0_58,
    n1232
  );


  buf
  g1204
  (
    n1268,
    n1231
  );


  not
  g1205
  (
    n1249,
    n1224
  );


  not
  g1206
  (
    n1257,
    n1225
  );


  not
  g1207
  (
    n1254,
    n1244
  );


  not
  g1208
  (
    n1262,
    n1239
  );


  buf
  g1209
  (
    n1253,
    n1221
  );


  buf
  g1210
  (
    n1272,
    n1248
  );


  not
  g1211
  (
    KeyWire_0_14,
    n1250
  );


  buf
  g1212
  (
    n1287,
    n1249
  );


  not
  g1213
  (
    n1292,
    n1250
  );


  not
  g1214
  (
    n1282,
    n1248
  );


  buf
  g1215
  (
    n1277,
    n1251
  );


  buf
  g1216
  (
    n1288,
    n1246
  );


  not
  g1217
  (
    KeyWire_0_20,
    n1249
  );


  buf
  g1218
  (
    n1289,
    n1249
  );


  not
  g1219
  (
    n1285,
    n1246
  );


  buf
  g1220
  (
    n1283,
    n1251
  );


  buf
  g1221
  (
    n1291,
    n1246
  );


  not
  g1222
  (
    n1280,
    n1247
  );


  not
  g1223
  (
    n1281,
    n1251
  );


  buf
  g1224
  (
    n1271,
    n1248
  );


  not
  g1225
  (
    n1278,
    n1247
  );


  not
  g1226
  (
    n1274,
    n1246
  );


  buf
  g1227
  (
    n1286,
    n1247
  );


  not
  g1228
  (
    n1279,
    n1248
  );


  buf
  g1229
  (
    n1284,
    n1249
  );


  not
  g1230
  (
    n1276,
    n1250
  );


  not
  g1231
  (
    KeyWire_0_35,
    n1250
  );


  xor
  g1232
  (
    n1273,
    n1244,
    n1247
  );


  buf
  g1233
  (
    n1372,
    n1269
  );


  buf
  g1234
  (
    n1361,
    n1283
  );


  not
  g1235
  (
    n1316,
    n1275
  );


  buf
  g1236
  (
    n1298,
    n1260
  );


  buf
  g1237
  (
    n1320,
    n1271
  );


  buf
  g1238
  (
    n1341,
    n1283
  );


  not
  g1239
  (
    n1326,
    n1265
  );


  buf
  g1240
  (
    n1324,
    n1179
  );


  buf
  g1241
  (
    n1371,
    n1178
  );


  not
  g1242
  (
    n1319,
    n1290
  );


  buf
  g1243
  (
    n1308,
    n1262
  );


  buf
  g1244
  (
    n1342,
    n1285
  );


  not
  g1245
  (
    n1367,
    n1256
  );


  not
  g1246
  (
    n1305,
    n1277
  );


  buf
  g1247
  (
    n1339,
    n1274
  );


  buf
  g1248
  (
    n1313,
    n1258
  );


  not
  g1249
  (
    n1358,
    n1270
  );


  buf
  g1250
  (
    n1381,
    n1253
  );


  buf
  g1251
  (
    n1302,
    n1270
  );


  not
  g1252
  (
    n1321,
    n1281
  );


  not
  g1253
  (
    n1345,
    n1264
  );


  buf
  g1254
  (
    n1347,
    n1275
  );


  buf
  g1255
  (
    n1380,
    n1273
  );


  buf
  g1256
  (
    n1333,
    n1268
  );


  not
  g1257
  (
    n1306,
    n1273
  );


  buf
  g1258
  (
    n1322,
    n1276
  );


  not
  g1259
  (
    n1354,
    n1268
  );


  buf
  g1260
  (
    n1310,
    n1284
  );


  buf
  g1261
  (
    n1353,
    n1275
  );


  buf
  g1262
  (
    n1351,
    n1280
  );


  buf
  g1263
  (
    n1373,
    n1180
  );


  not
  g1264
  (
    n1364,
    n1287
  );


  not
  g1265
  (
    n1295,
    n1180
  );


  not
  g1266
  (
    n1299,
    n1257
  );


  not
  g1267
  (
    n1370,
    n1253
  );


  not
  g1268
  (
    n1382,
    n1277
  );


  not
  g1269
  (
    n1348,
    n1179
  );


  buf
  g1270
  (
    n1365,
    n1262
  );


  not
  g1271
  (
    KeyWire_0_47,
    n1291
  );


  buf
  g1272
  (
    n1294,
    n1260
  );


  buf
  g1273
  (
    n1377,
    n1283
  );


  not
  g1274
  (
    n1343,
    n1266
  );


  buf
  g1275
  (
    n1314,
    n1177
  );


  not
  g1276
  (
    n1296,
    n1179
  );


  not
  g1277
  (
    n1357,
    n1276
  );


  not
  g1278
  (
    n1340,
    n1278
  );


  buf
  g1279
  (
    KeyWire_0_22,
    n1267
  );


  not
  g1280
  (
    n1335,
    n1261
  );


  not
  g1281
  (
    n1303,
    n1270
  );


  buf
  g1282
  (
    n1355,
    n1277
  );


  not
  g1283
  (
    n1301,
    n1252
  );


  buf
  g1284
  (
    n1384,
    n1259
  );


  buf
  g1285
  (
    n1366,
    n1267
  );


  buf
  g1286
  (
    n1300,
    n1268
  );


  buf
  g1287
  (
    n1315,
    n1261
  );


  buf
  g1288
  (
    n1329,
    n1253
  );


  buf
  g1289
  (
    n1359,
    n1262
  );


  buf
  g1290
  (
    n1325,
    n1287
  );


  buf
  g1291
  (
    n1312,
    n1282
  );


  not
  g1292
  (
    n1346,
    n1265
  );


  xor
  g1293
  (
    n1337,
    n1179,
    n534,
    n1282,
    n1271
  );


  or
  g1294
  (
    n1368,
    n1292,
    n1252,
    n1260,
    n1178
  );


  and
  g1295
  (
    n1328,
    n1283,
    n1274,
    n1291,
    n1288
  );


  and
  g1296
  (
    KeyWire_0_29,
    n1281,
    n1281,
    n1287,
    n1272
  );


  nor
  g1297
  (
    n1362,
    n1282,
    n1273,
    n1286,
    n1264
  );


  xor
  g1298
  (
    n1374,
    n1256,
    n1280,
    n1284
  );


  or
  g1299
  (
    n1307,
    n1264,
    n1259,
    n1266,
    n1279
  );


  nor
  g1300
  (
    n1323,
    n1289,
    n1263,
    n1287,
    n1290
  );


  or
  g1301
  (
    n1338,
    n1290,
    n1279,
    n1257,
    n1259
  );


  nor
  g1302
  (
    n1375,
    n1281,
    n1177,
    n1180
  );


  xnor
  g1303
  (
    n1383,
    n1252,
    n1269,
    n1285,
    n1280
  );


  nor
  g1304
  (
    n1332,
    n1275,
    n1267,
    n1285,
    n1254
  );


  nand
  g1305
  (
    n1297,
    n1282,
    n1265,
    n1251,
    n1285
  );


  and
  g1306
  (
    n1330,
    n1176,
    n1276,
    n1255,
    n1279
  );


  nor
  g1307
  (
    n1344,
    n1177,
    n1278,
    n1257,
    n1254
  );


  or
  g1308
  (
    n1369,
    n1258,
    n1178,
    n1261,
    n1292
  );


  nor
  g1309
  (
    n1349,
    n1269,
    n1258,
    n1291,
    n1256
  );


  nor
  g1310
  (
    n1376,
    n1289,
    n1255,
    n1265,
    n1268
  );


  or
  g1311
  (
    n1378,
    n533,
    n1266,
    n1276,
    n1263
  );


  xor
  g1312
  (
    n1363,
    n1279,
    n1272,
    n1291,
    n1254
  );


  or
  g1313
  (
    n1317,
    n1266,
    n1288,
    n1177,
    n1278
  );


  xnor
  g1314
  (
    n1334,
    n1267,
    n1288,
    n1272,
    n1269
  );


  and
  g1315
  (
    n1350,
    n1289,
    n1261,
    n1264,
    n1257
  );


  xnor
  g1316
  (
    n1311,
    n1178,
    n1176,
    n1278,
    n1259
  );


  and
  g1317
  (
    n1327,
    n1288,
    n1286,
    n1263,
    n1284
  );


  nand
  g1318
  (
    n1379,
    n1271,
    n1290,
    n1286,
    n1260
  );


  xnor
  g1319
  (
    n1356,
    n1280,
    n1255,
    n1176,
    n1256
  );


  nand
  g1320
  (
    n1360,
    n1176,
    n1274,
    n1258,
    n1262
  );


  or
  g1321
  (
    n1293,
    n1286,
    n1253,
    n1289,
    n1292
  );


  nor
  g1322
  (
    n1336,
    n1273,
    n535,
    n1252,
    n1263
  );


  nor
  g1323
  (
    n1304,
    n1271,
    n1272,
    n1277,
    n1255
  );


  or
  g1324
  (
    n1331,
    n1292,
    n1274,
    n1270,
    n1254
  );


  and
  g1325
  (
    n1402,
    n1311,
    n1309,
    n1338,
    n1335
  );


  nand
  g1326
  (
    n1392,
    n1316,
    n1354,
    n1377,
    n1340
  );


  nand
  g1327
  (
    n1391,
    n1297,
    n1327,
    n1345,
    n1370
  );


  nand
  g1328
  (
    n1414,
    n1378,
    n1343,
    n1306,
    n1295
  );


  xor
  g1329
  (
    n1411,
    n1331,
    n1320,
    n1376,
    n1365
  );


  nand
  g1330
  (
    n1409,
    n1300,
    n1321,
    n1296,
    n1307
  );


  nand
  g1331
  (
    n1408,
    n1374,
    n1372,
    n1366,
    n1371
  );


  nor
  g1332
  (
    n1396,
    n1378,
    n1379,
    n1374,
    n1357
  );


  or
  g1333
  (
    n1400,
    n1362,
    n1317,
    n1293,
    n1337
  );


  nor
  g1334
  (
    n1405,
    n1373,
    n1319,
    n1370,
    n1371
  );


  nor
  g1335
  (
    n1399,
    n1352,
    n537,
    n1330,
    n1318
  );


  or
  g1336
  (
    n1404,
    n1374,
    n1339,
    n1379,
    n1347
  );


  nor
  g1337
  (
    n1410,
    n1329,
    n1373,
    n1356,
    n1333
  );


  xor
  g1338
  (
    n1388,
    n1328,
    n1303,
    n1375,
    n1324
  );


  and
  g1339
  (
    n1393,
    n1301,
    n1302,
    n1379,
    n1370
  );


  and
  g1340
  (
    n1407,
    n1326,
    n1314,
    n1322,
    n1358
  );


  nand
  g1341
  (
    n1397,
    n1374,
    n1376,
    n1377
  );


  xnor
  g1342
  (
    n1389,
    n1349,
    n1378,
    n1336,
    n1373
  );


  nand
  g1343
  (
    n1385,
    n1315,
    n1313,
    n1363,
    n1308
  );


  nor
  g1344
  (
    n1403,
    n1359,
    n1325,
    n1376,
    n1377
  );


  xor
  g1345
  (
    n1401,
    n1342,
    n1370,
    n1305,
    n1323
  );


  nand
  g1346
  (
    n1413,
    n1334,
    n1375,
    n1371,
    n1355
  );


  nor
  g1347
  (
    n1390,
    n1310,
    n1344,
    n1368,
    n1351
  );


  and
  g1348
  (
    n1386,
    n1371,
    n1346,
    n1377,
    n1348
  );


  nand
  g1349
  (
    n1406,
    n1361,
    n1372,
    n538,
    n1353
  );


  nand
  g1350
  (
    n1398,
    n1299,
    n1294,
    n536,
    n1312
  );


  nand
  g1351
  (
    n1412,
    n1373,
    n1360,
    n1341,
    n1298
  );


  xnor
  g1352
  (
    n1395,
    n1304,
    n1367,
    n1375,
    n1372
  );


  and
  g1353
  (
    n1394,
    n1364,
    n1378,
    n1369,
    n1375
  );


  or
  g1354
  (
    n1387,
    n1332,
    n539,
    n1372,
    n1350
  );


  xnor
  g1355
  (
    n1417,
    n1381,
    n1381,
    n1382,
    n1405
  );


  or
  g1356
  (
    n1421,
    n1380,
    n1407,
    n1384
  );


  nand
  g1357
  (
    n1418,
    n1383,
    n1382,
    n1408,
    n1409
  );


  and
  g1358
  (
    n1415,
    n1381,
    n1379,
    n1403,
    n1380
  );


  and
  g1359
  (
    n1419,
    n1404,
    n1384,
    n1383,
    n1380
  );


  or
  g1360
  (
    n1416,
    n1382,
    n1381,
    n1383,
    n1406
  );


  and
  g1361
  (
    n1420,
    n1382,
    n1380,
    n1383,
    n1384
  );


  buf
  g1362
  (
    KeyWire_0_37,
    n1420
  );


  not
  g1363
  (
    n1422,
    n540
  );


  nand
  g1364
  (
    n1424,
    n1419,
    n1421
  );


  not
  g1365
  (
    n1427,
    n1051
  );


  buf
  g1366
  (
    n1425,
    n1423
  );


  buf
  g1367
  (
    n1431,
    n1424
  );


  not
  g1368
  (
    n1430,
    n1423
  );


  buf
  g1369
  (
    n1432,
    n542
  );


  not
  g1370
  (
    n1433,
    n1424
  );


  xor
  g1371
  (
    n1428,
    n1423,
    n1424
  );


  xor
  g1372
  (
    n1429,
    n1424,
    n1052,
    n1422
  );


  nand
  g1373
  (
    n1426,
    n541,
    n1423,
    n1051
  );


  buf
  g1374
  (
    n1440,
    n1428
  );


  not
  g1375
  (
    n1441,
    n1425
  );


  not
  g1376
  (
    n1439,
    n1425
  );


  not
  g1377
  (
    n1443,
    n545
  );


  not
  g1378
  (
    n1437,
    n544
  );


  buf
  g1379
  (
    n1436,
    n548
  );


  not
  g1380
  (
    n1438,
    n547
  );


  buf
  g1381
  (
    n1444,
    n1427
  );


  buf
  g1382
  (
    n1434,
    n1427
  );


  not
  g1383
  (
    n1445,
    n1428
  );


  and
  g1384
  (
    n1442,
    n1426,
    n543,
    n1427,
    n546
  );


  xnor
  g1385
  (
    n1435,
    n1427,
    n1426
  );


  xor
  g1386
  (
    n1450,
    n1433,
    n1435,
    n559,
    n572
  );


  nand
  g1387
  (
    KeyWire_0_33,
    n550,
    n1436,
    n555,
    n574
  );


  and
  g1388
  (
    n1453,
    n1436,
    n1428,
    n1430,
    n569
  );


  xor
  g1389
  (
    n1460,
    n1438,
    n1433,
    n567,
    n1434
  );


  nor
  g1390
  (
    n1451,
    n1438,
    n570,
    n576,
    n565
  );


  nor
  g1391
  (
    n1452,
    n1439,
    n1435,
    n1437,
    n1430
  );


  xor
  g1392
  (
    n1458,
    n1430,
    n556,
    n577,
    n558
  );


  xor
  g1393
  (
    n1448,
    n1429,
    n571,
    n1433,
    n568
  );


  nand
  g1394
  (
    n1446,
    n562,
    n1435,
    n552,
    n1433
  );


  nor
  g1395
  (
    n1447,
    n561,
    n553,
    n575,
    n554
  );


  or
  g1396
  (
    KeyWire_0_46,
    n1432,
    n566,
    n1438,
    n1431
  );


  and
  g1397
  (
    n1457,
    n1430,
    n1429,
    n564,
    n1431
  );


  nand
  g1398
  (
    n1462,
    n1436,
    n573,
    n1431,
    n1439
  );


  or
  g1399
  (
    n1461,
    n1438,
    n551,
    n1428,
    n1436
  );


  xor
  g1400
  (
    n1463,
    n1429,
    n549,
    n1434,
    n1437
  );


  xor
  g1401
  (
    n1456,
    n1432,
    n1432,
    n560,
    n578
  );


  and
  g1402
  (
    n1449,
    n1437,
    n1432,
    n1429,
    n557
  );


  xnor
  g1403
  (
    n1454,
    n563,
    n1431,
    n1435,
    n1437
  );


  or
  g1404
  (
    n1464,
    n1440,
    n1451,
    n1439
  );


  not
  g1405
  (
    n1465,
    n1464
  );


  not
  g1406
  (
    KeyWire_0_51,
    n1464
  );


  nand
  g1407
  (
    n1474,
    n597,
    n1465,
    n601,
    n595
  );


  nor
  g1408
  (
    KeyWire_0_61,
    n1466,
    n584,
    n585,
    n589
  );


  xnor
  g1409
  (
    KeyWire_0_8,
    n587,
    n588,
    n600,
    n582
  );


  and
  g1410
  (
    n1471,
    n599,
    n1466,
    n583,
    n596
  );


  or
  g1411
  (
    n1468,
    n580,
    n602,
    n1465
  );


  nor
  g1412
  (
    n1472,
    n593,
    n590,
    n586,
    n592
  );


  xor
  g1413
  (
    n1467,
    n1465,
    n591,
    n1466,
    n579
  );


  xor
  g1414
  (
    n1469,
    n598,
    n581,
    n594,
    n1466
  );


  buf
  g1415
  (
    n1476,
    n1440
  );


  not
  g1416
  (
    n1481,
    n604
  );


  buf
  g1417
  (
    n1486,
    n1472
  );


  buf
  g1418
  (
    n1479,
    n1441
  );


  not
  g1419
  (
    n1482,
    n1468
  );


  not
  g1420
  (
    n1478,
    n1441
  );


  buf
  g1421
  (
    n1483,
    n1469
  );


  nand
  g1422
  (
    n1475,
    n1469,
    n1472
  );


  or
  g1423
  (
    n1484,
    n610,
    n1471
  );


  nand
  g1424
  (
    n1485,
    n1440,
    n1471,
    n603
  );


  nor
  g1425
  (
    n1488,
    n1470,
    n1441,
    n1471
  );


  nand
  g1426
  (
    n1487,
    n1441,
    n1467,
    n607
  );


  or
  g1427
  (
    n1480,
    n608,
    n609,
    n1470
  );


  nor
  g1428
  (
    n1477,
    n1472,
    n605,
    n1440
  );


  nor
  g1429
  (
    n1489,
    n1468,
    n1472,
    n606
  );


  xor
  g1430
  (
    n1492,
    n1474,
    n1474,
    n1479,
    n1207
  );


  xor
  g1431
  (
    n1493,
    n1208,
    n1481,
    n1482
  );


  and
  g1432
  (
    n1501,
    n611,
    n1480,
    n1478,
    n1206
  );


  xnor
  g1433
  (
    n1500,
    n1213,
    n612,
    n1477,
    n614
  );


  nor
  g1434
  (
    n1496,
    n1481,
    n616,
    n1476,
    n1210
  );


  or
  g1435
  (
    n1490,
    n1212,
    n1479,
    n1473
  );


  or
  g1436
  (
    n1494,
    n1480,
    n1483,
    n1481,
    n613
  );


  nor
  g1437
  (
    n1499,
    n1482,
    n1478
  );


  xor
  g1438
  (
    n1498,
    n1214,
    n1473,
    n1474
  );


  or
  g1439
  (
    n1491,
    n1209,
    n1473,
    n615,
    n1480
  );


  nand
  g1440
  (
    n1495,
    n1479,
    n1475,
    n617,
    n1482
  );


  nor
  g1441
  (
    n1497,
    n1482,
    n1474,
    n1480,
    n1211
  );


  nor
  g1442
  (
    n1504,
    n618,
    n1484,
    n621,
    n627
  );


  and
  g1443
  (
    n1518,
    n1486,
    n1483,
    n1487,
    n631
  );


  and
  g1444
  (
    n1502,
    n1484,
    n1487,
    n622,
    n634
  );


  nand
  g1445
  (
    n1503,
    n1485,
    n1494,
    n1486,
    n630
  );


  xnor
  g1446
  (
    n1507,
    n641,
    n1494,
    n1492,
    n635
  );


  and
  g1447
  (
    n1515,
    n1486,
    n1485,
    n620,
    n1489
  );


  xnor
  g1448
  (
    n1516,
    n1490,
    n628,
    n1491,
    n629
  );


  xnor
  g1449
  (
    n1514,
    n1489,
    n1493,
    n640,
    n636
  );


  nand
  g1450
  (
    n1510,
    n1486,
    n1493,
    n1491,
    n1484
  );


  and
  g1451
  (
    n1512,
    n624,
    n1485,
    n1489,
    n1493
  );


  nor
  g1452
  (
    n1513,
    n626,
    n1488,
    n1491,
    n632
  );


  nor
  g1453
  (
    n1508,
    n619,
    n1491,
    n623,
    n1493
  );


  nor
  g1454
  (
    n1517,
    n1492,
    n1489,
    n633,
    n1488
  );


  or
  g1455
  (
    n1505,
    n639,
    n1487,
    n1492,
    n1483
  );


  xor
  g1456
  (
    n1509,
    n1494,
    n1484,
    n1492,
    n1488
  );


  xor
  g1457
  (
    n1511,
    n1490,
    n1483,
    n637,
    n638
  );


  nand
  g1458
  (
    n1506,
    n1487,
    n625,
    n1488,
    n1485
  );


  nand
  g1459
  (
    n1528,
    n1508,
    n1495,
    n1216,
    n1499
  );


  xor
  g1460
  (
    n1526,
    n1442,
    n1509,
    n1500
  );


  nand
  g1461
  (
    n1524,
    n1499,
    n646,
    n642,
    n1497
  );


  xnor
  g1462
  (
    n1519,
    n649,
    n1505,
    n1500,
    n1498
  );


  or
  g1463
  (
    n1523,
    n1499,
    n1216,
    n1497,
    n1501
  );


  nand
  g1464
  (
    n1525,
    n1497,
    n645,
    n1216,
    n1442
  );


  nor
  g1465
  (
    n1520,
    n653,
    n1512,
    n1518,
    n1501
  );


  or
  g1466
  (
    n1532,
    n1517,
    n1496,
    n1516,
    n1514
  );


  nand
  g1467
  (
    n1521,
    n1498,
    n648,
    n1495,
    n1496
  );


  nor
  g1468
  (
    n1531,
    n1511,
    n1442,
    n1494,
    n644
  );


  xnor
  g1469
  (
    KeyWire_0_0,
    n1502,
    n1499,
    n1215,
    n1504
  );


  xnor
  g1470
  (
    n1533,
    n1495,
    n1515,
    n1507,
    n650
  );


  and
  g1471
  (
    n1535,
    n1496,
    n1495,
    n1216,
    n652
  );


  nor
  g1472
  (
    n1522,
    n1442,
    n1217,
    n1500,
    n1510
  );


  xor
  g1473
  (
    n1527,
    n1503,
    n1496,
    n1497,
    n1501
  );


  xnor
  g1474
  (
    n1530,
    n651,
    n1501,
    n1498,
    n1506
  );


  xnor
  g1475
  (
    n1529,
    n647,
    n1498,
    n1513,
    n643
  );


  nor
  g1476
  (
    n1568,
    n1526,
    n1076,
    n1068,
    n1075
  );


  nand
  g1477
  (
    n1561,
    n1073,
    n1069,
    n1220,
    n1443
  );


  or
  g1478
  (
    n1550,
    n1054,
    n1533,
    n1411,
    n1070
  );


  xnor
  g1479
  (
    n1547,
    n1217,
    n1066,
    n1070,
    n1454
  );


  xor
  g1480
  (
    n1541,
    n1071,
    n1062,
    n1217,
    n1063
  );


  or
  g1481
  (
    n1553,
    n1071,
    n1218,
    n1245,
    n1059
  );


  xor
  g1482
  (
    n1570,
    n1452,
    n1062,
    n1055,
    n1065
  );


  nor
  g1483
  (
    KeyWire_0_12,
    n1534,
    n1059,
    n1057,
    n1075
  );


  nor
  g1484
  (
    n1548,
    n1525,
    n1067,
    n1531
  );


  and
  g1485
  (
    n1544,
    n1219,
    n1064,
    n1533,
    n1072
  );


  nand
  g1486
  (
    n1579,
    n1534,
    n1443,
    n1531,
    n1072
  );


  or
  g1487
  (
    n1536,
    n1219,
    n1074,
    n1453,
    n1066
  );


  xnor
  g1488
  (
    n1572,
    n1076,
    n1532,
    n1056,
    n1062
  );


  or
  g1489
  (
    n1569,
    n1074,
    n1067,
    n1071,
    n1056
  );


  nor
  g1490
  (
    n1567,
    n1063,
    n1535,
    n1520,
    n1410
  );


  and
  g1491
  (
    n1543,
    n1076,
    n1055,
    n1069,
    n1071
  );


  xnor
  g1492
  (
    n1552,
    n1534,
    n1068,
    n1075,
    n1523
  );


  xor
  g1493
  (
    n1557,
    n1065,
    n1217,
    n1058,
    n1073
  );


  xnor
  g1494
  (
    n1556,
    n1065,
    n1058,
    n1072,
    n1052
  );


  xor
  g1495
  (
    n1582,
    n1056,
    n1524,
    n1065,
    n1075
  );


  xnor
  g1496
  (
    n1551,
    n1444,
    n1070,
    n1063,
    n1074
  );


  xnor
  g1497
  (
    n1537,
    n1058,
    n1519,
    n1060,
    n1521
  );


  nor
  g1498
  (
    n1564,
    n1069,
    n1534,
    n1059,
    n1220
  );


  nand
  g1499
  (
    n1539,
    n1528,
    n1526,
    n1218,
    n1220
  );


  xnor
  g1500
  (
    n1563,
    n1529,
    n1443,
    n1060,
    n1528
  );


  xor
  g1501
  (
    n1566,
    n1064,
    n1523,
    n1052,
    n1520
  );


  xor
  g1502
  (
    n1583,
    n1460,
    n1070,
    n1532,
    n1057
  );


  xor
  g1503
  (
    n1554,
    n1522,
    n1218,
    n1463,
    n1525
  );


  and
  g1504
  (
    n1577,
    n1220,
    n1055,
    n1054,
    n1063
  );


  xor
  g1505
  (
    n1578,
    n1062,
    n1458,
    n1053,
    n1061
  );


  xor
  g1506
  (
    n1560,
    n1531,
    n1412,
    n1053,
    n1461
  );


  xor
  g1507
  (
    n1562,
    n1058,
    n1532,
    n1064,
    n1076
  );


  xnor
  g1508
  (
    n1538,
    n1527,
    n1530,
    n1061
  );


  xnor
  g1509
  (
    n1571,
    n1457,
    n1066,
    n1530,
    n1068
  );


  nand
  g1510
  (
    n1549,
    n1413,
    n1068,
    n1456,
    n1535
  );


  or
  g1511
  (
    n1575,
    n1077,
    n1064,
    n1060,
    n1529
  );


  and
  g1512
  (
    n1559,
    n1057,
    n1533,
    n1067,
    n1245
  );


  nor
  g1513
  (
    n1555,
    n1077,
    n1069,
    n1053,
    n1052
  );


  nand
  g1514
  (
    n1580,
    n1074,
    n1057,
    n1219,
    n1414
  );


  nand
  g1515
  (
    n1573,
    n1077,
    n1059,
    n1531,
    n1529
  );


  or
  g1516
  (
    n1546,
    n1073,
    n1072,
    n1245,
    n1524
  );


  nand
  g1517
  (
    n1558,
    n1219,
    n1054,
    n1533,
    n1530
  );


  xnor
  g1518
  (
    n1581,
    n1519,
    n1054,
    n1529,
    n1218
  );


  xor
  g1519
  (
    n1542,
    n1462,
    n1077,
    n1530,
    n1522
  );


  xor
  g1520
  (
    n1545,
    n1527,
    n1245,
    n1060,
    n1521
  );


  nor
  g1521
  (
    n1565,
    n1443,
    n1056,
    n1053,
    n1532
  );


  xnor
  g1522
  (
    n1540,
    n1535,
    n1535,
    n1459,
    n1455
  );


  or
  g1523
  (
    n1576,
    n1061,
    n1073,
    n1066,
    n1055
  );


  nor
  g1524
  (
    n1632,
    n1551,
    n1580,
    n673,
    n1577
  );


  nand
  g1525
  (
    n1666,
    n1563,
    n761,
    n680,
    n669
  );


  or
  g1526
  (
    n1620,
    n924,
    n778,
    n913,
    n857
  );


  nor
  g1527
  (
    n1594,
    n928,
    n756,
    n659,
    n884
  );


  xnor
  g1528
  (
    n1674,
    n832,
    n1547,
    n935,
    n929
  );


  and
  g1529
  (
    n1669,
    n840,
    n1573,
    n805,
    n1569
  );


  or
  g1530
  (
    n1658,
    n765,
    n793,
    n1576,
    n957
  );


  or
  g1531
  (
    n1608,
    n1579,
    n727,
    n1573,
    n743
  );


  and
  g1532
  (
    n1642,
    n1562,
    n949,
    n912,
    n871
  );


  and
  g1533
  (
    n1614,
    n767,
    n876,
    n730,
    n917
  );


  or
  g1534
  (
    n1659,
    n1559,
    n804,
    n1548,
    n702
  );


  or
  g1535
  (
    n1675,
    n844,
    n802,
    n1583,
    n916
  );


  and
  g1536
  (
    n1671,
    n1560,
    n1563,
    n1552,
    n867
  );


  and
  g1537
  (
    n1661,
    n794,
    n1539,
    n1569,
    n810
  );


  and
  g1538
  (
    n1681,
    n724,
    n1550,
    n751,
    n654
  );


  and
  g1539
  (
    n1588,
    n695,
    n1578,
    n839,
    n879
  );


  xnor
  g1540
  (
    n1627,
    n915,
    n656,
    n704,
    n1570
  );


  or
  g1541
  (
    n1663,
    n1554,
    n758,
    n1557,
    n1565
  );


  xor
  g1542
  (
    n1616,
    n954,
    n849,
    n880,
    n1545
  );


  xor
  g1543
  (
    n1684,
    n734,
    n864,
    n1577,
    n783
  );


  or
  g1544
  (
    n1667,
    n684,
    n1575,
    n1581,
    n790
  );


  and
  g1545
  (
    n1672,
    n759,
    n862,
    n747,
    n1574
  );


  nand
  g1546
  (
    n1634,
    n723,
    n1580,
    n1564,
    n1558
  );


  nand
  g1547
  (
    n1613,
    n814,
    n1549,
    n722,
    n893
  );


  xnor
  g1548
  (
    n1662,
    n947,
    n786,
    n655,
    n908
  );


  and
  g1549
  (
    n1585,
    n930,
    n887,
    n665,
    n803
  );


  and
  g1550
  (
    n1603,
    n815,
    n686,
    n666,
    n760
  );


  nor
  g1551
  (
    n1595,
    n869,
    n1543,
    n670,
    n657
  );


  xor
  g1552
  (
    n1601,
    n755,
    n881,
    n818,
    n773
  );


  xnor
  g1553
  (
    n1646,
    n796,
    n919,
    n827,
    n720
  );


  and
  g1554
  (
    n1618,
    n874,
    n945,
    n901,
    n1549
  );


  and
  g1555
  (
    n1677,
    n714,
    n865,
    n835,
    n750
  );


  nor
  g1556
  (
    n1640,
    n948,
    n774,
    n737,
    n719
  );


  and
  g1557
  (
    n1647,
    n1554,
    n958,
    n1561,
    n795
  );


  xor
  g1558
  (
    n1617,
    n944,
    n822,
    n784,
    n1582
  );


  nand
  g1559
  (
    n1685,
    n1546,
    n733,
    n1571,
    n781
  );


  xnor
  g1560
  (
    KeyWire_0_21,
    n863,
    n956,
    n850,
    n892
  );


  or
  g1561
  (
    n1605,
    n927,
    n757,
    n1548,
    n1557
  );


  or
  g1562
  (
    n1637,
    n726,
    n661,
    n891,
    n672
  );


  xnor
  g1563
  (
    n1679,
    n1550,
    n922,
    n698,
    n894
  );


  and
  g1564
  (
    n1660,
    n1582,
    n817,
    n842,
    n691
  );


  nor
  g1565
  (
    n1643,
    n667,
    n914,
    n699,
    n819
  );


  nand
  g1566
  (
    n1644,
    n888,
    n709,
    n951,
    n946
  );


  nand
  g1567
  (
    n1651,
    n838,
    n687,
    n1553,
    n889
  );


  and
  g1568
  (
    n1604,
    n713,
    n668,
    n799,
    n693
  );


  xor
  g1569
  (
    n1606,
    n921,
    n937,
    n748,
    n735
  );


  xor
  g1570
  (
    n1628,
    n675,
    n703,
    n739,
    n885
  );


  nand
  g1571
  (
    n1615,
    n866,
    n843,
    n1572,
    n658
  );


  and
  g1572
  (
    n1612,
    n1567,
    n1571,
    n872,
    n768
  );


  xor
  g1573
  (
    n1611,
    n728,
    n825,
    n725,
    n955
  );


  and
  g1574
  (
    n1623,
    n782,
    n1568,
    n707,
    n676
  );


  nor
  g1575
  (
    n1610,
    n746,
    n1541,
    n834,
    n706
  );


  nand
  g1576
  (
    n1591,
    n854,
    n823,
    n700,
    n877
  );


  xor
  g1577
  (
    n1597,
    n1543,
    n950,
    n859,
    n1582
  );


  nor
  g1578
  (
    n1590,
    n800,
    n736,
    n738,
    n1552
  );


  nor
  g1579
  (
    n1589,
    n1564,
    n1537,
    n712,
    n808
  );


  xnor
  g1580
  (
    n1635,
    n816,
    n780,
    n868,
    n1581
  );


  nor
  g1581
  (
    n1584,
    n1541,
    n788,
    n682,
    n1566
  );


  xnor
  g1582
  (
    n1586,
    n688,
    n932,
    n903,
    n811
  );


  nand
  g1583
  (
    n1607,
    n1542,
    n741,
    n846,
    n813
  );


  or
  g1584
  (
    n1592,
    n787,
    n1581,
    n911,
    n1562
  );


  nor
  g1585
  (
    n1596,
    n1578,
    n762,
    n775,
    n764
  );


  nand
  g1586
  (
    n1622,
    n1555,
    n807,
    n1537,
    n685
  );


  or
  g1587
  (
    n1680,
    n1547,
    n754,
    n1555,
    n926
  );


  and
  g1588
  (
    n1593,
    n934,
    n1568,
    n898,
    n836
  );


  or
  g1589
  (
    n1636,
    n671,
    n749,
    n940,
    n753
  );


  and
  g1590
  (
    n1670,
    n1582,
    n847,
    n718,
    n890
  );


  nand
  g1591
  (
    n1602,
    n900,
    n705,
    n824,
    n1572
  );


  nand
  g1592
  (
    n1676,
    n772,
    n769,
    n1581,
    n886
  );


  and
  g1593
  (
    n1625,
    n1583,
    n831,
    n906,
    n697
  );


  and
  g1594
  (
    n1599,
    n660,
    n896,
    n777,
    n883
  );


  xor
  g1595
  (
    n1648,
    n902,
    n875,
    n763,
    n1576
  );


  and
  g1596
  (
    n1657,
    n841,
    n745,
    n820,
    n662
  );


  or
  g1597
  (
    n1621,
    n1566,
    n853,
    n806,
    n740
  );


  nand
  g1598
  (
    KeyWire_0_5,
    n1583,
    n941,
    n1561,
    n785
  );


  nand
  g1599
  (
    n1630,
    n674,
    n1556,
    n1575,
    n766
  );


  or
  g1600
  (
    n1600,
    n920,
    n959,
    n791,
    n731
  );


  nand
  g1601
  (
    n1638,
    n861,
    n708,
    n721,
    n716
  );


  nand
  g1602
  (
    n1649,
    n694,
    n858,
    n936,
    n1538
  );


  nor
  g1603
  (
    n1633,
    n1545,
    n677,
    n878,
    n1538
  );


  nor
  g1604
  (
    n1587,
    n789,
    n678,
    n1536,
    n1544
  );


  nor
  g1605
  (
    n1653,
    n907,
    n942,
    n770,
    n870
  );


  xnor
  g1606
  (
    n1598,
    n939,
    n1553,
    n829,
    n1570
  );


  xor
  g1607
  (
    n1673,
    n692,
    n953,
    n873,
    n821
  );


  xnor
  g1608
  (
    n1650,
    n1574,
    n717,
    n715,
    n812
  );


  xnor
  g1609
  (
    n1619,
    n1579,
    n848,
    n1542,
    n679
  );


  and
  g1610
  (
    n1678,
    n744,
    n1560,
    n797,
    n1556
  );


  nand
  g1611
  (
    KeyWire_0_45,
    n904,
    n742,
    n683,
    n899
  );


  nor
  g1612
  (
    n1645,
    n711,
    n1567,
    n855,
    n845
  );


  nor
  g1613
  (
    n1641,
    n923,
    n938,
    n895,
    n1539
  );


  and
  g1614
  (
    n1652,
    n809,
    n1540,
    n1559,
    n1551
  );


  nand
  g1615
  (
    n1629,
    n689,
    n931,
    n779,
    n696
  );


  nand
  g1616
  (
    n1683,
    n1536,
    n952,
    n856,
    n828
  );


  nand
  g1617
  (
    n1668,
    n909,
    n830,
    n798,
    n1540
  );


  xor
  g1618
  (
    n1626,
    n1558,
    n826,
    n664,
    n943
  );


  nor
  g1619
  (
    n1682,
    n771,
    n833,
    n897,
    n851
  );


  and
  g1620
  (
    n1655,
    n1565,
    n752,
    n882,
    n792
  );


  nand
  g1621
  (
    n1665,
    n905,
    n933,
    n1544,
    n860
  );


  xor
  g1622
  (
    n1654,
    n852,
    n837,
    n729,
    n701
  );


  or
  g1623
  (
    n1664,
    n1546,
    n732,
    n801,
    n681
  );


  and
  g1624
  (
    n1631,
    n710,
    n910,
    n925,
    n1583
  );


  xor
  g1625
  (
    n1609,
    n690,
    n663,
    n776,
    n918
  );


  nand
  g1626
  (
    n1686,
    n1624,
    n1622,
    n1588,
    n1605
  );


  nand
  g1627
  (
    n1696,
    n1610,
    n1620,
    n1596,
    n1589
  );


  xnor
  g1628
  (
    n1697,
    n1632,
    n1630,
    n1614,
    n1617
  );


  xnor
  g1629
  (
    n1693,
    n1635,
    n1602,
    n1611,
    n1612
  );


  nor
  g1630
  (
    n1688,
    n1609,
    n1629,
    n1625,
    n1606
  );


  xnor
  g1631
  (
    KeyWire_0_34,
    n1627,
    n1598,
    n1615,
    n1616
  );


  nor
  g1632
  (
    n1694,
    n1628,
    n1590,
    n1618,
    n1599
  );


  xnor
  g1633
  (
    n1692,
    n1585,
    n1607,
    n1586,
    n1631
  );


  nand
  g1634
  (
    n1687,
    n1595,
    n1600,
    n1597,
    n1587
  );


  nand
  g1635
  (
    n1690,
    n1626,
    n1619,
    n1604,
    n1584
  );


  xnor
  g1636
  (
    n1689,
    n1613,
    n1608,
    n1592,
    n1591
  );


  and
  g1637
  (
    n1698,
    n1633,
    n1621,
    n1634,
    n1623
  );


  and
  g1638
  (
    n1691,
    n1593,
    n1594,
    n1601,
    n1603
  );


  nor
  g1639
  (
    n1699,
    n1698,
    n1637,
    n1636,
    n1638
  );


  nor
  g1640
  (
    n1703,
    n1640,
    n1641,
    n1650,
    n1699
  );


  xnor
  g1641
  (
    n1700,
    n1649,
    n1648,
    n1646,
    n1647
  );


  or
  g1642
  (
    n1701,
    n1645,
    n1639,
    n1699,
    n1644
  );


  xor
  g1643
  (
    n1702,
    n1699,
    n1699,
    n1643,
    n1642
  );


  xor
  g1644
  (
    n1711,
    n1657,
    n1651,
    n1445,
    n1661
  );


  or
  g1645
  (
    KeyWire_0_59,
    n1656,
    n1703,
    n1664,
    n1655
  );


  xor
  g1646
  (
    n1714,
    n1658,
    n1676,
    n1445,
    n1665
  );


  xor
  g1647
  (
    n1718,
    n1666,
    n1122,
    n1702,
    n1444
  );


  xor
  g1648
  (
    n1715,
    n1701,
    n1702,
    n1674,
    n1092
  );


  nor
  g1649
  (
    n1717,
    n1703,
    n1672,
    n1671,
    n250
  );


  or
  g1650
  (
    n1707,
    n1702,
    n1444,
    n1703,
    n1700
  );


  or
  g1651
  (
    n1710,
    n1662,
    n1675,
    n1673,
    n1670
  );


  nand
  g1652
  (
    n1706,
    n1660,
    n1445,
    n1701,
    n1669
  );


  nor
  g1653
  (
    n1712,
    n1652,
    n1092,
    n1703,
    n1093
  );


  nor
  g1654
  (
    n1719,
    n1700,
    n1654,
    n1701,
    n1092
  );


  xnor
  g1655
  (
    n1705,
    n1679,
    n1667,
    n1122,
    n1659
  );


  nand
  g1656
  (
    n1704,
    n1444,
    n1445,
    n1653,
    n1093
  );


  xor
  g1657
  (
    n1713,
    n1663,
    n1092,
    n1700,
    n1678
  );


  nand
  g1658
  (
    n1708,
    n1093,
    n1702,
    n1121,
    n1701
  );


  xor
  g1659
  (
    n1716,
    n1700,
    n1093,
    n1677,
    n1668
  );


  nand
  g1660
  (
    n1722,
    n1717,
    n1719,
    n1715
  );


  and
  g1661
  (
    n1727,
    n1717,
    n1714,
    n1718,
    n1705
  );


  xnor
  g1662
  (
    n1724,
    n1708,
    n1717,
    n1719
  );


  and
  g1663
  (
    n1723,
    n1714,
    n1718,
    n1716,
    n1683
  );


  nor
  g1664
  (
    n1720,
    n1716,
    n1712,
    n1704,
    n1713
  );


  xor
  g1665
  (
    n1726,
    n1685,
    n1707,
    n1714
  );


  xor
  g1666
  (
    n1721,
    n1684,
    n1682,
    n1715,
    n1710
  );


  nor
  g1667
  (
    n1725,
    n1715,
    n1716,
    n1718,
    n1711
  );


  xor
  g1668
  (
    n1728,
    n1716,
    n1717,
    n1718,
    n1709
  );


  and
  g1669
  (
    n1729,
    n1706,
    n1719,
    n1680,
    n1681
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1534,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n635,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1160,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n294,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n618,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n1624,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1110,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1172,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1470,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n75,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n963,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n78,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1574,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1031,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1275,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n925,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n188,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n476,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n519,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n120,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1290,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1656,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1309,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n907,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1011,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1132,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n504,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1000,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n259,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1352,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n610,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n442,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n60,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n1459,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n1695,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n1270,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n795,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n1423,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n959,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n370,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n330,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n470,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n811,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n92,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n935,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n1639,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n1455,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n1318,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n89,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n372,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n803,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n1466,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n1166,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n637,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n67,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n727,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n308,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n119,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n1261,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n1709,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n480,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n1473,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n354,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n912,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


