

module Stat_3000_323
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1385,
  n1389,
  n1396,
  n1409,
  n3023,
  n3026,
  n3021,
  n3032,
  n3019,
  n3031,
  n3020,
  n3017,
  n3025,
  n3012,
  n3013,
  n3011,
  n3015,
  n3027,
  n3018,
  n3030,
  n3029,
  n3008,
  n3022,
  n3009,
  n3028,
  n3005,
  n3010,
  n3024,
  n3016,
  n3014,
  n3006,
  n3007
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1385;output n1389;output n1396;output n1409;output n3023;output n3026;output n3021;output n3032;output n3019;output n3031;output n3020;output n3017;output n3025;output n3012;output n3013;output n3011;output n3015;output n3027;output n3018;output n3030;output n3029;output n3008;output n3022;output n3009;output n3028;output n3005;output n3010;output n3024;output n3016;output n3014;output n3006;output n3007;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1386;wire n1387;wire n1388;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n50,
    n3
  );


  buf
  g1
  (
    n39,
    n1
  );


  not
  g2
  (
    n40,
    n4
  );


  buf
  g3
  (
    n41,
    n1
  );


  not
  g4
  (
    n43,
    n3
  );


  not
  g5
  (
    n33,
    n2
  );


  buf
  g6
  (
    n37,
    n4
  );


  buf
  g7
  (
    n38,
    n2
  );


  not
  g8
  (
    n36,
    n5
  );


  not
  g9
  (
    n47,
    n4
  );


  buf
  g10
  (
    n48,
    n2
  );


  buf
  g11
  (
    n49,
    n2
  );


  buf
  g12
  (
    n34,
    n3
  );


  buf
  g13
  (
    n45,
    n5
  );


  not
  g14
  (
    n42,
    n1
  );


  buf
  g15
  (
    n44,
    n3
  );


  not
  g16
  (
    n46,
    n1
  );


  not
  g17
  (
    n35,
    n4
  );


  not
  g18
  (
    n79,
    n33
  );


  buf
  g19
  (
    n55,
    n46
  );


  not
  g20
  (
    n86,
    n39
  );


  not
  g21
  (
    n101,
    n45
  );


  not
  g22
  (
    KeyWire_0_30,
    n35
  );


  buf
  g23
  (
    n109,
    n47
  );


  buf
  g24
  (
    n65,
    n43
  );


  buf
  g25
  (
    n63,
    n44
  );


  buf
  g26
  (
    n56,
    n40
  );


  buf
  g27
  (
    n60,
    n34
  );


  buf
  g28
  (
    n66,
    n44
  );


  buf
  g29
  (
    n91,
    n38
  );


  buf
  g30
  (
    n104,
    n40
  );


  buf
  g31
  (
    n98,
    n45
  );


  buf
  g32
  (
    n88,
    n35
  );


  buf
  g33
  (
    n97,
    n46
  );


  buf
  g34
  (
    n95,
    n43
  );


  not
  g35
  (
    n96,
    n40
  );


  buf
  g36
  (
    n71,
    n38
  );


  not
  g37
  (
    n58,
    n43
  );


  buf
  g38
  (
    n80,
    n37
  );


  not
  g39
  (
    n73,
    n33
  );


  buf
  g40
  (
    n52,
    n41
  );


  not
  g41
  (
    n64,
    n42
  );


  buf
  g42
  (
    n84,
    n42
  );


  buf
  g43
  (
    n54,
    n42
  );


  not
  g44
  (
    n87,
    n33
  );


  buf
  g45
  (
    n107,
    n35
  );


  buf
  g46
  (
    n59,
    n34
  );


  not
  g47
  (
    n99,
    n44
  );


  not
  g48
  (
    n67,
    n46
  );


  not
  g49
  (
    n57,
    n42
  );


  not
  g50
  (
    n77,
    n36
  );


  not
  g51
  (
    n68,
    n38
  );


  not
  g52
  (
    n69,
    n47
  );


  buf
  g53
  (
    n89,
    n34
  );


  not
  g54
  (
    n81,
    n37
  );


  buf
  g55
  (
    n106,
    n43
  );


  buf
  g56
  (
    n53,
    n34
  );


  not
  g57
  (
    n72,
    n35
  );


  buf
  g58
  (
    n83,
    n37
  );


  not
  g59
  (
    n92,
    n46
  );


  buf
  g60
  (
    n105,
    n38
  );


  not
  g61
  (
    n103,
    n39
  );


  buf
  g62
  (
    n76,
    n44
  );


  buf
  g63
  (
    KeyWire_0_21,
    n33
  );


  not
  g64
  (
    n51,
    n37
  );


  not
  g65
  (
    n85,
    n41
  );


  buf
  g66
  (
    n75,
    n36
  );


  not
  g67
  (
    n102,
    n41
  );


  buf
  g68
  (
    n78,
    n40
  );


  not
  g69
  (
    n74,
    n45
  );


  not
  g70
  (
    n62,
    n39
  );


  not
  g71
  (
    n70,
    n36
  );


  not
  g72
  (
    n61,
    n36
  );


  not
  g73
  (
    n93,
    n41
  );


  not
  g74
  (
    n108,
    n45
  );


  not
  g75
  (
    n100,
    n47
  );


  not
  g76
  (
    n82,
    n39
  );


  buf
  g77
  (
    n145,
    n100
  );


  buf
  g78
  (
    n271,
    n81
  );


  not
  g79
  (
    n319,
    n63
  );


  not
  g80
  (
    n128,
    n87
  );


  buf
  g81
  (
    n321,
    n88
  );


  not
  g82
  (
    n167,
    n91
  );


  not
  g83
  (
    n229,
    n99
  );


  not
  g84
  (
    n154,
    n80
  );


  not
  g85
  (
    n205,
    n51
  );


  not
  g86
  (
    n182,
    n66
  );


  buf
  g87
  (
    n270,
    n93
  );


  buf
  g88
  (
    n156,
    n81
  );


  not
  g89
  (
    n215,
    n79
  );


  buf
  g90
  (
    n155,
    n97
  );


  not
  g91
  (
    n313,
    n56
  );


  buf
  g92
  (
    n117,
    n68
  );


  buf
  g93
  (
    n115,
    n56
  );


  buf
  g94
  (
    n111,
    n94
  );


  not
  g95
  (
    n246,
    n93
  );


  not
  g96
  (
    n317,
    n55
  );


  buf
  g97
  (
    n259,
    n86
  );


  buf
  g98
  (
    n293,
    n66
  );


  not
  g99
  (
    n204,
    n76
  );


  not
  g100
  (
    n170,
    n65
  );


  not
  g101
  (
    n168,
    n60
  );


  buf
  g102
  (
    n119,
    n54
  );


  not
  g103
  (
    n203,
    n92
  );


  buf
  g104
  (
    n193,
    n68
  );


  not
  g105
  (
    n227,
    n62
  );


  buf
  g106
  (
    n110,
    n63
  );


  buf
  g107
  (
    n242,
    n78
  );


  not
  g108
  (
    n268,
    n53
  );


  buf
  g109
  (
    n276,
    n100
  );


  not
  g110
  (
    n300,
    n95
  );


  buf
  g111
  (
    n269,
    n75
  );


  buf
  g112
  (
    n261,
    n84
  );


  not
  g113
  (
    n149,
    n94
  );


  not
  g114
  (
    n264,
    n90
  );


  buf
  g115
  (
    n189,
    n92
  );


  not
  g116
  (
    n281,
    n58
  );


  buf
  g117
  (
    n161,
    n61
  );


  buf
  g118
  (
    n134,
    n52
  );


  buf
  g119
  (
    n152,
    n70
  );


  buf
  g120
  (
    n195,
    n77
  );


  buf
  g121
  (
    n263,
    n74
  );


  buf
  g122
  (
    n310,
    n96
  );


  not
  g123
  (
    n126,
    n57
  );


  not
  g124
  (
    n158,
    n89
  );


  not
  g125
  (
    n290,
    n88
  );


  buf
  g126
  (
    n160,
    n69
  );


  buf
  g127
  (
    n234,
    n67
  );


  not
  g128
  (
    n295,
    n67
  );


  not
  g129
  (
    n179,
    n94
  );


  not
  g130
  (
    n129,
    n100
  );


  not
  g131
  (
    n267,
    n61
  );


  buf
  g132
  (
    n207,
    n90
  );


  not
  g133
  (
    n210,
    n55
  );


  not
  g134
  (
    n162,
    n57
  );


  buf
  g135
  (
    n188,
    n51
  );


  not
  g136
  (
    n127,
    n71
  );


  buf
  g137
  (
    n202,
    n61
  );


  buf
  g138
  (
    n151,
    n103
  );


  buf
  g139
  (
    n125,
    n69
  );


  not
  g140
  (
    n164,
    n83
  );


  buf
  g141
  (
    n294,
    n74
  );


  buf
  g142
  (
    n185,
    n54
  );


  not
  g143
  (
    n196,
    n103
  );


  buf
  g144
  (
    n183,
    n91
  );


  buf
  g145
  (
    n216,
    n83
  );


  not
  g146
  (
    n273,
    n76
  );


  buf
  g147
  (
    n178,
    n62
  );


  buf
  g148
  (
    n201,
    n79
  );


  buf
  g149
  (
    n173,
    n71
  );


  not
  g150
  (
    n275,
    n69
  );


  not
  g151
  (
    n212,
    n67
  );


  buf
  g152
  (
    n116,
    n69
  );


  not
  g153
  (
    n312,
    n101
  );


  buf
  g154
  (
    n118,
    n71
  );


  buf
  g155
  (
    n133,
    n80
  );


  buf
  g156
  (
    n251,
    n59
  );


  buf
  g157
  (
    n181,
    n78
  );


  not
  g158
  (
    n279,
    n64
  );


  not
  g159
  (
    n309,
    n73
  );


  not
  g160
  (
    n320,
    n72
  );


  not
  g161
  (
    n296,
    n91
  );


  not
  g162
  (
    n304,
    n98
  );


  not
  g163
  (
    n228,
    n81
  );


  not
  g164
  (
    n175,
    n99
  );


  buf
  g165
  (
    n123,
    n83
  );


  not
  g166
  (
    n214,
    n75
  );


  not
  g167
  (
    n138,
    n96
  );


  buf
  g168
  (
    n274,
    n97
  );


  buf
  g169
  (
    n157,
    n78
  );


  buf
  g170
  (
    n256,
    n77
  );


  not
  g171
  (
    n282,
    n57
  );


  not
  g172
  (
    n131,
    n65
  );


  buf
  g173
  (
    n209,
    n60
  );


  not
  g174
  (
    n236,
    n70
  );


  not
  g175
  (
    n114,
    n77
  );


  buf
  g176
  (
    n143,
    n75
  );


  buf
  g177
  (
    n146,
    n75
  );


  buf
  g178
  (
    n198,
    n91
  );


  buf
  g179
  (
    n140,
    n89
  );


  buf
  g180
  (
    n262,
    n56
  );


  not
  g181
  (
    n253,
    n53
  );


  buf
  g182
  (
    n306,
    n58
  );


  buf
  g183
  (
    n187,
    n76
  );


  buf
  g184
  (
    n177,
    n62
  );


  not
  g185
  (
    n169,
    n60
  );


  not
  g186
  (
    n283,
    n59
  );


  buf
  g187
  (
    n277,
    n70
  );


  not
  g188
  (
    n255,
    n87
  );


  buf
  g189
  (
    n112,
    n87
  );


  not
  g190
  (
    n221,
    n73
  );


  buf
  g191
  (
    n147,
    n102
  );


  buf
  g192
  (
    n244,
    n66
  );


  not
  g193
  (
    n176,
    n58
  );


  not
  g194
  (
    n284,
    n56
  );


  buf
  g195
  (
    n199,
    n90
  );


  not
  g196
  (
    n250,
    n55
  );


  not
  g197
  (
    n314,
    n53
  );


  buf
  g198
  (
    n297,
    n104
  );


  buf
  g199
  (
    n248,
    n102
  );


  buf
  g200
  (
    n211,
    n86
  );


  buf
  g201
  (
    n219,
    n52
  );


  buf
  g202
  (
    n184,
    n76
  );


  not
  g203
  (
    n142,
    n80
  );


  buf
  g204
  (
    n258,
    n67
  );


  not
  g205
  (
    n289,
    n95
  );


  not
  g206
  (
    n141,
    n58
  );


  buf
  g207
  (
    n163,
    n85
  );


  not
  g208
  (
    n322,
    n73
  );


  not
  g209
  (
    n132,
    n90
  );


  buf
  g210
  (
    n136,
    n53
  );


  not
  g211
  (
    n315,
    n103
  );


  buf
  g212
  (
    n311,
    n83
  );


  not
  g213
  (
    n124,
    n68
  );


  buf
  g214
  (
    n298,
    n64
  );


  not
  g215
  (
    n278,
    n84
  );


  buf
  g216
  (
    n324,
    n84
  );


  not
  g217
  (
    n208,
    n97
  );


  buf
  g218
  (
    n252,
    n59
  );


  not
  g219
  (
    n220,
    n96
  );


  buf
  g220
  (
    n194,
    n87
  );


  buf
  g221
  (
    n240,
    n94
  );


  not
  g222
  (
    n260,
    n104
  );


  not
  g223
  (
    n222,
    n95
  );


  buf
  g224
  (
    n245,
    n101
  );


  buf
  g225
  (
    n192,
    n70
  );


  not
  g226
  (
    n121,
    n98
  );


  not
  g227
  (
    n218,
    n68
  );


  buf
  g228
  (
    n303,
    n64
  );


  buf
  g229
  (
    n257,
    n93
  );


  not
  g230
  (
    n265,
    n98
  );


  buf
  g231
  (
    n206,
    n82
  );


  not
  g232
  (
    n190,
    n72
  );


  not
  g233
  (
    n225,
    n85
  );


  buf
  g234
  (
    n287,
    n51
  );


  not
  g235
  (
    n280,
    n99
  );


  buf
  g236
  (
    n137,
    n86
  );


  buf
  g237
  (
    n318,
    n61
  );


  not
  g238
  (
    n135,
    n72
  );


  buf
  g239
  (
    n230,
    n60
  );


  not
  g240
  (
    n166,
    n51
  );


  buf
  g241
  (
    n139,
    n55
  );


  buf
  g242
  (
    n226,
    n54
  );


  buf
  g243
  (
    n307,
    n100
  );


  not
  g244
  (
    n299,
    n72
  );


  buf
  g245
  (
    n316,
    n79
  );


  not
  g246
  (
    n171,
    n98
  );


  buf
  g247
  (
    n191,
    n71
  );


  buf
  g248
  (
    n197,
    n63
  );


  not
  g249
  (
    n217,
    n85
  );


  not
  g250
  (
    n302,
    n101
  );


  buf
  g251
  (
    n122,
    n74
  );


  not
  g252
  (
    n301,
    n73
  );


  not
  g253
  (
    n180,
    n79
  );


  not
  g254
  (
    n285,
    n88
  );


  buf
  g255
  (
    n231,
    n77
  );


  buf
  g256
  (
    n286,
    n81
  );


  buf
  g257
  (
    n150,
    n66
  );


  not
  g258
  (
    n144,
    n52
  );


  buf
  g259
  (
    n200,
    n102
  );


  buf
  g260
  (
    n305,
    n96
  );


  buf
  g261
  (
    n148,
    n82
  );


  buf
  g262
  (
    n254,
    n89
  );


  buf
  g263
  (
    n223,
    n85
  );


  buf
  g264
  (
    n174,
    n84
  );


  not
  g265
  (
    n249,
    n57
  );


  not
  g266
  (
    n292,
    n88
  );


  not
  g267
  (
    n241,
    n102
  );


  buf
  g268
  (
    n224,
    n99
  );


  buf
  g269
  (
    n247,
    n65
  );


  not
  g270
  (
    n266,
    n63
  );


  not
  g271
  (
    n172,
    n89
  );


  buf
  g272
  (
    n165,
    n78
  );


  not
  g273
  (
    n239,
    n82
  );


  buf
  g274
  (
    n243,
    n92
  );


  not
  g275
  (
    n291,
    n92
  );


  buf
  g276
  (
    n237,
    n59
  );


  not
  g277
  (
    n272,
    n62
  );


  buf
  g278
  (
    n288,
    n64
  );


  not
  g279
  (
    n153,
    n93
  );


  buf
  g280
  (
    n113,
    n101
  );


  buf
  g281
  (
    n159,
    n82
  );


  not
  g282
  (
    n130,
    n80
  );


  buf
  g283
  (
    n186,
    n52
  );


  buf
  g284
  (
    n233,
    n54
  );


  buf
  g285
  (
    n120,
    n104
  );


  buf
  g286
  (
    n238,
    n95
  );


  not
  g287
  (
    n232,
    n86
  );


  not
  g288
  (
    n213,
    n65
  );


  buf
  g289
  (
    n235,
    n97
  );


  not
  g290
  (
    n308,
    n74
  );


  buf
  g291
  (
    n323,
    n103
  );


  buf
  g292
  (
    n987,
    n258
  );


  not
  g293
  (
    n857,
    n148
  );


  buf
  g294
  (
    n365,
    n264
  );


  not
  g295
  (
    n679,
    n227
  );


  buf
  g296
  (
    n789,
    n194
  );


  not
  g297
  (
    n1069,
    n238
  );


  not
  g298
  (
    n1091,
    n114
  );


  not
  g299
  (
    n708,
    n182
  );


  buf
  g300
  (
    n573,
    n254
  );


  not
  g301
  (
    n681,
    n115
  );


  buf
  g302
  (
    n938,
    n151
  );


  not
  g303
  (
    n1119,
    n253
  );


  not
  g304
  (
    n771,
    n141
  );


  buf
  g305
  (
    n1080,
    n224
  );


  buf
  g306
  (
    n610,
    n180
  );


  not
  g307
  (
    n329,
    n136
  );


  buf
  g308
  (
    n1099,
    n260
  );


  buf
  g309
  (
    n812,
    n271
  );


  not
  g310
  (
    n492,
    n111
  );


  not
  g311
  (
    n523,
    n132
  );


  buf
  g312
  (
    n747,
    n171
  );


  not
  g313
  (
    n1117,
    n245
  );


  buf
  g314
  (
    n645,
    n165
  );


  not
  g315
  (
    n803,
    n235
  );


  buf
  g316
  (
    n452,
    n152
  );


  not
  g317
  (
    n764,
    n196
  );


  not
  g318
  (
    n1038,
    n248
  );


  not
  g319
  (
    n893,
    n162
  );


  buf
  g320
  (
    n548,
    n255
  );


  buf
  g321
  (
    n728,
    n203
  );


  buf
  g322
  (
    n382,
    n196
  );


  not
  g323
  (
    n1071,
    n307
  );


  not
  g324
  (
    n744,
    n142
  );


  not
  g325
  (
    n560,
    n316
  );


  buf
  g326
  (
    n528,
    n203
  );


  buf
  g327
  (
    n609,
    n114
  );


  buf
  g328
  (
    n978,
    n170
  );


  not
  g329
  (
    n831,
    n303
  );


  buf
  g330
  (
    n828,
    n176
  );


  buf
  g331
  (
    n1097,
    n187
  );


  not
  g332
  (
    n886,
    n131
  );


  buf
  g333
  (
    n643,
    n258
  );


  not
  g334
  (
    n897,
    n147
  );


  buf
  g335
  (
    n863,
    n298
  );


  buf
  g336
  (
    n770,
    n303
  );


  buf
  g337
  (
    n758,
    n188
  );


  buf
  g338
  (
    n425,
    n249
  );


  not
  g339
  (
    n468,
    n246
  );


  buf
  g340
  (
    n1116,
    n121
  );


  not
  g341
  (
    n343,
    n314
  );


  buf
  g342
  (
    n570,
    n275
  );


  not
  g343
  (
    n846,
    n159
  );


  not
  g344
  (
    n858,
    n130
  );


  not
  g345
  (
    n980,
    n238
  );


  not
  g346
  (
    n1008,
    n261
  );


  buf
  g347
  (
    n335,
    n229
  );


  not
  g348
  (
    n1017,
    n212
  );


  not
  g349
  (
    n504,
    n188
  );


  not
  g350
  (
    n402,
    n288
  );


  not
  g351
  (
    n1000,
    n220
  );


  not
  g352
  (
    n840,
    n151
  );


  buf
  g353
  (
    n765,
    n225
  );


  buf
  g354
  (
    n508,
    n182
  );


  not
  g355
  (
    n882,
    n266
  );


  buf
  g356
  (
    n493,
    n284
  );


  not
  g357
  (
    n775,
    n211
  );


  buf
  g358
  (
    n383,
    n204
  );


  buf
  g359
  (
    n370,
    n259
  );


  buf
  g360
  (
    n704,
    n170
  );


  not
  g361
  (
    n445,
    n168
  );


  not
  g362
  (
    n843,
    n218
  );


  not
  g363
  (
    n711,
    n193
  );


  not
  g364
  (
    n476,
    n317
  );


  buf
  g365
  (
    n838,
    n276
  );


  not
  g366
  (
    n735,
    n313
  );


  buf
  g367
  (
    n577,
    n188
  );


  not
  g368
  (
    n680,
    n202
  );


  buf
  g369
  (
    n371,
    n306
  );


  buf
  g370
  (
    n340,
    n168
  );


  buf
  g371
  (
    n617,
    n150
  );


  buf
  g372
  (
    n740,
    n191
  );


  not
  g373
  (
    n620,
    n137
  );


  not
  g374
  (
    n1075,
    n264
  );


  not
  g375
  (
    n821,
    n194
  );


  buf
  g376
  (
    n540,
    n208
  );


  buf
  g377
  (
    n1124,
    n174
  );


  buf
  g378
  (
    n602,
    n314
  );


  not
  g379
  (
    n794,
    n270
  );


  not
  g380
  (
    n347,
    n175
  );


  not
  g381
  (
    n443,
    n279
  );


  buf
  g382
  (
    n599,
    n201
  );


  buf
  g383
  (
    n1090,
    n147
  );


  not
  g384
  (
    n860,
    n238
  );


  not
  g385
  (
    n1024,
    n262
  );


  not
  g386
  (
    n554,
    n239
  );


  buf
  g387
  (
    n888,
    n192
  );


  not
  g388
  (
    n687,
    n180
  );


  not
  g389
  (
    n807,
    n234
  );


  buf
  g390
  (
    n885,
    n239
  );


  buf
  g391
  (
    n727,
    n125
  );


  buf
  g392
  (
    n1077,
    n138
  );


  not
  g393
  (
    n428,
    n225
  );


  buf
  g394
  (
    n899,
    n224
  );


  not
  g395
  (
    n342,
    n128
  );


  buf
  g396
  (
    n692,
    n308
  );


  not
  g397
  (
    n559,
    n204
  );


  not
  g398
  (
    n480,
    n237
  );


  not
  g399
  (
    n429,
    n115
  );


  not
  g400
  (
    n1003,
    n144
  );


  buf
  g401
  (
    n346,
    n304
  );


  buf
  g402
  (
    n1112,
    n142
  );


  not
  g403
  (
    n652,
    n273
  );


  not
  g404
  (
    n798,
    n253
  );


  buf
  g405
  (
    n940,
    n135
  );


  not
  g406
  (
    n823,
    n180
  );


  buf
  g407
  (
    n379,
    n259
  );


  buf
  g408
  (
    n677,
    n199
  );


  not
  g409
  (
    n1126,
    n126
  );


  buf
  g410
  (
    n816,
    n135
  );


  not
  g411
  (
    n871,
    n309
  );


  not
  g412
  (
    n1009,
    n302
  );


  not
  g413
  (
    n1131,
    n155
  );


  buf
  g414
  (
    n802,
    n251
  );


  not
  g415
  (
    n942,
    n191
  );


  not
  g416
  (
    n376,
    n296
  );


  buf
  g417
  (
    n1025,
    n128
  );


  not
  g418
  (
    n563,
    n237
  );


  not
  g419
  (
    n826,
    n218
  );


  buf
  g420
  (
    n939,
    n149
  );


  buf
  g421
  (
    n759,
    n211
  );


  not
  g422
  (
    n334,
    n240
  );


  buf
  g423
  (
    n467,
    n268
  );


  not
  g424
  (
    n396,
    n228
  );


  buf
  g425
  (
    n353,
    n215
  );


  buf
  g426
  (
    n869,
    n281
  );


  not
  g427
  (
    n776,
    n117
  );


  not
  g428
  (
    n964,
    n262
  );


  not
  g429
  (
    n403,
    n214
  );


  not
  g430
  (
    n588,
    n205
  );


  not
  g431
  (
    n1109,
    n279
  );


  buf
  g432
  (
    n394,
    n138
  );


  not
  g433
  (
    n1026,
    n296
  );


  buf
  g434
  (
    n567,
    n163
  );


  not
  g435
  (
    n1021,
    n256
  );


  not
  g436
  (
    n572,
    n310
  );


  not
  g437
  (
    n1018,
    n171
  );


  not
  g438
  (
    n457,
    n127
  );


  buf
  g439
  (
    n385,
    n177
  );


  not
  g440
  (
    n753,
    n291
  );


  buf
  g441
  (
    n597,
    n138
  );


  buf
  g442
  (
    n736,
    n312
  );


  buf
  g443
  (
    n1065,
    n167
  );


  buf
  g444
  (
    n731,
    n308
  );


  not
  g445
  (
    n539,
    n302
  );


  buf
  g446
  (
    n461,
    n182
  );


  buf
  g447
  (
    n666,
    n291
  );


  not
  g448
  (
    n688,
    n265
  );


  not
  g449
  (
    n739,
    n173
  );


  buf
  g450
  (
    n478,
    n135
  );


  not
  g451
  (
    n1121,
    n162
  );


  buf
  g452
  (
    n985,
    n118
  );


  buf
  g453
  (
    n1039,
    n113
  );


  not
  g454
  (
    n913,
    n164
  );


  buf
  g455
  (
    n326,
    n246
  );


  buf
  g456
  (
    n787,
    n155
  );


  buf
  g457
  (
    n700,
    n242
  );


  not
  g458
  (
    n583,
    n283
  );


  buf
  g459
  (
    n600,
    n223
  );


  not
  g460
  (
    n330,
    n254
  );


  buf
  g461
  (
    n788,
    n272
  );


  not
  g462
  (
    n1006,
    n297
  );


  not
  g463
  (
    n929,
    n185
  );


  not
  g464
  (
    n1015,
    n223
  );


  buf
  g465
  (
    n636,
    n203
  );


  not
  g466
  (
    n702,
    n110
  );


  buf
  g467
  (
    n1114,
    n188
  );


  buf
  g468
  (
    n818,
    n128
  );


  not
  g469
  (
    n780,
    n279
  );


  buf
  g470
  (
    n1082,
    n311
  );


  not
  g471
  (
    n782,
    n300
  );


  not
  g472
  (
    n1036,
    n134
  );


  not
  g473
  (
    n738,
    n206
  );


  buf
  g474
  (
    n797,
    n277
  );


  buf
  g475
  (
    n951,
    n248
  );


  buf
  g476
  (
    n390,
    n196
  );


  buf
  g477
  (
    n1125,
    n126
  );


  not
  g478
  (
    n530,
    n214
  );


  not
  g479
  (
    n533,
    n139
  );


  buf
  g480
  (
    n1047,
    n177
  );


  not
  g481
  (
    n368,
    n201
  );


  buf
  g482
  (
    n1103,
    n292
  );


  buf
  g483
  (
    n1014,
    n292
  );


  buf
  g484
  (
    n432,
    n214
  );


  buf
  g485
  (
    n465,
    n135
  );


  buf
  g486
  (
    n921,
    n293
  );


  not
  g487
  (
    n594,
    n185
  );


  buf
  g488
  (
    n462,
    n157
  );


  buf
  g489
  (
    n667,
    n311
  );


  buf
  g490
  (
    n935,
    n301
  );


  buf
  g491
  (
    n625,
    n279
  );


  buf
  g492
  (
    n1032,
    n216
  );


  not
  g493
  (
    n532,
    n160
  );


  buf
  g494
  (
    n853,
    n119
  );


  not
  g495
  (
    n686,
    n315
  );


  buf
  g496
  (
    n751,
    n287
  );


  buf
  g497
  (
    n348,
    n218
  );


  not
  g498
  (
    n502,
    n316
  );


  buf
  g499
  (
    n380,
    n142
  );


  not
  g500
  (
    n454,
    n204
  );


  not
  g501
  (
    n995,
    n249
  );


  not
  g502
  (
    n580,
    n234
  );


  not
  g503
  (
    n623,
    n210
  );


  not
  g504
  (
    n367,
    n130
  );


  buf
  g505
  (
    n809,
    n205
  );


  buf
  g506
  (
    n829,
    n268
  );


  buf
  g507
  (
    n796,
    n314
  );


  buf
  g508
  (
    n814,
    n131
  );


  buf
  g509
  (
    n579,
    n174
  );


  buf
  g510
  (
    n763,
    n290
  );


  not
  g511
  (
    n962,
    n307
  );


  buf
  g512
  (
    n684,
    n285
  );


  buf
  g513
  (
    n1138,
    n257
  );


  not
  g514
  (
    n416,
    n232
  );


  not
  g515
  (
    n608,
    n252
  );


  buf
  g516
  (
    n949,
    n220
  );


  not
  g517
  (
    n426,
    n241
  );


  not
  g518
  (
    n971,
    n247
  );


  not
  g519
  (
    n908,
    n129
  );


  not
  g520
  (
    n496,
    n158
  );


  buf
  g521
  (
    n477,
    n154
  );


  not
  g522
  (
    n820,
    n277
  );


  not
  g523
  (
    n694,
    n231
  );


  buf
  g524
  (
    n1105,
    n209
  );


  not
  g525
  (
    n344,
    n311
  );


  not
  g526
  (
    n527,
    n119
  );


  buf
  g527
  (
    n466,
    n298
  );


  not
  g528
  (
    n505,
    n161
  );


  not
  g529
  (
    n1133,
    n173
  );


  buf
  g530
  (
    n561,
    n275
  );


  not
  g531
  (
    n552,
    n271
  );


  not
  g532
  (
    n1023,
    n145
  );


  not
  g533
  (
    n892,
    n293
  );


  buf
  g534
  (
    n549,
    n280
  );


  buf
  g535
  (
    n358,
    n300
  );


  not
  g536
  (
    n1108,
    n136
  );


  not
  g537
  (
    n564,
    n286
  );


  not
  g538
  (
    n873,
    n138
  );


  not
  g539
  (
    n659,
    n232
  );


  buf
  g540
  (
    n413,
    n315
  );


  not
  g541
  (
    n363,
    n221
  );


  buf
  g542
  (
    n510,
    n213
  );


  buf
  g543
  (
    n864,
    n186
  );


  buf
  g544
  (
    n515,
    n259
  );


  not
  g545
  (
    n1056,
    n178
  );


  not
  g546
  (
    n1063,
    n161
  );


  buf
  g547
  (
    n841,
    n282
  );


  not
  g548
  (
    n474,
    n112
  );


  buf
  g549
  (
    n656,
    n295
  );


  not
  g550
  (
    n369,
    n197
  );


  not
  g551
  (
    n336,
    n139
  );


  not
  g552
  (
    n868,
    n149
  );


  buf
  g553
  (
    n859,
    n161
  );


  buf
  g554
  (
    n584,
    n286
  );


  buf
  g555
  (
    n745,
    n126
  );


  buf
  g556
  (
    n519,
    n117
  );


  buf
  g557
  (
    n494,
    n287
  );


  buf
  g558
  (
    n958,
    n129
  );


  not
  g559
  (
    n590,
    n171
  );


  not
  g560
  (
    n475,
    n151
  );


  not
  g561
  (
    n722,
    n131
  );


  not
  g562
  (
    n635,
    n119
  );


  buf
  g563
  (
    n619,
    n304
  );


  buf
  g564
  (
    n469,
    n281
  );


  buf
  g565
  (
    n655,
    n280
  );


  not
  g566
  (
    n663,
    n275
  );


  not
  g567
  (
    n726,
    n165
  );


  not
  g568
  (
    n960,
    n166
  );


  not
  g569
  (
    n889,
    n152
  );


  buf
  g570
  (
    n410,
    n197
  );


  not
  g571
  (
    n786,
    n298
  );


  buf
  g572
  (
    n910,
    n183
  );


  buf
  g573
  (
    n488,
    n317
  );


  buf
  g574
  (
    n836,
    n133
  );


  not
  g575
  (
    n989,
    n161
  );


  not
  g576
  (
    n984,
    n141
  );


  buf
  g577
  (
    n337,
    n125
  );


  buf
  g578
  (
    n341,
    n144
  );


  buf
  g579
  (
    n1074,
    n215
  );


  buf
  g580
  (
    n536,
    n226
  );


  not
  g581
  (
    n917,
    n276
  );


  buf
  g582
  (
    n1050,
    n191
  );


  not
  g583
  (
    n1081,
    n245
  );


  buf
  g584
  (
    n698,
    n189
  );


  buf
  g585
  (
    n447,
    n143
  );


  buf
  g586
  (
    n1113,
    n134
  );


  buf
  g587
  (
    n784,
    n273
  );


  not
  g588
  (
    n641,
    n113
  );


  not
  g589
  (
    n947,
    n122
  );


  buf
  g590
  (
    n781,
    n317
  );


  not
  g591
  (
    n723,
    n303
  );


  not
  g592
  (
    n783,
    n230
  );


  not
  g593
  (
    n500,
    n227
  );


  not
  g594
  (
    n934,
    n114
  );


  buf
  g595
  (
    n405,
    n274
  );


  not
  g596
  (
    n1048,
    n251
  );


  buf
  g597
  (
    n997,
    n310
  );


  buf
  g598
  (
    n966,
    n308
  );


  not
  g599
  (
    n999,
    n263
  );


  buf
  g600
  (
    n1052,
    n282
  );


  not
  g601
  (
    n415,
    n139
  );


  not
  g602
  (
    n364,
    n262
  );


  buf
  g603
  (
    n1106,
    n290
  );


  not
  g604
  (
    n695,
    n212
  );


  not
  g605
  (
    n844,
    n283
  );


  buf
  g606
  (
    n664,
    n303
  );


  not
  g607
  (
    n661,
    n196
  );


  not
  g608
  (
    n963,
    n284
  );


  not
  g609
  (
    n430,
    n190
  );


  buf
  g610
  (
    n395,
    n140
  );


  not
  g611
  (
    n1135,
    n121
  );


  buf
  g612
  (
    n785,
    n172
  );


  buf
  g613
  (
    n1051,
    n286
  );


  not
  g614
  (
    n433,
    n179
  );


  buf
  g615
  (
    n638,
    n155
  );


  not
  g616
  (
    n815,
    n179
  );


  not
  g617
  (
    n749,
    n163
  );


  not
  g618
  (
    n981,
    n288
  );


  buf
  g619
  (
    n557,
    n227
  );


  buf
  g620
  (
    n755,
    n284
  );


  buf
  g621
  (
    n808,
    n143
  );


  buf
  g622
  (
    n1079,
    n140
  );


  not
  g623
  (
    n362,
    n133
  );


  buf
  g624
  (
    n969,
    n263
  );


  buf
  g625
  (
    n1136,
    n221
  );


  not
  g626
  (
    n525,
    n224
  );


  buf
  g627
  (
    n613,
    n312
  );


  not
  g628
  (
    n644,
    n245
  );


  not
  g629
  (
    n642,
    n189
  );


  buf
  g630
  (
    n470,
    n299
  );


  not
  g631
  (
    n1022,
    n278
  );


  buf
  g632
  (
    n511,
    n291
  );


  buf
  g633
  (
    n925,
    n229
  );


  not
  g634
  (
    n451,
    n294
  );


  buf
  g635
  (
    n497,
    n185
  );


  not
  g636
  (
    n630,
    n236
  );


  buf
  g637
  (
    n1137,
    n256
  );


  not
  g638
  (
    n571,
    n163
  );


  not
  g639
  (
    n1029,
    n158
  );


  buf
  g640
  (
    n611,
    n207
  );


  not
  g641
  (
    n1076,
    n209
  );


  buf
  g642
  (
    n1033,
    n208
  );


  not
  g643
  (
    n1064,
    n124
  );


  buf
  g644
  (
    n598,
    n298
  );


  not
  g645
  (
    n839,
    n313
  );


  buf
  g646
  (
    n516,
    n176
  );


  buf
  g647
  (
    n710,
    n112
  );


  not
  g648
  (
    n556,
    n228
  );


  not
  g649
  (
    n1115,
    n182
  );


  buf
  g650
  (
    n1020,
    n134
  );


  not
  g651
  (
    n720,
    n115
  );


  buf
  g652
  (
    n982,
    n159
  );


  buf
  g653
  (
    n357,
    n124
  );


  not
  g654
  (
    n819,
    n252
  );


  buf
  g655
  (
    n631,
    n172
  );


  not
  g656
  (
    n481,
    n246
  );


  not
  g657
  (
    n628,
    n283
  );


  buf
  g658
  (
    n503,
    n145
  );


  buf
  g659
  (
    n526,
    n146
  );


  not
  g660
  (
    n1095,
    n236
  );


  buf
  g661
  (
    n325,
    n232
  );


  not
  g662
  (
    n778,
    n281
  );


  buf
  g663
  (
    n931,
    n202
  );


  buf
  g664
  (
    n414,
    n194
  );


  buf
  g665
  (
    n673,
    n120
  );


  not
  g666
  (
    n670,
    n274
  );


  not
  g667
  (
    n896,
    n167
  );


  not
  g668
  (
    n1041,
    n116
  );


  not
  g669
  (
    n994,
    n239
  );


  buf
  g670
  (
    n1093,
    n118
  );


  not
  g671
  (
    n845,
    n265
  );


  not
  g672
  (
    n769,
    n250
  );


  buf
  g673
  (
    n972,
    n185
  );


  not
  g674
  (
    KeyWire_0_10,
    n145
  );


  buf
  g675
  (
    n862,
    n220
  );


  not
  g676
  (
    n616,
    n241
  );


  not
  g677
  (
    n351,
    n195
  );


  not
  g678
  (
    n472,
    n251
  );


  buf
  g679
  (
    n1001,
    n146
  );


  not
  g680
  (
    n955,
    n306
  );


  not
  g681
  (
    n842,
    n301
  );


  not
  g682
  (
    n954,
    n313
  );


  buf
  g683
  (
    n520,
    n257
  );


  buf
  g684
  (
    n378,
    n277
  );


  buf
  g685
  (
    n861,
    n302
  );


  buf
  g686
  (
    n360,
    n176
  );


  buf
  g687
  (
    n944,
    n207
  );


  buf
  g688
  (
    n671,
    n236
  );


  not
  g689
  (
    n463,
    n270
  );


  not
  g690
  (
    n923,
    n122
  );


  buf
  g691
  (
    n707,
    n207
  );


  not
  g692
  (
    n1087,
    n193
  );


  buf
  g693
  (
    n400,
    n129
  );


  buf
  g694
  (
    n437,
    n301
  );


  not
  g695
  (
    n618,
    n187
  );


  not
  g696
  (
    n774,
    n133
  );


  not
  g697
  (
    n575,
    n189
  );


  not
  g698
  (
    n653,
    n261
  );


  not
  g699
  (
    n937,
    n219
  );


  buf
  g700
  (
    n874,
    n120
  );


  not
  g701
  (
    n509,
    n208
  );


  buf
  g702
  (
    n651,
    n205
  );


  not
  g703
  (
    n970,
    n215
  );


  buf
  g704
  (
    n976,
    n316
  );


  not
  g705
  (
    n959,
    n122
  );


  buf
  g706
  (
    n1054,
    n256
  );


  buf
  g707
  (
    n404,
    n272
  );


  buf
  g708
  (
    n800,
    n305
  );


  buf
  g709
  (
    n471,
    n314
  );


  not
  g710
  (
    n713,
    n271
  );


  not
  g711
  (
    n943,
    n159
  );


  buf
  g712
  (
    n894,
    n294
  );


  not
  g713
  (
    n489,
    n288
  );


  not
  g714
  (
    n660,
    n258
  );


  not
  g715
  (
    n696,
    n297
  );


  buf
  g716
  (
    n1092,
    n215
  );


  buf
  g717
  (
    n499,
    n257
  );


  buf
  g718
  (
    n453,
    n260
  );


  buf
  g719
  (
    n865,
    n151
  );


  not
  g720
  (
    n627,
    n167
  );


  not
  g721
  (
    n895,
    n168
  );


  not
  g722
  (
    n507,
    n285
  );


  not
  g723
  (
    n1016,
    n114
  );


  buf
  g724
  (
    n427,
    n221
  );


  not
  g725
  (
    n444,
    n289
  );


  not
  g726
  (
    n1059,
    n208
  );


  buf
  g727
  (
    n1012,
    n210
  );


  not
  g728
  (
    KeyWire_0_23,
    n117
  );


  not
  g729
  (
    n729,
    n184
  );


  buf
  g730
  (
    n373,
    n243
  );


  buf
  g731
  (
    n1046,
    n292
  );


  not
  g732
  (
    n1068,
    n192
  );


  not
  g733
  (
    n968,
    n305
  );


  not
  g734
  (
    n1060,
    n198
  );


  not
  g735
  (
    n1002,
    n170
  );


  not
  g736
  (
    n328,
    n210
  );


  not
  g737
  (
    n332,
    n250
  );


  buf
  g738
  (
    n408,
    n222
  );


  buf
  g739
  (
    n1055,
    n160
  );


  not
  g740
  (
    n914,
    n197
  );


  not
  g741
  (
    n629,
    n199
  );


  not
  g742
  (
    n333,
    n146
  );


  not
  g743
  (
    n904,
    n149
  );


  not
  g744
  (
    n715,
    n229
  );


  not
  g745
  (
    n535,
    n211
  );


  buf
  g746
  (
    n442,
    n269
  );


  not
  g747
  (
    n832,
    n244
  );


  buf
  g748
  (
    n456,
    n269
  );


  buf
  g749
  (
    n777,
    n309
  );


  buf
  g750
  (
    n361,
    n306
  );


  buf
  g751
  (
    n952,
    n174
  );


  buf
  g752
  (
    n512,
    n247
  );


  buf
  g753
  (
    n902,
    n164
  );


  buf
  g754
  (
    KeyWire_0_5,
    n157
  );


  not
  g755
  (
    n1031,
    n159
  );


  not
  g756
  (
    n640,
    n169
  );


  buf
  g757
  (
    n595,
    n235
  );


  buf
  g758
  (
    n867,
    n253
  );


  buf
  g759
  (
    n876,
    n190
  );


  not
  g760
  (
    n714,
    n287
  );


  buf
  g761
  (
    n440,
    n255
  );


  not
  g762
  (
    n1028,
    n149
  );


  not
  g763
  (
    n905,
    n214
  );


  buf
  g764
  (
    n534,
    n132
  );


  not
  g765
  (
    n654,
    n262
  );


  buf
  g766
  (
    n975,
    n266
  );


  not
  g767
  (
    n1037,
    n294
  );


  not
  g768
  (
    n596,
    n157
  );


  buf
  g769
  (
    n678,
    n254
  );


  not
  g770
  (
    n992,
    n137
  );


  not
  g771
  (
    n506,
    n212
  );


  not
  g772
  (
    n983,
    n237
  );


  not
  g773
  (
    n941,
    n252
  );


  not
  g774
  (
    n648,
    n141
  );


  buf
  g775
  (
    n1058,
    n255
  );


  not
  g776
  (
    n406,
    n200
  );


  not
  g777
  (
    n805,
    n123
  );


  not
  g778
  (
    n950,
    n209
  );


  buf
  g779
  (
    KeyWire_0_13,
    n156
  );


  not
  g780
  (
    n543,
    n115
  );


  not
  g781
  (
    n531,
    n150
  );


  buf
  g782
  (
    n898,
    n152
  );


  buf
  g783
  (
    n387,
    n139
  );


  buf
  g784
  (
    n912,
    n244
  );


  not
  g785
  (
    n375,
    n118
  );


  not
  g786
  (
    n870,
    n253
  );


  buf
  g787
  (
    n327,
    n162
  );


  not
  g788
  (
    n482,
    n256
  );


  buf
  g789
  (
    n381,
    n278
  );


  not
  g790
  (
    n606,
    n315
  );


  not
  g791
  (
    n901,
    n137
  );


  buf
  g792
  (
    n1085,
    n197
  );


  buf
  g793
  (
    n911,
    n297
  );


  buf
  g794
  (
    n725,
    n198
  );


  buf
  g795
  (
    n1088,
    n191
  );


  buf
  g796
  (
    n791,
    n178
  );


  buf
  g797
  (
    n790,
    n154
  );


  not
  g798
  (
    n1104,
    n211
  );


  not
  g799
  (
    n449,
    n110
  );


  not
  g800
  (
    n847,
    n202
  );


  not
  g801
  (
    n936,
    n285
  );


  buf
  g802
  (
    n1096,
    n243
  );


  buf
  g803
  (
    n485,
    n220
  );


  buf
  g804
  (
    n690,
    n150
  );


  not
  g805
  (
    n918,
    n261
  );


  not
  g806
  (
    n856,
    n157
  );


  buf
  g807
  (
    n574,
    n265
  );


  not
  g808
  (
    n439,
    n123
  );


  buf
  g809
  (
    n990,
    n189
  );


  not
  g810
  (
    n930,
    n156
  );


  not
  g811
  (
    n706,
    n148
  );


  not
  g812
  (
    n1120,
    n233
  );


  not
  g813
  (
    n883,
    n222
  );


  not
  g814
  (
    n338,
    n174
  );


  not
  g815
  (
    n719,
    n128
  );


  not
  g816
  (
    n479,
    n281
  );


  not
  g817
  (
    n547,
    n278
  );


  buf
  g818
  (
    n683,
    n192
  );


  buf
  g819
  (
    n906,
    n117
  );


  not
  g820
  (
    n1013,
    n190
  );


  buf
  g821
  (
    n890,
    n154
  );


  not
  g822
  (
    n647,
    n186
  );


  not
  g823
  (
    n401,
    n127
  );


  not
  g824
  (
    n919,
    n164
  );


  buf
  g825
  (
    n933,
    n187
  );


  buf
  g826
  (
    n1139,
    n267
  );


  not
  g827
  (
    n1007,
    n175
  );


  buf
  g828
  (
    n592,
    n270
  );


  buf
  g829
  (
    n1128,
    n153
  );


  not
  g830
  (
    n691,
    n267
  );


  buf
  g831
  (
    n422,
    n169
  );


  buf
  g832
  (
    n920,
    n153
  );


  buf
  g833
  (
    n372,
    n184
  );


  not
  g834
  (
    n483,
    n187
  );


  not
  g835
  (
    n1011,
    n147
  );


  not
  g836
  (
    n1132,
    n200
  );


  buf
  g837
  (
    n473,
    n222
  );


  not
  g838
  (
    n834,
    n152
  );


  not
  g839
  (
    n916,
    n181
  );


  buf
  g840
  (
    n657,
    n264
  );


  not
  g841
  (
    n682,
    n116
  );


  buf
  g842
  (
    n544,
    n316
  );


  buf
  g843
  (
    n953,
    n275
  );


  not
  g844
  (
    n374,
    n219
  );


  not
  g845
  (
    n1043,
    n226
  );


  buf
  g846
  (
    n779,
    n283
  );


  buf
  g847
  (
    n446,
    n230
  );


  buf
  g848
  (
    n709,
    n296
  );


  buf
  g849
  (
    n927,
    n295
  );


  not
  g850
  (
    n350,
    n183
  );


  not
  g851
  (
    n866,
    n127
  );


  not
  g852
  (
    n417,
    n295
  );


  not
  g853
  (
    n546,
    n244
  );


  buf
  g854
  (
    n551,
    n123
  );


  buf
  g855
  (
    n578,
    n310
  );


  buf
  g856
  (
    n754,
    n111
  );


  buf
  g857
  (
    n756,
    n291
  );


  buf
  g858
  (
    n946,
    n234
  );


  buf
  g859
  (
    n887,
    n305
  );


  buf
  g860
  (
    n1053,
    n274
  );


  buf
  g861
  (
    n676,
    n193
  );


  buf
  g862
  (
    n965,
    n217
  );


  not
  g863
  (
    n649,
    n186
  );


  not
  g864
  (
    n345,
    n312
  );


  buf
  g865
  (
    n881,
    n168
  );


  not
  g866
  (
    n748,
    n264
  );


  buf
  g867
  (
    n1035,
    n299
  );


  not
  g868
  (
    n674,
    n177
  );


  buf
  g869
  (
    n542,
    n218
  );


  buf
  g870
  (
    n903,
    n140
  );


  buf
  g871
  (
    n491,
    n200
  );


  not
  g872
  (
    n762,
    n141
  );


  not
  g873
  (
    KeyWire_0_19,
    n309
  );


  not
  g874
  (
    n604,
    n199
  );


  buf
  g875
  (
    n741,
    n198
  );


  buf
  g876
  (
    n793,
    n246
  );


  buf
  g877
  (
    KeyWire_0_4,
    n179
  );


  buf
  g878
  (
    n384,
    n136
  );


  not
  g879
  (
    n612,
    n180
  );


  buf
  g880
  (
    n1127,
    n235
  );


  buf
  g881
  (
    n835,
    n222
  );


  buf
  g882
  (
    n988,
    n302
  );


  buf
  g883
  (
    n772,
    n297
  );


  not
  g884
  (
    n993,
    n147
  );


  buf
  g885
  (
    n813,
    n129
  );


  buf
  g886
  (
    n880,
    n199
  );


  not
  g887
  (
    n558,
    n244
  );


  buf
  g888
  (
    n562,
    n233
  );


  not
  g889
  (
    n697,
    n178
  );


  not
  g890
  (
    n742,
    n263
  );


  buf
  g891
  (
    n998,
    n266
  );


  not
  g892
  (
    n730,
    n125
  );


  not
  g893
  (
    n900,
    n304
  );


  buf
  g894
  (
    n1101,
    n217
  );


  not
  g895
  (
    n411,
    n148
  );


  not
  g896
  (
    n435,
    n280
  );


  buf
  g897
  (
    n1122,
    n223
  );


  not
  g898
  (
    n650,
    n240
  );


  not
  g899
  (
    n622,
    n276
  );


  buf
  g900
  (
    n458,
    n242
  );


  not
  g901
  (
    n928,
    n293
  );


  buf
  g902
  (
    n1004,
    n252
  );


  not
  g903
  (
    n1005,
    n216
  );


  not
  g904
  (
    n412,
    n195
  );


  not
  g905
  (
    n801,
    n278
  );


  not
  g906
  (
    n601,
    n269
  );


  buf
  g907
  (
    KeyWire_0_15,
    n263
  );


  not
  g908
  (
    n537,
    n209
  );


  not
  g909
  (
    n665,
    n234
  );


  not
  g910
  (
    n915,
    n273
  );


  buf
  g911
  (
    n354,
    n167
  );


  buf
  g912
  (
    n716,
    n305
  );


  not
  g913
  (
    n424,
    n165
  );


  buf
  g914
  (
    n810,
    n312
  );


  buf
  g915
  (
    n977,
    n284
  );


  not
  g916
  (
    n1062,
    n267
  );


  buf
  g917
  (
    n621,
    n160
  );


  not
  g918
  (
    n852,
    n181
  );


  not
  g919
  (
    n624,
    n144
  );


  buf
  g920
  (
    n366,
    n130
  );


  not
  g921
  (
    n795,
    n265
  );


  not
  g922
  (
    n1098,
    n307
  );


  not
  g923
  (
    n926,
    n235
  );


  buf
  g924
  (
    n699,
    n124
  );


  buf
  g925
  (
    n830,
    n307
  );


  buf
  g926
  (
    n356,
    n204
  );


  not
  g927
  (
    n986,
    n169
  );


  not
  g928
  (
    n498,
    n120
  );


  buf
  g929
  (
    n974,
    n241
  );


  not
  g930
  (
    n399,
    n206
  );


  not
  g931
  (
    n331,
    n124
  );


  not
  g932
  (
    n589,
    n289
  );


  not
  g933
  (
    n1086,
    n247
  );


  not
  g934
  (
    n669,
    n146
  );


  not
  g935
  (
    n441,
    n166
  );


  not
  g936
  (
    n495,
    n287
  );


  not
  g937
  (
    n607,
    n155
  );


  not
  g938
  (
    n668,
    n296
  );


  not
  g939
  (
    n724,
    n274
  );


  not
  g940
  (
    n1083,
    n311
  );


  buf
  g941
  (
    n799,
    n172
  );


  buf
  g942
  (
    n945,
    n272
  );


  not
  g943
  (
    n359,
    n112
  );


  buf
  g944
  (
    n979,
    n170
  );


  not
  g945
  (
    n603,
    n200
  );


  not
  g946
  (
    n593,
    n132
  );


  not
  g947
  (
    n662,
    n111
  );


  buf
  g948
  (
    n701,
    n164
  );


  not
  g949
  (
    n1073,
    n260
  );


  not
  g950
  (
    n875,
    n217
  );


  buf
  g951
  (
    n1130,
    n171
  );


  buf
  g952
  (
    n484,
    n248
  );


  not
  g953
  (
    n851,
    n194
  );


  not
  g954
  (
    n431,
    n127
  );


  buf
  g955
  (
    n633,
    n294
  );


  buf
  g956
  (
    n639,
    n140
  );


  not
  g957
  (
    n513,
    n113
  );


  buf
  g958
  (
    n879,
    n158
  );


  buf
  g959
  (
    n389,
    n231
  );


  not
  g960
  (
    n397,
    n295
  );


  not
  g961
  (
    n732,
    n227
  );


  buf
  g962
  (
    n569,
    n300
  );


  not
  g963
  (
    n586,
    n186
  );


  buf
  g964
  (
    n450,
    n247
  );


  not
  g965
  (
    n689,
    n156
  );


  not
  g966
  (
    n817,
    n286
  );


  not
  g967
  (
    n568,
    n229
  );


  not
  g968
  (
    n1111,
    n271
  );


  not
  g969
  (
    n792,
    n110
  );


  buf
  g970
  (
    n1102,
    n217
  );


  not
  g971
  (
    n409,
    n230
  );


  not
  g972
  (
    n760,
    n242
  );


  buf
  g973
  (
    n518,
    n219
  );


  not
  g974
  (
    n718,
    n216
  );


  not
  g975
  (
    n811,
    n213
  );


  buf
  g976
  (
    n717,
    n116
  );


  buf
  g977
  (
    n566,
    n111
  );


  not
  g978
  (
    n884,
    n250
  );


  not
  g979
  (
    n632,
    n123
  );


  not
  g980
  (
    n448,
    n158
  );


  not
  g981
  (
    n398,
    n154
  );


  buf
  g982
  (
    n733,
    n315
  );


  not
  g983
  (
    n825,
    n184
  );


  not
  g984
  (
    n693,
    n118
  );


  not
  g985
  (
    n768,
    n162
  );


  not
  g986
  (
    n766,
    n219
  );


  not
  g987
  (
    n761,
    n132
  );


  buf
  g988
  (
    n486,
    n226
  );


  buf
  g989
  (
    n743,
    n165
  );


  buf
  g990
  (
    n737,
    n306
  );


  buf
  g991
  (
    KeyWire_0_2,
    n226
  );


  not
  g992
  (
    n646,
    n126
  );


  buf
  g993
  (
    n529,
    n206
  );


  buf
  g994
  (
    n521,
    n122
  );


  not
  g995
  (
    n541,
    n232
  );


  buf
  g996
  (
    n1010,
    n145
  );


  not
  g997
  (
    n996,
    n201
  );


  not
  g998
  (
    n922,
    n310
  );


  buf
  g999
  (
    n703,
    n156
  );


  buf
  g1000
  (
    n455,
    n290
  );


  buf
  g1001
  (
    n872,
    n131
  );


  buf
  g1002
  (
    n827,
    n137
  );


  buf
  g1003
  (
    n545,
    n285
  );


  buf
  g1004
  (
    n352,
    n221
  );


  not
  g1005
  (
    n877,
    n173
  );


  not
  g1006
  (
    n956,
    n134
  );


  not
  g1007
  (
    n634,
    n267
  );


  not
  g1008
  (
    n837,
    n181
  );


  not
  g1009
  (
    n850,
    n190
  );


  buf
  g1010
  (
    n459,
    n251
  );


  not
  g1011
  (
    n833,
    n121
  );


  buf
  g1012
  (
    n1107,
    n228
  );


  not
  g1013
  (
    n555,
    n304
  );


  buf
  g1014
  (
    n1044,
    n301
  );


  not
  g1015
  (
    n1134,
    n238
  );


  not
  g1016
  (
    n907,
    n268
  );


  buf
  g1017
  (
    n1123,
    n166
  );


  not
  g1018
  (
    n804,
    n272
  );


  not
  g1019
  (
    n576,
    n260
  );


  buf
  g1020
  (
    n750,
    n243
  );


  not
  g1021
  (
    n407,
    n300
  );


  buf
  g1022
  (
    n581,
    n258
  );


  buf
  g1023
  (
    n1084,
    n195
  );


  buf
  g1024
  (
    n1100,
    n110
  );


  buf
  g1025
  (
    n848,
    n276
  );


  buf
  g1026
  (
    n637,
    n233
  );


  not
  g1027
  (
    n434,
    n231
  );


  not
  g1028
  (
    n773,
    n160
  );


  not
  g1029
  (
    n1019,
    n290
  );


  not
  g1030
  (
    n392,
    n193
  );


  buf
  g1031
  (
    n1066,
    n293
  );


  not
  g1032
  (
    n672,
    n121
  );


  buf
  g1033
  (
    n932,
    n216
  );


  buf
  g1034
  (
    n1072,
    n228
  );


  not
  g1035
  (
    n582,
    n233
  );


  not
  g1036
  (
    n909,
    n225
  );


  not
  g1037
  (
    n757,
    n143
  );


  not
  g1038
  (
    n436,
    n254
  );


  buf
  g1039
  (
    n1030,
    n166
  );


  buf
  g1040
  (
    n605,
    n313
  );


  not
  g1041
  (
    n685,
    n239
  );


  buf
  g1042
  (
    n1040,
    n136
  );


  buf
  g1043
  (
    n420,
    n250
  );


  not
  g1044
  (
    n891,
    n242
  );


  buf
  g1045
  (
    n721,
    n143
  );


  buf
  g1046
  (
    n1042,
    n243
  );


  not
  g1047
  (
    n1110,
    n205
  );


  buf
  g1048
  (
    n1061,
    n270
  );


  not
  g1049
  (
    n524,
    n277
  );


  not
  g1050
  (
    n973,
    n184
  );


  buf
  g1051
  (
    n438,
    n308
  );


  buf
  g1052
  (
    KeyWire_0_26,
    n175
  );


  not
  g1053
  (
    n1067,
    n142
  );


  not
  g1054
  (
    n391,
    n273
  );


  not
  g1055
  (
    n1078,
    n266
  );


  buf
  g1056
  (
    n490,
    n203
  );


  not
  g1057
  (
    n501,
    n169
  );


  not
  g1058
  (
    n421,
    n201
  );


  not
  g1059
  (
    n854,
    n113
  );


  buf
  g1060
  (
    n538,
    n240
  );


  buf
  g1061
  (
    n1089,
    n183
  );


  buf
  g1062
  (
    n585,
    n181
  );


  buf
  g1063
  (
    n587,
    n249
  );


  not
  g1064
  (
    n822,
    n175
  );


  not
  g1065
  (
    n1045,
    n309
  );


  not
  g1066
  (
    n565,
    n240
  );


  buf
  g1067
  (
    n339,
    n150
  );


  not
  g1068
  (
    n1118,
    n248
  );


  buf
  g1069
  (
    n855,
    n213
  );


  not
  g1070
  (
    n878,
    n130
  );


  buf
  g1071
  (
    n615,
    n299
  );


  not
  g1072
  (
    n418,
    n230
  );


  buf
  g1073
  (
    n514,
    n225
  );


  buf
  g1074
  (
    n487,
    n269
  );


  buf
  g1075
  (
    n626,
    n236
  );


  buf
  g1076
  (
    n550,
    n245
  );


  buf
  g1077
  (
    n948,
    n288
  );


  buf
  g1078
  (
    n386,
    n176
  );


  not
  g1079
  (
    n460,
    n125
  );


  buf
  g1080
  (
    n658,
    n153
  );


  not
  g1081
  (
    n712,
    n317
  );


  buf
  g1082
  (
    n824,
    n299
  );


  not
  g1083
  (
    n746,
    n153
  );


  buf
  g1084
  (
    n961,
    n224
  );


  buf
  g1085
  (
    n675,
    n177
  );


  not
  g1086
  (
    n767,
    n231
  );


  not
  g1087
  (
    n1129,
    n210
  );


  not
  g1088
  (
    n1034,
    n212
  );


  buf
  g1089
  (
    n423,
    n195
  );


  buf
  g1090
  (
    n752,
    n179
  );


  not
  g1091
  (
    n991,
    n116
  );


  buf
  g1092
  (
    n377,
    n198
  );


  buf
  g1093
  (
    n1057,
    n257
  );


  not
  g1094
  (
    n517,
    n237
  );


  not
  g1095
  (
    n355,
    n119
  );


  not
  g1096
  (
    n1094,
    n163
  );


  not
  g1097
  (
    n806,
    n289
  );


  not
  g1098
  (
    n591,
    n178
  );


  not
  g1099
  (
    n967,
    n292
  );


  nand
  g1100
  (
    n705,
    n241,
    n192
  );


  nor
  g1101
  (
    n1027,
    n112,
    n207
  );


  or
  g1102
  (
    n957,
    n249,
    n261,
    n144,
    n282
  );


  nor
  g1103
  (
    n1070,
    n202,
    n133,
    n172,
    n289
  );


  xnor
  g1104
  (
    n553,
    n213,
    n255,
    n282,
    n120
  );


  or
  g1105
  (
    n849,
    n280,
    n173,
    n223,
    n259
  );


  nand
  g1106
  (
    n349,
    n268,
    n206,
    n148,
    n183
  );


  xor
  g1107
  (
    n1256,
    n640,
    n558,
    n533,
    n800
  );


  xor
  g1108
  (
    n1224,
    n507,
    n1102,
    n462,
    n851
  );


  and
  g1109
  (
    n1171,
    n483,
    n545,
    n1030,
    n386
  );


  and
  g1110
  (
    n1249,
    n352,
    n677,
    n1008,
    n982
  );


  xnor
  g1111
  (
    n1277,
    n540,
    n476,
    n642,
    n838
  );


  xnor
  g1112
  (
    n1306,
    n567,
    n826,
    n815,
    n1069
  );


  and
  g1113
  (
    n1156,
    n370,
    n784,
    n732,
    n983
  );


  xnor
  g1114
  (
    n1184,
    n820,
    n842,
    n853,
    n901
  );


  xor
  g1115
  (
    n1283,
    n753,
    n681,
    n612,
    n822
  );


  nand
  g1116
  (
    n1192,
    n963,
    n1087,
    n759,
    n442
  );


  xor
  g1117
  (
    n1259,
    n809,
    n895,
    n512,
    n931
  );


  nand
  g1118
  (
    n1189,
    n551,
    n745,
    n795,
    n1099
  );


  nor
  g1119
  (
    n1307,
    n936,
    n439,
    n868,
    n816
  );


  nand
  g1120
  (
    n1247,
    n773,
    n1010,
    n557,
    n930
  );


  and
  g1121
  (
    n1197,
    n750,
    n635,
    n423,
    n531
  );


  or
  g1122
  (
    n1239,
    n1015,
    n695,
    n768,
    n333
  );


  nand
  g1123
  (
    n1202,
    n463,
    n388,
    n879,
    n948
  );


  nor
  g1124
  (
    n1167,
    n814,
    n790,
    n690,
    n457
  );


  nor
  g1125
  (
    n1285,
    n398,
    n758,
    n541,
    n973
  );


  or
  g1126
  (
    n1294,
    n385,
    n698,
    n996,
    n906
  );


  xnor
  g1127
  (
    n1272,
    n1063,
    n657,
    n1045,
    n378
  );


  and
  g1128
  (
    n1203,
    n630,
    n1070,
    n513,
    n817
  );


  nand
  g1129
  (
    n1164,
    n847,
    n489,
    n871,
    n441
  );


  xor
  g1130
  (
    n1251,
    n669,
    n1072,
    n430,
    n468
  );


  nor
  g1131
  (
    n1289,
    n535,
    n726,
    n992,
    n966
  );


  nand
  g1132
  (
    n1291,
    n436,
    n775,
    n420,
    n629
  );


  nor
  g1133
  (
    n1245,
    n914,
    n849,
    n550,
    n371
  );


  and
  g1134
  (
    n1280,
    n549,
    n362,
    n818,
    n797
  );


  xnor
  g1135
  (
    n1241,
    n702,
    n782,
    n437,
    n583
  );


  nand
  g1136
  (
    n1205,
    n808,
    n325,
    n751,
    n350
  );


  nor
  g1137
  (
    n1158,
    n919,
    n345,
    n515,
    n353
  );


  nand
  g1138
  (
    n1297,
    n989,
    n903,
    n576,
    n860
  );


  xnor
  g1139
  (
    n1242,
    n1081,
    n834,
    n661,
    n670
  );


  nor
  g1140
  (
    n1264,
    n344,
    n869,
    n747,
    n343
  );


  xnor
  g1141
  (
    n1252,
    n696,
    n426,
    n984,
    n451
  );


  nand
  g1142
  (
    n1292,
    n943,
    n892,
    n380,
    n391
  );


  nand
  g1143
  (
    n1319,
    n571,
    n406,
    n1088,
    n332
  );


  xor
  g1144
  (
    n1270,
    n1033,
    n1056,
    n520,
    n968
  );


  xnor
  g1145
  (
    n1144,
    n662,
    n1096,
    n401,
    n418
  );


  xnor
  g1146
  (
    n1331,
    n446,
    n777,
    n337,
    n1024
  );


  nand
  g1147
  (
    n1255,
    n978,
    n918,
    n665,
    n947
  );


  xor
  g1148
  (
    n1322,
    n1020,
    n1057,
    n1003,
    n673
  );


  or
  g1149
  (
    n1181,
    n429,
    n1001,
    n921,
    n565
  );


  xor
  g1150
  (
    n1151,
    n884,
    n939,
    n461,
    n647
  );


  nor
  g1151
  (
    n1216,
    n360,
    n603,
    n588,
    n453
  );


  and
  g1152
  (
    n1260,
    n718,
    n574,
    n626,
    n606
  );


  xnor
  g1153
  (
    n1262,
    n465,
    n538,
    n503,
    n894
  );


  and
  g1154
  (
    n1198,
    n639,
    n1060,
    n664,
    n835
  );


  nand
  g1155
  (
    n1293,
    n445,
    n1038,
    n827,
    n1097
  );


  xor
  g1156
  (
    n1223,
    n659,
    n740,
    n688,
    n944
  );


  and
  g1157
  (
    KeyWire_0_0,
    n686,
    n706,
    n1034,
    n529
  );


  xor
  g1158
  (
    n1305,
    n631,
    n774,
    n393,
    n499
  );


  xnor
  g1159
  (
    n1316,
    n694,
    n585,
    n757,
    n472
  );


  xor
  g1160
  (
    n1195,
    n789,
    n743,
    n972,
    n1083
  );


  nand
  g1161
  (
    n1199,
    n500,
    n793,
    n922,
    n582
  );


  nor
  g1162
  (
    n1254,
    n709,
    n554,
    n544,
    n925
  );


  nand
  g1163
  (
    n1211,
    n564,
    n464,
    n475,
    n638
  );


  xor
  g1164
  (
    n1253,
    n1071,
    n794,
    n762,
    n598
  );


  nand
  g1165
  (
    n1302,
    n848,
    n942,
    n419,
    n712
  );


  nor
  g1166
  (
    n1178,
    n828,
    n813,
    n786,
    n605
  );


  xnor
  g1167
  (
    n1166,
    n552,
    n508,
    n769,
    n327
  );


  nand
  g1168
  (
    n1318,
    n1047,
    n372,
    n466,
    n637
  );


  xnor
  g1169
  (
    n1185,
    n701,
    n716,
    n1074,
    n594
  );


  nand
  g1170
  (
    n1175,
    n609,
    n447,
    n599,
    n619
  );


  nor
  g1171
  (
    n1244,
    n810,
    n608,
    n1029,
    n632
  );


  and
  g1172
  (
    n1250,
    n923,
    n699,
    n413,
    n411
  );


  or
  g1173
  (
    n1206,
    n843,
    n1027,
    n787,
    n514
  );


  or
  g1174
  (
    n1188,
    n364,
    n1086,
    n502,
    n870
  );


  xnor
  g1175
  (
    n1308,
    n953,
    n737,
    n749,
    n1077
  );


  xor
  g1176
  (
    n1311,
    n330,
    n691,
    n841,
    n358
  );


  xor
  g1177
  (
    n1142,
    n534,
    n591,
    n1002,
    n649
  );


  nor
  g1178
  (
    n1235,
    n1028,
    n524,
    n766,
    n952
  );


  and
  g1179
  (
    n1204,
    n1094,
    n799,
    n443,
    n334
  );


  and
  g1180
  (
    n1246,
    n897,
    n985,
    n1059,
    n575
  );


  nor
  g1181
  (
    n1296,
    n623,
    n404,
    n1100,
    n405
  );


  nor
  g1182
  (
    n1145,
    n700,
    n440,
    n1031,
    n1007
  );


  nor
  g1183
  (
    n1177,
    n748,
    n862,
    n528,
    n875
  );


  nor
  g1184
  (
    n1234,
    n738,
    n374,
    n744,
    n579
  );


  or
  g1185
  (
    n1238,
    n671,
    n891,
    n1025,
    n1032
  );


  or
  g1186
  (
    n1217,
    n491,
    n929,
    n880,
    n555
  );


  xor
  g1187
  (
    n1295,
    n850,
    n883,
    n467,
    n410
  );


  and
  g1188
  (
    n1230,
    n1090,
    n331,
    n480,
    n941
  );


  xor
  g1189
  (
    n1231,
    n1067,
    n368,
    n525,
    n909
  );


  or
  g1190
  (
    n1212,
    n846,
    n864,
    n381,
    n521
  );


  xor
  g1191
  (
    n1268,
    n627,
    n346,
    n487,
    n733
  );


  nor
  g1192
  (
    n1183,
    n348,
    n653,
    n924,
    n837
  );


  or
  g1193
  (
    n1169,
    n396,
    n804,
    n832,
    n422
  );


  xnor
  g1194
  (
    n1190,
    n980,
    n811,
    n361,
    n648
  );


  xnor
  g1195
  (
    n1159,
    n377,
    n902,
    n604,
    n542
  );


  nor
  g1196
  (
    n1174,
    n1040,
    n645,
    n363,
    n424
  );


  xnor
  g1197
  (
    n1141,
    n1017,
    n735,
    n537,
    n711
  );


  xnor
  g1198
  (
    n1222,
    n459,
    n1014,
    n824,
    n1098
  );


  nand
  g1199
  (
    n1172,
    n548,
    n741,
    n937,
    n651
  );


  xnor
  g1200
  (
    n1168,
    n729,
    n1064,
    n1011,
    n633
  );


  or
  g1201
  (
    n1213,
    n920,
    n482,
    n478,
    n428
  );


  nand
  g1202
  (
    n1271,
    n680,
    n1022,
    n610,
    n589
  );


  xor
  g1203
  (
    n1300,
    n357,
    n1079,
    n636,
    n584
  );


  and
  g1204
  (
    n1304,
    n960,
    n934,
    n383,
    n1051
  );


  xor
  g1205
  (
    n1312,
    n889,
    n369,
    n994,
    n679
  );


  or
  g1206
  (
    n1193,
    n1018,
    n339,
    n526,
    n618
  );


  xnor
  g1207
  (
    n1290,
    n407,
    n728,
    n867,
    n1021
  );


  or
  g1208
  (
    n1269,
    n833,
    n742,
    n964,
    n821
  );


  and
  g1209
  (
    n1329,
    n865,
    n493,
    n915,
    n427
  );


  xor
  g1210
  (
    n1328,
    n907,
    n975,
    n354,
    n456
  );


  nor
  g1211
  (
    n1314,
    n394,
    n704,
    n976,
    n561
  );


  nor
  g1212
  (
    n1276,
    n477,
    n416,
    n438,
    n1062
  );


  or
  g1213
  (
    n1310,
    n874,
    n1036,
    n615,
    n572
  );


  nand
  g1214
  (
    n1327,
    n580,
    n556,
    n779,
    n504
  );


  and
  g1215
  (
    n1320,
    n998,
    n559,
    n873,
    n1058
  );


  xor
  g1216
  (
    n1274,
    n1080,
    n1005,
    n519,
    n505
  );


  xor
  g1217
  (
    n1321,
    n641,
    n683,
    n855,
    n658
  );


  and
  g1218
  (
    n1179,
    n607,
    n1104,
    n628,
    n812
  );


  or
  g1219
  (
    n1303,
    n1082,
    n689,
    n595,
    n560
  );


  and
  g1220
  (
    n1149,
    n387,
    n896,
    n715,
    n460
  );


  xor
  g1221
  (
    n1209,
    n755,
    n736,
    n536,
    n425
  );


  or
  g1222
  (
    n1150,
    n625,
    n977,
    n484,
    n955
  );


  or
  g1223
  (
    n1143,
    n831,
    n1043,
    n634,
    n1055
  );


  and
  g1224
  (
    n1154,
    n490,
    n336,
    n592,
    n1095
  );


  and
  g1225
  (
    n1325,
    n783,
    n845,
    n375,
    n581
  );


  xnor
  g1226
  (
    n1218,
    n342,
    n938,
    n444,
    n965
  );


  xor
  g1227
  (
    n1258,
    n433,
    n1044,
    n1073,
    n1078
  );


  xor
  g1228
  (
    n1221,
    n928,
    n365,
    n703,
    n951
  );


  xnor
  g1229
  (
    n1180,
    n705,
    n993,
    n899,
    n667
  );


  or
  g1230
  (
    n1284,
    n359,
    n516,
    n933,
    n624
  );


  or
  g1231
  (
    n1176,
    n586,
    n876,
    n959,
    n373
  );


  nand
  g1232
  (
    n1146,
    n721,
    n780,
    n962,
    n448
  );


  or
  g1233
  (
    n1191,
    n771,
    n991,
    n553,
    n1023
  );


  and
  g1234
  (
    n1186,
    n971,
    n326,
    n518,
    n656
  );


  xnor
  g1235
  (
    n1240,
    n1101,
    n668,
    n912,
    n685
  );


  xor
  g1236
  (
    n1263,
    n1004,
    n1019,
    n1068,
    n997
  );


  and
  g1237
  (
    n1324,
    n593,
    n577,
    n796,
    n431
  );


  nand
  g1238
  (
    n1152,
    n935,
    n434,
    n678,
    n421
  );


  nand
  g1239
  (
    n1157,
    n693,
    n995,
    n587,
    n328
  );


  or
  g1240
  (
    n1214,
    n825,
    n1037,
    n458,
    n961
  );


  nor
  g1241
  (
    n1265,
    n829,
    n1091,
    n522,
    n1035
  );


  xnor
  g1242
  (
    n1232,
    n355,
    n1013,
    n1084,
    n496
  );


  nand
  g1243
  (
    n1279,
    n400,
    n990,
    n986,
    n517
  );


  and
  g1244
  (
    n1210,
    n954,
    n710,
    n886,
    n878
  );


  nor
  g1245
  (
    n1313,
    n616,
    n682,
    n798,
    n905
  );


  xnor
  g1246
  (
    n1317,
    n765,
    n772,
    n347,
    n946
  );


  nand
  g1247
  (
    n1153,
    n687,
    n1052,
    n852,
    n1076
  );


  and
  g1248
  (
    n1165,
    n644,
    n725,
    n408,
    n498
  );


  xnor
  g1249
  (
    n1227,
    n449,
    n562,
    n731,
    n547
  );


  and
  g1250
  (
    n1298,
    n958,
    n597,
    n940,
    n926
  );


  xnor
  g1251
  (
    n1309,
    n1075,
    n893,
    n614,
    n970
  );


  xor
  g1252
  (
    n1333,
    n707,
    n384,
    n674,
    n486
  );


  nor
  g1253
  (
    n1225,
    n746,
    n417,
    n546,
    n720
  );


  nand
  g1254
  (
    n1162,
    n470,
    n877,
    n435,
    n349
  );


  or
  g1255
  (
    n1160,
    n719,
    n807,
    n672,
    n511
  );


  nand
  g1256
  (
    n1170,
    n495,
    n887,
    n563,
    n969
  );


  and
  g1257
  (
    n1278,
    n1000,
    n454,
    n999,
    n613
  );


  nor
  g1258
  (
    n1323,
    n501,
    n979,
    n450,
    n739
  );


  and
  g1259
  (
    n1248,
    n568,
    n455,
    n338,
    n1093
  );


  nor
  g1260
  (
    n1330,
    n727,
    n830,
    n1085,
    n601
  );


  xnor
  g1261
  (
    n1299,
    n510,
    n340,
    n872,
    n1054
  );


  nor
  g1262
  (
    n1243,
    n335,
    n904,
    n366,
    n857
  );


  or
  g1263
  (
    n1233,
    n844,
    n945,
    n730,
    n432
  );


  and
  g1264
  (
    n1201,
    n494,
    n523,
    n932,
    n916
  );


  or
  g1265
  (
    n1301,
    n981,
    n770,
    n785,
    n646
  );


  nor
  g1266
  (
    n1208,
    n474,
    n1006,
    n471,
    n473
  );


  xnor
  g1267
  (
    n1287,
    n367,
    n761,
    n756,
    n600
  );


  nand
  g1268
  (
    n1187,
    n376,
    n1092,
    n570,
    n652
  );


  xor
  g1269
  (
    n1148,
    n697,
    n530,
    n776,
    n752
  );


  and
  g1270
  (
    n1163,
    n341,
    n1089,
    n910,
    n497
  );


  nor
  g1271
  (
    n1288,
    n734,
    n684,
    n402,
    n806
  );


  and
  g1272
  (
    n1326,
    n666,
    n379,
    n655,
    n650
  );


  nand
  g1273
  (
    n1273,
    n527,
    n861,
    n713,
    n805
  );


  or
  g1274
  (
    n1266,
    n967,
    n415,
    n890,
    n492
  );


  nand
  g1275
  (
    n1282,
    n792,
    n1041,
    n676,
    n596
  );


  nand
  g1276
  (
    n1173,
    n974,
    n488,
    n819,
    n590
  );


  and
  g1277
  (
    n1161,
    n708,
    n908,
    n356,
    n927
  );


  xnor
  g1278
  (
    n1236,
    n621,
    n692,
    n1050,
    n399
  );


  or
  g1279
  (
    n1267,
    n791,
    n617,
    n602,
    n573
  );


  or
  g1280
  (
    n1315,
    n760,
    n1042,
    n663,
    n900
  );


  xnor
  g1281
  (
    n1147,
    n1065,
    n885,
    n724,
    n764
  );


  xor
  g1282
  (
    n1194,
    n801,
    n485,
    n950,
    n452
  );


  or
  g1283
  (
    n1228,
    n802,
    n859,
    n1103,
    n506
  );


  nor
  g1284
  (
    n1237,
    n858,
    n566,
    n911,
    n1026
  );


  xor
  g1285
  (
    n1261,
    n479,
    n1016,
    n1049,
    n1012
  );


  or
  g1286
  (
    n1281,
    n409,
    n723,
    n763,
    n329
  );


  or
  g1287
  (
    n1207,
    n611,
    n389,
    n881,
    n622
  );


  xor
  g1288
  (
    n1226,
    n957,
    n1066,
    n392,
    n469
  );


  xor
  g1289
  (
    n1334,
    n532,
    n412,
    n882,
    n722
  );


  and
  g1290
  (
    n1332,
    n823,
    n839,
    n1053,
    n395
  );


  and
  g1291
  (
    n1196,
    n917,
    n569,
    n543,
    n539
  );


  nor
  g1292
  (
    n1200,
    n1046,
    n717,
    n866,
    n988
  );


  nand
  g1293
  (
    n1220,
    n987,
    n778,
    n888,
    n1009
  );


  xor
  g1294
  (
    n1286,
    n1039,
    n675,
    n660,
    n414
  );


  xor
  g1295
  (
    n1155,
    n643,
    n754,
    n781,
    n767
  );


  and
  g1296
  (
    n1219,
    n788,
    n382,
    n836,
    n956
  );


  and
  g1297
  (
    n1229,
    n856,
    n578,
    n481,
    n1061
  );


  xnor
  g1298
  (
    n1257,
    n1048,
    n854,
    n509,
    n863
  );


  xor
  g1299
  (
    n1140,
    n714,
    n351,
    n654,
    n898
  );


  or
  g1300
  (
    n1275,
    n397,
    n403,
    n390,
    n803
  );


  xnor
  g1301
  (
    n1182,
    n620,
    n913,
    n949,
    n840
  );


  buf
  g1302
  (
    n1337,
    n1146
  );


  not
  g1303
  (
    n1344,
    n1145
  );


  not
  g1304
  (
    n1345,
    n1150
  );


  buf
  g1305
  (
    n1348,
    n1141
  );


  not
  g1306
  (
    n1347,
    n1152
  );


  not
  g1307
  (
    n1336,
    n1149
  );


  buf
  g1308
  (
    n1346,
    n1156
  );


  not
  g1309
  (
    n1341,
    n1144
  );


  not
  g1310
  (
    n1342,
    n1158
  );


  buf
  g1311
  (
    n1343,
    n1155
  );


  buf
  g1312
  (
    n1339,
    n1142
  );


  xnor
  g1313
  (
    n1335,
    n1151,
    n1148,
    n1143
  );


  xnor
  g1314
  (
    n1338,
    n1159,
    n1153,
    n1140,
    n1157
  );


  or
  g1315
  (
    n1340,
    n1154,
    n1147,
    n1161,
    n1160
  );


  nand
  g1316
  (
    n1350,
    n1116,
    n319,
    n1339,
    n1113
  );


  nor
  g1317
  (
    n1353,
    n318,
    n1337,
    n1111
  );


  or
  g1318
  (
    n1358,
    n321,
    n1118,
    n320,
    n1338
  );


  xor
  g1319
  (
    n1352,
    n1105,
    n1338,
    n319,
    n1115
  );


  nand
  g1320
  (
    n1349,
    n1121,
    n1112,
    n319,
    n320
  );


  xnor
  g1321
  (
    n1356,
    n1109,
    n320,
    n1114,
    n1335
  );


  nor
  g1322
  (
    n1357,
    n1120,
    n1107,
    n1117,
    n319
  );


  or
  g1323
  (
    n1355,
    n1106,
    n1110,
    n1108,
    n1338
  );


  nor
  g1324
  (
    n1351,
    n1338,
    n318,
    n320
  );


  nor
  g1325
  (
    n1354,
    n1337,
    n318,
    n1119,
    n1336
  );


  not
  g1326
  (
    n1359,
    n1349
  );


  and
  g1327
  (
    n1361,
    n1170,
    n1163,
    n1162,
    n1167
  );


  xnor
  g1328
  (
    n1362,
    n1169,
    n1165,
    n1359,
    n1168
  );


  xor
  g1329
  (
    n1360,
    n1164,
    n1359,
    n1166
  );


  xor
  g1330
  (
    n1364,
    n1199,
    n1186,
    n1361,
    n1178
  );


  nor
  g1331
  (
    n1371,
    n1181,
    n1193,
    n1360,
    n1177
  );


  nand
  g1332
  (
    n1366,
    n1176,
    n1203,
    n1184,
    n1204
  );


  xor
  g1333
  (
    n1373,
    n1196,
    n1185,
    n1179,
    n1360
  );


  nor
  g1334
  (
    n1368,
    n1190,
    n1202,
    n1197,
    n1200
  );


  nand
  g1335
  (
    n1370,
    n1361,
    n1194,
    n1189,
    n1174
  );


  xor
  g1336
  (
    n1363,
    n1362,
    n1188,
    n1205,
    n1192
  );


  nand
  g1337
  (
    n1372,
    n1361,
    n1171,
    n1362,
    n1172
  );


  xnor
  g1338
  (
    n1369,
    n1362,
    n1180,
    n1173,
    n1360
  );


  xor
  g1339
  (
    n1367,
    n1175,
    n1183,
    n1182,
    n1187
  );


  nand
  g1340
  (
    n1365,
    n1362,
    n1360,
    n1361,
    n1191
  );


  or
  g1341
  (
    n1374,
    n1198,
    n1195,
    n1201,
    n1206
  );


  nand
  g1342
  (
    n1375,
    n1363,
    n6,
    n5
  );


  or
  g1343
  (
    n1377,
    n48,
    n1375,
    n49,
    n47
  );


  nand
  g1344
  (
    n1376,
    n1375,
    n48
  );


  xnor
  g1345
  (
    n1378,
    n109,
    n106,
    n108,
    n1376
  );


  nor
  g1346
  (
    n1380,
    n1376,
    n105,
    n1377
  );


  xor
  g1347
  (
    n1382,
    n104,
    n106,
    n108,
    n1377
  );


  xnor
  g1348
  (
    n1384,
    n109,
    n105,
    n107
  );


  nor
  g1349
  (
    n1383,
    n1377,
    n108,
    n107,
    n109
  );


  nor
  g1350
  (
    n1379,
    n1376,
    n106,
    n105
  );


  or
  g1351
  (
    n1381,
    n109,
    n1377,
    n107,
    n108
  );


  nand
  g1352
  (
    n1385,
    n324,
    n322,
    n323
  );


  nor
  g1353
  (
    n1388,
    n1382,
    n323,
    n1380
  );


  xor
  g1354
  (
    n1387,
    n321,
    n1379,
    n1381,
    n322
  );


  xor
  g1355
  (
    n1389,
    n324,
    n1378,
    n321
  );


  or
  g1356
  (
    n1386,
    n323,
    n324,
    n322
  );


  not
  g1357
  (
    n1392,
    n1123
  );


  xnor
  g1358
  (
    n1390,
    n1124,
    n1126,
    n1388
  );


  and
  g1359
  (
    n1391,
    n1389,
    n1122,
    n1125,
    n1387
  );


  xnor
  g1360
  (
    n1399,
    n1226,
    n1211,
    n1207,
    n1216
  );


  or
  g1361
  (
    n1401,
    n1232,
    n1224,
    n1208,
    n1218
  );


  or
  g1362
  (
    n1396,
    n1219,
    n1390,
    n1209,
    n1210
  );


  xnor
  g1363
  (
    n1400,
    n1214,
    n1391,
    n1215
  );


  nand
  g1364
  (
    n1395,
    n1390,
    n1227,
    n1391,
    n1221
  );


  xor
  g1365
  (
    n1397,
    n1213,
    n1217,
    n1231,
    n1228
  );


  nor
  g1366
  (
    n1393,
    n1229,
    n1212,
    n1223,
    n1233
  );


  and
  g1367
  (
    n1394,
    n1392,
    n1230,
    n1390
  );


  xor
  g1368
  (
    n1398,
    n1391,
    n1220,
    n1225,
    n1222
  );


  buf
  g1369
  (
    n1402,
    n1399
  );


  not
  g1370
  (
    n1403,
    n1398
  );


  buf
  g1371
  (
    n1407,
    n1395
  );


  buf
  g1372
  (
    n1406,
    n1396
  );


  not
  g1373
  (
    n1405,
    n1397
  );


  buf
  g1374
  (
    n1404,
    n1394
  );


  xnor
  g1375
  (
    n1408,
    n1236,
    n1238,
    n1402,
    n1355
  );


  and
  g1376
  (
    n1410,
    n1356,
    n1357,
    n1403,
    n1352
  );


  nand
  g1377
  (
    n1412,
    n1235,
    n1237,
    n1354,
    n1402
  );


  xnor
  g1378
  (
    n1411,
    n1353,
    n1234,
    n1402
  );


  and
  g1379
  (
    n1409,
    n1239,
    n1350,
    n1358,
    n1351
  );


  buf
  g1380
  (
    n1416,
    n1412
  );


  buf
  g1381
  (
    n1415,
    n1409
  );


  not
  g1382
  (
    n1413,
    n1411
  );


  not
  g1383
  (
    n1414,
    n1410
  );


  not
  g1384
  (
    n1417,
    n1244
  );


  not
  g1385
  (
    n1427,
    n1415
  );


  buf
  g1386
  (
    n1421,
    n1415
  );


  buf
  g1387
  (
    n1419,
    n1414
  );


  buf
  g1388
  (
    n1431,
    n1416
  );


  not
  g1389
  (
    n1418,
    n1416
  );


  buf
  g1390
  (
    n1422,
    n1250
  );


  not
  g1391
  (
    n1432,
    n1242
  );


  buf
  g1392
  (
    n1428,
    n1252
  );


  buf
  g1393
  (
    n1430,
    n1253
  );


  not
  g1394
  (
    n1429,
    n1243
  );


  nor
  g1395
  (
    n1425,
    n1415,
    n1254,
    n1414,
    n1245
  );


  xnor
  g1396
  (
    n1420,
    n1413,
    n1416,
    n1414
  );


  xor
  g1397
  (
    n1424,
    n1414,
    n1241,
    n1246,
    n1249
  );


  or
  g1398
  (
    n1426,
    n1240,
    n1413,
    n1248
  );


  xor
  g1399
  (
    n1423,
    n1247,
    n1415,
    n1413,
    n1251
  );


  not
  g1400
  (
    n1435,
    n1421
  );


  xor
  g1401
  (
    n1439,
    n1366,
    n1417,
    n1419,
    n1373
  );


  and
  g1402
  (
    n1438,
    n1367,
    n1365,
    n1366,
    n1368
  );


  xor
  g1403
  (
    n1449,
    n1371,
    n1374,
    n1364,
    n1370
  );


  nand
  g1404
  (
    n1441,
    n1369,
    n1369,
    n1368,
    n1364
  );


  or
  g1405
  (
    n1436,
    n1420,
    n1367,
    n1417,
    n1371
  );


  xnor
  g1406
  (
    n1444,
    n1417,
    n1373,
    n1365,
    n1418
  );


  xor
  g1407
  (
    n1448,
    n1371,
    n1364,
    n1419,
    n1417
  );


  xnor
  g1408
  (
    n1440,
    n1367,
    n1374,
    n1363,
    n1369
  );


  nor
  g1409
  (
    n1443,
    n1255,
    n1373,
    n1419
  );


  nor
  g1410
  (
    n1433,
    n1363,
    n1372,
    n1370,
    n1365
  );


  nor
  g1411
  (
    n1446,
    n1420,
    n1371,
    n1368,
    n1374
  );


  nand
  g1412
  (
    n1445,
    n1370,
    n1372,
    n1420,
    n1363
  );


  and
  g1413
  (
    n1447,
    n1367,
    n1418,
    n1372,
    n1373
  );


  nor
  g1414
  (
    n1442,
    n1418,
    n1370,
    n1369,
    n1368
  );


  nor
  g1415
  (
    n1437,
    n1420,
    n1364,
    n1365,
    n1366
  );


  nand
  g1416
  (
    n1434,
    n1372,
    n1374,
    n1418,
    n1366
  );


  and
  g1417
  (
    n1457,
    n1139,
    n1272,
    n1282,
    n1276
  );


  nor
  g1418
  (
    n1458,
    n1266,
    n1284,
    n1436
  );


  xor
  g1419
  (
    n1453,
    n1262,
    n1131,
    n1434,
    n1433
  );


  nand
  g1420
  (
    n1454,
    n1128,
    n1137,
    n1436,
    n1434
  );


  nand
  g1421
  (
    n1464,
    n1271,
    n1259,
    n1277,
    n1433
  );


  or
  g1422
  (
    n1459,
    n1136,
    n1435,
    n1127,
    n1132
  );


  and
  g1423
  (
    n1463,
    n1275,
    n1433,
    n1273,
    n1285
  );


  xnor
  g1424
  (
    n1456,
    n1267,
    n1129,
    n1286,
    n1134
  );


  nor
  g1425
  (
    n1452,
    n1133,
    n1281,
    n1274,
    n1264
  );


  and
  g1426
  (
    n1455,
    n1287,
    n1278,
    n1130,
    n1435
  );


  xor
  g1427
  (
    n1462,
    n1435,
    n1256,
    n1279,
    n1268
  );


  nor
  g1428
  (
    n1460,
    n1270,
    n1435,
    n1269,
    n1260
  );


  or
  g1429
  (
    n1450,
    n1433,
    n1138,
    n1280,
    n1263
  );


  xor
  g1430
  (
    n1461,
    n1434,
    n1261,
    n1283,
    n1265
  );


  xnor
  g1431
  (
    n1451,
    n1135,
    n1258,
    n1257,
    n1434
  );


  nand
  g1432
  (
    n1465,
    n1293,
    n1450,
    n1292,
    n1451
  );


  xor
  g1433
  (
    n1466,
    n1291,
    n1289,
    n1290,
    n1288
  );


  nor
  g1434
  (
    n1469,
    n1466,
    n1465,
    n1383,
    n1294
  );


  nand
  g1435
  (
    n1470,
    n1296,
    n1297,
    n1465,
    n1300
  );


  xor
  g1436
  (
    n1472,
    n1466,
    n1307,
    n1309,
    n1465
  );


  nor
  g1437
  (
    n1471,
    n1306,
    n1465,
    n1298,
    n1302
  );


  and
  g1438
  (
    n1468,
    n1304,
    n1301,
    n1305,
    n1308
  );


  or
  g1439
  (
    n1467,
    n1384,
    n1303,
    n1295,
    n1299
  );


  not
  g1440
  (
    n1480,
    n1346
  );


  buf
  g1441
  (
    n1485,
    n1346
  );


  buf
  g1442
  (
    n1488,
    n1343
  );


  buf
  g1443
  (
    n1487,
    n1469
  );


  not
  g1444
  (
    n1483,
    n1339
  );


  buf
  g1445
  (
    n1473,
    n1344
  );


  buf
  g1446
  (
    n1495,
    n1345
  );


  not
  g1447
  (
    n1493,
    n1347
  );


  not
  g1448
  (
    n1492,
    n1310
  );


  buf
  g1449
  (
    KeyWire_0_24,
    n1345
  );


  xnor
  g1450
  (
    n1490,
    n1342,
    n1348,
    n1341
  );


  xnor
  g1451
  (
    n1482,
    n1346,
    n1468,
    n1342
  );


  nor
  g1452
  (
    n1489,
    n1347,
    n1347,
    n1344,
    n1311
  );


  or
  g1453
  (
    n1478,
    n1341,
    n1470,
    n1345,
    n1467
  );


  nand
  g1454
  (
    n1477,
    n1342,
    n1340,
    n1346,
    n1472
  );


  nor
  g1455
  (
    n1486,
    n1472,
    n1344,
    n1468,
    n1467
  );


  xnor
  g1456
  (
    n1496,
    n1344,
    n1467,
    n1347,
    n1469
  );


  and
  g1457
  (
    n1475,
    n1470,
    n1345,
    n1341,
    n1340
  );


  xor
  g1458
  (
    n1474,
    n1339,
    n1471,
    n1467,
    n1343
  );


  or
  g1459
  (
    n1481,
    n1342,
    n1343,
    n1472
  );


  nand
  g1460
  (
    n1491,
    n1471,
    n1340,
    n1470,
    n1343
  );


  nand
  g1461
  (
    n1494,
    n1469,
    n1470,
    n1340,
    n1339
  );


  xnor
  g1462
  (
    n1479,
    n1348,
    n1471,
    n1341
  );


  and
  g1463
  (
    n1476,
    n1312,
    n1469,
    n1348,
    n1468
  );


  not
  g1464
  (
    n1539,
    n1482
  );


  buf
  g1465
  (
    n1556,
    n1473
  );


  not
  g1466
  (
    n1561,
    n1495
  );


  buf
  g1467
  (
    n1533,
    n1489
  );


  buf
  g1468
  (
    n1507,
    n1484
  );


  not
  g1469
  (
    n1528,
    n1494
  );


  not
  g1470
  (
    n1515,
    n1475
  );


  not
  g1471
  (
    n1529,
    n1475
  );


  buf
  g1472
  (
    n1564,
    n1457
  );


  not
  g1473
  (
    n1558,
    n1475
  );


  buf
  g1474
  (
    n1551,
    n1457
  );


  buf
  g1475
  (
    n1544,
    n1494
  );


  not
  g1476
  (
    n1572,
    n1488
  );


  buf
  g1477
  (
    n1583,
    n1488
  );


  not
  g1478
  (
    n1511,
    n1495
  );


  not
  g1479
  (
    n1549,
    n1496
  );


  not
  g1480
  (
    n1559,
    n1484
  );


  buf
  g1481
  (
    n1523,
    n1392
  );


  not
  g1482
  (
    n1504,
    n1492
  );


  buf
  g1483
  (
    n1568,
    n1478
  );


  not
  g1484
  (
    n1498,
    n1452
  );


  not
  g1485
  (
    n1554,
    n1392
  );


  not
  g1486
  (
    n1553,
    n1455
  );


  not
  g1487
  (
    n1542,
    n1485
  );


  buf
  g1488
  (
    n1503,
    n1488
  );


  not
  g1489
  (
    n1582,
    n1491
  );


  not
  g1490
  (
    n1545,
    n1487
  );


  buf
  g1491
  (
    n1508,
    n1477
  );


  buf
  g1492
  (
    n1532,
    n1474
  );


  not
  g1493
  (
    n1519,
    n1454
  );


  not
  g1494
  (
    n1500,
    n1473
  );


  not
  g1495
  (
    n1586,
    n1496
  );


  buf
  g1496
  (
    n1563,
    n1474
  );


  buf
  g1497
  (
    n1514,
    n1457
  );


  buf
  g1498
  (
    n1566,
    n1478
  );


  not
  g1499
  (
    n1527,
    n1487
  );


  not
  g1500
  (
    n1509,
    n1487
  );


  not
  g1501
  (
    n1587,
    n1490
  );


  not
  g1502
  (
    n1591,
    n1481
  );


  buf
  g1503
  (
    n1578,
    n1482
  );


  not
  g1504
  (
    n1524,
    n1480
  );


  not
  g1505
  (
    n1567,
    n1485
  );


  not
  g1506
  (
    n1522,
    n1477
  );


  not
  g1507
  (
    n1569,
    n1482
  );


  buf
  g1508
  (
    n1520,
    n1456
  );


  not
  g1509
  (
    n1534,
    n1493
  );


  not
  g1510
  (
    n1497,
    n1476
  );


  buf
  g1511
  (
    n1562,
    n1479
  );


  buf
  g1512
  (
    n1547,
    n1491
  );


  not
  g1513
  (
    n1525,
    n1479
  );


  not
  g1514
  (
    n1512,
    n1455
  );


  not
  g1515
  (
    n1555,
    n1483
  );


  buf
  g1516
  (
    n1576,
    n1491
  );


  not
  g1517
  (
    n1573,
    n1476
  );


  not
  g1518
  (
    n1537,
    n1474
  );


  not
  g1519
  (
    n1588,
    n1489
  );


  not
  g1520
  (
    n1536,
    n1456
  );


  not
  g1521
  (
    n1552,
    n1476
  );


  buf
  g1522
  (
    n1510,
    n1486
  );


  buf
  g1523
  (
    n1592,
    n1481
  );


  buf
  g1524
  (
    n1543,
    n1457
  );


  buf
  g1525
  (
    n1550,
    n1495
  );


  not
  g1526
  (
    n1506,
    n1478
  );


  buf
  g1527
  (
    n1584,
    n1481
  );


  buf
  g1528
  (
    n1548,
    n1479
  );


  not
  g1529
  (
    KeyWire_0_8,
    n1492
  );


  not
  g1530
  (
    n1560,
    n1488
  );


  not
  g1531
  (
    n1557,
    n1493
  );


  buf
  g1532
  (
    n1521,
    n1473
  );


  not
  g1533
  (
    n1535,
    n1494
  );


  not
  g1534
  (
    n1540,
    n1477
  );


  not
  g1535
  (
    n1570,
    n1487
  );


  buf
  g1536
  (
    n1574,
    n1478
  );


  not
  g1537
  (
    n1501,
    n1474
  );


  and
  g1538
  (
    n1546,
    n1480,
    n1384
  );


  or
  g1539
  (
    n1579,
    n1456,
    n1485
  );


  nor
  g1540
  (
    n1577,
    n1493,
    n1495
  );


  xnor
  g1541
  (
    n1502,
    n1489,
    n1482
  );


  nor
  g1542
  (
    n1518,
    n1458,
    n1454
  );


  nand
  g1543
  (
    n1590,
    n1484,
    n1486
  );


  xor
  g1544
  (
    n1575,
    n1483,
    n1491
  );


  nor
  g1545
  (
    n1530,
    n1492,
    n1477
  );


  and
  g1546
  (
    n1531,
    n1490,
    n1496
  );


  xnor
  g1547
  (
    n1516,
    n1455,
    n1490
  );


  nor
  g1548
  (
    n1581,
    n1480,
    n1392
  );


  and
  g1549
  (
    n1538,
    n1486,
    n1473
  );


  nor
  g1550
  (
    n1589,
    n1476,
    n1453
  );


  nand
  g1551
  (
    n1585,
    n1475,
    n1456
  );


  xor
  g1552
  (
    n1505,
    n1454,
    n1496
  );


  xnor
  g1553
  (
    n1499,
    n1493,
    n1483
  );


  and
  g1554
  (
    n1513,
    n1486,
    n1484
  );


  xor
  g1555
  (
    n1541,
    n1490,
    n1483
  );


  xnor
  g1556
  (
    n1517,
    n1494,
    n1458
  );


  xnor
  g1557
  (
    n1565,
    n1489,
    n1480
  );


  nand
  g1558
  (
    n1526,
    n1492,
    n1485
  );


  xor
  g1559
  (
    n1580,
    n1481,
    n1479
  );


  not
  g1560
  (
    n1895,
    n1549
  );


  not
  g1561
  (
    n1713,
    n1578
  );


  not
  g1562
  (
    n1644,
    n1522
  );


  buf
  g1563
  (
    n1839,
    n1520
  );


  buf
  g1564
  (
    n1798,
    n1545
  );


  not
  g1565
  (
    n1942,
    n1531
  );


  buf
  g1566
  (
    n1681,
    n1516
  );


  buf
  g1567
  (
    n1629,
    n1532
  );


  not
  g1568
  (
    n1807,
    n1543
  );


  buf
  g1569
  (
    n1675,
    n1458
  );


  not
  g1570
  (
    n1828,
    n1508
  );


  buf
  g1571
  (
    n1919,
    n1526
  );


  not
  g1572
  (
    n1750,
    n1527
  );


  buf
  g1573
  (
    n1599,
    n1554
  );


  buf
  g1574
  (
    n1617,
    n1550
  );


  not
  g1575
  (
    n1641,
    n1568
  );


  not
  g1576
  (
    n1834,
    n1511
  );


  not
  g1577
  (
    n1817,
    n1558
  );


  not
  g1578
  (
    n1647,
    n1553
  );


  buf
  g1579
  (
    n1646,
    n1576
  );


  buf
  g1580
  (
    n1862,
    n1553
  );


  not
  g1581
  (
    n1913,
    n1325
  );


  not
  g1582
  (
    n1855,
    n1538
  );


  not
  g1583
  (
    n1692,
    n1511
  );


  not
  g1584
  (
    n1931,
    n1556
  );


  not
  g1585
  (
    n1915,
    n1507
  );


  not
  g1586
  (
    n1593,
    n1513
  );


  buf
  g1587
  (
    n1604,
    n1572
  );


  buf
  g1588
  (
    n1718,
    n1534
  );


  buf
  g1589
  (
    n1687,
    n1518
  );


  buf
  g1590
  (
    n1638,
    n1524
  );


  buf
  g1591
  (
    n1914,
    n1519
  );


  not
  g1592
  (
    n1916,
    n1585
  );


  not
  g1593
  (
    n1694,
    n1540
  );


  not
  g1594
  (
    n1655,
    n1577
  );


  buf
  g1595
  (
    n1661,
    n1545
  );


  buf
  g1596
  (
    n1634,
    n1556
  );


  buf
  g1597
  (
    n1933,
    n1557
  );


  not
  g1598
  (
    n1753,
    n1574
  );


  buf
  g1599
  (
    n1632,
    n1507
  );


  buf
  g1600
  (
    n1899,
    n1577
  );


  buf
  g1601
  (
    n1596,
    n1550
  );


  buf
  g1602
  (
    n1875,
    n1567
  );


  buf
  g1603
  (
    n1935,
    n1544
  );


  not
  g1604
  (
    n1723,
    n1561
  );


  buf
  g1605
  (
    n1722,
    n1562
  );


  not
  g1606
  (
    n1643,
    n1314
  );


  buf
  g1607
  (
    n1921,
    n1528
  );


  buf
  g1608
  (
    n1946,
    n1460
  );


  not
  g1609
  (
    n1835,
    n1558
  );


  buf
  g1610
  (
    n1937,
    n1535
  );


  buf
  g1611
  (
    n1755,
    n1518
  );


  buf
  g1612
  (
    n1699,
    n1580
  );


  buf
  g1613
  (
    n1944,
    n1461
  );


  not
  g1614
  (
    n1806,
    n1568
  );


  not
  g1615
  (
    n1735,
    n1547
  );


  not
  g1616
  (
    n1633,
    n1500
  );


  buf
  g1617
  (
    n1668,
    n1316
  );


  buf
  g1618
  (
    n1748,
    n1546
  );


  buf
  g1619
  (
    n1702,
    n1560
  );


  buf
  g1620
  (
    n1866,
    n1565
  );


  not
  g1621
  (
    n1832,
    n1568
  );


  buf
  g1622
  (
    n1901,
    n1459
  );


  buf
  g1623
  (
    n1628,
    n1535
  );


  buf
  g1624
  (
    n1867,
    n1548
  );


  not
  g1625
  (
    n1793,
    n1503
  );


  buf
  g1626
  (
    n1622,
    n1542
  );


  not
  g1627
  (
    n1701,
    n1570
  );


  buf
  g1628
  (
    n1816,
    n1552
  );


  not
  g1629
  (
    n1686,
    n1525
  );


  buf
  g1630
  (
    n1877,
    n1463
  );


  not
  g1631
  (
    n1890,
    n1554
  );


  not
  g1632
  (
    n1613,
    n1528
  );


  buf
  g1633
  (
    n1665,
    n1575
  );


  not
  g1634
  (
    n1853,
    n1512
  );


  buf
  g1635
  (
    n1874,
    n1501
  );


  buf
  g1636
  (
    KeyWire_0_6,
    n1547
  );


  not
  g1637
  (
    n1651,
    n1567
  );


  not
  g1638
  (
    n1891,
    n1536
  );


  buf
  g1639
  (
    n1889,
    n1520
  );


  not
  g1640
  (
    n1873,
    n1538
  );


  not
  g1641
  (
    n1941,
    n1581
  );


  buf
  g1642
  (
    n1637,
    n1498
  );


  buf
  g1643
  (
    n1690,
    n1315
  );


  not
  g1644
  (
    n1685,
    n1558
  );


  not
  g1645
  (
    n1598,
    n1323
  );


  not
  g1646
  (
    n1905,
    n1499
  );


  not
  g1647
  (
    n1934,
    n1579
  );


  buf
  g1648
  (
    n1765,
    n1529
  );


  buf
  g1649
  (
    n1715,
    n1577
  );


  buf
  g1650
  (
    n1773,
    n1576
  );


  buf
  g1651
  (
    n1801,
    n1539
  );


  buf
  g1652
  (
    n1739,
    n1563
  );


  buf
  g1653
  (
    n1659,
    n1573
  );


  buf
  g1654
  (
    n1923,
    n1566
  );


  buf
  g1655
  (
    n1927,
    n1509
  );


  buf
  g1656
  (
    n1671,
    n1504
  );


  not
  g1657
  (
    n1908,
    n1497
  );


  buf
  g1658
  (
    n1782,
    n1511
  );


  buf
  g1659
  (
    n1707,
    n1527
  );


  buf
  g1660
  (
    n1597,
    n1546
  );


  not
  g1661
  (
    n1683,
    n1533
  );


  buf
  g1662
  (
    n1907,
    n1505
  );


  buf
  g1663
  (
    n1612,
    n1580
  );


  buf
  g1664
  (
    n1682,
    n1564
  );


  not
  g1665
  (
    n1814,
    n1561
  );


  not
  g1666
  (
    n1654,
    n1463
  );


  buf
  g1667
  (
    n1911,
    n1573
  );


  buf
  g1668
  (
    n1666,
    n1502
  );


  not
  g1669
  (
    n1872,
    n1549
  );


  not
  g1670
  (
    n1880,
    n1531
  );


  buf
  g1671
  (
    n1850,
    n1513
  );


  buf
  g1672
  (
    n1627,
    n1531
  );


  not
  g1673
  (
    n1887,
    n1566
  );


  buf
  g1674
  (
    n1805,
    n1499
  );


  buf
  g1675
  (
    n1714,
    n1512
  );


  not
  g1676
  (
    n1883,
    n1555
  );


  buf
  g1677
  (
    n1656,
    n1565
  );


  not
  g1678
  (
    n1840,
    n1571
  );


  not
  g1679
  (
    n1747,
    n1548
  );


  buf
  g1680
  (
    n1670,
    n1576
  );


  not
  g1681
  (
    n1838,
    n1584
  );


  buf
  g1682
  (
    n1885,
    n1552
  );


  not
  g1683
  (
    n1625,
    n1579
  );


  not
  g1684
  (
    n1712,
    n1517
  );


  buf
  g1685
  (
    n1772,
    n1459
  );


  buf
  g1686
  (
    n1710,
    n1508
  );


  not
  g1687
  (
    n1815,
    n1534
  );


  not
  g1688
  (
    n1876,
    n1569
  );


  buf
  g1689
  (
    n1930,
    n1530
  );


  not
  g1690
  (
    n1928,
    n1534
  );


  buf
  g1691
  (
    n1785,
    n1551
  );


  buf
  g1692
  (
    n1726,
    n1546
  );


  buf
  g1693
  (
    n1909,
    n1545
  );


  not
  g1694
  (
    n1878,
    n1460
  );


  buf
  g1695
  (
    n1653,
    n1526
  );


  not
  g1696
  (
    n1818,
    n1569
  );


  not
  g1697
  (
    n1757,
    n1585
  );


  buf
  g1698
  (
    n1938,
    n1332
  );


  not
  g1699
  (
    n1730,
    n1517
  );


  not
  g1700
  (
    n1809,
    n1568
  );


  not
  g1701
  (
    n1594,
    n1559
  );


  not
  g1702
  (
    n1775,
    n1519
  );


  not
  g1703
  (
    n1849,
    n1580
  );


  not
  g1704
  (
    n1679,
    n1584
  );


  buf
  g1705
  (
    n1879,
    n1541
  );


  not
  g1706
  (
    n1852,
    n1564
  );


  not
  g1707
  (
    n1871,
    n1329
  );


  buf
  g1708
  (
    n1920,
    n1526
  );


  not
  g1709
  (
    n1642,
    n1563
  );


  not
  g1710
  (
    n1733,
    n1509
  );


  buf
  g1711
  (
    n1897,
    n1573
  );


  not
  g1712
  (
    n1759,
    n1525
  );


  buf
  g1713
  (
    n1618,
    n1527
  );


  buf
  g1714
  (
    n1658,
    n1498
  );


  buf
  g1715
  (
    n1760,
    n1515
  );


  buf
  g1716
  (
    n1774,
    n1531
  );


  buf
  g1717
  (
    n1746,
    n1554
  );


  not
  g1718
  (
    n1904,
    n1514
  );


  not
  g1719
  (
    n1764,
    n1581
  );


  buf
  g1720
  (
    n1900,
    n1508
  );


  not
  g1721
  (
    n1940,
    n1505
  );


  not
  g1722
  (
    n1893,
    n1558
  );


  buf
  g1723
  (
    n1766,
    n1516
  );


  not
  g1724
  (
    n1886,
    n1400
  );


  not
  g1725
  (
    n1922,
    n1578
  );


  buf
  g1726
  (
    n1894,
    n1510
  );


  not
  g1727
  (
    n1619,
    n1503
  );


  not
  g1728
  (
    n1906,
    n1560
  );


  buf
  g1729
  (
    n1860,
    n1575
  );


  buf
  g1730
  (
    n1945,
    n1321
  );


  not
  g1731
  (
    n1822,
    n1501
  );


  not
  g1732
  (
    n1608,
    n1554
  );


  buf
  g1733
  (
    n1736,
    n1560
  );


  buf
  g1734
  (
    n1856,
    n1532
  );


  buf
  g1735
  (
    n1667,
    n1567
  );


  buf
  g1736
  (
    n1819,
    n1575
  );


  not
  g1737
  (
    n1721,
    n1511
  );


  not
  g1738
  (
    n1803,
    n1319
  );


  buf
  g1739
  (
    n1776,
    n1566
  );


  buf
  g1740
  (
    n1826,
    n1463
  );


  buf
  g1741
  (
    n1657,
    n1515
  );


  not
  g1742
  (
    n1607,
    n1317
  );


  not
  g1743
  (
    n1680,
    n1530
  );


  not
  g1744
  (
    n1851,
    n1572
  );


  not
  g1745
  (
    n1892,
    n1524
  );


  buf
  g1746
  (
    n1800,
    n1509
  );


  buf
  g1747
  (
    n1729,
    n1541
  );


  buf
  g1748
  (
    n1863,
    n1530
  );


  buf
  g1749
  (
    n1844,
    n1561
  );


  not
  g1750
  (
    n1770,
    n1566
  );


  not
  g1751
  (
    n1827,
    n1322
  );


  not
  g1752
  (
    n1903,
    n1549
  );


  buf
  g1753
  (
    n1859,
    n1550
  );


  not
  g1754
  (
    n1898,
    n1581
  );


  not
  g1755
  (
    n1868,
    n1561
  );


  not
  g1756
  (
    n1756,
    n1518
  );


  buf
  g1757
  (
    n1896,
    n1559
  );


  not
  g1758
  (
    n1724,
    n1510
  );


  buf
  g1759
  (
    n1857,
    n1562
  );


  buf
  g1760
  (
    KeyWire_0_3,
    n1536
  );


  not
  g1761
  (
    n1698,
    n1552
  );


  buf
  g1762
  (
    n1912,
    n1463
  );


  buf
  g1763
  (
    n1881,
    n1540
  );


  not
  g1764
  (
    n1663,
    n1528
  );


  buf
  g1765
  (
    n1623,
    n1553
  );


  buf
  g1766
  (
    n1674,
    n1461
  );


  buf
  g1767
  (
    n1652,
    n1544
  );


  not
  g1768
  (
    n1631,
    n1573
  );


  not
  g1769
  (
    n1791,
    n1517
  );


  not
  g1770
  (
    n1693,
    n1553
  );


  buf
  g1771
  (
    n1762,
    n1571
  );


  buf
  g1772
  (
    n1639,
    n1327
  );


  buf
  g1773
  (
    n1910,
    n1509
  );


  buf
  g1774
  (
    n1783,
    n1535
  );


  buf
  g1775
  (
    n1917,
    n1559
  );


  not
  g1776
  (
    n1741,
    n1522
  );


  buf
  g1777
  (
    n1595,
    n1462
  );


  not
  g1778
  (
    n1833,
    n1462
  );


  not
  g1779
  (
    n1810,
    n1574
  );


  not
  g1780
  (
    n1869,
    n1578
  );


  not
  g1781
  (
    n1734,
    n1540
  );


  buf
  g1782
  (
    n1700,
    n1582
  );


  not
  g1783
  (
    n1605,
    n1512
  );


  not
  g1784
  (
    n1697,
    n1548
  );


  not
  g1785
  (
    n1610,
    n1556
  );


  buf
  g1786
  (
    n1602,
    n1583
  );


  buf
  g1787
  (
    n1843,
    n1510
  );


  not
  g1788
  (
    n1794,
    n1533
  );


  buf
  g1789
  (
    n1708,
    n1536
  );


  not
  g1790
  (
    n1790,
    n1584
  );


  not
  g1791
  (
    n1813,
    n1460
  );


  buf
  g1792
  (
    n1695,
    n1503
  );


  not
  g1793
  (
    n1858,
    n1500
  );


  not
  g1794
  (
    n1751,
    n1550
  );


  not
  g1795
  (
    n1768,
    n1542
  );


  not
  g1796
  (
    n1796,
    n1523
  );


  not
  g1797
  (
    n1600,
    n1521
  );


  buf
  g1798
  (
    n1669,
    n1501
  );


  buf
  g1799
  (
    n1821,
    n1466
  );


  not
  g1800
  (
    n1609,
    n1543
  );


  not
  g1801
  (
    n1846,
    n1502
  );


  not
  g1802
  (
    n1672,
    n1557
  );


  buf
  g1803
  (
    n1703,
    n1581
  );


  not
  g1804
  (
    n1836,
    n1569
  );


  buf
  g1805
  (
    n1688,
    n1500
  );


  not
  g1806
  (
    n1924,
    n1580
  );


  buf
  g1807
  (
    n1728,
    n1570
  );


  buf
  g1808
  (
    KeyWire_0_9,
    n1579
  );


  buf
  g1809
  (
    n1635,
    n1520
  );


  not
  g1810
  (
    n1630,
    n1462
  );


  buf
  g1811
  (
    n1823,
    n1500
  );


  not
  g1812
  (
    n1740,
    n1549
  );


  buf
  g1813
  (
    n1926,
    n1498
  );


  buf
  g1814
  (
    n1706,
    n1584
  );


  buf
  g1815
  (
    n1673,
    n1497
  );


  buf
  g1816
  (
    n1788,
    n1502
  );


  not
  g1817
  (
    n1660,
    n1507
  );


  buf
  g1818
  (
    n1743,
    n1523
  );


  buf
  g1819
  (
    n1787,
    n1528
  );


  buf
  g1820
  (
    n1696,
    n1513
  );


  buf
  g1821
  (
    n1725,
    n1547
  );


  not
  g1822
  (
    n1731,
    n1540
  );


  buf
  g1823
  (
    n1689,
    n1564
  );


  buf
  g1824
  (
    n1779,
    n1577
  );


  not
  g1825
  (
    n1837,
    n1543
  );


  not
  g1826
  (
    n1615,
    n1506
  );


  buf
  g1827
  (
    n1749,
    n1535
  );


  buf
  g1828
  (
    n1704,
    n1331
  );


  not
  g1829
  (
    n1789,
    n1513
  );


  buf
  g1830
  (
    n1738,
    n1571
  );


  not
  g1831
  (
    n1611,
    n1565
  );


  buf
  g1832
  (
    n1888,
    n1330
  );


  not
  g1833
  (
    n1847,
    n1525
  );


  not
  g1834
  (
    n1830,
    n1582
  );


  not
  g1835
  (
    n1786,
    n1544
  );


  not
  g1836
  (
    n1603,
    n1537
  );


  not
  g1837
  (
    n1761,
    n1460
  );


  not
  g1838
  (
    n1781,
    n1514
  );


  not
  g1839
  (
    n1732,
    n1521
  );


  buf
  g1840
  (
    n1745,
    n1576
  );


  buf
  g1841
  (
    n1778,
    n1510
  );


  buf
  g1842
  (
    n1649,
    n1570
  );


  buf
  g1843
  (
    n1902,
    n1504
  );


  buf
  g1844
  (
    n1626,
    n1516
  );


  buf
  g1845
  (
    n1720,
    n1567
  );


  not
  g1846
  (
    n1829,
    n1521
  );


  buf
  g1847
  (
    n1936,
    n1542
  );


  buf
  g1848
  (
    n1754,
    n1541
  );


  buf
  g1849
  (
    n1716,
    n1541
  );


  not
  g1850
  (
    n1758,
    n1401
  );


  not
  g1851
  (
    n1705,
    n1506
  );


  buf
  g1852
  (
    n1767,
    n1506
  );


  buf
  g1853
  (
    n1865,
    n1514
  );


  not
  g1854
  (
    n1882,
    n1519
  );


  not
  g1855
  (
    n1691,
    n1326
  );


  buf
  g1856
  (
    n1709,
    n1548
  );


  not
  g1857
  (
    n1792,
    n1537
  );


  not
  g1858
  (
    n1645,
    n1505
  );


  buf
  g1859
  (
    n1820,
    n1459
  );


  buf
  g1860
  (
    n1744,
    n1514
  );


  buf
  g1861
  (
    n1808,
    n1582
  );


  buf
  g1862
  (
    KeyWire_0_31,
    n1530
  );


  buf
  g1863
  (
    n1648,
    n1538
  );


  buf
  g1864
  (
    n1664,
    n1571
  );


  not
  g1865
  (
    n1717,
    n1508
  );


  not
  g1866
  (
    n1662,
    n1519
  );


  not
  g1867
  (
    n1939,
    n1497
  );


  not
  g1868
  (
    n1918,
    n1570
  );


  not
  g1869
  (
    n1676,
    n1502
  );


  buf
  g1870
  (
    n1606,
    n1537
  );


  buf
  g1871
  (
    n1727,
    n1525
  );


  not
  g1872
  (
    n1684,
    n1499
  );


  buf
  g1873
  (
    n1802,
    n1520
  );


  not
  g1874
  (
    n1769,
    n1583
  );


  buf
  g1875
  (
    n1621,
    n1515
  );


  buf
  g1876
  (
    n1811,
    n1582
  );


  not
  g1877
  (
    n1884,
    n1526
  );


  not
  g1878
  (
    n1854,
    n1557
  );


  not
  g1879
  (
    n1825,
    n1515
  );


  not
  g1880
  (
    n1864,
    n1533
  );


  buf
  g1881
  (
    n1777,
    n1537
  );


  buf
  g1882
  (
    n1719,
    n1459
  );


  not
  g1883
  (
    n1799,
    n1328
  );


  not
  g1884
  (
    n1812,
    n1504
  );


  not
  g1885
  (
    n1848,
    n1527
  );


  buf
  g1886
  (
    n1737,
    n1507
  );


  not
  g1887
  (
    n1601,
    n1547
  );


  buf
  g1888
  (
    n1784,
    n1560
  );


  buf
  g1889
  (
    n1620,
    n1504
  );


  not
  g1890
  (
    n1870,
    n1574
  );


  buf
  g1891
  (
    n1842,
    n1522
  );


  buf
  g1892
  (
    n1742,
    n1461
  );


  buf
  g1893
  (
    n1929,
    n1461
  );


  not
  g1894
  (
    n1795,
    n1506
  );


  buf
  g1895
  (
    n1752,
    n1458
  );


  buf
  g1896
  (
    n1771,
    n1555
  );


  buf
  g1897
  (
    n1841,
    n1552
  );


  buf
  g1898
  (
    n1925,
    n1523
  );


  nor
  g1899
  (
    n1824,
    n1517,
    n1569,
    n1529,
    n1544
  );


  nor
  g1900
  (
    n1804,
    n1538,
    n1533,
    n1551,
    n1546
  );


  and
  g1901
  (
    n1616,
    n1320,
    n1574,
    n1555,
    n1578
  );


  or
  g1902
  (
    n1711,
    n1503,
    n1512,
    n1523,
    n1579
  );


  nor
  g1903
  (
    n1932,
    n1562,
    n1539,
    n1505,
    n1529
  );


  nand
  g1904
  (
    n1678,
    n1524,
    n1562,
    n1498,
    n1518
  );


  nand
  g1905
  (
    n1861,
    n1543,
    n1556,
    n1532,
    n1539
  );


  nor
  g1906
  (
    n1797,
    n1583,
    n1524,
    n1575,
    n1539
  );


  nand
  g1907
  (
    n1677,
    n1551,
    n1529,
    n1563,
    n1313
  );


  or
  g1908
  (
    n1640,
    n1572,
    n1462,
    n1497,
    n1583
  );


  or
  g1909
  (
    n1845,
    n1521,
    n1565,
    n1318,
    n1542
  );


  xnor
  g1910
  (
    n1831,
    n1516,
    n1551,
    n1324,
    n1559
  );


  xor
  g1911
  (
    n1763,
    n1534,
    n1555,
    n1545,
    n1557
  );


  xor
  g1912
  (
    n1614,
    n1532,
    n1536,
    n1522,
    n1564
  );


  or
  g1913
  (
    n1624,
    n1563,
    n1499,
    n1501,
    n1572
  );


  not
  g1914
  (
    n2391,
    n1691
  );


  not
  g1915
  (
    n2598,
    n1891
  );


  buf
  g1916
  (
    n2480,
    n1642
  );


  not
  g1917
  (
    n2639,
    n1742
  );


  not
  g1918
  (
    n1967,
    n1901
  );


  buf
  g1919
  (
    n2055,
    n1914
  );


  buf
  g1920
  (
    n2162,
    n1944
  );


  buf
  g1921
  (
    n2344,
    n1877
  );


  not
  g1922
  (
    n2352,
    n1804
  );


  buf
  g1923
  (
    n2507,
    n1743
  );


  not
  g1924
  (
    KeyWire_0_11,
    n1934
  );


  buf
  g1925
  (
    n2111,
    n1857
  );


  buf
  g1926
  (
    n2695,
    n1927
  );


  buf
  g1927
  (
    n2491,
    n1614
  );


  buf
  g1928
  (
    n2673,
    n1664
  );


  buf
  g1929
  (
    n2611,
    n1812
  );


  not
  g1930
  (
    n2478,
    n1779
  );


  buf
  g1931
  (
    n2363,
    n1648
  );


  not
  g1932
  (
    n1972,
    n1741
  );


  not
  g1933
  (
    n2202,
    n1810
  );


  not
  g1934
  (
    n1987,
    n1620
  );


  not
  g1935
  (
    n2585,
    n1818
  );


  buf
  g1936
  (
    n2136,
    n1618
  );


  not
  g1937
  (
    n2147,
    n1702
  );


  not
  g1938
  (
    n2153,
    n1658
  );


  not
  g1939
  (
    n2039,
    n1799
  );


  buf
  g1940
  (
    n2371,
    n1805
  );


  not
  g1941
  (
    n2261,
    n1861
  );


  not
  g1942
  (
    n2157,
    n1871
  );


  not
  g1943
  (
    n2472,
    n1888
  );


  buf
  g1944
  (
    n2453,
    n1877
  );


  buf
  g1945
  (
    n1957,
    n1690
  );


  not
  g1946
  (
    n2699,
    n1779
  );


  buf
  g1947
  (
    n2353,
    n1881
  );


  not
  g1948
  (
    n2434,
    n1928
  );


  not
  g1949
  (
    n2077,
    n1945
  );


  not
  g1950
  (
    n2316,
    n1622
  );


  not
  g1951
  (
    n2536,
    n1942
  );


  not
  g1952
  (
    KeyWire_0_20,
    n1754
  );


  not
  g1953
  (
    n2454,
    n1593
  );


  buf
  g1954
  (
    n2525,
    n1666
  );


  buf
  g1955
  (
    n2346,
    n1610
  );


  buf
  g1956
  (
    n2249,
    n1618
  );


  buf
  g1957
  (
    n1988,
    n1678
  );


  buf
  g1958
  (
    n2240,
    n1704
  );


  buf
  g1959
  (
    n2646,
    n1644
  );


  not
  g1960
  (
    n2469,
    n1680
  );


  not
  g1961
  (
    n2255,
    n1907
  );


  buf
  g1962
  (
    n2350,
    n1920
  );


  not
  g1963
  (
    n2022,
    n1797
  );


  not
  g1964
  (
    n2375,
    n1825
  );


  buf
  g1965
  (
    n2278,
    n1832
  );


  not
  g1966
  (
    n2592,
    n1910
  );


  not
  g1967
  (
    n2221,
    n1794
  );


  not
  g1968
  (
    n2268,
    n1766
  );


  not
  g1969
  (
    n2501,
    n1892
  );


  not
  g1970
  (
    n2382,
    n1732
  );


  not
  g1971
  (
    n1990,
    n1831
  );


  buf
  g1972
  (
    n2123,
    n1807
  );


  not
  g1973
  (
    n2170,
    n1617
  );


  buf
  g1974
  (
    n1981,
    n1798
  );


  buf
  g1975
  (
    n2277,
    n1634
  );


  buf
  g1976
  (
    n2050,
    n1924
  );


  not
  g1977
  (
    n2176,
    n1785
  );


  not
  g1978
  (
    n2446,
    n1618
  );


  not
  g1979
  (
    n2095,
    n1856
  );


  buf
  g1980
  (
    n2410,
    n1887
  );


  buf
  g1981
  (
    n2683,
    n1681
  );


  not
  g1982
  (
    n2625,
    n1887
  );


  not
  g1983
  (
    n2571,
    n1822
  );


  buf
  g1984
  (
    n2407,
    n1887
  );


  buf
  g1985
  (
    n2292,
    n1788
  );


  buf
  g1986
  (
    n2186,
    n1656
  );


  buf
  g1987
  (
    n2212,
    n1945
  );


  not
  g1988
  (
    n2440,
    n1631
  );


  buf
  g1989
  (
    n2655,
    n1726
  );


  not
  g1990
  (
    n2298,
    n1719
  );


  buf
  g1991
  (
    n2545,
    n1651
  );


  not
  g1992
  (
    n2564,
    n1744
  );


  not
  g1993
  (
    n2286,
    n1774
  );


  not
  g1994
  (
    n2297,
    n1694
  );


  not
  g1995
  (
    n2000,
    n1630
  );


  not
  g1996
  (
    n2066,
    n1703
  );


  not
  g1997
  (
    n2635,
    n1758
  );


  buf
  g1998
  (
    n2072,
    n1775
  );


  not
  g1999
  (
    n2531,
    n1932
  );


  not
  g2000
  (
    n2467,
    n1650
  );


  buf
  g2001
  (
    n2328,
    n1938
  );


  not
  g2002
  (
    n1971,
    n1698
  );


  buf
  g2003
  (
    n2075,
    n1742
  );


  buf
  g2004
  (
    n2216,
    n1852
  );


  buf
  g2005
  (
    n1991,
    n1865
  );


  buf
  g2006
  (
    n2489,
    n1617
  );


  not
  g2007
  (
    n2435,
    n1749
  );


  not
  g2008
  (
    n2465,
    n1911
  );


  buf
  g2009
  (
    n2518,
    n1933
  );


  buf
  g2010
  (
    n2456,
    n1711
  );


  not
  g2011
  (
    n2497,
    n1726
  );


  not
  g2012
  (
    n2019,
    n1823
  );


  not
  g2013
  (
    n2599,
    n1822
  );


  not
  g2014
  (
    n2348,
    n1796
  );


  buf
  g2015
  (
    n2442,
    n1945
  );


  buf
  g2016
  (
    n2423,
    n1636
  );


  not
  g2017
  (
    n2612,
    n1773
  );


  not
  g2018
  (
    n2396,
    n1896
  );


  buf
  g2019
  (
    n2134,
    n1822
  );


  not
  g2020
  (
    n2390,
    n1881
  );


  buf
  g2021
  (
    n2677,
    n1862
  );


  not
  g2022
  (
    n2025,
    n1597
  );


  not
  g2023
  (
    n2506,
    n1716
  );


  buf
  g2024
  (
    n2288,
    n1937
  );


  buf
  g2025
  (
    n2538,
    n1853
  );


  not
  g2026
  (
    n2533,
    n1675
  );


  buf
  g2027
  (
    n2400,
    n1609
  );


  buf
  g2028
  (
    n1986,
    n1790
  );


  not
  g2029
  (
    n2560,
    n1604
  );


  not
  g2030
  (
    n2237,
    n1805
  );


  buf
  g2031
  (
    n2345,
    n1869
  );


  not
  g2032
  (
    n2184,
    n1726
  );


  buf
  g2033
  (
    n2042,
    n1670
  );


  not
  g2034
  (
    n2339,
    n1801
  );


  not
  g2035
  (
    n2565,
    n1720
  );


  buf
  g2036
  (
    n2614,
    n1873
  );


  not
  g2037
  (
    n2559,
    n1917
  );


  buf
  g2038
  (
    n2033,
    n1855
  );


  not
  g2039
  (
    n2293,
    n1671
  );


  not
  g2040
  (
    n2693,
    n1717
  );


  buf
  g2041
  (
    n2492,
    n1604
  );


  buf
  g2042
  (
    n2351,
    n1632
  );


  not
  g2043
  (
    n2680,
    n1729
  );


  buf
  g2044
  (
    n2703,
    n1869
  );


  not
  g2045
  (
    n2265,
    n1928
  );


  not
  g2046
  (
    n2159,
    n1763
  );


  buf
  g2047
  (
    n2178,
    n1939
  );


  not
  g2048
  (
    n2318,
    n1714
  );


  not
  g2049
  (
    n2463,
    n1909
  );


  not
  g2050
  (
    n2018,
    n1597
  );


  buf
  g2051
  (
    n2575,
    n1816
  );


  not
  g2052
  (
    n2154,
    n1844
  );


  not
  g2053
  (
    n2577,
    n1615
  );


  not
  g2054
  (
    KeyWire_0_7,
    n1856
  );


  not
  g2055
  (
    n2160,
    n1905
  );


  not
  g2056
  (
    n2366,
    n1647
  );


  not
  g2057
  (
    n1949,
    n1704
  );


  buf
  g2058
  (
    n2607,
    n1911
  );


  not
  g2059
  (
    n2411,
    n1627
  );


  buf
  g2060
  (
    n2347,
    n1863
  );


  not
  g2061
  (
    n2670,
    n1903
  );


  not
  g2062
  (
    n2040,
    n1682
  );


  not
  g2063
  (
    n2010,
    n1876
  );


  not
  g2064
  (
    n2473,
    n1855
  );


  not
  g2065
  (
    n2096,
    n1661
  );


  buf
  g2066
  (
    n2498,
    n1765
  );


  buf
  g2067
  (
    n2364,
    n1811
  );


  not
  g2068
  (
    n2447,
    n1917
  );


  buf
  g2069
  (
    n2636,
    n1662
  );


  buf
  g2070
  (
    n2228,
    n1712
  );


  not
  g2071
  (
    n2105,
    n1602
  );


  not
  g2072
  (
    n2319,
    n1858
  );


  not
  g2073
  (
    n2030,
    n1842
  );


  not
  g2074
  (
    n2597,
    n1636
  );


  buf
  g2075
  (
    n2459,
    n1866
  );


  not
  g2076
  (
    n2628,
    n1761
  );


  not
  g2077
  (
    n1978,
    n1798
  );


  buf
  g2078
  (
    n2151,
    n1644
  );


  buf
  g2079
  (
    n2661,
    n1672
  );


  buf
  g2080
  (
    n1974,
    n1929
  );


  buf
  g2081
  (
    n2388,
    n1720
  );


  not
  g2082
  (
    n2398,
    n1700
  );


  not
  g2083
  (
    n2688,
    n1705
  );


  not
  g2084
  (
    n2649,
    n1403
  );


  not
  g2085
  (
    n2341,
    n1941
  );


  buf
  g2086
  (
    n2289,
    n1677
  );


  buf
  g2087
  (
    n2108,
    n1876
  );


  buf
  g2088
  (
    n2397,
    n1699
  );


  buf
  g2089
  (
    n2691,
    n1914
  );


  buf
  g2090
  (
    n2615,
    n1833
  );


  buf
  g2091
  (
    n2358,
    n1931
  );


  not
  g2092
  (
    n2320,
    n1865
  );


  not
  g2093
  (
    n2594,
    n1701
  );


  buf
  g2094
  (
    n2386,
    n1860
  );


  buf
  g2095
  (
    n1973,
    n1803
  );


  not
  g2096
  (
    n2572,
    n1728
  );


  buf
  g2097
  (
    n2372,
    n1628
  );


  not
  g2098
  (
    n1951,
    n1707
  );


  buf
  g2099
  (
    n2222,
    n1839
  );


  not
  g2100
  (
    n2083,
    n1778
  );


  buf
  g2101
  (
    n2168,
    n1826
  );


  not
  g2102
  (
    n2331,
    n1608
  );


  buf
  g2103
  (
    n2458,
    n1643
  );


  not
  g2104
  (
    n2449,
    n1880
  );


  buf
  g2105
  (
    n2455,
    n1664
  );


  not
  g2106
  (
    n2385,
    n1908
  );


  not
  g2107
  (
    n2191,
    n1609
  );


  not
  g2108
  (
    n2129,
    n1680
  );


  buf
  g2109
  (
    n2643,
    n1772
  );


  buf
  g2110
  (
    n2137,
    n1605
  );


  buf
  g2111
  (
    n2550,
    n1884
  );


  buf
  g2112
  (
    n2461,
    n1940
  );


  buf
  g2113
  (
    n2503,
    n1716
  );


  buf
  g2114
  (
    n1966,
    n1894
  );


  buf
  g2115
  (
    n2312,
    n1888
  );


  buf
  g2116
  (
    n2068,
    n1942
  );


  buf
  g2117
  (
    n2384,
    n1634
  );


  buf
  g2118
  (
    n2368,
    n1668
  );


  buf
  g2119
  (
    n2576,
    n1406
  );


  not
  g2120
  (
    n2563,
    n1835
  );


  not
  g2121
  (
    n2175,
    n1670
  );


  not
  g2122
  (
    n2477,
    n1913
  );


  buf
  g2123
  (
    n2054,
    n1829
  );


  not
  g2124
  (
    n2245,
    n1782
  );


  buf
  g2125
  (
    n2660,
    n1647
  );


  buf
  g2126
  (
    n2008,
    n1913
  );


  buf
  g2127
  (
    n2696,
    n1900
  );


  buf
  g2128
  (
    n2031,
    n1932
  );


  not
  g2129
  (
    n2052,
    n1867
  );


  buf
  g2130
  (
    KeyWire_0_17,
    n1680
  );


  not
  g2131
  (
    n2235,
    n1654
  );


  not
  g2132
  (
    n2187,
    n1784
  );


  buf
  g2133
  (
    n2193,
    n1755
  );


  not
  g2134
  (
    n2425,
    n1866
  );


  not
  g2135
  (
    n2413,
    n1758
  );


  buf
  g2136
  (
    n2326,
    n1602
  );


  not
  g2137
  (
    n2591,
    n1824
  );


  buf
  g2138
  (
    n2295,
    n1593
  );


  not
  g2139
  (
    n2279,
    n1405
  );


  buf
  g2140
  (
    n2437,
    n1858
  );


  not
  g2141
  (
    n2149,
    n1748
  );


  buf
  g2142
  (
    n2679,
    n1753
  );


  buf
  g2143
  (
    n2317,
    n1921
  );


  buf
  g2144
  (
    n2056,
    n1601
  );


  not
  g2145
  (
    n2618,
    n1602
  );


  buf
  g2146
  (
    n2511,
    n1750
  );


  not
  g2147
  (
    n2632,
    n1889
  );


  buf
  g2148
  (
    n2596,
    n1645
  );


  not
  g2149
  (
    n1999,
    n1946
  );


  buf
  g2150
  (
    n2698,
    n1812
  );


  not
  g2151
  (
    n2409,
    n1740
  );


  buf
  g2152
  (
    n2013,
    n1681
  );


  buf
  g2153
  (
    n2051,
    n1767
  );


  not
  g2154
  (
    n2307,
    n1846
  );


  buf
  g2155
  (
    n2354,
    n1883
  );


  buf
  g2156
  (
    n2158,
    n1631
  );


  buf
  g2157
  (
    n1968,
    n1663
  );


  buf
  g2158
  (
    n2462,
    n1941
  );


  not
  g2159
  (
    n2028,
    n1698
  );


  buf
  g2160
  (
    n2579,
    n1691
  );


  not
  g2161
  (
    n2260,
    n1853
  );


  buf
  g2162
  (
    n1996,
    n1735
  );


  buf
  g2163
  (
    n2543,
    n1851
  );


  not
  g2164
  (
    n2441,
    n1788
  );


  buf
  g2165
  (
    n2327,
    n1827
  );


  buf
  g2166
  (
    n2061,
    n1608
  );


  not
  g2167
  (
    n2091,
    n1755
  );


  buf
  g2168
  (
    n2547,
    n1621
  );


  not
  g2169
  (
    n2131,
    n1648
  );


  buf
  g2170
  (
    n2404,
    n1799
  );


  buf
  g2171
  (
    n2304,
    n1628
  );


  not
  g2172
  (
    n2405,
    n1792
  );


  not
  g2173
  (
    n2026,
    n1797
  );


  buf
  g2174
  (
    n1955,
    n1793
  );


  buf
  g2175
  (
    n2244,
    n1407
  );


  buf
  g2176
  (
    n2238,
    n1789
  );


  buf
  g2177
  (
    n2148,
    n1872
  );


  buf
  g2178
  (
    n2471,
    n1831
  );


  buf
  g2179
  (
    n2487,
    n1619
  );


  buf
  g2180
  (
    n2381,
    n1728
  );


  not
  g2181
  (
    n2183,
    n1406
  );


  not
  g2182
  (
    n2512,
    n1872
  );


  buf
  g2183
  (
    n2383,
    n1714
  );


  buf
  g2184
  (
    n2552,
    n1830
  );


  buf
  g2185
  (
    n2120,
    n1893
  );


  not
  g2186
  (
    n2637,
    n1762
  );


  not
  g2187
  (
    n2036,
    n1652
  );


  not
  g2188
  (
    n2225,
    n1900
  );


  buf
  g2189
  (
    n2089,
    n1706
  );


  not
  g2190
  (
    n2035,
    n1841
  );


  not
  g2191
  (
    n2692,
    n1907
  );


  buf
  g2192
  (
    n2024,
    n1643
  );


  not
  g2193
  (
    n2359,
    n1904
  );


  not
  g2194
  (
    n2638,
    n1819
  );


  not
  g2195
  (
    n2067,
    n1708
  );


  not
  g2196
  (
    n2064,
    n1757
  );


  not
  g2197
  (
    n2126,
    n1666
  );


  not
  g2198
  (
    n2570,
    n1808
  );


  not
  g2199
  (
    n2248,
    n1781
  );


  not
  g2200
  (
    n2627,
    n1717
  );


  buf
  g2201
  (
    n2082,
    n1731
  );


  buf
  g2202
  (
    n2601,
    n1684
  );


  buf
  g2203
  (
    n2156,
    n1595
  );


  not
  g2204
  (
    n1982,
    n1636
  );


  not
  g2205
  (
    n2644,
    n1676
  );


  not
  g2206
  (
    n2626,
    n1405
  );


  not
  g2207
  (
    n2623,
    n1821
  );


  buf
  g2208
  (
    n2011,
    n1745
  );


  buf
  g2209
  (
    n2513,
    n1815
  );


  not
  g2210
  (
    n2115,
    n1891
  );


  buf
  g2211
  (
    n2110,
    n1913
  );


  not
  g2212
  (
    n2648,
    n1603
  );


  not
  g2213
  (
    n2610,
    n1629
  );


  buf
  g2214
  (
    n2208,
    n1644
  );


  buf
  g2215
  (
    n2609,
    n1784
  );


  not
  g2216
  (
    n2284,
    n1787
  );


  buf
  g2217
  (
    n2500,
    n1776
  );


  buf
  g2218
  (
    n2392,
    n1796
  );


  buf
  g2219
  (
    n2488,
    n1875
  );


  not
  g2220
  (
    n2132,
    n1744
  );


  not
  g2221
  (
    n2047,
    n1872
  );


  not
  g2222
  (
    n2076,
    n1874
  );


  not
  g2223
  (
    n1964,
    n1791
  );


  buf
  g2224
  (
    n2164,
    n1727
  );


  buf
  g2225
  (
    n2349,
    n1630
  );


  not
  g2226
  (
    n2100,
    n1615
  );


  buf
  g2227
  (
    n2438,
    n1711
  );


  buf
  g2228
  (
    n2605,
    n1870
  );


  buf
  g2229
  (
    n2101,
    n1769
  );


  buf
  g2230
  (
    n2595,
    n1694
  );


  not
  g2231
  (
    n2686,
    n1617
  );


  buf
  g2232
  (
    n2195,
    n1406
  );


  not
  g2233
  (
    n2029,
    n1899
  );


  buf
  g2234
  (
    n2204,
    n1768
  );


  buf
  g2235
  (
    n2657,
    n1778
  );


  buf
  g2236
  (
    n2306,
    n1647
  );


  buf
  g2237
  (
    n2098,
    n1931
  );


  buf
  g2238
  (
    n2562,
    n1608
  );


  buf
  g2239
  (
    n2430,
    n1885
  );


  not
  g2240
  (
    n2189,
    n1693
  );


  not
  g2241
  (
    n2548,
    n1898
  );


  not
  g2242
  (
    n2106,
    n1857
  );


  not
  g2243
  (
    n2218,
    n1833
  );


  not
  g2244
  (
    n2509,
    n1868
  );


  not
  g2245
  (
    n2494,
    n1724
  );


  buf
  g2246
  (
    n2034,
    n1673
  );


  not
  g2247
  (
    n2012,
    n1840
  );


  buf
  g2248
  (
    n2074,
    n1618
  );


  not
  g2249
  (
    n2439,
    n1723
  );


  buf
  g2250
  (
    n2038,
    n1656
  );


  buf
  g2251
  (
    n2419,
    n1795
  );


  not
  g2252
  (
    n2043,
    n1683
  );


  not
  g2253
  (
    n2063,
    n1614
  );


  buf
  g2254
  (
    n2551,
    n1722
  );


  buf
  g2255
  (
    n2104,
    n1895
  );


  buf
  g2256
  (
    n2379,
    n1849
  );


  not
  g2257
  (
    n2311,
    n1657
  );


  not
  g2258
  (
    n2528,
    n1881
  );


  not
  g2259
  (
    n2694,
    n1847
  );


  buf
  g2260
  (
    n2418,
    n1686
  );


  not
  g2261
  (
    n2165,
    n1854
  );


  not
  g2262
  (
    n2269,
    n1729
  );


  buf
  g2263
  (
    n2124,
    n1883
  );


  buf
  g2264
  (
    n2333,
    n1918
  );


  not
  g2265
  (
    n2046,
    n1601
  );


  buf
  g2266
  (
    n1950,
    n1697
  );


  buf
  g2267
  (
    n2233,
    n1803
  );


  buf
  g2268
  (
    n2088,
    n1715
  );


  not
  g2269
  (
    n2116,
    n1651
  );


  not
  g2270
  (
    n2642,
    n1756
  );


  not
  g2271
  (
    n2044,
    n1747
  );


  not
  g2272
  (
    n1952,
    n1840
  );


  buf
  g2273
  (
    n2527,
    n1916
  );


  buf
  g2274
  (
    n2324,
    n1870
  );


  not
  g2275
  (
    n2338,
    n1615
  );


  not
  g2276
  (
    n2262,
    n1705
  );


  not
  g2277
  (
    n2583,
    n1665
  );


  buf
  g2278
  (
    n2514,
    n1684
  );


  not
  g2279
  (
    n2622,
    n1725
  );


  not
  g2280
  (
    n2181,
    n1884
  );


  not
  g2281
  (
    n2180,
    n1700
  );


  buf
  g2282
  (
    n2361,
    n1932
  );


  buf
  g2283
  (
    n2373,
    n1902
  );


  buf
  g2284
  (
    n2581,
    n1936
  );


  not
  g2285
  (
    n2522,
    n1825
  );


  buf
  g2286
  (
    n1995,
    n1771
  );


  not
  g2287
  (
    n2215,
    n1612
  );


  buf
  g2288
  (
    n2336,
    n1691
  );


  buf
  g2289
  (
    n2516,
    n1722
  );


  not
  g2290
  (
    n2697,
    n1783
  );


  not
  g2291
  (
    n2122,
    n1626
  );


  not
  g2292
  (
    n2675,
    n1739
  );


  not
  g2293
  (
    n1977,
    n1843
  );


  not
  g2294
  (
    n2272,
    n1657
  );


  not
  g2295
  (
    n2210,
    n1929
  );


  not
  g2296
  (
    n2460,
    n1629
  );


  not
  g2297
  (
    n2199,
    n1407
  );


  buf
  g2298
  (
    n2300,
    n1667
  );


  not
  g2299
  (
    n2532,
    n1744
  );


  buf
  g2300
  (
    n2079,
    n1675
  );


  buf
  g2301
  (
    n2001,
    n1934
  );


  buf
  g2302
  (
    n2285,
    n1757
  );


  not
  g2303
  (
    n2097,
    n1838
  );


  buf
  g2304
  (
    n2421,
    n1741
  );


  not
  g2305
  (
    n2429,
    n1638
  );


  not
  g2306
  (
    n2145,
    n1622
  );


  buf
  g2307
  (
    n2004,
    n1787
  );


  buf
  g2308
  (
    n2408,
    n1687
  );


  buf
  g2309
  (
    n1962,
    n1691
  );


  not
  g2310
  (
    n2201,
    n1834
  );


  buf
  g2311
  (
    n2378,
    n1905
  );


  not
  g2312
  (
    n2194,
    n1633
  );


  buf
  g2313
  (
    n2309,
    n1706
  );


  buf
  g2314
  (
    n2206,
    n1660
  );


  not
  g2315
  (
    n2656,
    n1837
  );


  not
  g2316
  (
    n2523,
    n1693
  );


  not
  g2317
  (
    n2588,
    n1407
  );


  not
  g2318
  (
    n2335,
    n1728
  );


  not
  g2319
  (
    n2236,
    n1938
  );


  buf
  g2320
  (
    n2602,
    n1695
  );


  buf
  g2321
  (
    n2534,
    n1926
  );


  buf
  g2322
  (
    n2377,
    n1651
  );


  not
  g2323
  (
    n2166,
    n1931
  );


  buf
  g2324
  (
    KeyWire_0_18,
    n1746
  );


  buf
  g2325
  (
    n2182,
    n1630
  );


  not
  g2326
  (
    n2048,
    n1827
  );


  buf
  g2327
  (
    KeyWire_0_27,
    n1899
  );


  buf
  g2328
  (
    n2422,
    n1751
  );


  not
  g2329
  (
    n1975,
    n1629
  );


  not
  g2330
  (
    n2299,
    n1688
  );


  not
  g2331
  (
    n2630,
    n1738
  );


  not
  g2332
  (
    n2252,
    n1624
  );


  not
  g2333
  (
    n2702,
    n1855
  );


  not
  g2334
  (
    n2253,
    n1860
  );


  buf
  g2335
  (
    n2606,
    n1665
  );


  buf
  g2336
  (
    n2426,
    n1881
  );


  buf
  g2337
  (
    n2229,
    n1785
  );


  buf
  g2338
  (
    n2073,
    n1673
  );


  not
  g2339
  (
    n2021,
    n1707
  );


  not
  g2340
  (
    n2578,
    n1650
  );


  buf
  g2341
  (
    n2332,
    n1821
  );


  buf
  g2342
  (
    n2394,
    n1747
  );


  buf
  g2343
  (
    n2483,
    n1797
  );


  not
  g2344
  (
    n2417,
    n1852
  );


  not
  g2345
  (
    n2259,
    n1681
  );


  buf
  g2346
  (
    n2109,
    n1610
  );


  not
  g2347
  (
    n2389,
    n1769
  );


  buf
  g2348
  (
    n2659,
    n1700
  );


  buf
  g2349
  (
    n2190,
    n1819
  );


  buf
  g2350
  (
    n2466,
    n1915
  );


  buf
  g2351
  (
    n2330,
    n1637
  );


  buf
  g2352
  (
    n2177,
    n1745
  );


  buf
  g2353
  (
    n2334,
    n1780
  );


  buf
  g2354
  (
    n2620,
    n1814
  );


  buf
  g2355
  (
    n2230,
    n1830
  );


  not
  g2356
  (
    n2555,
    n1640
  );


  buf
  g2357
  (
    n2682,
    n1600
  );


  buf
  g2358
  (
    n2321,
    n1659
  );


  not
  g2359
  (
    n1959,
    n1624
  );


  buf
  g2360
  (
    n2086,
    n1725
  );


  not
  g2361
  (
    n2380,
    n1860
  );


  buf
  g2362
  (
    n2016,
    n1334
  );


  not
  g2363
  (
    n2294,
    n1687
  );


  buf
  g2364
  (
    n2537,
    n1734
  );


  not
  g2365
  (
    n2475,
    n1766
  );


  not
  g2366
  (
    n2443,
    n1745
  );


  not
  g2367
  (
    n2486,
    n1627
  );


  not
  g2368
  (
    n2667,
    n1632
  );


  buf
  g2369
  (
    n2322,
    n1661
  );


  buf
  g2370
  (
    n2290,
    n1809
  );


  buf
  g2371
  (
    n2172,
    n1836
  );


  not
  g2372
  (
    n2340,
    n1752
  );


  not
  g2373
  (
    n2549,
    n1800
  );


  not
  g2374
  (
    n2653,
    n1800
  );


  not
  g2375
  (
    n2343,
    n1756
  );


  buf
  g2376
  (
    n2634,
    n1645
  );


  buf
  g2377
  (
    n2070,
    n1835
  );


  not
  g2378
  (
    n2573,
    n1938
  );


  buf
  g2379
  (
    n2274,
    n1901
  );


  buf
  g2380
  (
    n2701,
    n1816
  );


  not
  g2381
  (
    n2112,
    n1781
  );


  buf
  g2382
  (
    n2664,
    n1753
  );


  buf
  g2383
  (
    n2062,
    n1942
  );


  not
  g2384
  (
    n2167,
    n1708
  );


  buf
  g2385
  (
    n2556,
    n1845
  );


  not
  g2386
  (
    n2690,
    n1888
  );


  not
  g2387
  (
    n1956,
    n1873
  );


  not
  g2388
  (
    n2059,
    n1603
  );


  not
  g2389
  (
    n2546,
    n1679
  );


  buf
  g2390
  (
    n2017,
    n1811
  );


  not
  g2391
  (
    n2574,
    n1871
  );


  buf
  g2392
  (
    n2651,
    n1836
  );


  buf
  g2393
  (
    n2329,
    n1809
  );


  not
  g2394
  (
    n2291,
    n1935
  );


  buf
  g2395
  (
    n2569,
    n1800
  );


  buf
  g2396
  (
    n2428,
    n1595
  );


  not
  g2397
  (
    n2650,
    n1867
  );


  not
  g2398
  (
    n2142,
    n1645
  );


  buf
  g2399
  (
    n2496,
    n1613
  );


  not
  g2400
  (
    n1985,
    n1608
  );


  buf
  g2401
  (
    n1984,
    n1786
  );


  buf
  g2402
  (
    n2247,
    n1747
  );


  not
  g2403
  (
    n2401,
    n1777
  );


  buf
  g2404
  (
    n2213,
    n1863
  );


  buf
  g2405
  (
    n2687,
    n1752
  );


  not
  g2406
  (
    n2540,
    n1596
  );


  buf
  g2407
  (
    n2479,
    n1803
  );


  not
  g2408
  (
    n2313,
    n1730
  );


  not
  g2409
  (
    n2270,
    n1772
  );


  buf
  g2410
  (
    n2608,
    n1920
  );


  not
  g2411
  (
    n2517,
    n1842
  );


  not
  g2412
  (
    n2093,
    n1911
  );


  not
  g2413
  (
    n2530,
    n1765
  );


  buf
  g2414
  (
    n2355,
    n1669
  );


  not
  g2415
  (
    n2393,
    n1879
  );


  not
  g2416
  (
    n1980,
    n1657
  );


  buf
  g2417
  (
    n2027,
    n1774
  );


  not
  g2418
  (
    KeyWire_0_12,
    n1738
  );


  buf
  g2419
  (
    n2143,
    n1926
  );


  buf
  g2420
  (
    n2520,
    n1813
  );


  not
  g2421
  (
    n2631,
    n1856
  );


  buf
  g2422
  (
    n1993,
    n1653
  );


  buf
  g2423
  (
    n2662,
    n1914
  );


  buf
  g2424
  (
    n2266,
    n1884
  );


  not
  g2425
  (
    n2283,
    n1944
  );


  buf
  g2426
  (
    n2005,
    n1894
  );


  not
  g2427
  (
    n2529,
    n1649
  );


  buf
  g2428
  (
    n2071,
    n1654
  );


  buf
  g2429
  (
    n2406,
    n1612
  );


  buf
  g2430
  (
    n2604,
    n1690
  );


  buf
  g2431
  (
    n2205,
    n1783
  );


  buf
  g2432
  (
    n2203,
    n1775
  );


  not
  g2433
  (
    n2258,
    n1789
  );


  buf
  g2434
  (
    n2217,
    n1816
  );


  not
  g2435
  (
    n2658,
    n1658
  );


  buf
  g2436
  (
    n2669,
    n1920
  );


  not
  g2437
  (
    n2402,
    n1806
  );


  buf
  g2438
  (
    n2231,
    n1915
  );


  not
  g2439
  (
    n2414,
    n1731
  );


  not
  g2440
  (
    n2242,
    n1836
  );


  not
  g2441
  (
    n2541,
    n1797
  );


  not
  g2442
  (
    n2476,
    n1716
  );


  not
  g2443
  (
    n2271,
    n1717
  );


  nand
  g2444
  (
    n2174,
    n1601,
    n1759,
    n1623,
    n1749
  );


  or
  g2445
  (
    n2342,
    n1832,
    n1743,
    n1846,
    n1701
  );


  and
  g2446
  (
    n2495,
    n1786,
    n1865,
    n1667,
    n1895
  );


  xor
  g2447
  (
    n2633,
    n1939,
    n1837,
    n1808,
    n1621
  );


  xnor
  g2448
  (
    n2600,
    n1682,
    n1771,
    n1652,
    n1834
  );


  or
  g2449
  (
    n2399,
    n1333,
    n1653,
    n1687,
    n1858
  );


  xor
  g2450
  (
    n2510,
    n1611,
    n1776,
    n1742,
    n1730
  );


  nor
  g2451
  (
    n2301,
    n1662,
    n1624,
    n1666,
    n1838
  );


  xnor
  g2452
  (
    n2468,
    n1658,
    n1946,
    n1595,
    n1598
  );


  and
  g2453
  (
    n2499,
    n1864,
    n1829,
    n1685,
    n1596
  );


  xnor
  g2454
  (
    n2094,
    n1933,
    n1903,
    n1853,
    n1944
  );


  xnor
  g2455
  (
    n2121,
    n1652,
    n1776,
    n1602,
    n1625
  );


  xor
  g2456
  (
    n1961,
    n1814,
    n1695,
    n1699,
    n1859
  );


  xnor
  g2457
  (
    n2521,
    n1634,
    n1665,
    n1689,
    n1727
  );


  and
  g2458
  (
    n2356,
    n1850,
    n1900,
    n1741,
    n1765
  );


  xnor
  g2459
  (
    n1983,
    n1594,
    n1705,
    n1721,
    n1713
  );


  nor
  g2460
  (
    n2362,
    n1632,
    n1850,
    n1733,
    n1659
  );


  xor
  g2461
  (
    n2015,
    n1646,
    n1920,
    n1725,
    n1604
  );


  nor
  g2462
  (
    n2376,
    n1649,
    n1834,
    n1758,
    n1875
  );


  or
  g2463
  (
    n2424,
    n1760,
    n1647,
    n1875,
    n1791
  );


  and
  g2464
  (
    n2003,
    n1697,
    n1764,
    n1703,
    n1713
  );


  xor
  g2465
  (
    n2539,
    n1679,
    n1807,
    n1737,
    n1935
  );


  and
  g2466
  (
    n2085,
    n1763,
    n1828,
    n1823,
    n1734
  );


  nand
  g2467
  (
    n1976,
    n1923,
    n1666,
    n1616,
    n1715
  );


  and
  g2468
  (
    n2685,
    n1774,
    n1813,
    n1595,
    n1846
  );


  xnor
  g2469
  (
    n2369,
    n1711,
    n1650,
    n1686,
    n1641
  );


  or
  g2470
  (
    n2049,
    n1646,
    n1736,
    n1756,
    n1761
  );


  nor
  g2471
  (
    n2007,
    n1873,
    n1606,
    n1946,
    n1908
  );


  and
  g2472
  (
    n2117,
    n1767,
    n1724,
    n1739,
    n1708
  );


  xnor
  g2473
  (
    n2171,
    n1670,
    n1607,
    n1904,
    n1919
  );


  nor
  g2474
  (
    n2192,
    n1627,
    n1863,
    n1818,
    n1903
  );


  nor
  g2475
  (
    n2188,
    n1799,
    n1886,
    n1732,
    n1807
  );


  xnor
  g2476
  (
    n2065,
    n1835,
    n1868,
    n1762,
    n1736
  );


  and
  g2477
  (
    n2415,
    n1879,
    n1668,
    n1787,
    n1814
  );


  nor
  g2478
  (
    n2624,
    n1830,
    n1610,
    n1778,
    n1786
  );


  xnor
  g2479
  (
    n2568,
    n1847,
    n1607,
    n1639,
    n1629
  );


  or
  g2480
  (
    n2087,
    n1943,
    n1916,
    n1861,
    n1606
  );


  nand
  g2481
  (
    n2672,
    n1635,
    n1677,
    n1671,
    n1752
  );


  nor
  g2482
  (
    n2387,
    n1719,
    n1688,
    n1733,
    n1804
  );


  nor
  g2483
  (
    n2141,
    n1861,
    n1642,
    n1905,
    n1740
  );


  xnor
  g2484
  (
    n2209,
    n1721,
    n1876,
    n1886,
    n1894
  );


  nor
  g2485
  (
    n2224,
    n1895,
    n1759,
    n1775,
    n1838
  );


  nor
  g2486
  (
    n2515,
    n1619,
    n1844,
    n1936,
    n1823
  );


  xor
  g2487
  (
    n1965,
    n1840,
    n1827,
    n1613,
    n1915
  );


  xor
  g2488
  (
    n2603,
    n1803,
    n1684,
    n1621,
    n1914
  );


  xor
  g2489
  (
    n2053,
    n1936,
    n1646,
    n1930,
    n1599
  );


  and
  g2490
  (
    n2640,
    n1896,
    n1701,
    n1697,
    n1403
  );


  xnor
  g2491
  (
    n2619,
    n1825,
    n1922,
    n1639,
    n1759
  );


  xnor
  g2492
  (
    n2621,
    n1600,
    n1909,
    n1762,
    n1770
  );


  or
  g2493
  (
    n2102,
    n1609,
    n1638,
    n1750,
    n1727
  );


  xnor
  g2494
  (
    n1998,
    n1763,
    n1637,
    n1619,
    n1773
  );


  xor
  g2495
  (
    n2526,
    n1874,
    n1858,
    n1685,
    n1834
  );


  xor
  g2496
  (
    n2303,
    n1878,
    n1764,
    n1611,
    n1893
  );


  xnor
  g2497
  (
    n2395,
    n1805,
    n1856,
    n1944,
    n1788
  );


  xor
  g2498
  (
    n2586,
    n1731,
    n1466,
    n1845,
    n1671
  );


  nand
  g2499
  (
    n2535,
    n1946,
    n1777,
    n1669,
    n1737
  );


  nor
  g2500
  (
    n2474,
    n1633,
    n1717,
    n1908,
    n1777
  );


  xnor
  g2501
  (
    n2524,
    n1876,
    n1901,
    n1884,
    n1939
  );


  or
  g2502
  (
    n2561,
    n1912,
    n1801,
    n1904,
    n1883
  );


  and
  g2503
  (
    n2226,
    n1846,
    n1864,
    n1648,
    n1637
  );


  xnor
  g2504
  (
    n2613,
    n1848,
    n1714,
    n1706,
    n1927
  );


  or
  g2505
  (
    n2444,
    n1713,
    n1869,
    n1917,
    n1771
  );


  xnor
  g2506
  (
    n2367,
    n1643,
    n1927,
    n1600,
    n1639
  );


  nor
  g2507
  (
    n2590,
    n1868,
    n1866,
    n1643,
    n1929
  );


  xor
  g2508
  (
    n1960,
    n1883,
    n1787,
    n1593,
    n1734
  );


  xor
  g2509
  (
    n2427,
    n1712,
    n1605,
    n1847,
    n1663
  );


  xor
  g2510
  (
    n1958,
    n1721,
    n1620,
    n1631,
    n1845
  );


  xor
  g2511
  (
    n2276,
    n1906,
    n1781,
    n1625,
    n1718
  );


  xor
  g2512
  (
    n2629,
    n1748,
    n1890,
    n1736,
    n1675
  );


  xor
  g2513
  (
    n2684,
    n1700,
    n1922,
    n1754,
    n1673
  );


  xor
  g2514
  (
    n2567,
    n1822,
    n1623,
    n1687,
    n1886
  );


  and
  g2515
  (
    n2557,
    n1851,
    n1828,
    n1623,
    n1751
  );


  xnor
  g2516
  (
    n2584,
    n1673,
    n1871,
    n1789,
    n1804
  );


  nand
  g2517
  (
    n2457,
    n1820,
    n1889,
    n1857,
    n1940
  );


  nor
  g2518
  (
    n2150,
    n1612,
    n1710,
    n1916,
    n1942
  );


  nor
  g2519
  (
    n2370,
    n1740,
    n1795,
    n1828,
    n1930
  );


  nor
  g2520
  (
    n2254,
    n1806,
    n1840,
    n1709,
    n1719
  );


  nor
  g2521
  (
    n2357,
    n1640,
    n1686,
    n1681,
    n1854
  );


  xor
  g2522
  (
    n2374,
    n1654,
    n1739,
    n1857,
    n1664
  );


  xor
  g2523
  (
    n2310,
    n1805,
    n1807,
    n1695,
    n1658
  );


  xnor
  g2524
  (
    n1997,
    n1918,
    n1880,
    n1849,
    n1622
  );


  or
  g2525
  (
    n1947,
    n1601,
    n1661,
    n1897,
    n1918
  );


  or
  g2526
  (
    n2582,
    n1843,
    n1910,
    n1748,
    n1791
  );


  or
  g2527
  (
    n2239,
    n1810,
    n1793,
    n1851,
    n1772
  );


  and
  g2528
  (
    n2647,
    n1835,
    n1737,
    n1879,
    n1943
  );


  and
  g2529
  (
    n2544,
    n1785,
    n1751,
    n1620,
    n1896
  );


  xor
  g2530
  (
    n2365,
    n1862,
    n1839,
    n1749,
    n1616
  );


  xor
  g2531
  (
    n2092,
    n1746,
    n1937,
    n1878,
    n1877
  );


  and
  g2532
  (
    n2246,
    n1599,
    n1655,
    n1812,
    n1638
  );


  xnor
  g2533
  (
    n2198,
    n1769,
    n1781,
    n1702,
    n1743
  );


  or
  g2534
  (
    n2616,
    n1651,
    n1744,
    n1636,
    n1925
  );


  and
  g2535
  (
    n2433,
    n1925,
    n1848,
    n1926,
    n1626
  );


  xnor
  g2536
  (
    n2234,
    n1699,
    n1778,
    n1750,
    n1678
  );


  xor
  g2537
  (
    n2256,
    n1925,
    n1831,
    n1905,
    n1906
  );


  xnor
  g2538
  (
    n2482,
    n1599,
    n1701,
    n1826,
    n1827
  );


  and
  g2539
  (
    n2250,
    n1735,
    n1915,
    n1938,
    n1653
  );


  nand
  g2540
  (
    n2185,
    n1801,
    n1891,
    n1773,
    n1719
  );


  xnor
  g2541
  (
    n2470,
    n1849,
    n1922,
    n1897,
    n1847
  );


  or
  g2542
  (
    n2263,
    n1669,
    n1902,
    n1757,
    n1720
  );


  and
  g2543
  (
    n2589,
    n1890,
    n1764,
    n1613,
    n1696
  );


  nor
  g2544
  (
    n2700,
    n1820,
    n1646,
    n1908,
    n1882
  );


  xor
  g2545
  (
    n1963,
    n1712,
    n1780,
    n1850,
    n1937
  );


  and
  g2546
  (
    n2032,
    n1853,
    n1879,
    n1907,
    n1746
  );


  xor
  g2547
  (
    n2169,
    n1696,
    n1746,
    n1405,
    n1722
  );


  xnor
  g2548
  (
    n2125,
    n1707,
    n1819,
    n1685,
    n1702
  );


  xor
  g2549
  (
    n2323,
    n1817,
    n1690,
    n1596,
    n1407
  );


  or
  g2550
  (
    n2281,
    n1674,
    n1672,
    n1760,
    n1864
  );


  or
  g2551
  (
    n2666,
    n1771,
    n1728,
    n1692
  );


  nand
  g2552
  (
    n2305,
    n1718,
    n1641,
    n1404,
    n1659
  );


  or
  g2553
  (
    n2119,
    n1839,
    n1885,
    n1828,
    n1874
  );


  or
  g2554
  (
    n2689,
    n1767,
    n1760,
    n1684,
    n1813
  );


  or
  g2555
  (
    n2060,
    n1930,
    n1817,
    n1628,
    n1782
  );


  or
  g2556
  (
    n2668,
    n1812,
    n1929,
    n1894,
    n1722
  );


  or
  g2557
  (
    n2452,
    n1888,
    n1926,
    n1860,
    n1817
  );


  nand
  g2558
  (
    n2090,
    n1635,
    n1806,
    n1649,
    n1594
  );


  xnor
  g2559
  (
    n2251,
    n1849,
    n1655,
    n1832,
    n1598
  );


  nor
  g2560
  (
    n2275,
    n1909,
    n1760,
    n1842,
    n1864
  );


  or
  g2561
  (
    n2508,
    n1603,
    n1830,
    n1769,
    n1599
  );


  and
  g2562
  (
    n2128,
    n1910,
    n1594,
    n1707,
    n1705
  );


  or
  g2563
  (
    n2654,
    n1794,
    n1405,
    n1842,
    n1820
  );


  nand
  g2564
  (
    n2058,
    n1733,
    n1749,
    n1758,
    n1780
  );


  nand
  g2565
  (
    n2325,
    n1917,
    n1815,
    n1652,
    n1841
  );


  and
  g2566
  (
    n2566,
    n1837,
    n1663,
    n1713,
    n1924
  );


  xnor
  g2567
  (
    n2308,
    n1683,
    n1610,
    n1777,
    n1850
  );


  nand
  g2568
  (
    n2665,
    n1635,
    n1694,
    n1802,
    n1940
  );


  xnor
  g2569
  (
    n2179,
    n1877,
    n1818,
    n1754,
    n1824
  );


  nand
  g2570
  (
    n2554,
    n1770,
    n1660,
    n1924,
    n1671
  );


  xnor
  g2571
  (
    n2587,
    n1919,
    n1625,
    n1885,
    n1723
  );


  or
  g2572
  (
    n2416,
    n1913,
    n1804,
    n1936,
    n1679
  );


  xnor
  g2573
  (
    n2553,
    n1907,
    n1823,
    n1820,
    n1683
  );


  nand
  g2574
  (
    n2580,
    n1893,
    n1843,
    n1939,
    n1941
  );


  xor
  g2575
  (
    n2267,
    n1921,
    n1662,
    n1604,
    n1627
  );


  and
  g2576
  (
    n2214,
    n1641,
    n1882,
    n1817,
    n1716
  );


  or
  g2577
  (
    n1979,
    n1770,
    n1762,
    n1941,
    n1715
  );


  and
  g2578
  (
    n2403,
    n1770,
    n1833,
    n1650,
    n1895
  );


  nand
  g2579
  (
    n2243,
    n1644,
    n1912,
    n1754,
    n1753
  );


  xnor
  g2580
  (
    n2451,
    n1791,
    n1738,
    n1866,
    n1937
  );


  and
  g2581
  (
    n2264,
    n1775,
    n1755,
    n1678,
    n1854
  );


  nand
  g2582
  (
    n1969,
    n1680,
    n1788,
    n1845,
    n1922
  );


  and
  g2583
  (
    n2287,
    n1739,
    n1616,
    n1831,
    n1898
  );


  xor
  g2584
  (
    n1948,
    n1815,
    n1726,
    n1718,
    n1794
  );


  or
  g2585
  (
    n2484,
    n1755,
    n1648,
    n1790,
    n1873
  );


  and
  g2586
  (
    n2009,
    n1793,
    n1609,
    n1886,
    n1694
  );


  and
  g2587
  (
    n2152,
    n1620,
    n1782,
    n1676,
    n1792
  );


  or
  g2588
  (
    n2113,
    n1600,
    n1625,
    n1900,
    n1889
  );


  xor
  g2589
  (
    n1994,
    n1906,
    n1928,
    n1837,
    n1875
  );


  nor
  g2590
  (
    n2432,
    n1893,
    n1743,
    n1821,
    n1631
  );


  or
  g2591
  (
    n2671,
    n1930,
    n1611,
    n1638,
    n1852
  );


  xnor
  g2592
  (
    n2219,
    n1772,
    n1868,
    n1696,
    n1598
  );


  xnor
  g2593
  (
    n1970,
    n1752,
    n1689,
    n1668,
    n1899
  );


  xor
  g2594
  (
    n2504,
    n1829,
    n1814,
    n1909,
    n1656
  );


  nor
  g2595
  (
    n2080,
    n1645,
    n1709,
    n1747,
    n1832
  );


  nor
  g2596
  (
    n2241,
    n1742,
    n1698,
    n1833,
    n1616
  );


  nor
  g2597
  (
    n2130,
    n1720,
    n1733,
    n1672,
    n1736
  );


  xnor
  g2598
  (
    n2099,
    n1945,
    n1632,
    n1927,
    n1843
  );


  xor
  g2599
  (
    n2140,
    n1810,
    n1819,
    n1904,
    n1670
  );


  xnor
  g2600
  (
    n2197,
    n1912,
    n1821,
    n1765,
    n1679
  );


  nand
  g2601
  (
    n2542,
    n1715,
    n1614,
    n1911,
    n1675
  );


  and
  g2602
  (
    n2057,
    n1709,
    n1682,
    n1921,
    n1597
  );


  xor
  g2603
  (
    n2200,
    n1634,
    n1661,
    n1848,
    n1870
  );


  xor
  g2604
  (
    n2041,
    n1630,
    n1826,
    n1925,
    n1748
  );


  xor
  g2605
  (
    n2014,
    n1683,
    n1919,
    n1899,
    n1735
  );


  or
  g2606
  (
    n2139,
    n1789,
    n1923,
    n1859,
    n1891
  );


  and
  g2607
  (
    n2257,
    n1676,
    n1897,
    n1606,
    n1596
  );


  xnor
  g2608
  (
    n2505,
    n1621,
    n1698,
    n1626,
    n1839
  );


  nand
  g2609
  (
    n2114,
    n1934,
    n1810,
    n1708,
    n1703
  );


  or
  g2610
  (
    n2002,
    n1768,
    n1598,
    n1745,
    n1764
  );


  xnor
  g2611
  (
    n2135,
    n1808,
    n1799,
    n1593,
    n1714
  );


  or
  g2612
  (
    n2448,
    n1766,
    n1702,
    n1615,
    n1767
  );


  xor
  g2613
  (
    n2337,
    n1688,
    n1848,
    n1660,
    n1808
  );


  nand
  g2614
  (
    n2155,
    n1892,
    n1696,
    n1732,
    n1880
  );


  xor
  g2615
  (
    n2674,
    n1826,
    n1921,
    n1692,
    n1712
  );


  nor
  g2616
  (
    n2450,
    n1655,
    n1815,
    n1940,
    n1699
  );


  and
  g2617
  (
    n2273,
    n1784,
    n1718,
    n1607,
    n1935
  );


  and
  g2618
  (
    n2436,
    n1829,
    n1890,
    n1923,
    n1844
  );


  and
  g2619
  (
    n2211,
    n1607,
    n1795,
    n1741,
    n1783
  );


  nor
  g2620
  (
    n2314,
    n1674,
    n1725,
    n1933,
    n1619
  );


  or
  g2621
  (
    n2144,
    n1802,
    n1641,
    n1695,
    n1623
  );


  nor
  g2622
  (
    n2023,
    n1660,
    n1624,
    n1730,
    n1928
  );


  or
  g2623
  (
    n2207,
    n1792,
    n1809,
    n1932,
    n1796
  );


  nor
  g2624
  (
    n2118,
    n1723,
    n1710,
    n1867,
    n1859
  );


  or
  g2625
  (
    n2081,
    n1924,
    n1738,
    n1697,
    n1790
  );


  xnor
  g2626
  (
    n2431,
    n1677,
    n1774,
    n1811,
    n1597
  );


  nor
  g2627
  (
    n2652,
    n1865,
    n1796,
    n1882,
    n1613
  );


  xor
  g2628
  (
    n2280,
    n1903,
    n1662,
    n1790,
    n1813
  );


  nor
  g2629
  (
    n2412,
    n1626,
    n1653,
    n1943,
    n1740
  );


  xor
  g2630
  (
    n2045,
    n1657,
    n1750,
    n1403,
    n1756
  );


  or
  g2631
  (
    n2103,
    n1724,
    n1674,
    n1689
  );


  or
  g2632
  (
    n2663,
    n1664,
    n1779,
    n1686,
    n1836
  );


  xor
  g2633
  (
    n2681,
    n1800,
    n1795,
    n1863,
    n1874
  );


  and
  g2634
  (
    n2502,
    n1612,
    n1730,
    n1704,
    n1654
  );


  nand
  g2635
  (
    n2161,
    n1642,
    n1633,
    n1935,
    n1784
  );


  and
  g2636
  (
    n2302,
    n1706,
    n1406,
    n1751,
    n1676
  );


  xnor
  g2637
  (
    n2617,
    n1872,
    n1605,
    n1801,
    n1614
  );


  nand
  g2638
  (
    n2220,
    n1902,
    n1898,
    n1727,
    n1682
  );


  nor
  g2639
  (
    n2232,
    n1792,
    n1809,
    n1639,
    n1735
  );


  xor
  g2640
  (
    n2020,
    n1404,
    n1878,
    n1757,
    n1734
  );


  nor
  g2641
  (
    n2593,
    n1918,
    n1862,
    n1667,
    n1844
  );


  and
  g2642
  (
    n2481,
    n1768,
    n1878,
    n1889,
    n1818
  );


  or
  g2643
  (
    n2519,
    n1901,
    n1802,
    n1693,
    n1934
  );


  nor
  g2644
  (
    n1989,
    n1768,
    n1688,
    n1729,
    n1656
  );


  or
  g2645
  (
    n2678,
    n1773,
    n1711,
    n1692,
    n1933
  );


  nand
  g2646
  (
    n2490,
    n1721,
    n1729,
    n1731,
    n1892
  );


  xnor
  g2647
  (
    n2315,
    n1693,
    n1890,
    n1862,
    n1898
  );


  xor
  g2648
  (
    n1954,
    n1793,
    n1871,
    n1776,
    n1824
  );


  xor
  g2649
  (
    n2173,
    n1685,
    n1912,
    n1637,
    n1854
  );


  nor
  g2650
  (
    n2069,
    n1404,
    n1710,
    n1882,
    n1640
  );


  xor
  g2651
  (
    n2360,
    n1779,
    n1861,
    n1887,
    n1677
  );


  xnor
  g2652
  (
    n2127,
    n1761,
    n1923,
    n1816,
    n1690
  );


  xor
  g2653
  (
    n2282,
    n1709,
    n1906,
    n1880,
    n1902
  );


  or
  g2654
  (
    n2196,
    n1798,
    n1931,
    n1897,
    n1674
  );


  xor
  g2655
  (
    n2037,
    n1404,
    n1605,
    n1916,
    n1703
  );


  and
  g2656
  (
    n1953,
    n1855,
    n1611,
    n1640,
    n1867
  );


  nor
  g2657
  (
    n2078,
    n1655,
    n1841,
    n1806,
    n1943
  );


  or
  g2658
  (
    n2084,
    n1622,
    n1892,
    n1919,
    n1780
  );


  xnor
  g2659
  (
    n2445,
    n1824,
    n1724,
    n1732,
    n1763
  );


  and
  g2660
  (
    n2464,
    n1761,
    n1635,
    n1896,
    n1841
  );


  xnor
  g2661
  (
    n2133,
    n1669,
    n1870,
    n1838,
    n1628
  );


  and
  g2662
  (
    n2493,
    n1665,
    n1667,
    n1859,
    n1802
  );


  xnor
  g2663
  (
    n2296,
    n1617,
    n1633,
    n1798,
    n1851
  );


  nor
  g2664
  (
    n2558,
    n1678,
    n1885,
    n1782,
    n1594
  );


  xor
  g2665
  (
    n2485,
    n1603,
    n1737,
    n1794,
    n1825
  );


  xnor
  g2666
  (
    n1992,
    n1606,
    n1642,
    n1759,
    n1704
  );


  and
  g2667
  (
    n2146,
    n1852,
    n1785,
    n1783,
    n1766
  );


  or
  g2668
  (
    n2420,
    n1659,
    n1710,
    n1663,
    n1753
  );


  or
  g2669
  (
    n2641,
    n1811,
    n1869,
    n1786,
    n1910
  );


  nand
  g2670
  (
    n2645,
    n1668,
    n1723,
    n1649,
    n1672
  );


  nand
  g2671
  (
    n2774,
    n2662,
    n2661,
    n2392,
    n2639
  );


  xor
  g2672
  (
    n2833,
    n2336,
    n2675,
    n2428,
    n2423
  );


  xor
  g2673
  (
    n2708,
    n2257,
    n2185,
    n2261,
    n2457
  );


  xnor
  g2674
  (
    n2808,
    n1464,
    n2228,
    n2041,
    n1955
  );


  nor
  g2675
  (
    n2739,
    n2410,
    n2586,
    n2048,
    n2370
  );


  and
  g2676
  (
    n2725,
    n2262,
    n2439,
    n2074,
    n2326
  );


  and
  g2677
  (
    n2749,
    n1994,
    n2032,
    n2098,
    n2192
  );


  xnor
  g2678
  (
    n2784,
    n2095,
    n2462,
    n2176,
    n2210
  );


  xnor
  g2679
  (
    n2872,
    n2054,
    n2309,
    n2174,
    n1963
  );


  and
  g2680
  (
    n2705,
    n2397,
    n2629,
    n2282,
    n2212
  );


  nand
  g2681
  (
    n2712,
    n1986,
    n2444,
    n2345,
    n2484
  );


  nand
  g2682
  (
    n2895,
    n2502,
    n2250,
    n2243,
    n2209
  );


  xor
  g2683
  (
    KeyWire_0_25,
    n2355,
    n1586,
    n2574,
    n2623
  );


  and
  g2684
  (
    n2776,
    n1957,
    n2232,
    n1948,
    n2231
  );


  nand
  g2685
  (
    n2853,
    n2059,
    n2512,
    n2471,
    n2088
  );


  nor
  g2686
  (
    n2803,
    n2158,
    n2079,
    n2404,
    n2486
  );


  nor
  g2687
  (
    n2719,
    n2634,
    n2490,
    n2701,
    n1464
  );


  xnor
  g2688
  (
    n2817,
    n2476,
    n2686,
    n1969,
    n2625
  );


  and
  g2689
  (
    n2769,
    n2699,
    n2451,
    n2246,
    n1981
  );


  nand
  g2690
  (
    n2806,
    n2218,
    n2399,
    n2189,
    n2419
  );


  nor
  g2691
  (
    n2873,
    n2253,
    n2148,
    n2585,
    n2275
  );


  xor
  g2692
  (
    n2721,
    n2598,
    n2622,
    n2655,
    n2556
  );


  nor
  g2693
  (
    n2790,
    n2702,
    n2422,
    n2468,
    n2251
  );


  and
  g2694
  (
    n2802,
    n2518,
    n2456,
    n2010,
    n2413
  );


  xor
  g2695
  (
    n2877,
    n2371,
    n2296,
    n2260,
    n2416
  );


  xor
  g2696
  (
    n2723,
    n2269,
    n2455,
    n2299,
    n1995
  );


  xor
  g2697
  (
    n2846,
    n2443,
    n2684,
    n2138,
    n2614
  );


  xnor
  g2698
  (
    n2761,
    n2638,
    n2433,
    n2412,
    n2626
  );


  nor
  g2699
  (
    n2762,
    n2482,
    n2503,
    n2594,
    n2698
  );


  and
  g2700
  (
    n2869,
    n2303,
    n2459,
    n2115,
    n2267
  );


  nand
  g2701
  (
    n2830,
    n2328,
    n2018,
    n2526,
    n2449
  );


  and
  g2702
  (
    n2879,
    n2070,
    n2230,
    n2248,
    n2057
  );


  xnor
  g2703
  (
    n2842,
    n2333,
    n2234,
    n2665,
    n2297
  );


  or
  g2704
  (
    n2825,
    n2441,
    n2663,
    n2483,
    n2613
  );


  and
  g2705
  (
    n2747,
    n2164,
    n2124,
    n2086,
    n2601
  );


  xnor
  g2706
  (
    n2801,
    n2245,
    n2538,
    n2378,
    n1990
  );


  xor
  g2707
  (
    n2779,
    n2201,
    n2649,
    n2331,
    n2052
  );


  xor
  g2708
  (
    n2850,
    n2347,
    n2571,
    n1968,
    n2628
  );


  xor
  g2709
  (
    n2887,
    n2259,
    n2568,
    n2699,
    n2562
  );


  nor
  g2710
  (
    n2718,
    n2437,
    n1587,
    n2266,
    n2151
  );


  nand
  g2711
  (
    n2861,
    n2026,
    n2380,
    n2056,
    n2701
  );


  nand
  g2712
  (
    n2811,
    n2472,
    n2161,
    n2697,
    n2363
  );


  or
  g2713
  (
    n2840,
    n2017,
    n2335,
    n1977,
    n1966
  );


  xor
  g2714
  (
    n2709,
    n2159,
    n2188,
    n2353,
    n2035
  );


  xnor
  g2715
  (
    n2734,
    n2386,
    n2310,
    n2507,
    n2227
  );


  nor
  g2716
  (
    n2824,
    n2244,
    n2620,
    n2187,
    n2533
  );


  xor
  g2717
  (
    n2897,
    n2489,
    n2016,
    n2172,
    n2669
  );


  nand
  g2718
  (
    n2768,
    n2298,
    n1947,
    n2170,
    n2668
  );


  xnor
  g2719
  (
    n2793,
    n2401,
    n2315,
    n2178,
    n2678
  );


  xnor
  g2720
  (
    n2717,
    n2208,
    n2168,
    n2539,
    n2082
  );


  nor
  g2721
  (
    n2829,
    n2534,
    n2121,
    n2621,
    n2196
  );


  or
  g2722
  (
    n2795,
    n2285,
    n2249,
    n2136,
    n2063
  );


  xor
  g2723
  (
    n2868,
    n2013,
    n2368,
    n2465,
    n2195
  );


  or
  g2724
  (
    n2780,
    n1956,
    n2509,
    n2475,
    n2633
  );


  nand
  g2725
  (
    n2822,
    n2140,
    n2525,
    n1951,
    n2153
  );


  nand
  g2726
  (
    n2771,
    n2203,
    n2101,
    n2306,
    n2458
  );


  xor
  g2727
  (
    n2763,
    n2036,
    n2184,
    n2350,
    n2100
  );


  and
  g2728
  (
    n2820,
    n2434,
    n2332,
    n2608,
    n2144
  );


  or
  g2729
  (
    n2875,
    n2589,
    n2450,
    n2391,
    n2076
  );


  xnor
  g2730
  (
    n2890,
    n2008,
    n2143,
    n2308,
    n2690
  );


  nand
  g2731
  (
    n2819,
    n1958,
    n2666,
    n2006,
    n2582
  );


  nor
  g2732
  (
    n2744,
    n2390,
    n2104,
    n2454,
    n2223
  );


  nor
  g2733
  (
    n2816,
    n2356,
    n2181,
    n2011,
    n2654
  );


  nand
  g2734
  (
    n2810,
    n2190,
    n2557,
    n2432,
    n2569
  );


  nor
  g2735
  (
    n2798,
    n2674,
    n2109,
    n1964,
    n2039
  );


  xor
  g2736
  (
    n2727,
    n2570,
    n2300,
    n2116,
    n2519
  );


  or
  g2737
  (
    n2773,
    n2517,
    n2435,
    n2235,
    n2566
  );


  nor
  g2738
  (
    n2728,
    n2497,
    n1959,
    n2364,
    n2200
  );


  or
  g2739
  (
    n2745,
    n2087,
    n2068,
    n2580,
    n2119
  );


  and
  g2740
  (
    n2860,
    n2292,
    n2155,
    n2236,
    n2645
  );


  and
  g2741
  (
    n2854,
    n2213,
    n2049,
    n2421,
    n2438
  );


  or
  g2742
  (
    n2781,
    n2498,
    n2581,
    n2617,
    n2053
  );


  or
  g2743
  (
    n2792,
    n1979,
    n2263,
    n1973,
    n2521
  );


  xnor
  g2744
  (
    n2710,
    n2508,
    n2448,
    n2516,
    n2090
  );


  or
  g2745
  (
    n2716,
    n2703,
    n2286,
    n2609,
    n2376
  );


  or
  g2746
  (
    n2837,
    n2340,
    n2131,
    n2550,
    n2112
  );


  nand
  g2747
  (
    n2866,
    n2311,
    n2099,
    n2327,
    n1952
  );


  nand
  g2748
  (
    n2863,
    n2004,
    n2513,
    n2113,
    n2106
  );


  nand
  g2749
  (
    n2874,
    n2487,
    n2288,
    n2214,
    n2372
  );


  nor
  g2750
  (
    n2714,
    n2092,
    n2123,
    n2549,
    n2352
  );


  or
  g2751
  (
    n2736,
    n2691,
    n2660,
    n2061,
    n1586
  );


  and
  g2752
  (
    n2799,
    n2445,
    n2329,
    n2702,
    n2268
  );


  or
  g2753
  (
    n2794,
    n2426,
    n2491,
    n2648,
    n2229
  );


  xnor
  g2754
  (
    KeyWire_0_22,
    n2595,
    n2646,
    n2207,
    n2652
  );


  xnor
  g2755
  (
    n2889,
    n2393,
    n2351,
    n2069,
    n2276
  );


  xnor
  g2756
  (
    n2839,
    n2072,
    n2673,
    n2511,
    n2206
  );


  xnor
  g2757
  (
    n2892,
    n2077,
    n2256,
    n1974,
    n2478
  );


  xor
  g2758
  (
    n2729,
    n2657,
    n2480,
    n2405,
    n2653
  );


  nor
  g2759
  (
    n2730,
    n2545,
    n2182,
    n2702,
    n2024
  );


  xor
  g2760
  (
    n2775,
    n2563,
    n2081,
    n2224,
    n2414
  );


  xor
  g2761
  (
    n2843,
    n2682,
    n2107,
    n2211,
    n2611
  );


  and
  g2762
  (
    n2855,
    n2692,
    n1975,
    n2312,
    n2021
  );


  xnor
  g2763
  (
    n2807,
    n2398,
    n2567,
    n2463,
    n2552
  );


  and
  g2764
  (
    n2870,
    n2022,
    n2671,
    n2014,
    n2152
  );


  nor
  g2765
  (
    n2789,
    n2627,
    n2323,
    n2542,
    n2314
  );


  nor
  g2766
  (
    n2788,
    n2096,
    n2150,
    n2640,
    n2317
  );


  nor
  g2767
  (
    n2859,
    n2418,
    n2241,
    n2656,
    n2033
  );


  and
  g2768
  (
    n2847,
    n2546,
    n2066,
    n1464,
    n2344
  );


  nor
  g2769
  (
    n2876,
    n2252,
    n2409,
    n2280,
    n2377
  );


  xnor
  g2770
  (
    n2838,
    n2658,
    n2341,
    n2374,
    n2381
  );


  nor
  g2771
  (
    n2735,
    n2367,
    n2584,
    n2637,
    n2366
  );


  nor
  g2772
  (
    n2764,
    n2278,
    n2424,
    n2075,
    n2084
  );


  and
  g2773
  (
    n2885,
    n2167,
    n2301,
    n2305,
    n2264
  );


  and
  g2774
  (
    n2894,
    n2681,
    n1585,
    n2283,
    n1971
  );


  and
  g2775
  (
    n2791,
    n2596,
    n2643,
    n2202,
    n2129
  );


  xor
  g2776
  (
    n2858,
    n2293,
    n2003,
    n2064,
    n2703
  );


  xnor
  g2777
  (
    n2831,
    n2551,
    n1976,
    n2126,
    n2284
  );


  and
  g2778
  (
    n2898,
    n2067,
    n2334,
    n2590,
    n2670
  );


  xor
  g2779
  (
    n2759,
    n2179,
    n2051,
    n2149,
    n2142
  );


  xor
  g2780
  (
    n2884,
    n2388,
    n2034,
    n2700,
    n2474
  );


  or
  g2781
  (
    n2755,
    n2289,
    n2577,
    n2488,
    n2122
  );


  nand
  g2782
  (
    n2731,
    n2604,
    n2005,
    n2447,
    n2565
  );


  nor
  g2783
  (
    n2800,
    n2023,
    n2560,
    n2616,
    n2031
  );


  nor
  g2784
  (
    n2845,
    n2515,
    n2470,
    n2173,
    n2103
  );


  or
  g2785
  (
    n2782,
    n2233,
    n2685,
    n2644,
    n2226
  );


  or
  g2786
  (
    n2751,
    n2346,
    n2607,
    n2215,
    n2411
  );


  nor
  g2787
  (
    n2754,
    n2029,
    n2091,
    n2169,
    n2677
  );


  nor
  g2788
  (
    n2804,
    n2313,
    n2591,
    n2216,
    n2541
  );


  xor
  g2789
  (
    n2722,
    n2060,
    n2528,
    n2602,
    n2290
  );


  or
  g2790
  (
    n2821,
    n2558,
    n1978,
    n2651,
    n2429
  );


  nor
  g2791
  (
    n2886,
    n2400,
    n2544,
    n2572,
    n2680
  );


  nor
  g2792
  (
    n2765,
    n2045,
    n2177,
    n2019,
    n2171
  );


  nor
  g2793
  (
    n2888,
    n2009,
    n2495,
    n2073,
    n2242
  );


  xor
  g2794
  (
    n2881,
    n2078,
    n2117,
    n2385,
    n2265
  );


  or
  g2795
  (
    n2812,
    n2700,
    n1960,
    n2561,
    n2536
  );


  or
  g2796
  (
    n2772,
    n2324,
    n1993,
    n2320,
    n2436
  );


  xnor
  g2797
  (
    n2733,
    n2238,
    n2325,
    n1992,
    n2473
  );


  and
  g2798
  (
    n2720,
    n2632,
    n2615,
    n2531,
    n2559
  );


  xnor
  g2799
  (
    n2856,
    n2395,
    n2065,
    n2270,
    n2291
  );


  xnor
  g2800
  (
    n2748,
    n2461,
    n2025,
    n1988,
    n2132
  );


  xor
  g2801
  (
    n2741,
    n2403,
    n2453,
    n2287,
    n2357
  );


  xor
  g2802
  (
    n2737,
    n1587,
    n2348,
    n2481,
    n2120
  );


  nand
  g2803
  (
    n2743,
    n2071,
    n2683,
    n2688,
    n2575
  );


  or
  g2804
  (
    n2849,
    n1997,
    n2540,
    n2040,
    n1953
  );


  nand
  g2805
  (
    n2740,
    n1586,
    n2406,
    n2612,
    n2427
  );


  nand
  g2806
  (
    n2857,
    n2693,
    n2479,
    n2362,
    n2446
  );


  and
  g2807
  (
    n2797,
    n2619,
    n2452,
    n2493,
    n2030
  );


  nor
  g2808
  (
    n2834,
    n2672,
    n2631,
    n2321,
    n1989
  );


  xor
  g2809
  (
    n2809,
    n2137,
    n2330,
    n2699,
    n1983
  );


  and
  g2810
  (
    n2777,
    n2514,
    n2166,
    n2139,
    n2695
  );


  or
  g2811
  (
    n2750,
    n2012,
    n2219,
    n2277,
    n2105
  );


  xor
  g2812
  (
    n2848,
    n2553,
    n2543,
    n2094,
    n2373
  );


  nor
  g2813
  (
    n2832,
    n2379,
    n2440,
    n2430,
    n2204
  );


  or
  g2814
  (
    n2827,
    n2500,
    n2295,
    n2055,
    n2588
  );


  nand
  g2815
  (
    n2871,
    n2358,
    n2630,
    n2548,
    n2271
  );


  or
  g2816
  (
    n2767,
    n2186,
    n2191,
    n2038,
    n2349
  );


  or
  g2817
  (
    n2815,
    n2135,
    n2273,
    n2389,
    n1950
  );


  nand
  g2818
  (
    n2883,
    n2042,
    n2110,
    n2576,
    n2460
  );


  or
  g2819
  (
    n2805,
    n2494,
    n2027,
    n1996,
    n2647
  );


  and
  g2820
  (
    n2841,
    n2587,
    n2431,
    n1586,
    n1987
  );


  xor
  g2821
  (
    n2787,
    n2319,
    n2659,
    n2156,
    n2597
  );


  nor
  g2822
  (
    n2704,
    n2510,
    n2102,
    n2307,
    n2080
  );


  or
  g2823
  (
    n2785,
    n2700,
    n2599,
    n2592,
    n2467
  );


  xnor
  g2824
  (
    n2766,
    n2279,
    n2322,
    n2047,
    n2028
  );


  nor
  g2825
  (
    n2864,
    n2636,
    n2361,
    n1998,
    n1954
  );


  nand
  g2826
  (
    n2786,
    n2492,
    n2664,
    n1962,
    n2425
  );


  nor
  g2827
  (
    n2865,
    n2281,
    n2442,
    n2134,
    n2485
  );


  nor
  g2828
  (
    n2713,
    n2111,
    n2125,
    n2221,
    n2464
  );


  xor
  g2829
  (
    n2844,
    n2205,
    n2650,
    n1980,
    n2127
  );


  nand
  g2830
  (
    n2752,
    n2506,
    n2524,
    n2579,
    n2058
  );


  nand
  g2831
  (
    n2893,
    n2338,
    n2523,
    n2369,
    n2520
  );


  nand
  g2832
  (
    n2896,
    n2396,
    n2147,
    n1949,
    n1587
  );


  and
  g2833
  (
    n2756,
    n2505,
    n2239,
    n2583,
    n2618
  );


  xnor
  g2834
  (
    n2882,
    n2007,
    n2530,
    n2679,
    n2194
  );


  xor
  g2835
  (
    n2818,
    n2175,
    n2193,
    n2160,
    n2694
  );


  xnor
  g2836
  (
    n2770,
    n2703,
    n1965,
    n2605,
    n1970
  );


  xnor
  g2837
  (
    n2746,
    n2365,
    n2183,
    n2083,
    n2145
  );


  and
  g2838
  (
    n2778,
    n2154,
    n2118,
    n2339,
    n2294
  );


  nand
  g2839
  (
    n2880,
    n2222,
    n2220,
    n2407,
    n2408
  );


  nand
  g2840
  (
    n2813,
    n2532,
    n2255,
    n2600,
    n2217
  );


  nor
  g2841
  (
    n2828,
    n1999,
    n2635,
    n2108,
    n1585
  );


  xor
  g2842
  (
    n2826,
    n2573,
    n2676,
    n2337,
    n1967
  );


  xor
  g2843
  (
    n2814,
    n2387,
    n2130,
    n2527,
    n2163
  );


  nor
  g2844
  (
    n2796,
    n2529,
    n1464,
    n2247,
    n1984
  );


  nand
  g2845
  (
    n2706,
    n2199,
    n2420,
    n2272,
    n2062
  );


  xor
  g2846
  (
    n2823,
    n2302,
    n2044,
    n2624,
    n2258
  );


  or
  g2847
  (
    n2783,
    n2225,
    n2383,
    n2050,
    n2667
  );


  xnor
  g2848
  (
    n2836,
    n2354,
    n2237,
    n2696,
    n2146
  );


  xor
  g2849
  (
    n2724,
    n2180,
    n2157,
    n2555,
    n2496
  );


  nand
  g2850
  (
    n2891,
    n2043,
    n2384,
    n2522,
    n2318
  );


  xnor
  g2851
  (
    n2760,
    n2342,
    n2085,
    n2394,
    n2564
  );


  xor
  g2852
  (
    n2711,
    n2197,
    n2165,
    n2114,
    n1961
  );


  xor
  g2853
  (
    n2852,
    n2360,
    n2603,
    n2133,
    n2089
  );


  nand
  g2854
  (
    n2753,
    n2000,
    n2593,
    n2304,
    n2382
  );


  xnor
  g2855
  (
    n2757,
    n2547,
    n2687,
    n2578,
    n2046
  );


  or
  g2856
  (
    n2732,
    n2402,
    n2641,
    n2417,
    n2375
  );


  and
  g2857
  (
    n2726,
    n2316,
    n2343,
    n2469,
    n2606
  );


  or
  g2858
  (
    n2707,
    n2128,
    n2093,
    n1982,
    n2701
  );


  and
  g2859
  (
    n2758,
    n2642,
    n2415,
    n2141,
    n2162
  );


  or
  g2860
  (
    n2862,
    n2359,
    n2240,
    n2501,
    n2015
  );


  nand
  g2861
  (
    n2715,
    n2254,
    n2610,
    n1991,
    n2037
  );


  xnor
  g2862
  (
    n2851,
    n2537,
    n2504,
    n2020,
    n2002
  );


  nand
  g2863
  (
    n2835,
    n2689,
    n2477,
    n2499,
    n2535
  );


  and
  g2864
  (
    n2742,
    n1985,
    n2274,
    n2466,
    n1972
  );


  nand
  g2865
  (
    n2878,
    n2001,
    n2554,
    n2198,
    n2097
  );


  nor
  g2866
  (
    n2910,
    n2780,
    n2862,
    n2721,
    n2741
  );


  xnor
  g2867
  (
    n2938,
    n2818,
    n2821,
    n2819,
    n2884
  );


  xor
  g2868
  (
    n2929,
    n2742,
    n2766,
    n2772,
    n2723
  );


  or
  g2869
  (
    n2948,
    n2729,
    n2733,
    n2739,
    n2713
  );


  or
  g2870
  (
    n2933,
    n2858,
    n2710,
    n2761,
    n1591
  );


  nand
  g2871
  (
    n2908,
    n2894,
    n2730,
    n2783,
    n2715
  );


  or
  g2872
  (
    n2905,
    n2711,
    n2833,
    n2850,
    n2828
  );


  nor
  g2873
  (
    n2921,
    n2865,
    n2795,
    n2806,
    n2848
  );


  nor
  g2874
  (
    n2944,
    n2752,
    n2746,
    n2814,
    n2797
  );


  nand
  g2875
  (
    n2952,
    n2837,
    n2842,
    n2734,
    n1588
  );


  nand
  g2876
  (
    n2911,
    n2890,
    n2878,
    n2807,
    n2722
  );


  nand
  g2877
  (
    n2946,
    n2705,
    n2801,
    n2817,
    n2748
  );


  nor
  g2878
  (
    n2939,
    n2835,
    n2871,
    n2770,
    n2897
  );


  xor
  g2879
  (
    n2951,
    n2775,
    n2784,
    n2743,
    n2836
  );


  or
  g2880
  (
    n2932,
    n2829,
    n2843,
    n2876,
    n2892
  );


  or
  g2881
  (
    n2902,
    n2808,
    n2767,
    n1592,
    n2792
  );


  nand
  g2882
  (
    n2909,
    n2898,
    n2869,
    n2725,
    n2861
  );


  xor
  g2883
  (
    n2925,
    n2840,
    n2726,
    n2773,
    n2812
  );


  xor
  g2884
  (
    n2926,
    n2769,
    n2895,
    n1592,
    n2882
  );


  nor
  g2885
  (
    n2941,
    n2854,
    n2708,
    n2781,
    n2859
  );


  xnor
  g2886
  (
    n2900,
    n2872,
    n2896,
    n2738,
    n2802
  );


  or
  g2887
  (
    n2903,
    n2866,
    n2809,
    n2864,
    n2707
  );


  xor
  g2888
  (
    n2945,
    n2847,
    n2893,
    n2747,
    n2791
  );


  and
  g2889
  (
    n2942,
    n2724,
    n2716,
    n1590,
    n2778
  );


  and
  g2890
  (
    n2914,
    n2728,
    n2860,
    n2834,
    n2887
  );


  xor
  g2891
  (
    n2950,
    n2785,
    n2827,
    n2815,
    n2868
  );


  xor
  g2892
  (
    n2917,
    n2793,
    n2714,
    n2841,
    n2880
  );


  xor
  g2893
  (
    n2931,
    n2853,
    n1589,
    n2756,
    n2844
  );


  and
  g2894
  (
    KeyWire_0_28,
    n2765,
    n2790,
    n2857,
    n1590
  );


  or
  g2895
  (
    n2920,
    n2838,
    n2735,
    n2754,
    n2846
  );


  xor
  g2896
  (
    n2923,
    n2763,
    n2874,
    n2831,
    n2855
  );


  xor
  g2897
  (
    KeyWire_0_16,
    n2779,
    n2881,
    n2788,
    n2856
  );


  nor
  g2898
  (
    n2913,
    n2737,
    n2744,
    n2825,
    n2740
  );


  xor
  g2899
  (
    n2922,
    n2717,
    n2867,
    n2820,
    n2777
  );


  xor
  g2900
  (
    n2918,
    n2888,
    n2800,
    n2852,
    n1592
  );


  or
  g2901
  (
    n2901,
    n2851,
    n2719,
    n2863,
    n1589
  );


  nand
  g2902
  (
    n2937,
    n1591,
    n2839,
    n2811,
    n2706
  );


  or
  g2903
  (
    n2907,
    n2745,
    n2830,
    n2759,
    n2879
  );


  nor
  g2904
  (
    n2915,
    n2768,
    n2787,
    n2758,
    n1587
  );


  xor
  g2905
  (
    n2943,
    n2751,
    n2822,
    n2891,
    n2755
  );


  xnor
  g2906
  (
    n2927,
    n1589,
    n2762,
    n2823,
    n2877
  );


  xnor
  g2907
  (
    n2919,
    n2776,
    n1590,
    n2720,
    n2794
  );


  nor
  g2908
  (
    n2947,
    n2750,
    n2774,
    n2883,
    n2870
  );


  or
  g2909
  (
    n2906,
    n2718,
    n2798,
    n2889,
    n2816
  );


  xor
  g2910
  (
    n2935,
    n1588,
    n2712,
    n2885,
    n2771
  );


  xor
  g2911
  (
    n2904,
    n2796,
    n2886,
    n2826,
    n2786
  );


  and
  g2912
  (
    n2916,
    n2704,
    n2709,
    n2805,
    n2727
  );


  xor
  g2913
  (
    n2899,
    n2813,
    n2731,
    n2804,
    n1588
  );


  or
  g2914
  (
    n2924,
    n1592,
    n2873,
    n2757,
    n2753
  );


  xnor
  g2915
  (
    n2912,
    n2824,
    n2845,
    n2760,
    n1589
  );


  or
  g2916
  (
    n2928,
    n2875,
    n2803,
    n1590,
    n1591
  );


  and
  g2917
  (
    n2934,
    n2799,
    n2782,
    n2810,
    n2789
  );


  and
  g2918
  (
    n2949,
    n2749,
    n2736,
    n1591,
    n2832
  );


  and
  g2919
  (
    n2930,
    n2849,
    n2732,
    n2764,
    n1588
  );


  or
  g2920
  (
    n2988,
    n6,
    n2946,
    n9,
    n24
  );


  or
  g2921
  (
    n2992,
    n15,
    n2932,
    n2948,
    n20
  );


  xor
  g2922
  (
    n2996,
    n1430,
    n19,
    n2933,
    n1429
  );


  xor
  g2923
  (
    n2953,
    n1426,
    n2926,
    n2925,
    n1424
  );


  xnor
  g2924
  (
    n2991,
    n24,
    n2952,
    n10
  );


  or
  g2925
  (
    n2969,
    n2931,
    n26,
    n24,
    n2918
  );


  and
  g2926
  (
    n2956,
    n22,
    n22,
    n29,
    n1422
  );


  xnor
  g2927
  (
    n2975,
    n1421,
    n2908,
    n9,
    n19
  );


  nor
  g2928
  (
    n2990,
    n24,
    n18,
    n2899,
    n7
  );


  xnor
  g2929
  (
    n2978,
    n30,
    n29,
    n2950,
    n2912
  );


  nor
  g2930
  (
    n2994,
    n2945,
    n25,
    n26,
    n10
  );


  xnor
  g2931
  (
    n2974,
    n2938,
    n31,
    n2935,
    n1424
  );


  xor
  g2932
  (
    n2986,
    n17,
    n1423,
    n1422,
    n2907
  );


  nor
  g2933
  (
    n2984,
    n1430,
    n18,
    n2941,
    n1426
  );


  nand
  g2934
  (
    n2995,
    n2947,
    n27,
    n30,
    n17
  );


  and
  g2935
  (
    n2976,
    n1428,
    n25,
    n28,
    n2903
  );


  and
  g2936
  (
    n3002,
    n1427,
    n11,
    n30,
    n2927
  );


  xnor
  g2937
  (
    n2957,
    n19,
    n14,
    n2934,
    n16
  );


  or
  g2938
  (
    n2965,
    n1429,
    n2920,
    n26,
    n1432
  );


  xnor
  g2939
  (
    n2985,
    n8,
    n14,
    n2914,
    n1431
  );


  nor
  g2940
  (
    n2958,
    n31,
    n1427,
    n15
  );


  or
  g2941
  (
    n2962,
    n32,
    n23,
    n28,
    n2905
  );


  and
  g2942
  (
    n2981,
    n32,
    n18,
    n2944,
    n1421
  );


  and
  g2943
  (
    n2967,
    n2915,
    n27,
    n2929,
    n32
  );


  xnor
  g2944
  (
    n2989,
    n30,
    n1431,
    n2913,
    n10
  );


  and
  g2945
  (
    n2959,
    n1429,
    n2911,
    n17,
    n2943
  );


  xor
  g2946
  (
    n2968,
    n18,
    n8,
    n21,
    n1424
  );


  or
  g2947
  (
    n2971,
    n2951,
    n6,
    n32,
    n14
  );


  or
  g2948
  (
    n2993,
    n26,
    n16,
    n21,
    n1430
  );


  or
  g2949
  (
    n2961,
    n1425,
    n1428,
    n14,
    n7
  );


  or
  g2950
  (
    n2960,
    n2937,
    n7,
    n1431,
    n2921
  );


  or
  g2951
  (
    n3004,
    n20,
    n1422,
    n2939,
    n2904
  );


  nor
  g2952
  (
    n2955,
    n2949,
    n25,
    n2930,
    n6
  );


  xnor
  g2953
  (
    n2972,
    n13,
    n2902,
    n17,
    n23
  );


  xnor
  g2954
  (
    n2980,
    n2917,
    n12,
    n1423
  );


  xnor
  g2955
  (
    n2966,
    n2906,
    n22,
    n2942,
    n1431
  );


  nor
  g2956
  (
    n2977,
    n9,
    n2916,
    n21,
    n1432
  );


  xnor
  g2957
  (
    n2970,
    n31,
    n1422,
    n2923,
    n1423
  );


  and
  g2958
  (
    n2997,
    n1427,
    n12,
    n8,
    n9
  );


  and
  g2959
  (
    KeyWire_0_29,
    n8,
    n13,
    n11,
    n1423
  );


  or
  g2960
  (
    n2979,
    n2928,
    n1432,
    n2909,
    n2900
  );


  xor
  g2961
  (
    n2964,
    n13,
    n11,
    n1430,
    n27
  );


  and
  g2962
  (
    n2987,
    n2936,
    n25,
    n1425,
    n2901
  );


  nor
  g2963
  (
    n2983,
    n2940,
    n29,
    n20,
    n2910
  );


  xnor
  g2964
  (
    n3001,
    n1426,
    n22,
    n2922,
    n28
  );


  xnor
  g2965
  (
    n2998,
    n16,
    n23,
    n1429
  );


  nor
  g2966
  (
    n2982,
    n28,
    n16,
    n20,
    n2924
  );


  xnor
  g2967
  (
    n3000,
    n31,
    n1421,
    n15,
    n1428
  );


  xnor
  g2968
  (
    n2954,
    n1427,
    n1426,
    n7,
    n21
  );


  nor
  g2969
  (
    n3003,
    n13,
    n1424,
    n1428,
    n1425
  );


  xor
  g2970
  (
    n2963,
    n1425,
    n11,
    n29,
    n2919
  );


  or
  g2971
  (
    n2999,
    n27,
    n19,
    n12,
    n1432
  );


  nor
  g2972
  (
    n3007,
    n1449,
    n1445,
    n2981,
    n2965
  );


  nand
  g2973
  (
    n3013,
    n1437,
    n2956,
    n1439,
    n1440
  );


  nor
  g2974
  (
    n3032,
    n2983,
    n49,
    n3002,
    n2955
  );


  nor
  g2975
  (
    n3020,
    n2969,
    n1445,
    n3000,
    n1439
  );


  xor
  g2976
  (
    n3008,
    n1438,
    n1440,
    n2963,
    n1445
  );


  xor
  g2977
  (
    n3005,
    n2967,
    n2973,
    n1449,
    n1444
  );


  and
  g2978
  (
    KeyWire_0_14,
    n2977,
    n1439,
    n1446,
    n2993
  );


  and
  g2979
  (
    n3006,
    n2954,
    n2961,
    n2979,
    n1437
  );


  or
  g2980
  (
    n3009,
    n1436,
    n1447,
    n2953
  );


  xnor
  g2981
  (
    n3011,
    n1438,
    n1442,
    n3003,
    n2966
  );


  nand
  g2982
  (
    n3024,
    n1440,
    n1445,
    n2999,
    n1444
  );


  nor
  g2983
  (
    n3014,
    n2957,
    n2997,
    n2959,
    n1449
  );


  xor
  g2984
  (
    n3017,
    n1437,
    n3001,
    n1442,
    n2972
  );


  and
  g2985
  (
    n3019,
    n2991,
    n1443,
    n2990,
    n1447
  );


  xor
  g2986
  (
    n3018,
    n3004,
    n2971,
    n2975,
    n2992
  );


  xnor
  g2987
  (
    n3031,
    n2995,
    n49,
    n1439,
    n2996
  );


  and
  g2988
  (
    n3016,
    n1446,
    n2970,
    n1448,
    n1441
  );


  xnor
  g2989
  (
    n3029,
    n1437,
    n2962,
    n1441,
    n1447
  );


  xnor
  g2990
  (
    n3010,
    n1444,
    n2985,
    n2989,
    n50
  );


  xor
  g2991
  (
    n3030,
    n1446,
    n2982,
    n1438,
    n1449
  );


  xnor
  g2992
  (
    KeyWire_0_1,
    n50,
    n1442,
    n1448,
    n1441
  );


  xnor
  g2993
  (
    n3023,
    n2976,
    n2978,
    n2980,
    n1448
  );


  or
  g2994
  (
    n3026,
    n2968,
    n2960,
    n1444,
    n2998
  );


  or
  g2995
  (
    n3022,
    n1442,
    n1448,
    n2988,
    n2987
  );


  xor
  g2996
  (
    n3012,
    n2986,
    n1446,
    n1443,
    n2994
  );


  xor
  g2997
  (
    n3021,
    n50,
    n50,
    n1443,
    n1441
  );


  xor
  g2998
  (
    n3028,
    n1438,
    n1440,
    n2974,
    n2984
  );


  nor
  g2999
  (
    n3015,
    n2964,
    n49,
    n2958,
    n1443
  );


  xnor
  KeyGate_0_0
  (
    n1215,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n3025,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n522,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1650,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n388,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n1049,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1636,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n2107,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1571,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1943,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n734,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n2138,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n2227,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n393,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n3027,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n614,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n2940,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n2223,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n2676,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n464,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n2163,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n90,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n2738,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n924,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1484,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n2867,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n419,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n2006,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n2936,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n2973,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n94,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1780,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


