// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1057_14_11 written by SynthGen on 2021/05/24 19:42:16
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1057_14_11 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19,
 n771, n1065, n1076, n1074, n1071, n1070, n1067, n1069,
 n1075, n1073, n1061, n1057, n1064, n1068, n1072, n1058,
 n1066, n1055, n1056, n1063, n1062, n1059, n1060);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19;

output n771, n1065, n1076, n1074, n1071, n1070, n1067, n1069,
 n1075, n1073, n1061, n1057, n1064, n1068, n1072, n1058,
 n1066, n1055, n1056, n1063, n1062, n1059, n1060;

wire n20, n21, n22, n23, n24, n25, n26, n27,
 n28, n29, n30, n31, n32, n33, n34, n35,
 n36, n37, n38, n39, n40, n41, n42, n43,
 n44, n45, n46, n47, n48, n49, n50, n51,
 n52, n53, n54, n55, n56, n57, n58, n59,
 n60, n61, n62, n63, n64, n65, n66, n67,
 n68, n69, n70, n71, n72, n73, n74, n75,
 n76, n77, n78, n79, n80, n81, n82, n83,
 n84, n85, n86, n87, n88, n89, n90, n91,
 n92, n93, n94, n95, n96, n97, n98, n99,
 n100, n101, n102, n103, n104, n105, n106, n107,
 n108, n109, n110, n111, n112, n113, n114, n115,
 n116, n117, n118, n119, n120, n121, n122, n123,
 n124, n125, n126, n127, n128, n129, n130, n131,
 n132, n133, n134, n135, n136, n137, n138, n139,
 n140, n141, n142, n143, n144, n145, n146, n147,
 n148, n149, n150, n151, n152, n153, n154, n155,
 n156, n157, n158, n159, n160, n161, n162, n163,
 n164, n165, n166, n167, n168, n169, n170, n171,
 n172, n173, n174, n175, n176, n177, n178, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n189, n190, n191, n192, n193, n194, n195,
 n196, n197, n198, n199, n200, n201, n202, n203,
 n204, n205, n206, n207, n208, n209, n210, n211,
 n212, n213, n214, n215, n216, n217, n218, n219,
 n220, n221, n222, n223, n224, n225, n226, n227,
 n228, n229, n230, n231, n232, n233, n234, n235,
 n236, n237, n238, n239, n240, n241, n242, n243,
 n244, n245, n246, n247, n248, n249, n250, n251,
 n252, n253, n254, n255, n256, n257, n258, n259,
 n260, n261, n262, n263, n264, n265, n266, n267,
 n268, n269, n270, n271, n272, n273, n274, n275,
 n276, n277, n278, n279, n280, n281, n282, n283,
 n284, n285, n286, n287, n288, n289, n290, n291,
 n292, n293, n294, n295, n296, n297, n298, n299,
 n300, n301, n302, n303, n304, n305, n306, n307,
 n308, n309, n310, n311, n312, n313, n314, n315,
 n316, n317, n318, n319, n320, n321, n322, n323,
 n324, n325, n326, n327, n328, n329, n330, n331,
 n332, n333, n334, n335, n336, n337, n338, n339,
 n340, n341, n342, n343, n344, n345, n346, n347,
 n348, n349, n350, n351, n352, n353, n354, n355,
 n356, n357, n358, n359, n360, n361, n362, n363,
 n364, n365, n366, n367, n368, n369, n370, n371,
 n372, n373, n374, n375, n376, n377, n378, n379,
 n380, n381, n382, n383, n384, n385, n386, n387,
 n388, n389, n390, n391, n392, n393, n394, n395,
 n396, n397, n398, n399, n400, n401, n402, n403,
 n404, n405, n406, n407, n408, n409, n410, n411,
 n412, n413, n414, n415, n416, n417, n418, n419,
 n420, n421, n422, n423, n424, n425, n426, n427,
 n428, n429, n430, n431, n432, n433, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n634, n635,
 n636, n637, n638, n639, n640, n641, n642, n643,
 n644, n645, n646, n647, n648, n649, n650, n651,
 n652, n653, n654, n655, n656, n657, n658, n659,
 n660, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685, n686, n687, n688, n689, n690, n691,
 n692, n693, n694, n695, n696, n697, n698, n699,
 n700, n701, n702, n703, n704, n705, n706, n707,
 n708, n709, n710, n711, n712, n713, n714, n715,
 n716, n717, n718, n719, n720, n721, n722, n723,
 n724, n725, n726, n727, n728, n729, n730, n731,
 n732, n733, n734, n735, n736, n737, n738, n739,
 n740, n741, n742, n743, n744, n745, n746, n747,
 n748, n749, n750, n751, n752, n753, n754, n755,
 n756, n757, n758, n759, n760, n761, n762, n763,
 n764, n765, n766, n767, n768, n769, n770, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n865, n866, n867, n868,
 n869, n870, n871, n872, n873, n874, n875, n876,
 n877, n878, n879, n880, n881, n882, n883, n884,
 n885, n886, n887, n888, n889, n890, n891, n892,
 n893, n894, n895, n896, n897, n898, n899, n900,
 n901, n902, n903, n904, n905, n906, n907, n908,
 n909, n910, n911, n912, n913, n914, n915, n916,
 n917, n918, n919, n920, n921, n922, n923, n924,
 n925, n926, n927, n928, n929, n930, n931, n932,
 n933, n934, n935, n936, n937, n938, n939, n940,
 n941, n942, n943, n944, n945, n946, n947, n948,
 n949, n950, n951, n952, n953, n954, n955, n956,
 n957, n958, n959, n960, n961, n962, n963, n964,
 n965, n966, n967, n968, n969, n970, n971, n972,
 n973, n974, n975, n976, n977, n978, n979, n980,
 n981, n982, n983, n984, n985, n986, n987, n988,
 n989, n990, n991, n992, n993, n994, n995, n996,
 n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
 n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
 n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
 n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
 n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
 n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
 n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
 n1053, n1054;

buf  g0 (n90, n11);
not  g1 (n93, n8);
not  g2 (n79, n4);
not  g3 (n53, n13);
buf  g4 (n49, n10);
not  g5 (n77, n18);
buf  g6 (n70, n15);
not  g7 (n33, n12);
buf  g8 (n60, n9);
not  g9 (n34, n5);
buf  g10 (n78, n14);
buf  g11 (n65, n19);
buf  g12 (n21, n16);
not  g13 (n61, n19);
not  g14 (n75, n19);
buf  g15 (n26, n14);
buf  g16 (n32, n4);
buf  g17 (n86, n5);
not  g18 (n76, n8);
not  g19 (n43, n1);
buf  g20 (n48, n13);
not  g21 (n30, n14);
not  g22 (n41, n15);
buf  g23 (n91, n3);
not  g24 (n50, n15);
buf  g25 (n51, n7);
not  g26 (n67, n12);
not  g27 (n58, n1);
buf  g28 (n69, n2);
not  g29 (n22, n13);
not  g30 (n94, n7);
buf  g31 (n52, n7);
not  g32 (n27, n18);
not  g33 (n42, n4);
buf  g34 (n59, n3);
buf  g35 (n84, n4);
not  g36 (n71, n8);
not  g37 (n56, n6);
buf  g38 (n82, n12);
not  g39 (n20, n11);
buf  g40 (n39, n8);
not  g41 (n57, n6);
buf  g42 (n92, n2);
buf  g43 (n38, n17);
buf  g44 (n73, n9);
not  g45 (n68, n7);
not  g46 (n87, n17);
buf  g47 (n54, n1);
buf  g48 (n95, n19);
buf  g49 (n64, n2);
not  g50 (n72, n6);
not  g51 (n83, n15);
not  g52 (n31, n14);
not  g53 (n88, n6);
not  g54 (n40, n16);
buf  g55 (n74, n1);
buf  g56 (n89, n9);
not  g57 (n36, n3);
buf  g58 (n37, n17);
buf  g59 (n25, n5);
buf  g60 (n47, n16);
buf  g61 (n62, n17);
not  g62 (n44, n10);
buf  g63 (n24, n18);
not  g64 (n63, n5);
buf  g65 (n45, n18);
not  g66 (n29, n10);
not  g67 (n23, n16);
buf  g68 (n35, n12);
not  g69 (n46, n11);
not  g70 (n28, n2);
buf  g71 (n66, n10);
buf  g72 (n81, n13);
buf  g73 (n55, n9);
not  g74 (n85, n11);
not  g75 (n80, n3);
buf  g76 (n322, n56);
not  g77 (n366, n91);
buf  g78 (n265, n23);
not  g79 (n299, n41);
not  g80 (n237, n22);
buf  g81 (n104, n47);
buf  g82 (n157, n33);
not  g83 (n128, n68);
not  g84 (n107, n57);
buf  g85 (n148, n93);
buf  g86 (n315, n89);
not  g87 (n217, n50);
not  g88 (n290, n53);
not  g89 (n206, n57);
not  g90 (n369, n80);
buf  g91 (n150, n46);
not  g92 (n133, n42);
not  g93 (n121, n32);
not  g94 (n342, n94);
not  g95 (n240, n28);
buf  g96 (n296, n90);
not  g97 (n362, n56);
buf  g98 (n295, n49);
not  g99 (n102, n22);
buf  g100 (n360, n20);
buf  g101 (n142, n72);
not  g102 (n226, n30);
buf  g103 (n147, n59);
not  g104 (n208, n24);
not  g105 (n381, n89);
not  g106 (n307, n56);
buf  g107 (n215, n77);
buf  g108 (n389, n32);
buf  g109 (n123, n83);
not  g110 (n251, n21);
not  g111 (n122, n73);
not  g112 (n168, n47);
not  g113 (n309, n48);
not  g114 (n340, n82);
buf  g115 (n98, n73);
not  g116 (n328, n75);
buf  g117 (n184, n28);
not  g118 (n269, n80);
not  g119 (n278, n34);
buf  g120 (n117, n85);
not  g121 (n187, n83);
buf  g122 (n285, n27);
not  g123 (n384, n36);
not  g124 (n140, n39);
not  g125 (n195, n44);
not  g126 (n186, n63);
buf  g127 (n247, n52);
not  g128 (n266, n64);
not  g129 (n308, n51);
buf  g130 (n363, n84);
not  g131 (n116, n90);
buf  g132 (n234, n44);
buf  g133 (n352, n89);
not  g134 (n270, n26);
not  g135 (n317, n55);
not  g136 (n106, n88);
buf  g137 (n244, n40);
buf  g138 (n219, n91);
buf  g139 (n159, n60);
buf  g140 (n382, n41);
not  g141 (n292, n36);
not  g142 (n203, n69);
not  g143 (n262, n75);
buf  g144 (n174, n33);
not  g145 (n141, n30);
not  g146 (n127, n45);
not  g147 (n232, n48);
not  g148 (n139, n93);
buf  g149 (n282, n39);
not  g150 (n109, n58);
not  g151 (n151, n63);
buf  g152 (n349, n74);
buf  g153 (n199, n38);
buf  g154 (n257, n61);
buf  g155 (n129, n94);
not  g156 (n275, n47);
buf  g157 (n385, n63);
buf  g158 (n331, n62);
not  g159 (n394, n57);
buf  g160 (n119, n49);
buf  g161 (n396, n80);
not  g162 (n332, n62);
buf  g163 (n303, n77);
not  g164 (n231, n25);
buf  g165 (n306, n45);
not  g166 (n281, n71);
not  g167 (n143, n23);
not  g168 (n388, n92);
not  g169 (n361, n54);
not  g170 (n101, n31);
not  g171 (n166, n71);
buf  g172 (n372, n34);
buf  g173 (n393, n61);
buf  g174 (n209, n42);
not  g175 (n132, n70);
buf  g176 (n334, n92);
not  g177 (n387, n58);
buf  g178 (n204, n84);
not  g179 (n347, n29);
not  g180 (n351, n52);
buf  g181 (n239, n54);
buf  g182 (n355, n79);
not  g183 (n200, n58);
not  g184 (n326, n25);
not  g185 (n254, n38);
not  g186 (n249, n52);
buf  g187 (n344, n55);
not  g188 (n310, n73);
not  g189 (n259, n45);
not  g190 (n210, n90);
buf  g191 (n377, n70);
buf  g192 (n304, n83);
not  g193 (n131, n42);
not  g194 (n300, n71);
buf  g195 (n325, n35);
buf  g196 (n96, n54);
buf  g197 (n291, n87);
buf  g198 (n346, n66);
buf  g199 (n162, n43);
buf  g200 (n341, n93);
not  g201 (n316, n64);
buf  g202 (n323, n82);
buf  g203 (n177, n46);
not  g204 (n164, n53);
not  g205 (n336, n88);
not  g206 (n379, n35);
not  g207 (n190, n29);
not  g208 (n124, n74);
buf  g209 (n179, n30);
buf  g210 (n343, n94);
not  g211 (n213, n61);
not  g212 (n156, n67);
buf  g213 (n192, n69);
not  g214 (n223, n42);
not  g215 (n176, n20);
not  g216 (n233, n38);
buf  g217 (n264, n46);
buf  g218 (n335, n84);
buf  g219 (n197, n67);
buf  g220 (n145, n86);
not  g221 (n297, n81);
buf  g222 (n161, n91);
buf  g223 (n294, n23);
not  g224 (n312, n55);
not  g225 (n155, n66);
not  g226 (n365, n34);
buf  g227 (n238, n81);
buf  g228 (n110, n70);
buf  g229 (n392, n21);
not  g230 (n178, n31);
not  g231 (n152, n50);
not  g232 (n271, n80);
not  g233 (n327, n55);
buf  g234 (n284, n34);
buf  g235 (n373, n35);
buf  g236 (n207, n47);
not  g237 (n134, n86);
not  g238 (n380, n60);
buf  g239 (n391, n37);
not  g240 (n277, n29);
not  g241 (n293, n95);
buf  g242 (n205, n51);
buf  g243 (n321, n72);
buf  g244 (n286, n78);
buf  g245 (n170, n60);
buf  g246 (n337, n85);
not  g247 (n339, n86);
not  g248 (n202, n58);
not  g249 (n144, n85);
buf  g250 (n256, n25);
not  g251 (n149, n71);
not  g252 (n263, n78);
buf  g253 (n158, n33);
buf  g254 (n198, n88);
not  g255 (n287, n75);
not  g256 (n242, n76);
buf  g257 (n398, n65);
buf  g258 (n279, n95);
buf  g259 (n189, n72);
not  g260 (n246, n43);
not  g261 (n105, n24);
not  g262 (n350, n84);
buf  g263 (n111, n29);
buf  g264 (n320, n62);
not  g265 (n274, n41);
buf  g266 (n248, n92);
not  g267 (n114, n76);
buf  g268 (n193, n40);
buf  g269 (n333, n93);
not  g270 (n224, n36);
buf  g271 (n188, n37);
not  g272 (n367, n50);
not  g273 (n358, n75);
buf  g274 (n97, n59);
buf  g275 (n301, n57);
buf  g276 (n314, n59);
buf  g277 (n253, n65);
buf  g278 (n125, n78);
buf  g279 (n163, n61);
not  g280 (n115, n67);
buf  g281 (n108, n28);
buf  g282 (n368, n33);
buf  g283 (n180, n30);
buf  g284 (n216, n21);
not  g285 (n130, n50);
not  g286 (n330, n24);
not  g287 (n260, n73);
not  g288 (n126, n54);
buf  g289 (n99, n65);
buf  g290 (n235, n82);
buf  g291 (n222, n69);
buf  g292 (n250, n68);
not  g293 (n298, n83);
not  g294 (n305, n40);
not  g295 (n374, n22);
buf  g296 (n230, n79);
buf  g297 (n169, n81);
not  g298 (n338, n78);
not  g299 (n364, n68);
buf  g300 (n112, n74);
not  g301 (n243, n43);
not  g302 (n218, n67);
buf  g303 (n345, n25);
not  g304 (n329, n32);
not  g305 (n245, n26);
not  g306 (n182, n36);
not  g307 (n252, n76);
not  g308 (n241, n51);
buf  g309 (n185, n45);
buf  g310 (n227, n90);
buf  g311 (n319, n81);
buf  g312 (n288, n31);
not  g313 (n376, n53);
buf  g314 (n181, n87);
buf  g315 (n214, n38);
buf  g316 (n370, n27);
buf  g317 (n354, n27);
buf  g318 (n153, n74);
buf  g319 (n280, n79);
not  g320 (n258, n92);
not  g321 (n318, n77);
not  g322 (n302, n49);
buf  g323 (n118, n64);
not  g324 (n255, n39);
buf  g325 (n113, n64);
buf  g326 (n103, n56);
buf  g327 (n220, n39);
not  g328 (n324, n89);
buf  g329 (n378, n20);
buf  g330 (n383, n35);
not  g331 (n160, n77);
buf  g332 (n313, n52);
not  g333 (n191, n66);
buf  g334 (n283, n70);
buf  g335 (n356, n59);
not  g336 (n136, n79);
buf  g337 (n268, n63);
not  g338 (n261, n23);
buf  g339 (n276, n37);
not  g340 (n311, n46);
not  g341 (n375, n49);
buf  g342 (n289, n21);
buf  g343 (n173, n48);
buf  g344 (n175, n69);
not  g345 (n194, n82);
buf  g346 (n267, n87);
not  g347 (n183, n60);
not  g348 (n236, n62);
buf  g349 (n167, n22);
buf  g350 (n390, n26);
not  g351 (n100, n40);
not  g352 (n353, n88);
not  g353 (n212, n72);
buf  g354 (n154, n24);
buf  g355 (n357, n43);
buf  g356 (n371, n65);
not  g357 (n135, n20);
buf  g358 (n172, n27);
not  g359 (n171, n41);
not  g360 (n273, n76);
buf  g361 (n397, n86);
not  g362 (n348, n95);
not  g363 (n211, n28);
buf  g364 (n146, n44);
buf  g365 (n225, n94);
not  g366 (n138, n44);
buf  g367 (n395, n37);
buf  g368 (n386, n87);
buf  g369 (n137, n53);
buf  g370 (n120, n31);
not  g371 (n229, n85);
buf  g372 (n359, n66);
not  g373 (n221, n32);
not  g374 (n272, n48);
not  g375 (n196, n68);
buf  g376 (n165, n26);
buf  g377 (n228, n51);
buf  g378 (n201, n91);
buf  g379 (n624, n299);
not  g380 (n580, n357);
not  g381 (n556, n391);
buf  g382 (n412, n333);
not  g383 (n546, n376);
buf  g384 (n420, n313);
buf  g385 (n692, n215);
buf  g386 (n621, n191);
not  g387 (n493, n97);
not  g388 (n726, n380);
not  g389 (n471, n358);
not  g390 (n419, n369);
not  g391 (n442, n370);
not  g392 (n399, n390);
buf  g393 (n633, n221);
buf  g394 (n522, n253);
not  g395 (n504, n106);
not  g396 (n694, n201);
not  g397 (n429, n380);
not  g398 (n541, n133);
buf  g399 (n464, n199);
not  g400 (n590, n305);
buf  g401 (n611, n236);
buf  g402 (n698, n331);
buf  g403 (n720, n352);
not  g404 (n618, n359);
buf  g405 (n413, n357);
not  g406 (n647, n352);
not  g407 (n655, n372);
buf  g408 (n502, n185);
buf  g409 (n542, n183);
buf  g410 (n450, n225);
not  g411 (n607, n143);
not  g412 (n482, n208);
buf  g413 (n461, n390);
buf  g414 (n718, n272);
buf  g415 (n729, n322);
not  g416 (n747, n373);
buf  g417 (n595, n279);
not  g418 (n717, n368);
buf  g419 (n731, n114);
buf  g420 (n660, n344);
not  g421 (n734, n351);
not  g422 (n416, n149);
buf  g423 (n564, n275);
not  g424 (n439, n101);
not  g425 (n634, n388);
buf  g426 (n544, n323);
buf  g427 (n437, n381);
buf  g428 (n689, n379);
not  g429 (n638, n285);
not  g430 (n481, n338);
not  g431 (n579, n281);
not  g432 (n536, n301);
buf  g433 (n631, n232);
not  g434 (n679, n391);
buf  g435 (n555, n138);
not  g436 (n661, n386);
buf  g437 (n581, n240);
not  g438 (n497, n246);
not  g439 (n530, n242);
not  g440 (n748, n354);
buf  g441 (n709, n342);
buf  g442 (n714, n359);
not  g443 (n430, n227);
buf  g444 (n737, n355);
not  g445 (n742, n361);
buf  g446 (n405, n375);
buf  g447 (n623, n388);
not  g448 (n514, n283);
buf  g449 (n699, n269);
buf  g450 (n575, n344);
not  g451 (n697, n117);
not  g452 (n646, n142);
not  g453 (n553, n200);
buf  g454 (n677, n147);
buf  g455 (n500, n145);
not  g456 (n417, n366);
buf  g457 (n423, n336);
buf  g458 (n670, n156);
buf  g459 (n507, n315);
buf  g460 (n441, n312);
not  g461 (n418, n166);
not  g462 (n715, n367);
not  g463 (n627, n186);
buf  g464 (n604, n198);
buf  g465 (n733, n338);
not  g466 (n577, n298);
not  g467 (n512, n123);
not  g468 (n434, n377);
not  g469 (n616, n254);
buf  g470 (n691, n274);
buf  g471 (n465, n357);
not  g472 (n613, n118);
buf  g473 (n445, n293);
buf  g474 (n549, n360);
buf  g475 (n448, n165);
not  g476 (n738, n104);
buf  g477 (n444, n126);
not  g478 (n603, n245);
buf  g479 (n723, n169);
buf  g480 (n470, n328);
not  g481 (n548, n243);
buf  g482 (n711, n390);
buf  g483 (n705, n140);
not  g484 (n727, n187);
not  g485 (n440, n181);
buf  g486 (n532, n152);
buf  g487 (n523, n360);
buf  g488 (n732, n369);
buf  g489 (n710, n192);
buf  g490 (n740, n116);
not  g491 (n642, n334);
buf  g492 (n659, n353);
buf  g493 (n678, n220);
not  g494 (n400, n105);
not  g495 (n456, n378);
buf  g496 (n645, n373);
buf  g497 (n712, n290);
not  g498 (n650, n150);
buf  g499 (n432, n125);
not  g500 (n612, n174);
not  g501 (n680, n99);
not  g502 (n508, n136);
buf  g503 (n449, n258);
buf  g504 (n630, n334);
buf  g505 (n510, n311);
buf  g506 (n498, n259);
buf  g507 (n495, n160);
buf  g508 (n436, n226);
buf  g509 (n672, n154);
buf  g510 (n540, n383);
buf  g511 (n640, n379);
not  g512 (n473, n110);
not  g513 (n695, n155);
not  g514 (n704, n261);
not  g515 (n414, n196);
buf  g516 (n489, n251);
buf  g517 (n597, n282);
not  g518 (n629, n324);
not  g519 (n501, n341);
buf  g520 (n518, n300);
buf  g521 (n739, n354);
not  g522 (n703, n108);
buf  g523 (n681, n264);
not  g524 (n584, n382);
buf  g525 (n469, n375);
not  g526 (n422, n205);
buf  g527 (n520, n332);
buf  g528 (n525, n129);
not  g529 (n455, n249);
buf  g530 (n503, n379);
buf  g531 (n639, n276);
not  g532 (n543, n350);
buf  g533 (n499, n361);
not  g534 (n620, n308);
buf  g535 (n665, n364);
buf  g536 (n528, n347);
not  g537 (n632, n332);
not  g538 (n606, n351);
buf  g539 (n466, n389);
buf  g540 (n459, n137);
not  g541 (n669, n378);
buf  g542 (n708, n189);
buf  g543 (n526, n350);
not  g544 (n609, n153);
not  g545 (n447, n250);
buf  g546 (n568, n273);
not  g547 (n566, n384);
buf  g548 (n599, n223);
not  g549 (n651, n139);
not  g550 (n683, n386);
not  g551 (n668, n376);
not  g552 (n676, n372);
not  g553 (n690, n134);
buf  g554 (n460, n381);
buf  g555 (n454, n387);
buf  g556 (n458, n361);
buf  g557 (n602, n268);
buf  g558 (n664, n260);
not  g559 (n467, n348);
not  g560 (n476, n288);
buf  g561 (n598, n96);
not  g562 (n558, n204);
not  g563 (n741, n121);
buf  g564 (n527, n190);
buf  g565 (n744, n325);
not  g566 (n538, n148);
not  g567 (n474, n157);
not  g568 (n594, n228);
buf  g569 (n673, n381);
buf  g570 (n657, n337);
buf  g571 (n516, n385);
buf  g572 (n517, n144);
buf  g573 (n625, n321);
buf  g574 (n614, n314);
not  g575 (n636, n202);
not  g576 (n529, n341);
not  g577 (n656, n267);
not  g578 (n666, n329);
not  g579 (n452, n365);
buf  g580 (n574, n368);
not  g581 (n728, n241);
not  g582 (n572, n318);
buf  g583 (n571, n359);
buf  g584 (n674, n257);
buf  g585 (n589, n178);
buf  g586 (n648, n280);
buf  g587 (n426, n353);
not  g588 (n610, n319);
buf  g589 (n537, n384);
buf  g590 (n750, n320);
not  g591 (n688, n331);
buf  g592 (n685, n349);
not  g593 (n539, n327);
not  g594 (n496, n211);
buf  g595 (n684, n231);
not  g596 (n488, n238);
not  g597 (n535, n107);
not  g598 (n743, n307);
buf  g599 (n506, n385);
buf  g600 (n573, n214);
buf  g601 (n494, n162);
not  g602 (n479, n366);
buf  g603 (n588, n369);
buf  g604 (n578, n224);
not  g605 (n463, n376);
not  g606 (n401, n353);
not  g607 (n706, n367);
buf  g608 (n561, n203);
not  g609 (n424, n374);
not  g610 (n600, n336);
buf  g611 (n722, n248);
buf  g612 (n713, n366);
buf  g613 (n736, n335);
buf  g614 (n428, n349);
not  g615 (n560, n339);
buf  g616 (n457, n387);
not  g617 (n730, n306);
not  g618 (n567, n286);
buf  g619 (n505, n291);
not  g620 (n485, n345);
not  g621 (n586, n380);
not  g622 (n487, n345);
not  g623 (n591, n363);
not  g624 (n408, n364);
buf  g625 (n702, n218);
not  g626 (n596, n180);
buf  g627 (n663, n158);
not  g628 (n582, n230);
buf  g629 (n626, n141);
not  g630 (n545, n330);
buf  g631 (n643, n164);
not  g632 (n745, n216);
not  g633 (n667, n115);
buf  g634 (n622, n333);
not  g635 (n484, n170);
not  g636 (n653, n98);
not  g637 (n721, n206);
not  g638 (n480, n175);
buf  g639 (n521, n302);
not  g640 (n477, n168);
buf  g641 (n403, n335);
buf  g642 (n707, n340);
not  g643 (n451, n365);
not  g644 (n701, n256);
buf  g645 (n601, n356);
not  g646 (n415, n365);
not  g647 (n511, n348);
buf  g648 (n411, n102);
buf  g649 (n402, n383);
buf  g650 (n443, n356);
not  g651 (n431, n292);
not  g652 (n686, n316);
buf  g653 (n565, n362);
buf  g654 (n554, n284);
not  g655 (n483, n351);
not  g656 (n658, n130);
not  g657 (n746, n378);
buf  g658 (n519, n161);
not  g659 (n749, n239);
not  g660 (n559, n119);
buf  g661 (n587, n207);
not  g662 (n700, n382);
not  g663 (n409, n159);
not  g664 (n682, n194);
buf  g665 (n433, n271);
buf  g666 (n592, n358);
not  g667 (n628, n343);
not  g668 (n421, n128);
not  g669 (n675, n382);
buf  g670 (n593, n263);
buf  g671 (n513, n339);
not  g672 (n550, n362);
not  g673 (n492, n103);
not  g674 (n583, n184);
not  g675 (n515, n247);
buf  g676 (n427, n213);
not  g677 (n478, n372);
not  g678 (n534, n296);
not  g679 (n615, n167);
buf  g680 (n608, n289);
not  g681 (n425, n352);
not  g682 (n435, n370);
not  g683 (n562, n131);
buf  g684 (n491, n265);
not  g685 (n662, n360);
buf  g686 (n570, n368);
not  g687 (n547, n132);
buf  g688 (n475, n337);
not  g689 (n533, n217);
not  g690 (n453, n355);
buf  g691 (n637, n244);
buf  g692 (n563, n347);
not  g693 (n644, n277);
buf  g694 (n641, n358);
buf  g695 (n649, n188);
not  g696 (n605, n342);
not  g697 (n531, n356);
not  g698 (n407, n177);
not  g699 (n719, n210);
not  g700 (n585, n252);
not  g701 (n509, n171);
buf  g702 (n410, n349);
not  g703 (n524, n287);
buf  g704 (n490, n255);
not  g705 (n652, n163);
buf  g706 (n635, n383);
not  g707 (n735, n363);
not  g708 (n619, n303);
buf  g709 (n557, n377);
not  g710 (n406, n384);
buf  g711 (n671, n135);
buf  g712 (n486, n309);
not  g713 (n472, n237);
buf  g714 (n654, n374);
or   g715 (n462, n389, n295, n355, n127);
nand g716 (n438, n151, n362, n179, n233);
xnor g717 (n468, n120, n367, n386, n310);
and  g718 (n446, n219, n350, n370, n304);
and  g719 (n693, n377, n374, n270, n266);
and  g720 (n687, n262, n375, n193, n173);
nor  g721 (n552, n278, n209, n124, n195);
or   g722 (n569, n387, n234, n172, n389);
nand g723 (n404, n112, n176, n348, n297);
xnor g724 (n725, n222, n182, n326, n294);
xnor g725 (n617, n122, n100, n146, n235);
nand g726 (n696, n113, n197, n346, n317);
xnor g727 (n716, n373, n371, n111, n346);
nand g728 (n576, n371, n385, n212, n363);
nand g729 (n724, n229, n109, n388, n340);
nand g730 (n551, n364, n343, n354, n371);
xnor g731 (n754, n433, n480, n439, n502);
and  g732 (n760, n469, n495, n478, n421);
and  g733 (n767, n509, n526, n504, n527);
nor  g734 (n777, n416, n473, n459, n520);
nand g735 (n753, n529, n420, n506, n419);
nor  g736 (n765, n496, n524, n413, n431);
nand g737 (n758, n513, n514, n485, n501);
or   g738 (n771, n487, n425, n445, n522);
and  g739 (n768, n517, n458, n424, n508);
xnor g740 (n751, n484, n400, n523, n452);
and  g741 (n757, n482, n438, n455, n410);
and  g742 (n772, n449, n494, n491, n462);
xnor g743 (n755, n446, n476, n401, n479);
xnor g744 (n759, n407, n515, n481, n429);
and  g745 (n761, n486, n456, n464, n411);
or   g746 (n781, n519, n525, n500, n426);
xor  g747 (n778, n471, n403, n448, n460);
xor  g748 (n773, n530, n470, n477, n443);
nor  g749 (n775, n488, n434, n518, n512);
nand g750 (n756, n427, n467, n493, n475);
nor  g751 (n769, n447, n503, n505, n441);
and  g752 (n776, n414, n440, n406, n490);
xor  g753 (n766, n450, n428, n474, n528);
nor  g754 (n752, n489, n498, n417, n451);
nand g755 (n770, n453, n466, n454, n497);
nand g756 (n779, n408, n405, n442, n510);
nor  g757 (n782, n444, n507, n492, n465);
xor  g758 (n774, n472, n511, n432, n483);
or   g759 (n783, n516, n415, n521, n499);
nor  g760 (n763, n436, n461, n422, n457);
nand g761 (n762, n463, n430, n399, n412);
and  g762 (n764, n423, n468, n402, n418);
and  g763 (n780, n409, n435, n437, n404);
or   g764 (n812, n553, n545, n591, n574);
xor  g765 (n796, n609, n758, n778, n589);
nand g766 (n802, n606, n623, n780, n611);
or   g767 (n787, n766, n603, n575, n626);
and  g768 (n785, n586, n578, n579, n563);
xnor g769 (n795, n543, n617, n776, n584);
and  g770 (n814, n752, n595, n567, n583);
xor  g771 (n804, n544, n767, n756, n592);
and  g772 (n811, n775, n624, n546, n548);
or   g773 (n792, n618, n601, n533, n572);
nand g774 (n808, n566, n772, n612, n588);
xnor g775 (n789, n620, n764, n607, n569);
xnor g776 (n784, n759, n549, n762, n757);
or   g777 (n810, n550, n782, n777, n753);
xnor g778 (n809, n577, n593, n604, n568);
or   g779 (n800, n608, n561, n783, n538);
and  g780 (n801, n769, n770, n570, n536);
xor  g781 (n807, n754, n555, n779, n773);
xnor g782 (n815, n594, n587, n547, n534);
xnor g783 (n793, n613, n616, n560, n576);
nand g784 (n813, n597, n622, n571, n581);
xor  g785 (n794, n539, n556, n541, n559);
xor  g786 (n788, n552, n771, n573, n535);
nand g787 (n803, n781, n557, n760, n619);
and  g788 (n805, n598, n554, n537, n602);
nand g789 (n786, n605, n551, n614, n585);
and  g790 (n799, n540, n564, n558, n582);
nand g791 (n790, n768, n755, n531, n625);
and  g792 (n791, n600, n532, n580, n763);
and  g793 (n797, n774, n621, n761, n610);
or   g794 (n806, n565, n562, n615, n599);
or   g795 (n798, n542, n765, n596, n590);
buf  g796 (n843, n805);
buf  g797 (n830, n798);
buf  g798 (n838, n788);
buf  g799 (n850, n800);
not  g800 (n840, n801);
buf  g801 (n837, n804);
not  g802 (n819, n796);
not  g803 (n845, n802);
buf  g804 (n853, n789);
not  g805 (n820, n802);
buf  g806 (n832, n786);
buf  g807 (n839, n800);
buf  g808 (n821, n794);
not  g809 (n855, n808);
buf  g810 (n828, n805);
not  g811 (n856, n790);
buf  g812 (n834, n801);
buf  g813 (n844, n795);
not  g814 (n859, n797);
not  g815 (n842, n806);
not  g816 (n816, n796);
buf  g817 (n846, n810);
buf  g818 (n848, n786);
not  g819 (n825, n804);
xor  g820 (n818, n795, n793, n785, n807);
nor  g821 (n857, n798, n786, n791, n803);
xor  g822 (n824, n791, n788, n809);
xor  g823 (n854, n809, n787, n784, n803);
or   g824 (n858, n794, n794, n801, n807);
and  g825 (n831, n785, n806, n791, n810);
nor  g826 (n827, n802, n806, n795, n797);
xor  g827 (n860, n790, n788, n784, n792);
or   g828 (n836, n808, n799, n798, n793);
nand g829 (n823, n806, n785, n810, n790);
xnor g830 (n849, n785, n796, n789, n791);
nor  g831 (n841, n804, n809, n801, n786);
or   g832 (n822, n803, n799, n794, n792);
xnor g833 (n829, n792, n784, n807);
xnor g834 (n852, n800, n799, n808, n789);
and  g835 (n833, n793, n803, n799, n804);
or   g836 (n835, n807, n805, n810, n797);
xnor g837 (n847, n805, n798, n787, n808);
or   g838 (n817, n797, n790, n787, n792);
xnor g839 (n826, n802, n809, n796, n793);
nor  g840 (n851, n787, n789, n800, n795);
not  g841 (n864, n832);
buf  g842 (n867, n824);
not  g843 (n874, n823);
buf  g844 (n876, n825);
buf  g845 (n879, n826);
not  g846 (n877, n828);
not  g847 (n875, n817);
buf  g848 (n863, n822);
not  g849 (n861, n835);
not  g850 (n873, n819);
not  g851 (n880, n818);
not  g852 (n868, n827);
buf  g853 (n870, n820);
not  g854 (n865, n829);
buf  g855 (n878, n830);
buf  g856 (n866, n834);
buf  g857 (n871, n831);
not  g858 (n872, n816);
not  g859 (n862, n833);
buf  g860 (n869, n821);
not  g861 (n882, n868);
buf  g862 (n886, n874);
buf  g863 (n895, n866);
not  g864 (n893, n863);
buf  g865 (n897, n870);
buf  g866 (n898, n864);
buf  g867 (n883, n873);
buf  g868 (n885, n873);
not  g869 (n892, n861);
not  g870 (n894, n870);
not  g871 (n896, n869);
buf  g872 (n884, n867);
not  g873 (n881, n862);
not  g874 (n888, n872);
not  g875 (n887, n872);
not  g876 (n890, n871);
not  g877 (n891, n865);
not  g878 (n889, n871);
not  g879 (n938, n896);
buf  g880 (n950, n889);
not  g881 (n932, n875);
not  g882 (n934, n883);
not  g883 (n918, n885);
not  g884 (n926, n889);
buf  g885 (n953, n892);
buf  g886 (n928, n893);
buf  g887 (n946, n890);
not  g888 (n903, n887);
buf  g889 (n941, n886);
not  g890 (n900, n886);
buf  g891 (n925, n883);
buf  g892 (n930, n887);
buf  g893 (n921, n893);
not  g894 (n949, n897);
not  g895 (n937, n891);
not  g896 (n924, n898);
not  g897 (n913, n888);
buf  g898 (n951, n882);
buf  g899 (n919, n882);
buf  g900 (n907, n888);
not  g901 (n948, n881);
not  g902 (n911, n893);
buf  g903 (n909, n881);
buf  g904 (n929, n874);
buf  g905 (n905, n886);
buf  g906 (n935, n895);
not  g907 (n923, n885);
not  g908 (n943, n897);
not  g909 (n942, n890);
not  g910 (n917, n876);
buf  g911 (n899, n889);
not  g912 (n933, n892);
buf  g913 (n939, n884);
not  g914 (n904, n896);
buf  g915 (n947, n875);
not  g916 (n902, n898);
buf  g917 (n944, n876);
not  g918 (n914, n891);
not  g919 (n927, n898);
buf  g920 (n922, n887);
not  g921 (n931, n895);
buf  g922 (n952, n894);
buf  g923 (n912, n882);
not  g924 (n915, n888);
not  g925 (n910, n894);
buf  g926 (n936, n892);
buf  g927 (n906, n884);
not  g928 (n901, n896);
buf  g929 (n908, n895);
buf  g930 (n916, n885);
not  g931 (n945, n894);
nand g932 (n940, n890, n891, n881);
xor  g933 (n920, n897, n884, n898, n883);
nand g934 (n967, n926, n919, n904, n910);
and  g935 (n964, n928, n918, n906, n923);
and  g936 (n957, n916, n917, n926, n902);
xor  g937 (n954, n911, n907, n913, n899);
and  g938 (n960, n914, n927, n916, n929);
xor  g939 (n956, n904, n900, n905, n920);
xor  g940 (n965, n899, n925, n908, n906);
or   g941 (n966, n907, n925, n914, n931);
and  g942 (n955, n932, n902, n912, n901);
xor  g943 (n970, n910, n920, n931, n919);
and  g944 (n963, n915, n913, n927, n912);
nand g945 (n968, n930, n930, n909, n911);
nor  g946 (n962, n900, n903, n915, n917);
nand g947 (n958, n932, n901, n928, n929);
xnor g948 (n961, n905, n918, n903, n921);
nand g949 (n969, n909, n921, n923, n922);
or   g950 (n959, n908, n924, n922);
buf  g951 (n971, n957);
buf  g952 (n974, n954);
not  g953 (n972, n955);
not  g954 (n973, n956);
xnor g955 (n975, n971, n971, n967, n974);
xnor g956 (n985, n391, n966, n396, n965);
and  g957 (n983, n973, n974, n971, n878);
xor  g958 (n981, n974, n960, n392);
xor  g959 (n990, n973, n974, n395, n971);
xnor g960 (n988, n393, n972, n395);
nand g961 (n984, n812, n392, n972, n393);
xor  g962 (n980, n393, n878, n812, n811);
xor  g963 (n978, n972, n630, n629, n811);
and  g964 (n987, n812, n877, n811, n933);
xnor g965 (n989, n962, n396, n973, n395);
nand g966 (n982, n877, n961, n964, n969);
nand g967 (n977, n631, n879, n394, n811);
or   g968 (n986, n394, n973, n963, n397);
xor  g969 (n976, n959, n968, n396, n958);
xor  g970 (n979, n970, n628, n394, n627);
or   g971 (n1050, n648, n989, n710, n979);
xnor g972 (n1022, n977, n983, n666, n684);
or   g973 (n1026, n698, n688, n879, n686);
xor  g974 (n1006, n661, n851, n986, n978);
and  g975 (n998, n669, n697, n683, n646);
and  g976 (n1008, n939, n986, n95, n815);
nor  g977 (n1023, n691, n938, n981, n934);
and  g978 (n1018, n744, n815, n681, n814);
xnor g979 (n1054, n651, n977, n838, n983);
or   g980 (n1005, n741, n937, n846, n702);
nor  g981 (n1011, n813, n990, n842, n978);
or   g982 (n992, n935, n654, n855, n976);
and  g983 (n1035, n397, n985, n662, n841);
and  g984 (n1028, n655, n987, n849, n978);
nor  g985 (n1048, n658, n656, n732, n843);
nand g986 (n1027, n986, n815, n975, n671);
and  g987 (n1000, n712, n984, n728, n689);
nand g988 (n1030, n736, n980, n636, n988);
or   g989 (n1047, n659, n660, n981, n976);
xnor g990 (n1036, n982, n944, n813, n977);
nand g991 (n1031, n679, n813, n853, n990);
xnor g992 (n1024, n943, n632, n694, n980);
xnor g993 (n994, n937, n717, n680, n747);
nand g994 (n999, n750, n701, n734, n722);
or   g995 (n1034, n715, n976, n941, n668);
xor  g996 (n1044, n936, n988, n721, n985);
nor  g997 (n1039, n638, n735, n719, n738);
nand g998 (n1051, n985, n707, n645, n814);
and  g999 (n1012, n988, n685, n979, n672);
xor  g1000 (n1052, n975, n398, n649);
nand g1001 (n1014, n637, n983, n844, n988);
nand g1002 (n995, n980, n731, n982, n700);
xor  g1003 (n1025, n814, n852, n644, n714);
or   g1004 (n1032, n989, n639, n837, n749);
nor  g1005 (n1010, n979, n980, n984, n812);
nand g1006 (n1017, n858, n946, n641, n720);
or   g1007 (n1019, n941, n942, n705, n981);
and  g1008 (n1045, n938, n746, n989, n990);
or   g1009 (n1021, n984, n836, n982, n675);
nor  g1010 (n1049, n987, n860, n989, n737);
and  g1011 (n1002, n730, n667, n983, n703);
xnor g1012 (n997, n665, n944, n742, n642);
and  g1013 (n1038, n945, n985, n723, n740);
xor  g1014 (n993, n936, n946, n633, n945);
or   g1015 (n1029, n690, n942, n978, n848);
nor  g1016 (n1037, n673, n854, n724, n981);
nand g1017 (n1003, n711, n934, n856, n634);
xnor g1018 (n1013, n696, n726, n814, n713);
or   g1019 (n1033, n975, n682, n397, n987);
xnor g1020 (n1041, n725, n743, n990, n933);
xor  g1021 (n1040, n940, n745, n739, n706);
or   g1022 (n996, n678, n815, n845, n733);
nor  g1023 (n1020, n704, n687, n670, n748);
and  g1024 (n1016, n813, n664, n943, n709);
xor  g1025 (n1009, n699, n940, n986, n663);
xnor g1026 (n1053, n946, n643, n987, n653);
xor  g1027 (n1046, n939, n647, n859, n979);
and  g1028 (n1007, n635, n976, n984, n982);
nand g1029 (n991, n657, n716, n729, n727);
or   g1030 (n1043, n708, n650, n695, n975);
nor  g1031 (n1015, n718, n839, n935, n847);
xor  g1032 (n1004, n677, n676, n693, n850);
xor  g1033 (n1001, n857, n674, n652, n692);
and  g1034 (n1042, n840, n640, n977, n945);
xor  g1035 (n1058, n1023, n948, n1008, n1028);
nor  g1036 (n1060, n1038, n1053, n999, n1045);
nor  g1037 (n1057, n1009, n947, n1043, n1046);
and  g1038 (n1070, n992, n1037, n951, n952);
and  g1039 (n1073, n1001, n1027, n1050, n1051);
nor  g1040 (n1066, n1035, n947, n998, n948);
xnor g1041 (n1076, n1014, n1021, n1026, n1025);
xor  g1042 (n1065, n1042, n949, n1017, n1034);
xor  g1043 (n1072, n948, n950, n1012);
nor  g1044 (n1067, n1039, n398, n952, n1004);
or   g1045 (n1055, n1054, n949, n1030, n996);
nand g1046 (n1064, n952, n949, n953, n1011);
xor  g1047 (n1063, n880, n1016, n1013, n1019);
xnor g1048 (n1075, n1036, n1010, n1040, n947);
nor  g1049 (n1061, n1031, n1033, n1006, n1000);
or   g1050 (n1059, n953, n880, n994, n1015);
or   g1051 (n1068, n1022, n1032, n1020, n995);
or   g1052 (n1074, n1049, n1005, n1041, n1024);
nand g1053 (n1071, n1029, n1048, n953, n1018);
and  g1054 (n1069, n1047, n993, n1044, n1002);
xor  g1055 (n1062, n950, n951, n997);
nand g1056 (n1056, n1003, n1052, n1007, n991);
endmodule
