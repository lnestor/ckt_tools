

module Stat_183_517
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n122,
  n171,
  n124,
  n178,
  n160,
  n125,
  n165,
  n177,
  n130,
  n208,
  n204,
  n192,
  n199,
  n203,
  n205,
  n198,
  n200,
  n197,
  n201,
  n195,
  n196,
  n209,
  n194,
  n207,
  n206,
  n202,
  n193,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;
  output n122;output n171;output n124;output n178;output n160;output n125;output n165;output n177;output n130;output n208;output n204;output n192;output n199;output n203;output n205;output n198;output n200;output n197;output n201;output n195;output n196;output n209;output n194;output n207;output n206;output n202;output n193;
  wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n123;wire n126;wire n127;wire n128;wire n129;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n161;wire n162;wire n163;wire n164;wire n166;wire n167;wire n168;wire n169;wire n170;wire n172;wire n173;wire n174;wire n175;wire n176;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n54,
    n8
  );


  not
  g1
  (
    n61,
    n23
  );


  not
  g2
  (
    n64,
    n10
  );


  buf
  g3
  (
    n72,
    n1
  );


  buf
  g4
  (
    n28,
    n17
  );


  not
  g5
  (
    n73,
    n9
  );


  not
  g6
  (
    n80,
    n14
  );


  not
  g7
  (
    n91,
    n8
  );


  buf
  g8
  (
    n77,
    n4
  );


  buf
  g9
  (
    n79,
    n19
  );


  buf
  g10
  (
    n56,
    n10
  );


  not
  g11
  (
    n57,
    n11
  );


  buf
  g12
  (
    n47,
    n19
  );


  not
  g13
  (
    n50,
    n7
  );


  not
  g14
  (
    n37,
    n5
  );


  buf
  g15
  (
    n90,
    n20
  );


  not
  g16
  (
    n41,
    n4
  );


  not
  g17
  (
    n97,
    n23
  );


  not
  g18
  (
    n55,
    n7
  );


  not
  g19
  (
    n86,
    n12
  );


  not
  g20
  (
    n30,
    n3
  );


  buf
  g21
  (
    n84,
    n1
  );


  not
  g22
  (
    n70,
    n9
  );


  not
  g23
  (
    n78,
    n20
  );


  buf
  g24
  (
    n66,
    n13
  );


  not
  g25
  (
    n69,
    n14
  );


  not
  g26
  (
    n71,
    n22
  );


  buf
  g27
  (
    n32,
    n24
  );


  not
  g28
  (
    n58,
    n6
  );


  buf
  g29
  (
    n53,
    n20
  );


  not
  g30
  (
    n42,
    n2
  );


  buf
  g31
  (
    n76,
    n11
  );


  buf
  g32
  (
    n49,
    n3
  );


  buf
  g33
  (
    n83,
    n16
  );


  not
  g34
  (
    n92,
    n17
  );


  not
  g35
  (
    n40,
    n22
  );


  not
  g36
  (
    n38,
    n11
  );


  buf
  g37
  (
    n59,
    n6
  );


  buf
  g38
  (
    n33,
    n2
  );


  buf
  g39
  (
    n63,
    n5
  );


  not
  g40
  (
    n62,
    n8
  );


  not
  g41
  (
    n36,
    n14
  );


  buf
  g42
  (
    n96,
    n15
  );


  buf
  g43
  (
    n87,
    n21
  );


  not
  g44
  (
    n39,
    n1
  );


  not
  g45
  (
    n29,
    n6
  );


  not
  g46
  (
    n68,
    n5
  );


  not
  g47
  (
    n27,
    n13
  );


  not
  g48
  (
    n44,
    n13
  );


  buf
  g49
  (
    n74,
    n18
  );


  buf
  g50
  (
    n88,
    n10
  );


  buf
  g51
  (
    n34,
    n7
  );


  buf
  g52
  (
    n45,
    n3
  );


  buf
  g53
  (
    n43,
    n4
  );


  buf
  g54
  (
    n60,
    n9
  );


  not
  g55
  (
    n51,
    n18
  );


  not
  g56
  (
    n35,
    n15
  );


  buf
  g57
  (
    n48,
    n17
  );


  buf
  g58
  (
    n52,
    n16
  );


  not
  g59
  (
    n67,
    n23
  );


  buf
  g60
  (
    n75,
    n16
  );


  buf
  g61
  (
    n95,
    n18
  );


  buf
  g62
  (
    n89,
    n15
  );


  buf
  g63
  (
    n82,
    n12
  );


  not
  g64
  (
    n98,
    n21
  );


  buf
  g65
  (
    n81,
    n12
  );


  buf
  g66
  (
    n31,
    n24
  );


  buf
  g67
  (
    n46,
    n2
  );


  not
  g68
  (
    n65,
    n22
  );


  not
  g69
  (
    n94,
    n21
  );


  not
  g70
  (
    n93,
    n24
  );


  buf
  g71
  (
    n85,
    n19
  );


  not
  g72
  (
    n109,
    n30
  );


  not
  g73
  (
    n110,
    n29
  );


  not
  g74
  (
    n111,
    n33
  );


  buf
  g75
  (
    n106,
    n34
  );


  buf
  g76
  (
    n115,
    n31
  );


  not
  g77
  (
    n118,
    n26
  );


  not
  g78
  (
    n108,
    n28
  );


  buf
  g79
  (
    n119,
    n27
  );


  not
  g80
  (
    n114,
    n25
  );


  not
  g81
  (
    n107,
    n30
  );


  not
  g82
  (
    n99,
    n26
  );


  buf
  g83
  (
    n105,
    n26
  );


  buf
  g84
  (
    n102,
    n29
  );


  buf
  g85
  (
    n120,
    n25
  );


  buf
  g86
  (
    n100,
    n31
  );


  not
  g87
  (
    n104,
    n32
  );


  buf
  g88
  (
    n101,
    n27
  );


  buf
  g89
  (
    n117,
    n31
  );


  buf
  g90
  (
    n103,
    n33
  );


  buf
  g91
  (
    n112,
    n32
  );


  xnor
  g92
  (
    n116,
    n30,
    n27,
    n32,
    n28
  );


  nor
  g93
  (
    n113,
    n33,
    n28,
    n25,
    n29
  );


  and
  g94
  (
    n128,
    n49,
    n116,
    n95
  );


  or
  g95
  (
    n142,
    n42,
    n94,
    n113,
    n107
  );


  or
  g96
  (
    n160,
    n51,
    n69,
    n100,
    n60
  );


  or
  g97
  (
    n138,
    n83,
    n60,
    n79,
    n42
  );


  xnor
  g98
  (
    n149,
    n61,
    n66,
    n79,
    n56
  );


  nor
  g99
  (
    n147,
    n79,
    n94,
    n103,
    n73
  );


  and
  g100
  (
    n151,
    n82,
    n86,
    n109,
    n93
  );


  nor
  g101
  (
    n137,
    n50,
    n72,
    n41,
    n45
  );


  xor
  g102
  (
    n124,
    n51,
    n55,
    n57,
    n117
  );


  nand
  g103
  (
    n179,
    n104,
    n108,
    n77,
    n41
  );


  nand
  g104
  (
    n126,
    n72,
    n54,
    n53,
    n47
  );


  nor
  g105
  (
    n184,
    n43,
    n48,
    n40,
    n117
  );


  and
  g106
  (
    n182,
    n62,
    n80,
    n53,
    n82
  );


  xnor
  g107
  (
    n158,
    n113,
    n85,
    n64,
    n115
  );


  xor
  g108
  (
    n125,
    n36,
    n72,
    n78,
    n89
  );


  or
  g109
  (
    n134,
    n81,
    n82,
    n69,
    n84
  );


  xor
  g110
  (
    n172,
    n46,
    n114,
    n115,
    n108
  );


  or
  g111
  (
    n122,
    n77,
    n68,
    n80,
    n78
  );


  and
  g112
  (
    n139,
    n50,
    n43,
    n99,
    n68
  );


  and
  g113
  (
    n157,
    n93,
    n110,
    n100,
    n92
  );


  nand
  g114
  (
    n135,
    n87,
    n88,
    n71,
    n99
  );


  or
  g115
  (
    n156,
    n86,
    n111,
    n87,
    n73
  );


  and
  g116
  (
    AntiSAT_key_wire,
    n96,
    n76,
    n36,
    n52
  );


  nor
  g117
  (
    n171,
    n100,
    n38,
    n92,
    n34
  );


  xor
  g118
  (
    n153,
    n112,
    n93,
    n47,
    n89
  );


  or
  g119
  (
    n175,
    n103,
    n58,
    n88,
    n85
  );


  xnor
  g120
  (
    n166,
    n112,
    n96,
    n75,
    n99
  );


  or
  g121
  (
    n162,
    n83,
    n49,
    n67,
    n35
  );


  xnor
  g122
  (
    n155,
    n101,
    n84,
    n60,
    n61
  );


  or
  g123
  (
    n145,
    n103,
    n53,
    n106,
    n49
  );


  nand
  g124
  (
    n130,
    n59,
    n54,
    n62,
    n104
  );


  nand
  g125
  (
    n144,
    n106,
    n107,
    n105,
    n114
  );


  nor
  g126
  (
    n133,
    n78,
    n120,
    n70,
    n59
  );


  xnor
  g127
  (
    n127,
    n68,
    n57,
    n46,
    n64
  );


  xnor
  g128
  (
    n165,
    n35,
    n67,
    n76,
    n91
  );


  nor
  g129
  (
    n164,
    n111,
    n39,
    n63,
    n44
  );


  xor
  g130
  (
    n123,
    n112,
    n88,
    n44,
    n38
  );


  and
  g131
  (
    n152,
    n81,
    n71,
    n111,
    n65
  );


  nor
  g132
  (
    n163,
    n74,
    n66,
    n118,
    n51
  );


  xor
  g133
  (
    n169,
    n90,
    n90,
    n39,
    n84
  );


  nor
  g134
  (
    n143,
    n59,
    n104,
    n118,
    n63
  );


  nor
  g135
  (
    n140,
    n108,
    n62,
    n113,
    n52
  );


  xnor
  g136
  (
    n183,
    n97,
    n87,
    n55,
    n98
  );


  nor
  g137
  (
    n180,
    n58,
    n63,
    n119,
    n55
  );


  nand
  g138
  (
    n129,
    n44,
    n95,
    n98,
    n97
  );


  xor
  g139
  (
    n141,
    n102,
    n75,
    n71,
    n45
  );


  nand
  g140
  (
    n181,
    n74,
    n80,
    n118,
    n101
  );


  xor
  g141
  (
    n168,
    n102,
    n95,
    n61,
    n40
  );


  or
  g142
  (
    n121,
    n36,
    n57,
    n109,
    n120
  );


  xnor
  g143
  (
    n185,
    n90,
    n86,
    n47,
    n117
  );


  nor
  g144
  (
    n136,
    n83,
    n56,
    n75,
    n98
  );


  xnor
  g145
  (
    n131,
    n119,
    n74,
    n39,
    n69
  );


  xor
  g146
  (
    n177,
    n64,
    n35,
    n38,
    n34
  );


  xor
  g147
  (
    n148,
    n107,
    n102,
    n37,
    n65
  );


  and
  g148
  (
    n176,
    n54,
    n94,
    n45,
    n89
  );


  xor
  g149
  (
    n173,
    n48,
    n110,
    n81
  );


  or
  g150
  (
    n170,
    n76,
    n97,
    n92,
    n109
  );


  or
  g151
  (
    n146,
    n91,
    n105,
    n66,
    n40
  );


  and
  g152
  (
    n174,
    n46,
    n37,
    n65,
    n77
  );


  nand
  g153
  (
    n159,
    n67,
    n50,
    n115,
    n91
  );


  and
  g154
  (
    n132,
    n114,
    n73,
    n116,
    n96
  );


  or
  g155
  (
    n154,
    n58,
    n42,
    n119,
    n56
  );


  or
  g156
  (
    n161,
    n101,
    n37,
    n70,
    n106
  );


  nand
  g157
  (
    n150,
    n85,
    n105,
    n48,
    n52
  );


  nand
  g158
  (
    n167,
    n41,
    n116,
    n70,
    n43
  );


  buf
  g159
  (
    n191,
    n131
  );


  buf
  g160
  (
    n186,
    n132
  );


  buf
  g161
  (
    n190,
    n120
  );


  not
  g162
  (
    n189,
    n134
  );


  buf
  g163
  (
    n188,
    n133
  );


  or
  g164
  (
    n187,
    n135,
    n130
  );


  nor
  g165
  (
    n206,
    n139,
    n164,
    n150,
    n191
  );


  nand
  g166
  (
    n208,
    n190,
    n143,
    n159,
    n191
  );


  xor
  g167
  (
    n195,
    n187,
    n187,
    n144,
    n178
  );


  xor
  g168
  (
    n200,
    n176,
    n188,
    n163,
    n160
  );


  or
  g169
  (
    n194,
    n165,
    n138,
    n167,
    n181
  );


  xnor
  g170
  (
    n198,
    n166,
    n189,
    n171,
    n186
  );


  nor
  g171
  (
    n207,
    n172,
    n157,
    n151,
    n174
  );


  or
  g172
  (
    n209,
    n190,
    n191,
    n185,
    n155
  );


  nor
  g173
  (
    n205,
    n187,
    n145,
    n190,
    n149
  );


  or
  g174
  (
    n201,
    n189,
    n185,
    n175,
    n156
  );


  xor
  g175
  (
    n202,
    n148,
    n184,
    n146
  );


  or
  g176
  (
    n203,
    n140,
    n185,
    n162,
    n137
  );


  nand
  g177
  (
    n197,
    n184,
    n189,
    n186,
    n153
  );


  nor
  g178
  (
    n192,
    n173,
    n169,
    n186,
    n161
  );


  xor
  g179
  (
    n196,
    n188,
    n136,
    n147,
    n177
  );


  xor
  g180
  (
    n204,
    n179,
    n142,
    n141,
    n154
  );


  or
  g181
  (
    n199,
    n158,
    n182,
    n170,
    n152
  );


  nor
  g182
  (
    n193,
    n168,
    n188,
    n183,
    n180
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_0,
    keyIn_0_26,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_1,
    keyIn_0_27,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_2,
    keyIn_0_28,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_3,
    keyIn_0_29,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_4,
    keyIn_0_30,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_5,
    keyIn_0_31,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_6,
    keyIn_0_32,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_7,
    keyIn_0_33,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_8,
    keyIn_0_34,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_9,
    keyIn_0_35,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_10,
    keyIn_0_36,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_11,
    keyIn_0_37,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_12,
    keyIn_0_38,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_13,
    keyIn_0_39,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_14,
    keyIn_0_40,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_15,
    keyIn_0_41,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_16,
    keyIn_0_42,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_17,
    keyIn_0_43,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_18,
    keyIn_0_44,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_19,
    keyIn_0_45,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_20,
    keyIn_0_46,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_21,
    keyIn_0_47,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_22,
    keyIn_0_48,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_23,
    keyIn_0_49,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_24,
    keyIn_0_50,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_25,
    keyIn_0_51,
    n26
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n178,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

