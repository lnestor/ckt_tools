// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_311 written by SynthGen on 2021/04/05 11:23:41
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_311 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n892, n886, n877, n890, n870, n880, n872, n884,
 n871, n883, n881, n869, n891, n873, n887, n882,
 n866, n1953, n2028, n2023, n2022, n2020, n2027, n2031,
 n2029, n2025, n2030, n2021, n2019, n2026, n2032, n2024);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n892, n886, n877, n890, n870, n880, n872, n884,
 n871, n883, n881, n869, n891, n873, n887, n882,
 n866, n1953, n2028, n2023, n2022, n2020, n2027, n2031,
 n2029, n2025, n2030, n2021, n2019, n2026, n2032, n2024;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n867, n868, n874, n875, n876, n878, n879,
 n885, n888, n889, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
 n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
 n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
 n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
 n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
 n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
 n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
 n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
 n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
 n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
 n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
 n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
 n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
 n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
 n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
 n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
 n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
 n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
 n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
 n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
 n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
 n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
 n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
 n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
 n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
 n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
 n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
 n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
 n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
 n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
 n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
 n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
 n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
 n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
 n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
 n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
 n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
 n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
 n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
 n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
 n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
 n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
 n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
 n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
 n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
 n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
 n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
 n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
 n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
 n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
 n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
 n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
 n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
 n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
 n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
 n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
 n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
 n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
 n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
 n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
 n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
 n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
 n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
 n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
 n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
 n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
 n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
 n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
 n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
 n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
 n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
 n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
 n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
 n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
 n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
 n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
 n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
 n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
 n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
 n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
 n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
 n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
 n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
 n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
 n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
 n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
 n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
 n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
 n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
 n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
 n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
 n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
 n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
 n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
 n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
 n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
 n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
 n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
 n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
 n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
 n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
 n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
 n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
 n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
 n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
 n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
 n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
 n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
 n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
 n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
 n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
 n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
 n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
 n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018;

buf  g0 (n61, n24);
buf  g1 (n52, n20);
buf  g2 (n143, n29);
not  g3 (n50, n18);
not  g4 (n56, n9);
buf  g5 (n126, n19);
not  g6 (n131, n29);
not  g7 (n39, n13);
buf  g8 (n93, n11);
buf  g9 (n70, n25);
not  g10 (n103, n31);
buf  g11 (n65, n12);
not  g12 (n62, n7);
not  g13 (n134, n27);
not  g14 (n66, n23);
buf  g15 (n35, n27);
not  g16 (n105, n7);
buf  g17 (n40, n18);
not  g18 (n112, n7);
buf  g19 (n140, n30);
buf  g20 (n33, n3);
not  g21 (n94, n1);
buf  g22 (n67, n22);
not  g23 (n37, n19);
buf  g24 (n92, n20);
not  g25 (n108, n30);
not  g26 (n144, n13);
not  g27 (n88, n16);
not  g28 (n129, n3);
not  g29 (n46, n15);
buf  g30 (n136, n25);
buf  g31 (n47, n6);
buf  g32 (n45, n12);
not  g33 (n49, n7);
buf  g34 (n118, n9);
buf  g35 (n121, n29);
not  g36 (n34, n28);
not  g37 (n78, n13);
not  g38 (n132, n13);
buf  g39 (n122, n28);
not  g40 (n135, n26);
buf  g41 (n97, n23);
buf  g42 (n74, n8);
buf  g43 (n128, n26);
not  g44 (n130, n4);
buf  g45 (n58, n1);
buf  g46 (n107, n17);
buf  g47 (n53, n14);
buf  g48 (n63, n17);
buf  g49 (n96, n6);
buf  g50 (n42, n21);
not  g51 (n113, n8);
buf  g52 (n119, n15);
not  g53 (n44, n29);
not  g54 (n87, n11);
buf  g55 (n84, n5);
not  g56 (n55, n3);
not  g57 (n137, n5);
not  g58 (n139, n9);
buf  g59 (n141, n27);
not  g60 (n138, n23);
buf  g61 (n100, n8);
buf  g62 (n101, n14);
not  g63 (n69, n2);
not  g64 (n77, n26);
not  g65 (n115, n24);
not  g66 (n83, n20);
not  g67 (n89, n18);
buf  g68 (n81, n1);
buf  g69 (n124, n16);
buf  g70 (n57, n24);
not  g71 (n82, n22);
not  g72 (n111, n26);
not  g73 (n99, n2);
not  g74 (n106, n12);
buf  g75 (n114, n4);
not  g76 (n117, n9);
buf  g77 (n68, n23);
buf  g78 (n120, n10);
not  g79 (n38, n14);
not  g80 (n133, n16);
not  g81 (n95, n19);
buf  g82 (n125, n18);
not  g83 (n147, n25);
not  g84 (n64, n10);
buf  g85 (n109, n28);
not  g86 (n54, n10);
buf  g87 (n60, n17);
buf  g88 (n91, n22);
buf  g89 (n80, n8);
buf  g90 (n59, n21);
not  g91 (n98, n4);
buf  g92 (n127, n5);
not  g93 (n110, n21);
buf  g94 (n48, n11);
not  g95 (n43, n21);
not  g96 (n145, n30);
buf  g97 (n142, n6);
not  g98 (n51, n22);
not  g99 (n72, n14);
not  g100 (n148, n30);
not  g101 (n79, n16);
not  g102 (n90, n6);
not  g103 (n123, n24);
buf  g104 (n86, n2);
not  g105 (n75, n28);
buf  g106 (n102, n17);
not  g107 (n73, n27);
not  g108 (n85, n12);
buf  g109 (n41, n15);
buf  g110 (n116, n11);
not  g111 (n76, n25);
buf  g112 (n104, n15);
not  g113 (n71, n19);
not  g114 (n146, n20);
buf  g115 (n36, n10);
not  g116 (n446, n98);
buf  g117 (n292, n48);
not  g118 (n387, n85);
not  g119 (n463, n35);
not  g120 (n383, n66);
buf  g121 (n343, n111);
not  g122 (n376, n48);
not  g123 (n169, n97);
buf  g124 (n166, n72);
not  g125 (n335, n88);
not  g126 (n431, n49);
buf  g127 (n175, n36);
not  g128 (n185, n44);
not  g129 (n274, n49);
not  g130 (n237, n91);
buf  g131 (n219, n113);
buf  g132 (n440, n42);
not  g133 (n295, n68);
not  g134 (n331, n92);
buf  g135 (n277, n54);
not  g136 (n281, n87);
not  g137 (n485, n114);
buf  g138 (n260, n94);
not  g139 (n241, n73);
buf  g140 (n452, n37);
not  g141 (n242, n79);
not  g142 (n300, n92);
buf  g143 (n430, n52);
buf  g144 (n276, n87);
buf  g145 (n438, n89);
buf  g146 (n416, n101);
not  g147 (n244, n45);
not  g148 (n384, n101);
buf  g149 (n428, n104);
not  g150 (n195, n69);
buf  g151 (n330, n82);
buf  g152 (n378, n86);
not  g153 (n153, n68);
buf  g154 (n163, n58);
buf  g155 (n196, n65);
not  g156 (n471, n112);
not  g157 (n298, n60);
buf  g158 (n389, n74);
not  g159 (n417, n112);
not  g160 (n272, n41);
not  g161 (n412, n68);
buf  g162 (n315, n104);
not  g163 (n204, n50);
buf  g164 (n225, n116);
buf  g165 (n290, n117);
buf  g166 (n210, n84);
buf  g167 (n309, n100);
not  g168 (n443, n90);
not  g169 (n406, n63);
not  g170 (n371, n72);
not  g171 (n402, n77);
buf  g172 (n350, n114);
buf  g173 (n296, n77);
buf  g174 (n477, n44);
buf  g175 (n271, n85);
buf  g176 (n338, n108);
buf  g177 (n181, n65);
buf  g178 (n340, n89);
buf  g179 (n474, n115);
buf  g180 (n313, n71);
not  g181 (n191, n37);
buf  g182 (n388, n50);
buf  g183 (n461, n68);
buf  g184 (n421, n93);
not  g185 (n304, n38);
not  g186 (n324, n106);
buf  g187 (n186, n70);
buf  g188 (n256, n73);
not  g189 (n162, n66);
buf  g190 (n483, n106);
not  g191 (n265, n88);
buf  g192 (n280, n89);
not  g193 (n258, n33);
not  g194 (n359, n70);
not  g195 (n426, n115);
buf  g196 (n355, n110);
buf  g197 (n167, n52);
buf  g198 (n165, n39);
buf  g199 (n467, n64);
buf  g200 (n328, n83);
not  g201 (n423, n56);
not  g202 (n158, n77);
not  g203 (n351, n71);
not  g204 (n202, n56);
buf  g205 (n332, n51);
buf  g206 (n220, n74);
not  g207 (n170, n66);
not  g208 (n369, n95);
not  g209 (n187, n111);
not  g210 (n222, n85);
buf  g211 (n236, n38);
not  g212 (n311, n35);
not  g213 (n490, n98);
not  g214 (n229, n57);
not  g215 (n278, n102);
not  g216 (n156, n104);
buf  g217 (n245, n81);
buf  g218 (n396, n49);
not  g219 (n329, n62);
not  g220 (n414, n97);
not  g221 (n447, n95);
buf  g222 (n385, n106);
buf  g223 (n390, n90);
not  g224 (n294, n54);
not  g225 (n234, n62);
buf  g226 (n442, n96);
not  g227 (n363, n34);
not  g228 (n424, n67);
not  g229 (n221, n33);
not  g230 (n445, n39);
buf  g231 (n218, n61);
not  g232 (n200, n62);
not  g233 (n183, n72);
not  g234 (n392, n69);
not  g235 (n365, n80);
not  g236 (n456, n100);
buf  g237 (n382, n105);
buf  g238 (n320, n39);
not  g239 (n429, n38);
buf  g240 (n246, n64);
not  g241 (n238, n115);
not  g242 (n268, n60);
not  g243 (n286, n54);
not  g244 (n302, n113);
not  g245 (n386, n34);
buf  g246 (n336, n116);
not  g247 (n345, n112);
not  g248 (n160, n47);
not  g249 (n251, n63);
not  g250 (n151, n41);
buf  g251 (n189, n53);
buf  g252 (n168, n55);
not  g253 (n287, n61);
not  g254 (n283, n61);
not  g255 (n341, n73);
buf  g256 (n269, n35);
not  g257 (n481, n41);
buf  g258 (n157, n72);
buf  g259 (n472, n39);
not  g260 (n205, n99);
buf  g261 (n449, n116);
buf  g262 (n319, n107);
not  g263 (n325, n60);
not  g264 (n337, n90);
buf  g265 (n487, n61);
not  g266 (n259, n69);
not  g267 (n391, n75);
not  g268 (n398, n55);
not  g269 (n179, n103);
not  g270 (n413, n76);
buf  g271 (n275, n94);
not  g272 (n357, n96);
not  g273 (n354, n52);
not  g274 (n239, n76);
not  g275 (n451, n65);
not  g276 (n240, n59);
buf  g277 (n203, n44);
buf  g278 (n489, n46);
not  g279 (n444, n97);
not  g280 (n448, n40);
not  g281 (n310, n55);
not  g282 (n347, n107);
not  g283 (n194, n101);
not  g284 (n235, n93);
not  g285 (n326, n63);
buf  g286 (n373, n94);
buf  g287 (n411, n91);
buf  g288 (n314, n73);
not  g289 (n291, n64);
not  g290 (n334, n104);
buf  g291 (n395, n64);
not  g292 (n257, n99);
buf  g293 (n217, n46);
buf  g294 (n261, n52);
buf  g295 (n409, n118);
not  g296 (n255, n98);
buf  g297 (n422, n110);
not  g298 (n484, n91);
buf  g299 (n214, n37);
not  g300 (n273, n92);
not  g301 (n228, n83);
not  g302 (n152, n109);
buf  g303 (n394, n38);
not  g304 (n420, n96);
not  g305 (n410, n51);
not  g306 (n178, n99);
not  g307 (n397, n80);
not  g308 (n342, n54);
buf  g309 (n208, n53);
not  g310 (n233, n117);
buf  g311 (n486, n76);
not  g312 (n379, n93);
buf  g313 (n209, n114);
buf  g314 (n358, n78);
buf  g315 (n321, n111);
buf  g316 (n375, n33);
buf  g317 (n457, n50);
not  g318 (n348, n71);
buf  g319 (n279, n60);
not  g320 (n333, n92);
not  g321 (n466, n70);
not  g322 (n403, n67);
buf  g323 (n212, n108);
buf  g324 (n380, n95);
not  g325 (n254, n46);
buf  g326 (n437, n43);
buf  g327 (n289, n35);
buf  g328 (n312, n70);
buf  g329 (n188, n99);
buf  g330 (n197, n115);
buf  g331 (n364, n100);
buf  g332 (n404, n67);
buf  g333 (n308, n106);
buf  g334 (n473, n59);
not  g335 (n339, n102);
buf  g336 (n370, n65);
buf  g337 (n253, n78);
buf  g338 (n267, n34);
buf  g339 (n482, n109);
buf  g340 (n478, n77);
buf  g341 (n182, n48);
buf  g342 (n177, n57);
not  g343 (n206, n86);
not  g344 (n207, n113);
not  g345 (n401, n82);
buf  g346 (n159, n84);
buf  g347 (n353, n66);
buf  g348 (n262, n43);
buf  g349 (n465, n105);
not  g350 (n322, n78);
buf  g351 (n476, n59);
buf  g352 (n367, n83);
buf  g353 (n434, n85);
buf  g354 (n211, n102);
not  g355 (n480, n103);
not  g356 (n264, n105);
not  g357 (n180, n78);
buf  g358 (n366, n58);
not  g359 (n469, n80);
not  g360 (n393, n40);
buf  g361 (n432, n86);
not  g362 (n154, n76);
not  g363 (n293, n91);
buf  g364 (n149, n107);
not  g365 (n226, n113);
not  g366 (n468, n88);
not  g367 (n305, n87);
buf  g368 (n352, n79);
buf  g369 (n303, n58);
not  g370 (n318, n59);
not  g371 (n462, n40);
not  g372 (n356, n43);
buf  g373 (n323, n51);
not  g374 (n361, n41);
not  g375 (n231, n40);
not  g376 (n427, n67);
not  g377 (n285, n56);
buf  g378 (n435, n44);
not  g379 (n150, n58);
buf  g380 (n266, n82);
not  g381 (n458, n79);
not  g382 (n450, n57);
buf  g383 (n176, n80);
not  g384 (n299, n101);
buf  g385 (n232, n88);
buf  g386 (n263, n87);
buf  g387 (n199, n57);
buf  g388 (n174, n75);
buf  g389 (n190, n84);
buf  g390 (n297, n74);
buf  g391 (n164, n84);
not  g392 (n243, n69);
buf  g393 (n455, n42);
buf  g394 (n368, n33);
not  g395 (n247, n117);
buf  g396 (n439, n111);
buf  g397 (n216, n48);
not  g398 (n327, n45);
not  g399 (n193, n96);
not  g400 (n400, n110);
buf  g401 (n184, n36);
buf  g402 (n415, n83);
buf  g403 (n374, n117);
not  g404 (n282, n36);
buf  g405 (n192, n98);
buf  g406 (n418, n79);
not  g407 (n230, n51);
buf  g408 (n201, n108);
buf  g409 (n213, n36);
buf  g410 (n307, n100);
not  g411 (n464, n102);
buf  g412 (n407, n103);
buf  g413 (n284, n93);
buf  g414 (n316, n97);
buf  g415 (n408, n45);
not  g416 (n173, n55);
buf  g417 (n249, n81);
not  g418 (n362, n47);
not  g419 (n215, n43);
buf  g420 (n224, n49);
not  g421 (n317, n90);
not  g422 (n453, n103);
not  g423 (n475, n86);
not  g424 (n288, n109);
buf  g425 (n433, n89);
not  g426 (n372, n114);
not  g427 (n399, n105);
buf  g428 (n155, n74);
not  g429 (n425, n53);
buf  g430 (n470, n116);
buf  g431 (n248, n63);
buf  g432 (n360, n81);
buf  g433 (n301, n118);
not  g434 (n223, n108);
buf  g435 (n381, n62);
not  g436 (n488, n95);
not  g437 (n171, n109);
not  g438 (n270, n45);
not  g439 (n227, n46);
not  g440 (n454, n110);
buf  g441 (n349, n42);
not  g442 (n436, n50);
buf  g443 (n479, n81);
not  g444 (n198, n42);
buf  g445 (n344, n37);
buf  g446 (n419, n71);
not  g447 (n306, n75);
not  g448 (n161, n47);
buf  g449 (n252, n56);
not  g450 (n346, n107);
not  g451 (n441, n112);
not  g452 (n405, n94);
not  g453 (n172, n47);
not  g454 (n460, n53);
buf  g455 (n459, n34);
not  g456 (n377, n82);
not  g457 (n250, n75);
buf  g458 (n733, n289);
buf  g459 (n575, n410);
not  g460 (n594, n402);
not  g461 (n516, n463);
not  g462 (n623, n207);
buf  g463 (n504, n231);
buf  g464 (n546, n279);
not  g465 (n551, n309);
not  g466 (n672, n130);
buf  g467 (n579, n165);
not  g468 (n835, n418);
not  g469 (n804, n328);
buf  g470 (n653, n194);
not  g471 (n659, n402);
nor  g472 (n669, n176, n126, n311);
nand g473 (n513, n128, n405, n457, n390);
or   g474 (n693, n227, n296, n418, n123);
xnor g475 (n825, n392, n378, n454, n443);
nand g476 (n592, n365, n374, n123, n342);
xnor g477 (n599, n379, n347, n415, n307);
nor  g478 (n701, n431, n399, n345, n448);
and  g479 (n529, n364, n263, n273, n217);
or   g480 (n823, n250, n423, n449, n317);
xor  g481 (n614, n243, n185, n222);
nand g482 (n637, n354, n280, n306, n409);
nand g483 (n617, n191, n142, n366, n160);
and  g484 (n729, n437, n351, n320, n173);
nand g485 (n814, n184, n292, n275, n437);
and  g486 (n709, n319, n410, n364, n421);
nor  g487 (n522, n295, n137, n315, n455);
nand g488 (n569, n250, n188, n285, n284);
xnor g489 (n827, n150, n243, n184, n219);
xnor g490 (n536, n357, n324, n318, n287);
and  g491 (n773, n211, n189, n456, n438);
and  g492 (n567, n333, n215, n442, n163);
and  g493 (n717, n369, n178, n459, n157);
or   g494 (n721, n162, n372, n390, n376);
xor  g495 (n616, n240, n340, n439, n453);
and  g496 (n683, n275, n191, n452, n264);
nor  g497 (n707, n127, n328, n318, n383);
xor  g498 (n784, n119, n337, n359, n238);
and  g499 (n615, n135, n385, n198, n159);
and  g500 (n754, n237, n237, n138, n290);
nor  g501 (n788, n360, n128, n219, n427);
nor  g502 (n743, n197, n327, n408, n236);
and  g503 (n571, n284, n204, n308, n235);
nor  g504 (n620, n258, n198, n323, n281);
and  g505 (n787, n310, n371, n386, n425);
nand g506 (n570, n454, n318, n333, n194);
nand g507 (n770, n374, n195, n142, n332);
xnor g508 (n526, n264, n316, n393, n372);
or   g509 (n532, n351, n141, n275, n211);
nand g510 (n728, n261, n225, n449, n424);
nand g511 (n818, n290, n234, n356, n179);
nand g512 (n587, n234, n282, n176);
xor  g513 (n657, n157, n184, n457, n188);
xor  g514 (n673, n170, n165, n127, n432);
or   g515 (n793, n314, n181, n174, n198);
nand g516 (n760, n441, n328, n370, n353);
and  g517 (n766, n229, n344, n345, n442);
nand g518 (n745, n216, n444, n355, n323);
and  g519 (n639, n316, n143, n420, n336);
nor  g520 (n635, n153, n119, n461, n267);
nand g521 (n552, n406, n457, n318, n411);
or   g522 (n736, n245, n426, n371, n374);
xnor g523 (n803, n317, n261, n395, n170);
nand g524 (n660, n288, n224, n451, n363);
xor  g525 (n514, n139, n397, n272, n136);
xor  g526 (n842, n426, n256, n189, n201);
and  g527 (n578, n460, n358, n298, n151);
nand g528 (n649, n302, n356, n369, n403);
nand g529 (n624, n422, n245, n300, n215);
xor  g530 (n663, n451, n316, n245, n186);
nor  g531 (n506, n408, n163, n140, n173);
xnor g532 (n491, n254, n269, n443, n382);
xnor g533 (n824, n214, n136, n352, n181);
or   g534 (n661, n226, n226, n258, n425);
and  g535 (n613, n298, n158, n341, n230);
xor  g536 (n518, n217, n393, n435, n200);
nor  g537 (n610, n387, n459, n211, n413);
nand g538 (n727, n240, n259, n249, n357);
xor  g539 (n688, n385, n369, n163, n306);
xor  g540 (n495, n187, n131, n448, n168);
nand g541 (n682, n444, n436, n311, n297);
or   g542 (n550, n461, n181, n367, n334);
nor  g543 (n791, n263, n128, n347, n305);
xnor g544 (n515, n429, n445, n122, n359);
xnor g545 (n609, n127, n283, n321, n217);
and  g546 (n805, n439, n438, n128, n252);
nor  g547 (n564, n186, n391, n201, n250);
and  g548 (n723, n334, n294, n420, n207);
nand g549 (n598, n149, n371, n377, n429);
and  g550 (n815, n382, n229, n396, n418);
and  g551 (n519, n327, n120, n313, n345);
and  g552 (n811, n400, n160, n152);
xnor g553 (n744, n405, n313, n400, n459);
xnor g554 (n801, n139, n459, n264, n460);
nand g555 (n679, n305, n338, n381, n375);
and  g556 (n535, n450, n405, n169, n232);
nand g557 (n528, n252, n143, n140, n441);
xnor g558 (n580, n219, n223, n398, n379);
and  g559 (n530, n417, n322, n131, n151);
or   g560 (n658, n337, n430, n413, n278);
and  g561 (n525, n319, n298, n237, n150);
xor  g562 (n700, n194, n289, n173, n221);
xor  g563 (n675, n291, n453, n266, n153);
xor  g564 (n554, n372, n121, n203, n355);
and  g565 (n618, n224, n260, n390, n174);
nand g566 (n666, n263, n363, n376, n321);
nand g567 (n588, n379, n156, n266, n376);
and  g568 (n605, n270, n416, n401, n463);
or   g569 (n668, n320, n299, n350, n272);
and  g570 (n544, n319, n416, n387, n126);
or   g571 (n769, n388, n346, n368, n389);
xnor g572 (n708, n248, n269, n320, n296);
or   g573 (n547, n229, n368, n389, n167);
xor  g574 (n549, n449, n347, n161, n215);
and  g575 (n589, n202, n361, n253, n404);
and  g576 (n566, n431, n291, n362, n283);
and  g577 (n630, n182, n154, n407, n163);
nand g578 (n507, n243, n296, n378, n452);
nand g579 (n795, n174, n299, n213, n232);
nor  g580 (n565, n196, n274, n187, n289);
xor  g581 (n493, n461, n204, n230, n450);
xnor g582 (n828, n150, n434, n346, n212);
nor  g583 (n636, n412, n134, n439, n301);
and  g584 (n541, n152, n206, n351, n155);
and  g585 (n762, n352, n120, n341, n382);
xnor g586 (n687, n303, n187, n140, n449);
xnor g587 (n799, n236, n388, n189, n363);
xor  g588 (n591, n122, n404, n217, n222);
or   g589 (n523, n252, n322, n422, n291);
or   g590 (n832, n370, n360, n129, n440);
nand g591 (n511, n279, n339, n314, n286);
nor  g592 (n557, n266, n435, n279, n228);
xnor g593 (n582, n402, n244, n255, n311);
nand g594 (n713, n280, n190, n357, n287);
and  g595 (n667, n407, n218, n221, n377);
and  g596 (n711, n268, n313, n336, n462);
and  g597 (n619, n342, n303, n204, n247);
nand g598 (n771, n141, n285, n200, n359);
xor  g599 (n735, n338, n192, n406, n314);
or   g600 (n689, n118, n423, n246, n260);
xor  g601 (n696, n229, n430, n325, n349);
and  g602 (n739, n200, n271, n144, n391);
xor  g603 (n524, n219, n171, n391, n142);
xor  g604 (n782, n189, n282, n187, n417);
xor  g605 (n819, n193, n237, n225, n197);
xnor g606 (n656, n133, n232, n284, n412);
xnor g607 (n662, n394, n253, n170, n368);
xnor g608 (n652, n243, n132, n302, n195);
nor  g609 (n645, n268, n227, n425, n166);
nand g610 (n840, n144, n415, n262, n276);
and  g611 (n545, n440, n438, n166, n124);
xnor g612 (n562, n337, n168, n336, n210);
or   g613 (n703, n339, n373, n392, n435);
nor  g614 (n521, n433, n335, n201, n209);
or   g615 (n698, n216, n423, n279, n383);
nor  g616 (n633, n350, n261, n445, n253);
and  g617 (n642, n155, n238, n314, n276);
nor  g618 (n671, n215, n218, n278, n349);
or   g619 (n500, n142, n188, n307, n248);
xor  g620 (n681, n131, n406, n185, n329);
nand g621 (n759, n292, n418, n207, n428);
nand g622 (n830, n285, n305, n458, n380);
xnor g623 (n699, n348, n190, n233, n331);
and  g624 (n563, n366, n358, n143, n132);
xnor g625 (n680, n119, n233, n230, n201);
xor  g626 (n691, n133, n289, n386, n188);
and  g627 (n765, n427, n293, n316, n436);
xnor g628 (n593, n393, n387, n450, n180);
and  g629 (n806, n137, n294, n267, n446);
nand g630 (n737, n307, n420, n228, n421);
nand g631 (n749, n424, n456, n249, n395);
xnor g632 (n585, n342, n238, n358, n183);
nor  g633 (n790, n356, n406, n265, n330);
xor  g634 (n738, n277, n247, n137, n203);
nor  g635 (n752, n234, n305, n399, n304);
or   g636 (n651, n259, n296, n138, n199);
xnor g637 (n779, n306, n145, n401, n235);
xnor g638 (n692, n422, n274, n239, n151);
xnor g639 (n503, n281, n361, n440, n400);
nand g640 (n785, n267, n455, n249, n248);
nand g641 (n542, n177, n274, n303, n162);
and  g642 (n494, n401, n149, n389, n276);
xnor g643 (n750, n231, n213, n355, n170);
and  g644 (n686, n343, n433, n425, n302);
xnor g645 (n628, n233, n417, n414, n180);
xor  g646 (n600, n335, n412, n210, n132);
or   g647 (n757, n384, n202, n339, n319);
nor  g648 (n724, n443, n178, n144, n411);
nor  g649 (n556, n227, n295, n446, n152);
nor  g650 (n577, n438, n277, n445, n169);
nand g651 (n809, n285, n356, n302, n138);
nand g652 (n626, n192, n136, n159, n221);
xnor g653 (n670, n360, n327, n220, n136);
xor  g654 (n751, n254, n365, n336, n157);
nor  g655 (n621, n323, n268, n368, n446);
and  g656 (n798, n190, n197, n378, n431);
nand g657 (n706, n282, n326, n392, n145);
and  g658 (n810, n442, n258, n447, n451);
nor  g659 (n820, n390, n123, n154, n360);
nor  g660 (n634, n294, n396, n301, n175);
nor  g661 (n789, n329, n309, n444, n455);
or   g662 (n539, n304, n265, n164, n172);
or   g663 (n627, n426, n135, n242, n140);
and  g664 (n641, n199, n165, n378, n206);
xor  g665 (n838, n286, n387, n416, n220);
nor  g666 (n796, n269, n408, n162, n153);
xnor g667 (n677, n317, n295, n236, n332);
and  g668 (n829, n263, n343, n240, n130);
xnor g669 (n761, n386, n315, n311, n177);
xnor g670 (n568, n164, n251, n185, n376);
or   g671 (n697, n396, n177, n432, n191);
nor  g672 (n548, n179, n431, n380, n423);
nand g673 (n501, n242, n195, n340, n450);
nor  g674 (n678, n238, n380, n293, n176);
nor  g675 (n802, n297, n435, n426, n456);
or   g676 (n543, n324, n172, n458, n270);
nand g677 (n538, n228, n404, n299, n150);
and  g678 (n684, n299, n278, n403, n375);
nor  g679 (n622, n358, n329, n132, n137);
nor  g680 (n775, n224, n326, n381, n421);
xnor g681 (n643, n239, n331, n246, n380);
and  g682 (n772, n462, n312, n382, n164);
and  g683 (n517, n166, n354, n208, n452);
or   g684 (n734, n300, n199, n192, n256);
xor  g685 (n647, n151, n121, n347, n286);
nor  g686 (n822, n171, n153, n265, n428);
nor  g687 (n755, n293, n182, n350, n255);
and  g688 (n590, n275, n271, n283, n396);
or   g689 (n774, n362, n144, n260, n127);
or   g690 (n581, n287, n309, n308, n220);
nor  g691 (n715, n301, n264, n257, n134);
nor  g692 (n797, n191, n421, n135, n366);
xor  g693 (n502, n444, n304, n303, n167);
and  g694 (n595, n411, n443, n227, n448);
nor  g695 (n586, n291, n436, n241, n442);
xnor g696 (n654, n205, n175, n255, n218);
xnor g697 (n740, n301, n209, n258, n414);
nor  g698 (n821, n293, n331, n326, n129);
xnor g699 (n718, n274, n413, n174, n180);
xor  g700 (n836, n175, n181, n462, n411);
and  g701 (n533, n412, n131, n461, n306);
nand g702 (n510, n246, n397, n434, n367);
and  g703 (n674, n122, n119, n143, n460);
nor  g704 (n492, n394, n139, n255, n428);
nor  g705 (n572, n185, n300, n216, n434);
xnor g706 (n531, n180, n308, n122, n254);
nor  g707 (n534, n231, n224, n353, n197);
xor  g708 (n690, n251, n310, n177, n343);
nor  g709 (n527, n451, n196, n292, n322);
nor  g710 (n640, n400, n226, n337, n329);
nor  g711 (n625, n300, n212, n354, n343);
xnor g712 (n509, n242, n398, n183, n440);
xor  g713 (n747, n424, n458, n355, n262);
nand g714 (n753, n365, n298, n159, n161);
nor  g715 (n608, n167, n156, n335, n130);
or   g716 (n748, n214, n330, n223, n362);
nor  g717 (n646, n193, n322, n377);
or   g718 (n732, n138, n182, n341, n348);
nor  g719 (n596, n383, n272, n453, n164);
nor  g720 (n722, n231, n371, n359, n269);
nand g721 (n758, n346, n447, n179, n169);
or   g722 (n720, n251, n364, n385, n367);
and  g723 (n574, n419, n309, n134, n233);
xnor g724 (n655, n208, n384, n325, n157);
or   g725 (n555, n235, n453, n141, n308);
nand g726 (n781, n253, n324, n391, n272);
xor  g727 (n611, n121, n340, n433, n152);
and  g728 (n560, n344, n349, n433, n333);
xnor g729 (n764, n247, n288, n419);
nand g730 (n712, n161, n245, n198, n430);
and  g731 (n583, n381, n210, n256, n211);
xnor g732 (n710, n458, n385, n464, n193);
xor  g733 (n606, n402, n405, n196, n214);
and  g734 (n794, n234, n203, n373, n429);
xor  g735 (n508, n280, n206, n168, n395);
nand g736 (n792, n236, n447, n248, n249);
or   g737 (n839, n434, n124, n246, n325);
and  g738 (n786, n394, n221, n125, n213);
xnor g739 (n714, n223, n171, n257, n375);
nor  g740 (n597, n353, n313, n158, n321);
nand g741 (n837, n126, n262, n348, n195);
xor  g742 (n576, n184, n398, n222, n339);
xnor g743 (n780, n410, n183, n186, n407);
nor  g744 (n665, n439, n284, n280, n134);
xor  g745 (n612, n330, n327, n403, n125);
nor  g746 (n632, n244, n352, n315, n172);
xnor g747 (n741, n341, n230, n190, n204);
xor  g748 (n763, n383, n205, n266, n323);
xor  g749 (n843, n178, n139, n363, n398);
xnor g750 (n498, n273, n209, n457, n365);
nor  g751 (n584, n235, n123, n321, n373);
xnor g752 (n685, n239, n155, n388, n214);
xnor g753 (n631, n397, n463, n349, n270);
nand g754 (n812, n312, n294, n257, n125);
and  g755 (n676, n283, n118, n361, n352);
nor  g756 (n834, n166, n307, n448, n346);
or   g757 (n813, n158, n437, n415, n121);
nor  g758 (n704, n392, n129, n428);
and  g759 (n520, n460, n193, n455, n281);
xnor g760 (n831, n397, n270, n427);
xnor g761 (n817, n202, n286, n271, n209);
nor  g762 (n731, n162, n159, n141, n218);
nand g763 (n730, n432, n277, n344, n192);
xnor g764 (n756, n429, n273, n216, n342);
nand g765 (n768, n384, n331, n401, n315);
nand g766 (n783, n364, n271, n292, n223);
nor  g767 (n650, n367, n208, n145, n415);
xor  g768 (n629, n332, n156, n297, n247);
nand g769 (n702, n165, n374, n437, n179);
nor  g770 (n499, n244, n409, n447, n175);
or   g771 (n833, n194, n454, n261, n370);
xor  g772 (n776, n333, n332, n133, n203);
xnor g773 (n694, n196, n155, n372, n254);
or   g774 (n644, n259, n420, n220, n265);
nor  g775 (n767, n357, n369, n171, n409);
xnor g776 (n559, n176, n242, n154, n133);
and  g777 (n725, n256, n225, n407, n317);
nand g778 (n726, n335, n403, n430, n172);
xnor g779 (n777, n169, n257, n158, n324);
nor  g780 (n778, n202, n240, n445, n409);
xor  g781 (n601, n239, n441, n334, n379);
xnor g782 (n603, n416, n161, n232, n168);
xnor g783 (n496, n373, n205, n199, n226);
xor  g784 (n540, n208, n393, n320, n399);
nand g785 (n695, n381, n395, n375, n135);
nor  g786 (n742, n250, n419, n212, n326);
or   g787 (n841, n340, n278, n334, n251);
xor  g788 (n573, n344, n312, n244, n384);
xor  g789 (n561, n210, n160, n124, n297);
or   g790 (n719, n178, n173, n432, n441);
xor  g791 (n602, n312, n125, n213, n281);
nor  g792 (n553, n345, n295, n354, n462);
or   g793 (n558, n205, n225, n328, n304);
xor  g794 (n807, n290, n414, n241, n386);
nor  g795 (n648, n463, n273, n353, n351);
nor  g796 (n607, n424, n130, n241, n389);
and  g797 (n826, n370, n446, n252, n408);
xor  g798 (n800, n456, n212, n413, n330);
nor  g799 (n664, n149, n350, n325, n419);
nand g800 (n705, n156, n200, n338, n120);
and  g801 (n746, n366, n126, n267, n186);
xor  g802 (n497, n404, n436, n277, n310);
nand g803 (n808, n290, n454, n259, n452);
xnor g804 (n816, n120, n417, n414, n348);
nand g805 (n604, n228, n310, n394, n422);
and  g806 (n512, n207, n287, n268, n399);
and  g807 (n537, n260, n167, n288, n241);
or   g808 (n505, n182, n124, n338, n410);
nand g809 (n716, n262, n276, n183, n388);
and  g810 (n638, n154, n362, n206, n361);
not  g811 (n846, n495);
not  g812 (n854, n493);
not  g813 (n853, n492);
not  g814 (n855, n147);
not  g815 (n848, n496);
buf  g816 (n852, n494);
and  g817 (n850, n146, n145);
xnor g818 (n845, n146, n146, n492, n491);
nand g819 (n851, n494, n146, n491);
or   g820 (n849, n494, n495, n491, n493);
xnor g821 (n847, n493, n495, n494, n147);
nand g822 (n844, n492, n492, n493, n495);
buf  g823 (n857, n844);
not  g824 (n856, n844);
or   g825 (n865, n496, n501, n499, n857);
xnor g826 (n864, n857, n497, n500, n501);
nor  g827 (n862, n856, n498, n499);
xnor g828 (n859, n502, n501, n857, n856);
and  g829 (n863, n497, n499, n857, n500);
nor  g830 (n860, n497, n499, n501, n496);
or   g831 (n861, n500, n497, n498);
nor  g832 (n858, n500, n856, n496);
nand g833 (n869, n863, n466, n862, n470);
nor  g834 (n880, n477, n480, n861, n482);
nor  g835 (n876, n465, n476, n472);
xor  g836 (n885, n474, n479, n470, n859);
xnor g837 (n867, n860, n844, n476, n467);
and  g838 (n878, n859, n477, n863, n464);
xnor g839 (n870, n466, n465, n481, n464);
xnor g840 (n872, n478, n473, n845, n468);
and  g841 (n881, n469, n478, n473, n863);
xnor g842 (n891, n474, n860, n479, n862);
and  g843 (n879, n471, n475, n858, n478);
and  g844 (n887, n481, n468, n861, n471);
xor  g845 (n888, n480, n858, n470, n859);
and  g846 (n875, n863, n469, n478);
or   g847 (n877, n467, n858, n862, n469);
nand g848 (n874, n481, n468, n472, n473);
nor  g849 (n882, n466, n480, n471, n864);
xnor g850 (n883, n846, n465, n482, n858);
and  g851 (n889, n859, n477, n860, n861);
or   g852 (n884, n845, n475, n481, n476);
xnor g853 (n868, n864, n482, n475, n474);
nor  g854 (n890, n466, n482, n479, n477);
xor  g855 (n886, n861, n471, n845, n480);
xor  g856 (n871, n472, n475, n465, n470);
nor  g857 (n866, n479, n472, n860, n464);
nor  g858 (n892, n473, n474, n467);
or   g859 (n873, n862, n468, n845, n864);
xor  g860 (n893, n504, n502, n503);
nand g861 (n896, n886, n883, n503, n502);
nand g862 (n895, n505, n503, n884, n504);
or   g863 (n894, n885, n504, n502);
xor  g864 (n911, n507, n895, n511, n847);
and  g865 (n898, n893, n509, n505, n510);
xnor g866 (n900, n508, n513, n864, n846);
or   g867 (n906, n893, n512, n894);
xor  g868 (n901, n509, n508, n506, n896);
nand g869 (n910, n511, n847, n512, n846);
and  g870 (n899, n508, n507, n505, n895);
and  g871 (n897, n894, n896, n847, n506);
or   g872 (n907, n846, n894, n847);
and  g873 (n905, n509, n506, n514, n513);
or   g874 (n909, n510, n893, n512, n895);
nor  g875 (n902, n513, n895, n509, n507);
nor  g876 (n908, n893, n896, n505, n510);
and  g877 (n903, n511, n510, n508, n507);
xnor g878 (n904, n514, n513, n511, n506);
or   g879 (n916, n515, n517, n514);
xnor g880 (n917, n515, n518, n899);
nand g881 (n912, n901, n515, n516, n902);
nand g882 (n915, n515, n516, n900, n518);
xnor g883 (n914, n517, n516, n518, n898);
nor  g884 (n913, n517, n897, n516, n514);
not  g885 (n919, n915);
not  g886 (n918, n913);
buf  g887 (n920, n914);
not  g888 (n921, n915);
not  g889 (n922, n919);
not  g890 (n932, n907);
buf  g891 (n928, n921);
not  g892 (n924, n918);
buf  g893 (n923, n848);
buf  g894 (n936, n920);
or   g895 (n930, n904, n865);
nor  g896 (n933, n908, n920);
or   g897 (n935, n849, n918, n865, n919);
nor  g898 (n934, n921, n919, n848, n905);
xor  g899 (n931, n887, n889, n920, n921);
nor  g900 (n925, n910, n888, n849, n918);
xnor g901 (n926, n919, n918, n850, n849);
nor  g902 (n927, n890, n909, n891, n921);
xor  g903 (n937, n920, n906, n865, n850);
or   g904 (n929, n849, n903, n848);
buf  g905 (n941, n923);
not  g906 (n939, n922);
not  g907 (n940, n922);
buf  g908 (n942, n922);
not  g909 (n938, n923);
xnor g910 (n943, n922, n519, n916);
not  g911 (n946, n911);
not  g912 (n958, n923);
buf  g913 (n947, n943);
buf  g914 (n957, n850);
buf  g915 (n952, n939);
buf  g916 (n955, n924);
not  g917 (n950, n943);
not  g918 (n949, n519);
not  g919 (n954, n940);
not  g920 (n948, n938);
buf  g921 (n951, n940);
nand g922 (n944, n520, n942, n943);
nand g923 (n953, n911, n923, n942, n943);
nand g924 (n956, n939, n942, n941);
nand g925 (n945, n924, n519, n942);
nor  g926 (n961, n927, n945, n924, n926);
xor  g927 (n959, n928, n944, n926);
nor  g928 (n963, n944, n925, n927);
and  g929 (n960, n924, n925, n927);
xnor g930 (n962, n926, n944, n927);
nor  g931 (n968, n961, n865, n948, n960);
nand g932 (n969, n962, n950, n951);
and  g933 (n967, n947, n916, n946, n960);
xor  g934 (n966, n950, n945, n949, n962);
nor  g935 (n964, n950, n948, n961, n949);
nand g936 (n972, n945, n946, n948, n949);
nand g937 (n965, n951, n945, n946);
xor  g938 (n970, n959, n947, n963);
and  g939 (n971, n949, n947, n948);
not  g940 (n981, n968);
buf  g941 (n978, n967);
not  g942 (n974, n970);
not  g943 (n983, n929);
not  g944 (n982, n969);
not  g945 (n980, n970);
not  g946 (n984, n928);
buf  g947 (n979, n929);
not  g948 (n976, n964);
buf  g949 (n977, n971);
or   g950 (n975, n968, n965, n969, n966);
xnor g951 (n973, n929, n967, n928);
nor  g952 (n985, n929, n973);
xnor g953 (n986, n951, n985, n952);
nand g954 (n987, n985, n951, n520);
nand g955 (n988, n523, n973, n987, n520);
xnor g956 (n989, n987, n522, n523);
nor  g957 (n990, n973, n522, n986, n521);
or   g958 (n992, n986, n521, n987);
xor  g959 (n991, n523, n521, n522);
xnor g960 (n993, n486, n988, n990, n485);
nor  g961 (n1010, n990, n483, n992, n991);
and  g962 (n1002, n486, n853, n483, n992);
nand g963 (n1006, n992, n524, n852, n952);
xnor g964 (n1007, n989, n954, n953, n486);
and  g965 (n995, n988, n525, n524);
or   g966 (n998, n991, n972, n483, n851);
nand g967 (n999, n991, n990, n852, n954);
nor  g968 (n1004, n954, n991, n483, n525);
nand g969 (n996, n992, n972, n484, n853);
nor  g970 (n1003, n851, n989, n853, n525);
nor  g971 (n1008, n955, n955, n852, n953);
xor  g972 (n1001, n989, n988, n485, n851);
xnor g973 (n1000, n990, n851, n486, n954);
nor  g974 (n994, n484, n526, n485, n524);
nor  g975 (n1005, n484, n526, n953, n853);
nand g976 (n1009, n953, n952, n971, n485);
nor  g977 (n997, n852, n524, n850, n484);
nand g978 (n1014, n527, n529, n993);
or   g979 (n1012, n529, n526, n993);
nand g980 (n1011, n994, n528, n526);
and  g981 (n1013, n993, n528, n530, n527);
xnor g982 (n1015, n528, n527, n529);
buf  g983 (n1019, n1012);
buf  g984 (n1017, n1012);
not  g985 (n1022, n1011);
buf  g986 (n1020, n1011);
buf  g987 (n1016, n1013);
buf  g988 (n1024, n1011);
buf  g989 (n1023, n1011);
not  g990 (n1025, n1012);
not  g991 (n1018, n1013);
not  g992 (n1021, n1012);
xor  g993 (n1060, n981, n1018, n973, n1023);
xor  g994 (n1036, n981, n855, n930, n999);
or   g995 (n1050, n530, n1024, n930, n892);
or   g996 (n1044, n1022, n999, n933, n1019);
nor  g997 (n1032, n996, n855, n931);
xnor g998 (n1042, n1022, n975, n1021, n1025);
xnor g999 (n1045, n1025, n1023, n958);
xnor g1000 (n1029, n1001, n1000, n977, n998);
xor  g1001 (n1039, n1022, n979, n1002, n1020);
xor  g1002 (n1049, n958, n531, n1018, n1021);
or   g1003 (n1048, n930, n957, n1017, n532);
nand g1004 (n1038, n854, n995, n974, n1016);
xnor g1005 (n1056, n1023, n933, n995, n1024);
nor  g1006 (n1055, n994, n981, n1021, n1016);
nand g1007 (n1062, n979, n976, n1021, n1000);
nand g1008 (n1059, n956, n854, n955, n979);
or   g1009 (n1026, n974, n956, n996);
xor  g1010 (n1065, n1024, n1025, n1018, n531);
nand g1011 (n1061, n1020, n1024, n854, n979);
xnor g1012 (n1052, n932, n1017, n976, n854);
xor  g1013 (n1040, n982, n931, n932, n955);
nand g1014 (n1027, n933, n855, n996, n1000);
and  g1015 (n1033, n1020, n995, n994, n1022);
xor  g1016 (n1053, n999, n999, n930, n980);
nor  g1017 (n1051, n996, n530, n974, n531);
and  g1018 (n1030, n998, n978, n1016, n1019);
nand g1019 (n1046, n980, n975, n997, n994);
xnor g1020 (n1054, n1001, n956, n1017, n976);
nor  g1021 (n1063, n958, n934, n998, n957);
xnor g1022 (n1047, n1018, n980, n977, n997);
xnor g1023 (n1058, n933, n1000, n980, n995);
xnor g1024 (n1043, n975, n997, n532, n982);
nor  g1025 (n1064, n1001, n1017, n977, n533);
nand g1026 (n1037, n530, n531, n1020, n982);
and  g1027 (n1041, n855, n977, n532, n978);
or   g1028 (n1035, n1025, n932, n974);
or   g1029 (n1028, n978, n1019, n998, n1001);
or   g1030 (n1031, n997, n976, n978, n981);
nand g1031 (n1034, n1019, n957, n931, n975);
xnor g1032 (n1057, n957, n1016, n532, n958);
xnor g1033 (n1132, n626, n579, n561, n615);
nor  g1034 (n1190, n594, n629, n628, n566);
or   g1035 (n1177, n592, n1033, n553, n620);
xnor g1036 (n1102, n549, n567, n1064, n1036);
nor  g1037 (n1166, n628, n1063, n590, n1014);
xnor g1038 (n1208, n650, n1026, n541, n619);
xor  g1039 (n1113, n533, n646, n540, n1061);
and  g1040 (n1117, n1034, n577, n580, n1055);
and  g1041 (n1187, n643, n554, n577, n589);
nor  g1042 (n1186, n1030, n624, n646, n1028);
xor  g1043 (n1211, n620, n623, n595, n597);
xor  g1044 (n1179, n1043, n1047, n600, n599);
xor  g1045 (n1076, n1047, n543, n1043, n1044);
and  g1046 (n1189, n1032, n583, n1061, n636);
xor  g1047 (n1141, n626, n568, n566, n585);
nor  g1048 (n1171, n617, n639, n583, n550);
or   g1049 (n1140, n534, n589, n598, n1063);
and  g1050 (n1180, n1041, n577, n636, n641);
xor  g1051 (n1134, n643, n1059, n594, n631);
nor  g1052 (n1108, n638, n622, n572, n551);
and  g1053 (n1198, n536, n571, n1062, n1057);
nor  g1054 (n1195, n627, n535, n583, n602);
nand g1055 (n1105, n621, n552, n605);
xnor g1056 (n1178, n633, n582, n646, n1042);
and  g1057 (n1082, n586, n643, n648, n1028);
nand g1058 (n1212, n610, n564, n635, n585);
xor  g1059 (n1191, n645, n534, n567, n1035);
or   g1060 (n1217, n572, n1063, n555, n595);
xnor g1061 (n1072, n584, n535, n591, n574);
nor  g1062 (n1090, n1030, n563, n1038, n568);
nand g1063 (n1078, n581, n649, n611, n637);
xor  g1064 (n1183, n1059, n613, n1036, n600);
nor  g1065 (n1074, n627, n543, n1053, n592);
and  g1066 (n1207, n587, n1063, n584, n1052);
and  g1067 (n1147, n574, n1052, n606, n578);
nor  g1068 (n1167, n632, n1048, n600, n619);
nor  g1069 (n1160, n563, n555, n595, n621);
nand g1070 (n1094, n630, n1057, n1031, n538);
nor  g1071 (n1158, n1026, n590, n606, n638);
nand g1072 (n1081, n596, n983, n577, n555);
nor  g1073 (n1069, n982, n544, n576, n627);
or   g1074 (n1223, n614, n590, n1039, n559);
xnor g1075 (n1083, n648, n617, n1036, n643);
xor  g1076 (n1116, n1013, n618, n1064, n1033);
xnor g1077 (n1123, n1058, n1064, n588, n642);
xnor g1078 (n1193, n1039, n556, n575, n1035);
and  g1079 (n1219, n625, n568, n615, n1058);
xnor g1080 (n1203, n544, n603, n606, n632);
nor  g1081 (n1168, n1048, n605, n580, n564);
nand g1082 (n1104, n605, n639, n1037, n549);
xnor g1083 (n1096, n1050, n565, n1028, n597);
nand g1084 (n1111, n1031, n1053, n1027, n576);
or   g1085 (n1201, n600, n570, n611, n1041);
nand g1086 (n1097, n541, n557, n1059, n1046);
or   g1087 (n1086, n571, n536, n1026, n579);
nor  g1088 (n1109, n641, n558, n618, n648);
nand g1089 (n1070, n588, n597, n1051, n573);
or   g1090 (n1080, n571, n591, n597, n544);
nand g1091 (n1133, n623, n585, n596, n603);
and  g1092 (n1143, n1047, n612, n616, n618);
nand g1093 (n1126, n604, n645, n633, n649);
or   g1094 (n1206, n539, n1034, n595, n583);
xnor g1095 (n1200, n1065, n602, n1064, n537);
or   g1096 (n1192, n564, n543, n1037, n558);
and  g1097 (n1176, n593, n533, n549, n608);
or   g1098 (n1066, n609, n551, n1052, n1040);
or   g1099 (n1152, n1046, n615, n562, n645);
and  g1100 (n1071, n1034, n983, n601, n630);
xor  g1101 (n1087, n579, n561, n637, n567);
xor  g1102 (n1222, n560, n1054, n645, n650);
or   g1103 (n1121, n574, n1044, n538, n613);
xnor g1104 (n1079, n602, n539, n584, n618);
nor  g1105 (n1091, n544, n1027, n647, n598);
and  g1106 (n1225, n555, n550, n537, n566);
nor  g1107 (n1196, n1050, n1035, n548, n617);
or   g1108 (n1088, n1055, n538, n599, n1035);
nand g1109 (n1202, n536, n622, n533, n1043);
xor  g1110 (n1153, n1040, n559, n610, n1061);
nor  g1111 (n1095, n1028, n1040, n1041, n1045);
xor  g1112 (n1101, n545, n559, n1031, n622);
and  g1113 (n1213, n539, n542, n1014);
xor  g1114 (n1214, n1029, n564, n625, n575);
or   g1115 (n1172, n983, n546, n1058, n642);
or   g1116 (n1130, n568, n623, n647, n586);
or   g1117 (n1098, n1037, n1014, n586, n546);
and  g1118 (n1077, n641, n628, n581, n629);
nand g1119 (n1136, n553, n552, n649, n579);
xor  g1120 (n1085, n570, n538, n569, n1039);
and  g1121 (n1159, n562, n634, n609, n607);
or   g1122 (n1120, n1049, n630, n1048, n626);
nor  g1123 (n1182, n601, n614, n615, n619);
xnor g1124 (n1115, n984, n554, n644, n563);
nand g1125 (n1119, n553, n566, n638, n1049);
nor  g1126 (n1110, n593, n598, n1044, n535);
xnor g1127 (n1092, n1034, n1065, n644, n587);
xor  g1128 (n1164, n545, n541, n1049, n638);
xnor g1129 (n1199, n640, n1057, n548, n1038);
nand g1130 (n1138, n560, n644, n610, n604);
nand g1131 (n1156, n606, n570, n599, n1056);
xor  g1132 (n1100, n649, n619, n610, n546);
xnor g1133 (n1181, n648, n547, n554, n562);
or   g1134 (n1220, n537, n616, n621, n634);
and  g1135 (n1129, n536, n1060, n1045, n594);
nor  g1136 (n1224, n644, n631, n614, n635);
and  g1137 (n1089, n558, n572, n1056, n588);
nand g1138 (n1154, n624, n636, n574, n569);
xor  g1139 (n1197, n551, n1043, n603, n642);
and  g1140 (n1099, n633, n573, n545, n604);
nand g1141 (n1209, n563, n983, n560, n559);
xor  g1142 (n1163, n557, n635, n592, n625);
nand g1143 (n1075, n565, n628, n560, n1058);
or   g1144 (n1205, n575, n588, n591, n1050);
nor  g1145 (n1204, n534, n1039, n1054, n1046);
and  g1146 (n1218, n541, n552, n1030, n569);
or   g1147 (n1073, n556, n624, n547, n551);
or   g1148 (n1107, n1062, n621, n585, n608);
nor  g1149 (n1174, n591, n1030, n625, n1029);
nor  g1150 (n1103, n1045, n612, n594, n578);
xor  g1151 (n1106, n548, n608, n590, n547);
nor  g1152 (n1165, n1033, n601, n1051, n1061);
and  g1153 (n1145, n1053, n540, n1032, n640);
xor  g1154 (n1142, n534, n1065, n1056, n582);
nand g1155 (n1149, n626, n586, n1050, n578);
nor  g1156 (n1148, n604, n554, n647, n587);
nand g1157 (n1114, n1040, n1054, n1038, n631);
xnor g1158 (n1068, n570, n1013, n1047, n1060);
xor  g1159 (n1215, n1051, n569, n624, n1045);
nor  g1160 (n1124, n633, n1046, n640, n607);
and  g1161 (n1210, n539, n632, n1029, n614);
xor  g1162 (n1162, n616, n593, n634);
xor  g1163 (n1150, n576, n608, n1036, n646);
nor  g1164 (n1137, n580, n542, n1056, n556);
nand g1165 (n1146, n1060, n596, n553, n545);
nor  g1166 (n1131, n1049, n601, n1053, n578);
nand g1167 (n1194, n612, n582, n1062, n639);
nand g1168 (n1184, n589, n1065, n609, n622);
xor  g1169 (n1157, n581, n557, n641, n1060);
xor  g1170 (n1175, n1052, n1062, n613, n598);
xor  g1171 (n1155, n587, n548, n635, n1027);
and  g1172 (n1161, n582, n1026, n639, n556);
and  g1173 (n1170, n567, n617, n640, n565);
nor  g1174 (n1173, n1037, n636, n596, n607);
nand g1175 (n1144, n573, n543, n642, n613);
nand g1176 (n1169, n557, n1054, n647, n542);
xor  g1177 (n1216, n1042, n571, n581, n609);
and  g1178 (n1188, n620, n630, n552, n623);
nor  g1179 (n1093, n1032, n561, n1027, n607);
nand g1180 (n1122, n540, n562, n637, n1041);
xnor g1181 (n1067, n572, n629, n627, n573);
and  g1182 (n1151, n592, n611, n1044, n1048);
xnor g1183 (n1118, n589, n580, n602, n561);
nor  g1184 (n1139, n565, n550, n603, n549);
and  g1185 (n1125, n1038, n599, n1031, n540);
xnor g1186 (n1128, n1029, n1032, n558, n1057);
or   g1187 (n1135, n1055, n550, n584, n612);
and  g1188 (n1084, n616, n547, n632, n1059);
nand g1189 (n1127, n593, n546, n537, n575);
nor  g1190 (n1221, n576, n1051, n637, n1033);
xor  g1191 (n1112, n620, n631, n1042, n535);
nand g1192 (n1185, n611, n1055, n629, n1042);
buf  g1193 (n1316, n1090);
nor  g1194 (n1273, n1125, n1004, n1148, n1167);
xor  g1195 (n1305, n1145, n1163, n1157, n1138);
nor  g1196 (n1302, n1107, n1141, n1156, n1115);
xnor g1197 (n1262, n1173, n1119, n1176, n1136);
nand g1198 (n1301, n1141, n1175, n1131, n1125);
nand g1199 (n1279, n1077, n1173, n1106, n1005);
xnor g1200 (n1339, n1098, n1002, n1140, n1183);
and  g1201 (n1315, n937, n1180, n1096, n1112);
and  g1202 (n1296, n1148, n1070, n1143, n1134);
or   g1203 (n1360, n1086, n1153, n1143, n1145);
and  g1204 (n1270, n1080, n1153, n1167, n1083);
xnor g1205 (n1240, n1068, n1098, n1114, n1095);
nor  g1206 (n1234, n1126, n1072, n1087, n1170);
xor  g1207 (n1300, n1184, n1141, n1079, n1144);
nand g1208 (n1338, n1111, n1149, n1123, n1182);
xnor g1209 (n1285, n1132, n1005, n1181, n1155);
xor  g1210 (n1310, n1179, n1138, n651, n1078);
nor  g1211 (n1352, n1106, n1148, n1083, n1072);
xnor g1212 (n1344, n1083, n1181, n1087, n1102);
xnor g1213 (n1243, n1099, n1124, n935, n1111);
and  g1214 (n1246, n935, n1158, n1005, n1160);
or   g1215 (n1331, n1172, n1089, n1140, n1125);
nand g1216 (n1256, n1113, n1073, n1142, n1162);
xor  g1217 (n1321, n1166, n1185, n1089, n1076);
or   g1218 (n1238, n1103, n1181, n1154, n1010);
nand g1219 (n1319, n1118, n1007, n1176, n1159);
nor  g1220 (n1280, n1101, n1074, n1153, n1069);
or   g1221 (n1332, n1118, n1093, n1128, n1117);
xor  g1222 (n1269, n1086, n1104, n1068, n1174);
xnor g1223 (n1288, n1168, n1163, n1113, n1104);
nor  g1224 (n1231, n1097, n1154, n1098, n1089);
or   g1225 (n1320, n1073, n1099, n1002, n1104);
xnor g1226 (n1295, n1178, n1133, n1107, n934);
nor  g1227 (n1325, n652, n1138, n1172, n1105);
nand g1228 (n1260, n1112, n1120, n1184, n1178);
nand g1229 (n1244, n1117, n1082, n1120, n1173);
or   g1230 (n1329, n1159, n1183, n1116, n1142);
nand g1231 (n1347, n1082, n1143, n1066, n1115);
or   g1232 (n1290, n1129, n1174, n1086, n1156);
nand g1233 (n1228, n1110, n1183, n1138, n1100);
xnor g1234 (n1335, n1140, n1080, n1114, n1177);
and  g1235 (n1277, n1133, n1152, n1173, n1135);
xor  g1236 (n1237, n1094, n1073, n1147, n1137);
nand g1237 (n1275, n1132, n1175, n1135, n1078);
and  g1238 (n1272, n1125, n1171, n1110, n1127);
xor  g1239 (n1333, n1109, n1110, n1162, n1123);
or   g1240 (n1309, n1144, n1185, n1102, n937);
nand g1241 (n1343, n1097, n1003, n1160, n1112);
or   g1242 (n1322, n1124, n1180, n1127, n1179);
nand g1243 (n1304, n1159, n1115, n1161, n1153);
or   g1244 (n1266, n1091, n1164, n1069, n1093);
or   g1245 (n1247, n1131, n1120, n1091, n1006);
xnor g1246 (n1251, n1166, n1136, n1112, n652);
nand g1247 (n1351, n1004, n1077, n1009, n1161);
xnor g1248 (n1263, n1146, n1128, n1168, n1157);
xor  g1249 (n1233, n1009, n1121, n1094, n1171);
or   g1250 (n1291, n1072, n1102, n1085);
xnor g1251 (n1307, n1096, n1150, n1007, n1161);
and  g1252 (n1271, n1130, n1123, n1088, n1167);
nor  g1253 (n1337, n1148, n1079, n935, n1074);
and  g1254 (n1357, n1069, n1149, n1113, n1123);
nor  g1255 (n1254, n1067, n1151, n1164, n1106);
nand g1256 (n1283, n1139, n1068, n1119, n1135);
nor  g1257 (n1226, n1103, n1120, n1006, n1132);
nand g1258 (n1232, n1099, n1111, n1119, n1133);
xor  g1259 (n1249, n1094, n1071, n1119, n1155);
xor  g1260 (n1359, n1091, n1092, n1166, n1003);
xor  g1261 (n1230, n1085, n1166, n1122, n1150);
nor  g1262 (n1278, n1151, n1006, n1134, n1146);
or   g1263 (n1354, n1115, n1156, n1005, n1144);
and  g1264 (n1350, n937, n936, n1086, n1091);
nor  g1265 (n1340, n1186, n1126, n1010, n1142);
nand g1266 (n1252, n1163, n1108, n1146, n1179);
or   g1267 (n1314, n1117, n1164, n1137, n1067);
xnor g1268 (n1242, n1150, n1097, n1139, n1146);
or   g1269 (n1348, n1070, n1010, n1143, n1109);
nor  g1270 (n1346, n1176, n1067, n934, n1170);
and  g1271 (n1324, n1003, n917, n1007, n1172);
nand g1272 (n1236, n1095, n1157, n1078, n1177);
and  g1273 (n1265, n650, n1155, n1008, n1088);
nand g1274 (n1361, n1075, n650, n1182, n1087);
and  g1275 (n1345, n1080, n1110, n1002, n1089);
xnor g1276 (n1358, n1082, n1073, n1128, n1066);
nor  g1277 (n1289, n1163, n1136, n1066, n1124);
nor  g1278 (n1286, n1066, n1128, n651, n1183);
nor  g1279 (n1239, n1152, n1095, n1116, n1177);
nor  g1280 (n1284, n1114, n1004, n1116, n1177);
nand g1281 (n1330, n1075, n1184, n1084, n1150);
nor  g1282 (n1313, n1130, n1105, n1118, n1077);
xnor g1283 (n1274, n1084, n1116, n1076, n1137);
nor  g1284 (n1312, n1127, n1081, n1090, n1170);
nand g1285 (n1258, n1152, n1165, n1092, n1080);
nand g1286 (n1299, n1109, n1147, n652, n1136);
or   g1287 (n1298, n1105, n1126, n1129, n1006);
nor  g1288 (n1327, n1165, n1100, n1180, n936);
nand g1289 (n1318, n1145, n1097, n935, n1176);
nand g1290 (n1227, n1092, n1100, n1185, n1008);
nand g1291 (n1276, n1149, n1101, n1157, n1121);
nand g1292 (n1326, n1104, n1167, n1132, n1168);
xor  g1293 (n1336, n1094, n1181, n1141, n1071);
nand g1294 (n1323, n1103, n1084, n1008, n1168);
or   g1295 (n1341, n1078, n1008, n651, n1079);
and  g1296 (n1334, n1071, n1129, n1079, n1170);
nand g1297 (n1306, n1131, n1130, n1108, n1178);
or   g1298 (n1297, n1135, n1144, n1122, n1121);
xor  g1299 (n1287, n1169, n1075, n1149, n1070);
and  g1300 (n1267, n1004, n1175, n1172, n1165);
and  g1301 (n1248, n1105, n1070, n1162, n1185);
nand g1302 (n1342, n1130, n1169, n1122, n1108);
and  g1303 (n1235, n1109, n1075, n1152, n1118);
xor  g1304 (n1253, n1142, n1139, n1129, n1154);
xor  g1305 (n1241, n1090, n1133, n1147, n936);
xor  g1306 (n1250, n1074, n1147, n1140, n1082);
xor  g1307 (n1311, n1111, n917, n1067, n936);
and  g1308 (n1261, n1117, n1159, n1179, n1093);
xor  g1309 (n1294, n1081, n1180, n1162, n1093);
nand g1310 (n1293, n1174, n1009, n1158, n1077);
xnor g1311 (n1259, n1154, n1076, n1161);
xor  g1312 (n1281, n1092, n1099, n1100, n1158);
xnor g1313 (n1264, n1081, n1124, n1178, n1088);
or   g1314 (n1356, n1101, n1083, n1113, n1102);
xor  g1315 (n1257, n1098, n1160, n1169, n1175);
nand g1316 (n1255, n1139, n1010, n1085, n1088);
xor  g1317 (n1292, n1107, n1156, n1072, n1122);
nor  g1318 (n1268, n1007, n1069, n1127, n1169);
and  g1319 (n1282, n934, n1174, n1103, n1160);
or   g1320 (n1303, n1095, n1090, n1151, n651);
xor  g1321 (n1328, n1151, n1074, n1096);
and  g1322 (n1349, n1126, n1009, n1155, n1068);
xnor g1323 (n1353, n1114, n1171, n1134);
nor  g1324 (n1245, n1158, n1101, n1107, n1165);
or   g1325 (n1229, n1182, n1071, n1164, n1003);
or   g1326 (n1317, n1145, n1087, n1108, n1106);
xnor g1327 (n1355, n1171, n1084, n1131, n1182);
and  g1328 (n1308, n1184, n1137, n1121, n1081);
and  g1329 (n1677, n1292, n717, n780, n1360);
xnor g1330 (n1493, n1223, n1259, n1245, n728);
or   g1331 (n1590, n786, n695, n1293, n1283);
and  g1332 (n1514, n1345, n1253, n753);
and  g1333 (n1520, n682, n828, n1191, n1310);
nand g1334 (n1592, n837, n1253, n697, n1265);
xor  g1335 (n1704, n1318, n739, n1252, n662);
and  g1336 (n1474, n715, n1346, n1289, n1360);
or   g1337 (n1699, n715, n1243, n1221, n812);
xor  g1338 (n1568, n676, n832, n662, n1314);
xnor g1339 (n1503, n655, n1323, n839, n1297);
nand g1340 (n1484, n827, n1243, n1322, n1213);
or   g1341 (n1475, n712, n782, n490, n1230);
and  g1342 (n1695, n840, n749, n832, n1298);
or   g1343 (n1429, n1226, n801, n1237, n1015);
xor  g1344 (n1521, n774, n670, n747, n1342);
xor  g1345 (n1727, n1276, n1347, n1241, n1295);
nand g1346 (n1606, n1285, n1277, n821, n1219);
nor  g1347 (n1389, n790, n761, n742, n1236);
xor  g1348 (n1731, n826, n1339, n1343, n1313);
xor  g1349 (n1670, n792, n1236, n1298, n751);
and  g1350 (n1630, n1314, n694, n1223, n771);
xnor g1351 (n1644, n1208, n729, n1237, n673);
or   g1352 (n1496, n1214, n1192, n757, n843);
xor  g1353 (n1689, n726, n1251, n736, n1352);
nor  g1354 (n1382, n1187, n1361, n1291, n689);
nor  g1355 (n1435, n719, n1329, n1296, n807);
xor  g1356 (n1684, n1239, n1262, n705, n822);
xnor g1357 (n1585, n699, n746, n689, n1242);
xnor g1358 (n1694, n811, n836, n1199, n1222);
nand g1359 (n1528, n1198, n1209, n710, n1317);
nand g1360 (n1519, n811, n841, n1331, n742);
nor  g1361 (n1634, n1305, n1335, n1256, n699);
nor  g1362 (n1525, n1330, n838, n666, n671);
and  g1363 (n1579, n811, n727, n825, n1294);
and  g1364 (n1556, n767, n825, n812, n1194);
nand g1365 (n1529, n1250, n753, n1356, n729);
xor  g1366 (n1413, n1223, n715, n769, n694);
nand g1367 (n1444, n1202, n795, n685, n1217);
xor  g1368 (n1646, n1243, n817, n839, n1214);
xor  g1369 (n1708, n681, n743, n1211, n816);
xnor g1370 (n1460, n808, n740, n1263, n697);
xnor g1371 (n1669, n1322, n658, n653, n762);
xnor g1372 (n1485, n1205, n771, n1194, n674);
nand g1373 (n1655, n1276, n707, n1271, n1351);
or   g1374 (n1392, n734, n1300, n1257, n758);
and  g1375 (n1407, n1267, n1270, n745, n1315);
or   g1376 (n1645, n728, n770, n691, n725);
and  g1377 (n1406, n685, n770, n714, n814);
xor  g1378 (n1458, n837, n677, n1299, n1272);
nor  g1379 (n1553, n758, n793, n832, n764);
and  g1380 (n1540, n775, n1261, n782, n700);
nand g1381 (n1633, n1316, n822, n716, n756);
xnor g1382 (n1650, n819, n718, n1329, n1288);
xor  g1383 (n1602, n788, n789, n719, n1204);
xor  g1384 (n1608, n1312, n669, n1309, n819);
nand g1385 (n1533, n750, n1306, n653, n746);
or   g1386 (n1618, n1314, n700, n682, n669);
nor  g1387 (n1656, n768, n808, n1352, n1343);
or   g1388 (n1397, n738, n1259, n658, n777);
nor  g1389 (n1623, n656, n788, n800, n781);
xor  g1390 (n1654, n840, n824, n723, n843);
or   g1391 (n1719, n841, n712, n835, n1238);
nor  g1392 (n1467, n766, n1230, n1228, n1212);
or   g1393 (n1643, n752, n785, n666, n1329);
and  g1394 (n1723, n686, n1198, n1328, n1215);
nand g1395 (n1405, n1339, n693, n1233, n783);
or   g1396 (n1648, n825, n1304, n1300, n732);
or   g1397 (n1594, n800, n1215, n791, n1210);
xnor g1398 (n1588, n789, n661, n1188, n1272);
and  g1399 (n1398, n1265, n1335, n1250, n697);
or   g1400 (n1378, n663, n711, n817, n1190);
and  g1401 (n1721, n784, n748, n1228, n1015);
xor  g1402 (n1614, n1247, n754, n752, n787);
nor  g1403 (n1536, n820, n785, n698, n702);
nor  g1404 (n1679, n705, n1345, n841, n1210);
or   g1405 (n1619, n1239, n765, n489, n784);
or   g1406 (n1470, n1313, n688, n810, n1321);
nand g1407 (n1627, n1326, n713, n687, n830);
xor  g1408 (n1472, n1246, n684, n823, n820);
or   g1409 (n1576, n811, n722, n784, n740);
xnor g1410 (n1542, n726, n1271, n829, n1356);
xnor g1411 (n1483, n1333, n675, n1225, n1275);
or   g1412 (n1551, n802, n1261, n1298, n754);
xnor g1413 (n1587, n1205, n665, n682, n1288);
xnor g1414 (n1544, n1212, n1189, n1304, n700);
xnor g1415 (n1701, n488, n769, n1218, n1246);
xnor g1416 (n1543, n721, n734, n722, n688);
xor  g1417 (n1605, n756, n1340, n757, n1195);
xnor g1418 (n1687, n767, n1330, n1259, n828);
nor  g1419 (n1675, n1291, n786, n1359, n838);
nor  g1420 (n1658, n668, n777, n1347, n797);
and  g1421 (n1370, n1222, n684, n693, n718);
xnor g1422 (n1686, n1244, n827, n1230, n661);
or   g1423 (n1638, n1246, n1328, n690, n1292);
xor  g1424 (n1548, n1336, n1206, n657, n1352);
xnor g1425 (n1499, n1310, n1284, n774, n1290);
xor  g1426 (n1577, n1268, n1247, n808, n1319);
or   g1427 (n1570, n1342, n1261, n827, n725);
or   g1428 (n1511, n764, n831, n694, n984);
nand g1429 (n1416, n666, n1276, n831, n1309);
nand g1430 (n1452, n1212, n794, n737, n1331);
nor  g1431 (n1598, n817, n786, n698, n1234);
nand g1432 (n1404, n761, n703, n1238, n693);
nor  g1433 (n1364, n675, n829, n984, n1349);
nand g1434 (n1437, n803, n1332, n1233, n1301);
xor  g1435 (n1522, n1272, n1278, n719, n816);
xnor g1436 (n1698, n1189, n1225, n663, n743);
xnor g1437 (n1620, n694, n824, n1359, n829);
and  g1438 (n1418, n759, n666, n821, n766);
xor  g1439 (n1597, n1262, n1269, n746, n833);
xnor g1440 (n1479, n744, n734, n671, n790);
nand g1441 (n1586, n1322, n738, n1355, n670);
nor  g1442 (n1705, n660, n1288, n793, n1293);
and  g1443 (n1509, n785, n683, n723, n1345);
nand g1444 (n1412, n784, n775, n1353, n701);
nor  g1445 (n1569, n760, n1188, n1189, n732);
nor  g1446 (n1534, n1326, n1264, n487, n1245);
nand g1447 (n1440, n705, n679, n1341, n737);
and  g1448 (n1402, n488, n1346, n805, n757);
nand g1449 (n1447, n653, n724, n1280, n1318);
xor  g1450 (n1660, n1295, n1353, n813, n669);
xnor g1451 (n1446, n1324, n1265, n744, n755);
nor  g1452 (n1510, n793, n1348, n1259, n1263);
nor  g1453 (n1545, n1268, n1357, n779, n1348);
nor  g1454 (n1393, n728, n730, n1192, n720);
and  g1455 (n1451, n695, n1357, n805, n781);
nor  g1456 (n1575, n748, n772, n832, n823);
or   g1457 (n1517, n1291, n1280, n1279, n1338);
and  g1458 (n1601, n1323, n1324, n1215, n1286);
nor  g1459 (n1417, n680, n1341, n655, n1317);
nand g1460 (n1729, n654, n711, n751, n817);
nor  g1461 (n1672, n1260, n1337, n745, n1319);
or   g1462 (n1367, n800, n896, n1300, n1282);
or   g1463 (n1603, n1270, n682, n1320, n757);
xnor g1464 (n1450, n1313, n683, n767, n1273);
nand g1465 (n1631, n1278, n1320, n1318, n708);
xnor g1466 (n1647, n1313, n833, n842, n1202);
nand g1467 (n1464, n1316, n1301, n1312, n733);
or   g1468 (n1527, n779, n751, n790, n1206);
and  g1469 (n1507, n741, n1193, n831, n730);
nor  g1470 (n1371, n679, n1255, n1196, n658);
nor  g1471 (n1730, n1306, n1334, n1200, n798);
nand g1472 (n1461, n1197, n690, n1258, n704);
xor  g1473 (n1414, n794, n1337, n778, n834);
nand g1474 (n1408, n1322, n668, n1273, n755);
and  g1475 (n1506, n487, n838, n737, n1245);
or   g1476 (n1366, n1189, n731, n1219, n1355);
nand g1477 (n1425, n685, n729, n1253, n1267);
nor  g1478 (n1681, n1309, n701, n731, n1228);
xor  g1479 (n1637, n1264, n692, n748, n767);
or   g1480 (n1693, n1346, n684, n707, n1249);
xor  g1481 (n1494, n1204, n684, n1226, n1208);
xnor g1482 (n1428, n760, n659, n1211, n713);
xnor g1483 (n1573, n779, n1274, n683, n1333);
xnor g1484 (n1682, n673, n1257, n1213, n1305);
and  g1485 (n1615, n762, n1354, n1269, n1200);
or   g1486 (n1571, n1249, n735, n721, n716);
or   g1487 (n1700, n656, n700, n1321, n1344);
nor  g1488 (n1652, n1266, n1290, n809, n713);
xor  g1489 (n1728, n1300, n782, n803, n796);
or   g1490 (n1487, n1015, n1266, n1358, n1279);
xnor g1491 (n1668, n1342, n764, n1209, n1273);
nand g1492 (n1369, n679, n687, n1301, n790);
xnor g1493 (n1385, n763, n1250, n830, n490);
nand g1494 (n1726, n1187, n796, n1326, n724);
or   g1495 (n1430, n731, n702, n1224, n1306);
xnor g1496 (n1733, n1257, n1351, n688, n1251);
and  g1497 (n1667, n765, n1349, n1186, n1341);
xor  g1498 (n1635, n487, n803, n1336, n701);
and  g1499 (n1365, n768, n1345, n667, n1361);
and  g1500 (n1566, n724, n766, n1262, n754);
nand g1501 (n1690, n1281, n733, n1214, n739);
nand g1502 (n1535, n1227, n664, n1336, n1190);
nor  g1503 (n1531, n1240, n840, n796, n1354);
xor  g1504 (n1489, n661, n1229, n821, n760);
nand g1505 (n1439, n1015, n671, n805, n1197);
and  g1506 (n1478, n823, n1239, n1207, n768);
xnor g1507 (n1426, n1279, n1245, n1327, n1305);
xnor g1508 (n1607, n717, n662, n1197, n1254);
or   g1509 (n1593, n764, n1316, n1284, n781);
nand g1510 (n1639, n1188, n1337, n691, n1232);
nor  g1511 (n1659, n1295, n1252, n772, n686);
xor  g1512 (n1488, n816, n714, n1200, n806);
nor  g1513 (n1578, n812, n1266, n1303, n783);
nand g1514 (n1717, n691, n656, n487, n1271);
nor  g1515 (n1703, n667, n1267, n775, n1359);
xor  g1516 (n1716, n788, n1254, n798, n1355);
xor  g1517 (n1554, n842, n1204, n1237, n1235);
xnor g1518 (n1589, n1324, n795, n820, n815);
or   g1519 (n1604, n1344, n1351, n696, n804);
or   g1520 (n1626, n680, n1200, n1190, n1214);
and  g1521 (n1560, n1283, n678, n813, n1250);
xnor g1522 (n1676, n1273, n704, n819, n1340);
xnor g1523 (n1581, n697, n814, n1211, n1303);
xor  g1524 (n1713, n1279, n1354, n676, n1233);
nor  g1525 (n1410, n1334, n1341, n1207, n1221);
nand g1526 (n1584, n1223, n787, n1298, n1340);
nand g1527 (n1383, n1204, n1283, n1311, n1336);
xnor g1528 (n1495, n704, n667, n1242, n791);
nand g1529 (n1558, n1275, n712, n1284, n722);
nand g1530 (n1486, n802, n1206, n773, n775);
nor  g1531 (n1424, n681, n743, n696, n1263);
or   g1532 (n1420, n734, n719, n1217, n1357);
nand g1533 (n1629, n830, n1344, n747, n820);
nand g1534 (n1471, n1201, n1270, n723, n668);
nor  g1535 (n1664, n674, n704, n756, n1251);
nor  g1536 (n1436, n681, n1231, n1307, n736);
nand g1537 (n1691, n1350, n1248, n672, n1278);
and  g1538 (n1688, n1358, n1229, n1203, n1343);
xor  g1539 (n1621, n1307, n1218, n818, n799);
nor  g1540 (n1583, n680, n1260, n725, n747);
nor  g1541 (n1710, n1330, n1240, n1309, n828);
xnor g1542 (n1657, n1216, n1227, n840, n665);
nand g1543 (n1438, n810, n692, n1335, n1277);
xor  g1544 (n1375, n1220, n778, n706, n745);
or   g1545 (n1415, n1256, n1316, n1339, n675);
xor  g1546 (n1482, n1194, n741, n674, n1246);
and  g1547 (n1711, n1358, n1014, n1352, n489);
xnor g1548 (n1546, n1343, n827, n1335, n751);
and  g1549 (n1674, n685, n804, n670, n1257);
nand g1550 (n1476, n814, n676, n669, n1281);
or   g1551 (n1555, n766, n1206, n692, n1315);
nor  g1552 (n1539, n1210, n1190, n1290, n753);
or   g1553 (n1409, n1297, n1293, n759, n1347);
xor  g1554 (n1666, n1216, n749, n792, n1220);
nor  g1555 (n1411, n776, n758, n797, n843);
xor  g1556 (n1481, n673, n772, n1198, n1238);
nand g1557 (n1538, n1251, n1216, n1338, n1287);
xnor g1558 (n1616, n801, n824, n655, n1310);
and  g1559 (n1395, n1249, n1238, n1265, n663);
xor  g1560 (n1724, n1235, n1291, n752, n836);
xor  g1561 (n1683, n1353, n842, n714, n1191);
nor  g1562 (n1463, n716, n787, n1207, n1296);
or   g1563 (n1491, n1262, n703, n1296, n802);
and  g1564 (n1649, n1229, n709, n809, n813);
xor  g1565 (n1697, n1258, n777, n1244, n733);
xor  g1566 (n1500, n664, n1285, n1318, n1210);
xor  g1567 (n1427, n706, n789, n1353, n777);
nor  g1568 (n1718, n708, n1361, n1241, n687);
or   g1569 (n1445, n765, n821, n1289, n710);
or   g1570 (n1610, n802, n742, n1264, n1234);
or   g1571 (n1492, n1270, n1202, n735, n773);
nand g1572 (n1609, n703, n1269, n1264, n695);
xnor g1573 (n1595, n726, n657, n793, n1195);
or   g1574 (n1612, n1302, n774, n792, n1339);
nand g1575 (n1391, n661, n1268, n1360, n665);
or   g1576 (n1526, n1281, n1317, n756, n720);
and  g1577 (n1377, n740, n818, n769, n1232);
nand g1578 (n1562, n1234, n668, n712, n672);
nand g1579 (n1421, n689, n1222, n1358, n815);
xnor g1580 (n1530, n683, n654, n678, n1327);
and  g1581 (n1455, n1325, n1299, n776, n652);
nor  g1582 (n1665, n698, n1218, n701, n1306);
xor  g1583 (n1696, n842, n1356, n1319, n1354);
and  g1584 (n1640, n676, n717, n800, n1348);
nand g1585 (n1663, n804, n776, n720, n664);
and  g1586 (n1565, n809, n688, n1243, n1271);
nor  g1587 (n1399, n681, n680, n738, n798);
xnor g1588 (n1448, n1274, n689, n745, n657);
xor  g1589 (n1532, n1256, n1227, n797, n664);
and  g1590 (n1473, n1227, n825, n488, n782);
and  g1591 (n1707, n736, n843, n779, n1292);
xnor g1592 (n1559, n1221, n788, n1195, n1202);
xnor g1593 (n1734, n1280, n1289, n1216, n806);
and  g1594 (n1422, n1274, n1293, n806, n1326);
nor  g1595 (n1680, n1194, n490, n770);
and  g1596 (n1722, n809, n1187, n1272, n769);
xor  g1597 (n1591, n1290, n1237, n1292, n1320);
and  g1598 (n1574, n1218, n1258, n660, n1360);
xnor g1599 (n1714, n717, n1230, n801, n658);
xor  g1600 (n1561, n709, n686, n1355, n1208);
xor  g1601 (n1466, n781, n686, n813, n1304);
or   g1602 (n1403, n727, n765, n1331, n1330);
nor  g1603 (n1547, n1209, n829, n1356, n1207);
and  g1604 (n1596, n1323, n1317, n1242, n1307);
and  g1605 (n1502, n1247, n692, n1235, n815);
xnor g1606 (n1564, n831, n671, n1225, n1198);
or   g1607 (n1431, n1213, n834, n736, n1242);
nand g1608 (n1501, n1331, n739, n699, n797);
nor  g1609 (n1661, n750, n806, n678, n1221);
xor  g1610 (n1396, n796, n1303, n1219, n780);
or   g1611 (n1376, n1302, n1342, n1308, n1255);
xnor g1612 (n1512, n1338, n1220, n742, n1361);
xor  g1613 (n1394, n1233, n1226, n794, n1299);
xnor g1614 (n1362, n1299, n758, n761, n702);
xor  g1615 (n1456, n677, n1308, n799, n1333);
and  g1616 (n1613, n741, n1241, n1192, n794);
xnor g1617 (n1379, n750, n783, n1209, n1320);
xnor g1618 (n1720, n753, n1308, n743, n1254);
or   g1619 (n1384, n1319, n728, n708, n1303);
xor  g1620 (n1572, n698, n1277, n823, n709);
xor  g1621 (n1386, n659, n1276, n706, n1327);
or   g1622 (n1523, n1211, n747, n1261, n1240);
xnor g1623 (n1625, n1311, n1195, n1334, n763);
xor  g1624 (n1557, n1307, n761, n1289, n677);
nand g1625 (n1580, n699, n718, n801, n1247);
xor  g1626 (n1628, n750, n1208, n789, n1285);
or   g1627 (n1490, n662, n1260, n760, n706);
nand g1628 (n1480, n812, n828, n1197, n780);
and  g1629 (n1636, n1196, n726, n759, n837);
or   g1630 (n1537, n1296, n984, n792, n763);
xnor g1631 (n1725, n716, n1283, n1328, n804);
xor  g1632 (n1515, n741, n1332, n720, n1359);
or   g1633 (n1454, n836, n763, n835, n670);
xnor g1634 (n1433, n655, n1192, n772, n1231);
xor  g1635 (n1715, n732, n696, n1252);
and  g1636 (n1541, n679, n749, n1349, n1278);
xor  g1637 (n1390, n837, n771, n749, n488);
nor  g1638 (n1453, n799, n1249, n1350, n1281);
xor  g1639 (n1441, n1229, n778, n1324, n1203);
or   g1640 (n1401, n773, n1241, n791, n1191);
nand g1641 (n1374, n1301, n1255, n1236, n814);
or   g1642 (n1400, n776, n657, n1351, n1255);
nand g1643 (n1468, n755, n773, n1269, n729);
nor  g1644 (n1600, n818, n1282, n762, n1201);
nand g1645 (n1732, n740, n826, n1302, n707);
xnor g1646 (n1465, n1325, n731, n834, n822);
nor  g1647 (n1692, n687, n1228, n783, n1268);
or   g1648 (n1550, n1275, n1327, n836, n1232);
nand g1649 (n1443, n762, n1333, n1196, n818);
xnor g1650 (n1653, n1193, n1315, n1267, n1295);
nor  g1651 (n1624, n656, n1256, n834, n780);
or   g1652 (n1516, n799, n1311, n1334, n727);
or   g1653 (n1552, n702, n755, n703, n1286);
xor  g1654 (n1671, n725, n833, n1205, n711);
xnor g1655 (n1380, n1323, n1344, n1263, n1350);
nand g1656 (n1504, n774, n739, n1315, n1328);
xnor g1657 (n1449, n748, n1224, n1220, n1287);
nand g1658 (n1513, n710, n1325, n1347, n816);
xnor g1659 (n1432, n1340, n665, n1314, n770);
nor  g1660 (n1419, n1231, n795, n489, n807);
xor  g1661 (n1622, n1280, n839, n744, n659);
nand g1662 (n1368, n693, n1205, n815, n826);
xor  g1663 (n1388, n1244, n798, n715, n691);
xor  g1664 (n1524, n1203, n709, n1248, n1297);
xnor g1665 (n1372, n1346, n1294, n1235, n673);
nand g1666 (n1709, n737, n730, n1321, n654);
and  g1667 (n1706, n839, n659, n1349, n723);
or   g1668 (n1678, n1284, n1199, n1203, n1286);
nand g1669 (n1632, n718, n1285, n1287, n1244);
nand g1670 (n1673, n1224, n678, n830, n1282);
xor  g1671 (n1563, n1286, n660, n1186, n1321);
or   g1672 (n1505, n791, n1287, n1338, n1305);
xnor g1673 (n1423, n1329, n835, n1258, n771);
xnor g1674 (n1642, n1325, n653, n824, n1248);
or   g1675 (n1387, n835, n1191, n1288, n690);
xor  g1676 (n1442, n1224, n1332, n744, n785);
and  g1677 (n1498, n1188, n1294, n710, n807);
xnor g1678 (n1381, n795, n1240, n677, n1231);
and  g1679 (n1582, n778, n1196, n1217);
nor  g1680 (n1497, n730, n1310, n805, n768);
or   g1681 (n1477, n695, n674, n489, n711);
xnor g1682 (n1702, n1187, n833, n752, n1357);
xor  g1683 (n1549, n663, n660, n1236, n1277);
xnor g1684 (n1712, n714, n1201, n810, n786);
xnor g1685 (n1459, n1212, n721, n1332, n808);
nand g1686 (n1567, n1201, n735, n721, n1311);
or   g1687 (n1508, n838, n707, n675, n705);
xor  g1688 (n1611, n759, n1337, n654, n722);
nand g1689 (n1685, n1213, n1199, n696, n1282);
or   g1690 (n1363, n733, n1274, n819, n1266);
nor  g1691 (n1434, n1215, n1239, n1302, n672);
xnor g1692 (n1662, n708, n1304, n826, n1294);
nor  g1693 (n1373, n667, n1225, n787, n803);
xnor g1694 (n1518, n1219, n810, n724, n754);
xnor g1695 (n1641, n738, n1193, n1348, n1312);
xor  g1696 (n1651, n1254, n1312, n690, n746);
nor  g1697 (n1457, n1308, n735, n1222, n1248);
or   g1698 (n1617, n1199, n732, n822, n672);
and  g1699 (n1462, n1193, n1350, n1260, n1297);
nor  g1700 (n1469, n727, n1186, n1232, n713);
or   g1701 (n1599, n841, n1234, n1275, n807);
xnor g1702 (n1901, n1721, n1545, n1553, n1717);
nand g1703 (n1891, n1638, n1501, n1632, n1424);
nand g1704 (n1831, n1394, n1660, n1435, n1649);
nand g1705 (n1922, n1630, n1664, n1556, n1384);
xor  g1706 (n1929, n1730, n1622, n1665, n1643);
nand g1707 (n1907, n1674, n1632, n1424, n1543);
nor  g1708 (n1939, n1633, n1451, n1453, n1720);
xor  g1709 (n1777, n1492, n1416, n1641, n1387);
nand g1710 (n1743, n1418, n1579, n1440, n1386);
xnor g1711 (n1747, n1500, n1619, n148, n1493);
and  g1712 (n1857, n1515, n1410, n1507, n1477);
nand g1713 (n1832, n1487, n1460, n1596, n1591);
or   g1714 (n1790, n1636, n1372, n1590, n1415);
or   g1715 (n1821, n1698, n1418, n1400, n1438);
or   g1716 (n1896, n1557, n1587, n1699, n1459);
xnor g1717 (n1823, n1550, n1584, n1512, n1399);
xor  g1718 (n1859, n1386, n1598, n1649, n1609);
xor  g1719 (n1841, n1643, n1366, n1499, n1635);
nand g1720 (n1925, n1458, n1396, n1522, n1619);
nor  g1721 (n1858, n1678, n1701, n1415, n1516);
nor  g1722 (n1885, n1363, n1669, n1454, n1492);
or   g1723 (n1931, n1373, n1392, n1696, n1442);
or   g1724 (n1883, n1677, n1365, n1595, n1490);
or   g1725 (n1869, n1711, n1661, n1589, n1726);
nor  g1726 (n1873, n1468, n1497, n1607, n1517);
nor  g1727 (n1765, n1568, n1731, n1684, n1608);
and  g1728 (n1872, n1700, n1476, n1363, n1527);
nand g1729 (n1795, n1687, n1521, n1395, n1462);
nand g1730 (n1906, n1378, n1484, n1623, n1503);
or   g1731 (n1825, n1715, n1392, n1618, n1641);
and  g1732 (n1888, n1729, n1449, n1557, n1486);
xor  g1733 (n1882, n1441, n1388, n1685, n1372);
xor  g1734 (n1877, n1729, n1601, n1597, n1697);
xnor g1735 (n1932, n1672, n1465, n1376, n1658);
and  g1736 (n1820, n1611, n1429, n1455, n1644);
xnor g1737 (n1785, n1514, n1651, n1606, n1555);
nand g1738 (n1921, n1369, n1627, n1658, n1642);
xor  g1739 (n1833, n1437, n1634, n1534, n1652);
and  g1740 (n1917, n1645, n1670, n1380, n1639);
or   g1741 (n1770, n1620, n1434, n1382, n1423);
or   g1742 (n1934, n1460, n1605, n1681, n1524);
xnor g1743 (n1937, n1693, n1399, n1649, n1527);
and  g1744 (n1861, n1693, n1576, n1701, n1385);
or   g1745 (n1766, n1447, n1463, n1488, n1600);
nor  g1746 (n1864, n1519, n1398, n1544, n1564);
nand g1747 (n1830, n1474, n1521, n1431, n1432);
xor  g1748 (n1868, n1540, n1725, n1549, n1525);
xor  g1749 (n1920, n1433, n1570, n1412, n1502);
or   g1750 (n1912, n1439, n1713, n1539, n1663);
or   g1751 (n1769, n1678, n1377, n1592, n1468);
nor  g1752 (n1783, n1593, n1715, n1532, n1498);
xnor g1753 (n1893, n1510, n1518, n1708, n1678);
xnor g1754 (n1835, n1421, n1669, n1504, n1637);
or   g1755 (n1918, n1600, n1438, n1572, n1554);
and  g1756 (n1749, n1490, n1587, n1531, n1564);
and  g1757 (n1737, n1469, n1730, n1461, n1725);
or   g1758 (n1863, n1670, n1730, n1709, n1429);
xor  g1759 (n1940, n1463, n1441, n1653, n1425);
nor  g1760 (n1881, n1481, n1727, n1596, n1419);
or   g1761 (n1806, n1406, n1411, n1627, n1696);
nand g1762 (n1875, n1494, n1543, n1544, n1698);
xor  g1763 (n1776, n1548, n1456, n1417, n1554);
xor  g1764 (n1812, n1546, n1653, n1471, n1639);
xor  g1765 (n1780, n1542, n1512, n1686, n1690);
nand g1766 (n1816, n1571, n1484, n1476, n1560);
xnor g1767 (n1928, n1452, n1407, n1640, n1657);
or   g1768 (n1764, n1691, n1598, n1647, n1398);
or   g1769 (n1930, n1673, n1660, n1653, n1644);
xnor g1770 (n1786, n1538, n1668, n1594, n1676);
and  g1771 (n1935, n1505, n1532, n1546, n1537);
xor  g1772 (n1916, n1690, n1621, n1614, n1535);
nor  g1773 (n1754, n1648, n1426, n1697, n1671);
xor  g1774 (n1814, n1613, n1378, n1430, n1731);
nand g1775 (n1760, n1699, n1401, n1466, n1505);
or   g1776 (n1767, n1573, n1622, n1663, n1448);
nand g1777 (n1839, n1394, n1533, n1615, n1497);
xor  g1778 (n1779, n1475, n1461, n1584, n1482);
xor  g1779 (n1902, n1666, n1448, n1602, n1705);
or   g1780 (n1889, n1721, n1561, n1666, n1665);
nor  g1781 (n1746, n1577, n1430, n1595, n1605);
and  g1782 (n1851, n1530, n1582, n1370, n1520);
or   g1783 (n1813, n1526, n1703, n1674, n1523);
xor  g1784 (n1761, n1650, n1624, n1694, n1464);
xnor g1785 (n1897, n1691, n1621, n1562, n1609);
and  g1786 (n1850, n1513, n1422, n1580, n1453);
nand g1787 (n1910, n1528, n1408, n1610, n1680);
xor  g1788 (n1755, n1370, n1716, n1379);
xnor g1789 (n1871, n1633, n1411, n1642, n1625);
and  g1790 (n1890, n1570, n1679, n1626, n1648);
xnor g1791 (n1810, n1723, n1433, n1722, n1443);
xnor g1792 (n1900, n1599, n1593, n1470, n1629);
xnor g1793 (n1750, n1671, n1390, n1432, n1391);
nand g1794 (n1852, n1726, n1585, n1385, n1685);
nand g1795 (n1738, n1393, n1673, n1575, n1531);
or   g1796 (n1751, n1727, n1686, n1585, n1575);
nor  g1797 (n1775, n1533, n1455, n1501, n1526);
nand g1798 (n1778, n1374, n1643, n1634, n1608);
or   g1799 (n1845, n1603, n1637, n1467, n1402);
nor  g1800 (n1919, n1661, n1620, n1555, n1566);
nand g1801 (n1848, n1508, n1683, n1402, n1631);
or   g1802 (n1745, n1556, n1642, n1450, n1569);
and  g1803 (n1854, n1458, n1442, n1732, n1590);
nand g1804 (n1809, n1478, n1657, n1517, n1494);
xnor g1805 (n1791, n1695, n1375, n1405, n1439);
nand g1806 (n1773, n1698, n1446, n1478, n1450);
and  g1807 (n1846, n1654, n1679, n1423, n1387);
nor  g1808 (n1826, n1686, n1616, n1567, n1664);
xnor g1809 (n1894, n1718, n1537, n1528, n1367);
nand g1810 (n1739, n1727, n1507, n1456, n1731);
xor  g1811 (n1899, n1647, n1539, n1547, n1617);
xor  g1812 (n1753, n1656, n1702, n1565, n1722);
nor  g1813 (n1886, n1706, n1662, n1612, n1444);
nor  g1814 (n1815, n1413, n1583, n1700, n1524);
xor  g1815 (n1879, n1541, n1445, n1364, n1707);
xor  g1816 (n1756, n1371, n1683, n1519, n1389);
or   g1817 (n1774, n1631, n1676, n1691, n1396);
nand g1818 (n1834, n1467, n1509, n1733, n1431);
or   g1819 (n1862, n1628, n1655, n1509, n1495);
nor  g1820 (n1838, n1688, n1713, n1413, n1664);
or   g1821 (n1926, n1578, n1707, n1724, n1733);
or   g1822 (n1874, n1583, n1542, n1475, n1651);
xnor g1823 (n1741, n1452, n1669, n1503, n1723);
and  g1824 (n1803, n1706, n1491, n1551, n1661);
xor  g1825 (n1938, n1485, n1606, n1684, n1734);
or   g1826 (n1849, n1639, n1474, n1709, n1529);
xnor g1827 (n1933, n1658, n1485, n1719, n1705);
xnor g1828 (n1805, n1690, n1558, n1692, n1728);
xor  g1829 (n1837, n1733, n1373, n1689, n1688);
nor  g1830 (n1911, n1426, n1561, n1487, n1685);
xor  g1831 (n1811, n1479, n1362, n1414, n1705);
xor  g1832 (n1742, n1592, n937, n1529, n1571);
and  g1833 (n1772, n1435, n1672, n1550, n1563);
nand g1834 (n1793, n1405, n1629, n1486, n1628);
nor  g1835 (n1818, n1607, n1420, n1572, n1688);
or   g1836 (n1822, n1717, n1687, n1397, n1470);
nand g1837 (n1752, n1708, n1651, n1623, n1511);
and  g1838 (n1909, n1383, n1672, n1696, n1367);
and  g1839 (n1903, n1481, n1580, n1417, n1626);
xnor g1840 (n1799, n1680, n1675, n1559, n1654);
xnor g1841 (n1904, n1506, n1703, n1719, n1720);
or   g1842 (n1927, n1601, n1428, n1650, n1454);
xnor g1843 (n1840, n1712, n1469, n1710, n1728);
xor  g1844 (n1807, n1662, n1711, n1582, n1420);
nand g1845 (n1788, n1638, n1610, n1404, n1687);
nor  g1846 (n1943, n1547, n1446, n1704, n1694);
or   g1847 (n1853, n1641, n1617, n1545, n1440);
xor  g1848 (n1876, n1701, n1520, n1702, n1562);
xor  g1849 (n1923, n1668, n1573, n1489, n1436);
xor  g1850 (n1844, n1732, n1675, n1574, n1551);
xor  g1851 (n1787, n1568, n1714, n1578, n1389);
or   g1852 (n1798, n1612, n1427, n1722, n1645);
or   g1853 (n1794, n1491, n1714, n1436, n1449);
and  g1854 (n1781, n1563, n1704, n1522, n1644);
xnor g1855 (n1792, n1381, n1383, n1646, n1483);
xor  g1856 (n1836, n1496, n1660, n1703, n1376);
and  g1857 (n1842, n1699, n1422, n1530, n1707);
xor  g1858 (n1913, n1684, n1498, n1393, n1419);
and  g1859 (n1796, n1591, n1566, n1719, n1510);
nor  g1860 (n1887, n1677, n1645, n1680, n1514);
xor  g1861 (n1736, n1710, n1427, n1683, n1681);
xor  g1862 (n1915, n1525, n1368, n1364, n1715);
xor  g1863 (n1941, n147, n1692, n1388, n1451);
nor  g1864 (n1735, n1586, n1709, n1681, n1700);
and  g1865 (n1829, n1716, n1473, n1695, n1708);
and  g1866 (n1784, n1535, n1734, n1613, n1671);
and  g1867 (n1768, n1506, n1380, n1630, n1362);
xor  g1868 (n1936, n1720, n1552, n1646, n1724);
and  g1869 (n1867, n1646, n1656, n1712, n1473);
xnor g1870 (n1797, n1553, n1508, n1636, n1504);
nor  g1871 (n1771, n1513, n1523, n1710, n1511);
nor  g1872 (n1945, n1594, n1689, n1447, n1377);
xor  g1873 (n1880, n1652, n1403, n1589, n1410);
nor  g1874 (n1740, n1647, n1697, n1721, n1657);
xor  g1875 (n1944, n1640, n1462, n1464, n1725);
nand g1876 (n1748, n1637, n1611, n1712, n1635);
nor  g1877 (n1924, n1650, n1665, n1471, n1540);
xnor g1878 (n1870, n1662, n1673, n1412, n1401);
nor  g1879 (n1800, n1659, n1404, n1729, n1586);
and  g1880 (n1801, n1604, n1579, n1444, n1655);
xnor g1881 (n1855, n1384, n1655, n1652, n1569);
nor  g1882 (n1819, n1407, n1479, n1574, n1567);
and  g1883 (n1824, n1483, n1616, n148, n1718);
nor  g1884 (n1762, n1654, n1638, n1443, n1682);
and  g1885 (n1757, n1603, n1472, n1576, n1552);
and  g1886 (n1843, n1714, n1706, n1676, n1499);
xor  g1887 (n1860, n1548, n1732, n1488, n1711);
nor  g1888 (n1856, n1395, n1675, n1391, n1480);
and  g1889 (n1942, n1482, n1472, n1400, n1693);
or   g1890 (n1828, n1434, n1480, n1581);
nand g1891 (n1895, n1397, n1659, n1489, n1677);
xnor g1892 (n1865, n1445, n1718, n1602, n1694);
xnor g1893 (n1808, n1559, n1409, n1667, n1516);
nor  g1894 (n1789, n1428, n1459, n1382, n1536);
and  g1895 (n1905, n1663, n1541, n1577, n1495);
nor  g1896 (n1763, n1375, n1534, n1403, n1648);
and  g1897 (n1866, n1502, n1549, n1695, n1518);
and  g1898 (n1892, n1437, n1659, n1416, n1724);
nand g1899 (n1946, n1682, n147, n1666, n1565);
or   g1900 (n1744, n1366, n1728, n1515, n1618);
nand g1901 (n1759, n1682, n1624, n1406, n1702);
xor  g1902 (n1908, n1667, n1692, n1689, n1538);
and  g1903 (n1782, n1599, n1408, n1588, n1381);
and  g1904 (n1847, n1558, n1704, n1425, n1604);
xnor g1905 (n1804, n1597, n1588, n1457, n1496);
nand g1906 (n1827, n1614, n1466, n1723, n1379);
or   g1907 (n1914, n1368, n1560, n1500, n1409);
nand g1908 (n1758, n1625, n1726, n1713, n1457);
xnor g1909 (n1884, n1674, n1615, n1365, n1493);
nand g1910 (n1817, n1421, n1465, n1679, n1390);
and  g1911 (n1802, n1656, n1374, n1668, n1670);
xnor g1912 (n1898, n1667, n1371, n1717, n1414);
xnor g1913 (n1878, n1369, n1536, n1477, n1640);
nor  g1914 (n1962, n1774, n1736);
nand g1915 (n1952, n1765, n1773, n1748, n1789);
and  g1916 (n1957, n1794, n1762, n1788, n1784);
nand g1917 (n1955, n1780, n1778, n1792, n1783);
xnor g1918 (n1958, n1777, n1735, n1745, n1766);
nand g1919 (n1953, n1739, n1767, n1781, n1772);
xnor g1920 (n1959, n1790, n1741, n1787, n1760);
nand g1921 (n1954, n1779, n1768, n1743, n1755);
and  g1922 (n1947, n1749, n1763, n1756, n1795);
nor  g1923 (n1956, n1737, n1770, n1751, n1791);
xnor g1924 (n1950, n1793, n1744, n1771, n1776);
nand g1925 (n1951, n1764, n1769, n1786, n1747);
xor  g1926 (n1961, n1758, n1738, n1742, n1757);
xnor g1927 (n1960, n1759, n1746, n1752, n1754);
xnor g1928 (n1949, n1761, n1796, n1785, n1740);
nor  g1929 (n1948, n1782, n1750, n1753, n1775);
and  g1930 (n1971, n1894, n1812, n1961, n1841);
xor  g1931 (n2008, n1959, n1958, n1940);
and  g1932 (n1963, n1844, n1955, n1822, n1905);
nand g1933 (n1989, n1956, n1957, n1814, n32);
nor  g1934 (n1997, n1874, n1823, n1956, n1961);
nor  g1935 (n2000, n1926, n1940, n1939, n1924);
nor  g1936 (n1984, n1886, n1847, n1951, n1911);
nand g1937 (n1992, n1956, n1831, n1888, n1959);
xnor g1938 (n1968, n1914, n1806, n1908, n1933);
xor  g1939 (n1973, n1931, n1798, n1856, n1862);
nor  g1940 (n1974, n1954, n1938, n1951, n1960);
or   g1941 (n1996, n1945, n1827, n1901, n1937);
and  g1942 (n1980, n1870, n1896, n1839, n32);
nand g1943 (n1981, n1849, n1953, n1734, n1958);
or   g1944 (n2013, n1962, n1957, n1951, n148);
xnor g1945 (n2002, n1880, n1962, n1939, n1868);
nand g1946 (n1977, n1900, n1799, n1819, n1854);
or   g1947 (n2007, n1941, n1800, n1953, n1928);
or   g1948 (n1969, n31, n1950, n1804, n1955);
nor  g1949 (n1976, n1865, n1957, n1930, n1892);
xnor g1950 (n2018, n1863, n31, n1871, n1867);
or   g1951 (n2017, n1866, n1912, n1801, n1835);
or   g1952 (n2012, n1815, n1920, n1813, n1953);
xnor g1953 (n1965, n1932, n1950, n1942, n1952);
nand g1954 (n1988, n1898, n1845, n1927, n1837);
or   g1955 (n1986, n1954, n1936, n1913, n1891);
xor  g1956 (n2001, n1873, n1949, n1848, n1842);
xnor g1957 (n1998, n32, n1959, n1952, n1948);
xnor g1958 (n2006, n1950, n1910, n1917, n1810);
or   g1959 (n1987, n1805, n1923, n1859, n32);
xor  g1960 (n2004, n1944, n1952, n1828, n1878);
nor  g1961 (n1970, n1961, n1958, n1904, n1885);
xor  g1962 (n2009, n1941, n1889, n1851, n1949);
nor  g1963 (n1979, n1960, n1809, n1834, n1943);
xor  g1964 (n1978, n1949, n1853, n1893, n1852);
xor  g1965 (n2010, n148, n1947, n31, n1820);
nor  g1966 (n1985, n1925, n1816, n1959, n1869);
nand g1967 (n1983, n1843, n1846, n1922, n1811);
nor  g1968 (n2003, n1947, n1855, n1955, n1879);
xor  g1969 (n1975, n1946, n1954, n1919);
xor  g1970 (n1972, n1961, n1836, n1887, n1877);
xor  g1971 (n2005, n1860, n1817, n1829, n1909);
xor  g1972 (n1991, n1872, n1882, n1883, n1915);
xor  g1973 (n1982, n1861, n1962, n1832, n1956);
and  g1974 (n1990, n1942, n1876, n1934, n1826);
and  g1975 (n2011, n1962, n1825, n1821, n1857);
or   g1976 (n2014, n1875, n1858, n1921, n1797);
or   g1977 (n2016, n1960, n1895, n1808, n1902);
nand g1978 (n1964, n1803, n1944, n1864, n1903);
or   g1979 (n1993, n1906, n1929, n1918, n1960);
or   g1980 (n1966, n1884, n1943, n1840, n1890);
and  g1981 (n2015, n1907, n1850, n1802, n1838);
nor  g1982 (n1967, n1948, n1833, n1946, n1935);
and  g1983 (n1994, n1916, n1945, n1948, n1957);
xnor g1984 (n1999, n1807, n1955, n1830, n1897);
xor  g1985 (n1995, n1824, n1881, n1899, n1818);
xnor g1986 (n2032, n1996, n2004, n2017, n1973);
xor  g1987 (n2019, n2007, n2008, n1989, n1991);
nand g1988 (n2029, n1966, n1987, n1975, n1985);
nor  g1989 (n2025, n1971, n2012, n2003, n1992);
xor  g1990 (n2027, n2000, n1969, n2016, n2002);
nor  g1991 (n2020, n2013, n1983, n1986, n2005);
or   g1992 (n2030, n1984, n1974, n1978, n2001);
nand g1993 (n2021, n2009, n1993, n1964, n1970);
nor  g1994 (n2022, n1980, n1994, n1995, n2011);
xnor g1995 (n2028, n1967, n1972, n2014, n2015);
nor  g1996 (n2026, n1968, n1997, n1981, n1965);
nor  g1997 (n2023, n1979, n1998, n1976, n1977);
or   g1998 (n2024, n2010, n1990, n1988, n2018);
nand g1999 (n2031, n2006, n1982, n1963, n1999);
endmodule
