

module Stat_128_636
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n144,
  n135,
  n134,
  n129,
  n126,
  n147,
  n138,
  n136,
  n139,
  n140,
  n125,
  n137,
  n146,
  n142,
  n132,
  n127,
  n130,
  n143,
  n145,
  n133,
  n141,
  n148,
  n131,
  n128
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n144;output n135;output n134;output n129;output n126;output n147;output n138;output n136;output n139;output n140;output n125;output n137;output n146;output n142;output n132;output n127;output n130;output n143;output n145;output n133;output n141;output n148;output n131;output n128;
  wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    KeyWire_0_11,
    n2
  );


  buf
  g1
  (
    n25,
    n3
  );


  not
  g2
  (
    KeyWire_0_16,
    n1
  );


  buf
  g3
  (
    KeyWire_0_63,
    n4
  );


  buf
  g4
  (
    n23,
    n2
  );


  not
  g5
  (
    n22,
    n1
  );


  buf
  g6
  (
    KeyWire_0_29,
    n3
  );


  not
  g7
  (
    KeyWire_0_0,
    n27
  );


  buf
  g8
  (
    KeyWire_0_42,
    n21
  );


  buf
  g9
  (
    n32,
    n22
  );


  buf
  g10
  (
    n47,
    n25
  );


  buf
  g11
  (
    KeyWire_0_4,
    n25
  );


  buf
  g12
  (
    KeyWire_0_59,
    n24
  );


  not
  g13
  (
    KeyWire_0_28,
    n26
  );


  not
  g14
  (
    KeyWire_0_58,
    n22
  );


  not
  g15
  (
    n33,
    n22
  );


  not
  g16
  (
    n38,
    n24
  );


  not
  g17
  (
    n35,
    n26
  );


  buf
  g18
  (
    KeyWire_0_49,
    n27
  );


  not
  g19
  (
    n28,
    n27
  );


  buf
  g20
  (
    n52,
    n26
  );


  not
  g21
  (
    KeyWire_0_51,
    n25
  );


  not
  g22
  (
    KeyWire_0_40,
    n25
  );


  not
  g23
  (
    n42,
    n23
  );


  not
  g24
  (
    KeyWire_0_2,
    n26
  );


  buf
  g25
  (
    n37,
    n24
  );


  buf
  g26
  (
    KeyWire_0_36,
    n21
  );


  buf
  g27
  (
    n36,
    n24
  );


  buf
  g28
  (
    KeyWire_0_1,
    n21
  );


  not
  g29
  (
    n39,
    n23
  );


  not
  g30
  (
    KeyWire_0_12,
    n21
  );


  buf
  g31
  (
    n40,
    n23
  );


  not
  g32
  (
    n54,
    n23
  );


  not
  g33
  (
    n53,
    n22
  );


  not
  g34
  (
    KeyWire_0_15,
    n18
  );


  buf
  g35
  (
    KeyWire_0_54,
    n6
  );


  not
  g36
  (
    KeyWire_0_38,
    n41
  );


  buf
  g37
  (
    KeyWire_0_41,
    n39
  );


  not
  g38
  (
    n61,
    n44
  );


  not
  g39
  (
    KeyWire_0_22,
    n6
  );


  not
  g40
  (
    n82,
    n14
  );


  buf
  g41
  (
    n59,
    n43
  );


  buf
  g42
  (
    KeyWire_0_37,
    n37
  );


  buf
  g43
  (
    KeyWire_0_55,
    n15
  );


  not
  g44
  (
    n68,
    n40
  );


  buf
  g45
  (
    n76,
    n42
  );


  not
  g46
  (
    KeyWire_0_34,
    n13
  );


  buf
  g47
  (
    KeyWire_0_56,
    n41
  );


  not
  g48
  (
    KeyWire_0_17,
    n33
  );


  not
  g49
  (
    n100,
    n29
  );


  not
  g50
  (
    KeyWire_0_13,
    n36
  );


  buf
  g51
  (
    n74,
    n33
  );


  not
  g52
  (
    n99,
    n11
  );


  buf
  g53
  (
    n86,
    n38
  );


  buf
  g54
  (
    KeyWire_0_44,
    n18
  );


  buf
  g55
  (
    KeyWire_0_24,
    n28
  );


  nand
  g56
  (
    KeyWire_0_27,
    n5,
    n31,
    n36
  );


  nand
  g57
  (
    n95,
    n35,
    n32,
    n31,
    n14
  );


  nor
  g58
  (
    n85,
    n19,
    n17,
    n20,
    n13
  );


  xor
  g59
  (
    n102,
    n47,
    n29,
    n39,
    n35
  );


  xor
  g60
  (
    KeyWire_0_18,
    n19,
    n42,
    n28,
    n46
  );


  nor
  g61
  (
    n84,
    n48,
    n10,
    n40,
    n39
  );


  nor
  g62
  (
    n90,
    n34,
    n37,
    n45,
    n42
  );


  nand
  g63
  (
    n94,
    n11,
    n29,
    n12,
    n30
  );


  nand
  g64
  (
    KeyWire_0_30,
    n35,
    n34,
    n20,
    n33
  );


  nor
  g65
  (
    KeyWire_0_5,
    n16,
    n46,
    n32,
    n13
  );


  nor
  g66
  (
    KeyWire_0_35,
    n18,
    n11,
    n43,
    n19
  );


  and
  g67
  (
    KeyWire_0_46,
    n43,
    n20,
    n34,
    n9
  );


  xor
  g68
  (
    KeyWire_0_7,
    n17,
    n15,
    n16,
    n31
  );


  or
  g69
  (
    KeyWire_0_61,
    n10,
    n12,
    n7,
    n17
  );


  and
  g70
  (
    KeyWire_0_10,
    n14,
    n36,
    n37,
    n43
  );


  or
  g71
  (
    n93,
    n8,
    n45,
    n35
  );


  xnor
  g72
  (
    n77,
    n20,
    n10,
    n41,
    n44
  );


  and
  g73
  (
    n87,
    n17,
    n28,
    n44,
    n46
  );


  and
  g74
  (
    n97,
    n39,
    n15,
    n47,
    n13
  );


  or
  g75
  (
    n72,
    n48,
    n29,
    n47,
    n30
  );


  nand
  g76
  (
    n56,
    n12,
    n34,
    n28,
    n41
  );


  nand
  g77
  (
    KeyWire_0_53,
    n31,
    n8,
    n14,
    n5
  );


  or
  g78
  (
    n67,
    n33,
    n46,
    n10,
    n36
  );


  nand
  g79
  (
    n104,
    n7,
    n40,
    n16,
    n19
  );


  xnor
  g80
  (
    n75,
    n45,
    n18,
    n32,
    n4
  );


  xnor
  g81
  (
    KeyWire_0_43,
    n40,
    n38,
    n37,
    n11
  );


  xnor
  g82
  (
    KeyWire_0_21,
    n12,
    n16,
    n30,
    n42
  );


  nor
  g83
  (
    n60,
    n47,
    n38,
    n30
  );


  nor
  g84
  (
    KeyWire_0_62,
    n15,
    n9,
    n32,
    n44
  );


  xor
  g85
  (
    KeyWire_0_39,
    n62,
    n57,
    n63,
    n64
  );


  or
  g86
  (
    n107,
    n59,
    n66,
    n56,
    n61
  );


  xor
  g87
  (
    n112,
    n65,
    n60,
    n66,
    n67
  );


  xor
  g88
  (
    n109,
    n58,
    n60,
    n65,
    n55
  );


  xor
  g89
  (
    KeyWire_0_14,
    n57,
    n62,
    n63,
    n59
  );


  xor
  g90
  (
    n106,
    n67,
    n27,
    n68
  );


  nor
  g91
  (
    n111,
    n58,
    n64,
    n56,
    n61
  );


  and
  g92
  (
    KeyWire_0_60,
    n73,
    n52,
    n109,
    n53
  );


  or
  g93
  (
    n119,
    n108,
    n50,
    n72,
    n71
  );


  or
  g94
  (
    n113,
    n49,
    n110,
    n71,
    n112
  );


  xor
  g95
  (
    n114,
    n54,
    n111,
    n69
  );


  nand
  g96
  (
    KeyWire_0_32,
    n51,
    n50,
    n49,
    n112
  );


  nand
  g97
  (
    n118,
    n69,
    n54,
    n109
  );


  and
  g98
  (
    KeyWire_0_57,
    n51,
    n51,
    n50,
    n52
  );


  or
  g99
  (
    n122,
    n73,
    n106,
    n52
  );


  or
  g100
  (
    n116,
    n72,
    n53,
    n70
  );


  xor
  g101
  (
    n123,
    n53,
    n48,
    n70
  );


  xor
  g102
  (
    KeyWire_0_20,
    n110,
    n50,
    n49
  );


  and
  g103
  (
    n121,
    n107,
    n108,
    n51,
    n54
  );


  xnor
  g104
  (
    KeyWire_0_26,
    n122,
    n82,
    n116,
    n93
  );


  nand
  g105
  (
    n141,
    n94,
    n93,
    n102,
    n75
  );


  nand
  g106
  (
    KeyWire_0_25,
    n105,
    n123,
    n82,
    n79
  );


  nor
  g107
  (
    KeyWire_0_9,
    n119,
    n118,
    n122,
    n124
  );


  or
  g108
  (
    n131,
    n115,
    n92,
    n90,
    n75
  );


  or
  g109
  (
    n138,
    n85,
    n84,
    n102,
    n78
  );


  nor
  g110
  (
    KeyWire_0_3,
    n83,
    n89,
    n74,
    n120
  );


  xor
  g111
  (
    n136,
    n105,
    n114,
    n85,
    n79
  );


  xor
  g112
  (
    KeyWire_0_19,
    n78,
    n101,
    n99,
    n94
  );


  nand
  g113
  (
    KeyWire_0_47,
    n102,
    n102,
    n77,
    n97
  );


  xor
  g114
  (
    KeyWire_0_45,
    n99,
    n89,
    n86,
    n123
  );


  nor
  g115
  (
    KeyWire_0_31,
    n81,
    n103,
    n105,
    n95
  );


  and
  g116
  (
    n134,
    n100,
    n83,
    n98,
    n116
  );


  nand
  g117
  (
    KeyWire_0_23,
    n114,
    n80,
    n103,
    n124
  );


  xor
  g118
  (
    n132,
    n96,
    n96,
    n119,
    n100
  );


  nand
  g119
  (
    n128,
    n117,
    n92,
    n86,
    n113
  );


  nand
  g120
  (
    KeyWire_0_50,
    n74,
    n76,
    n103,
    n95
  );


  and
  g121
  (
    KeyWire_0_48,
    n91,
    n77,
    n120,
    n115
  );


  and
  g122
  (
    n125,
    n121,
    n104
  );


  nand
  g123
  (
    n127,
    n81,
    n113,
    n117,
    n87
  );


  or
  g124
  (
    KeyWire_0_6,
    n84,
    n97,
    n118,
    n76
  );


  or
  g125
  (
    KeyWire_0_52,
    n101,
    n88,
    n104
  );


  xnor
  g126
  (
    KeyWire_0_8,
    n121,
    n103,
    n98,
    n105
  );


  or
  g127
  (
    KeyWire_0_33,
    n91,
    n87,
    n90,
    n80
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n41,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n44,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n48,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n145,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n31,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n88,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n137,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n103,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n144,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n148,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n81,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n24,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n45,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n65,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n110,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n80,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n27,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n83,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n101,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n129,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n117,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n57,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n64,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n126,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n92,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n130,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n147,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n89,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n34,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n26,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n71,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n133,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n120,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n139,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n70,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n63,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n46,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n79,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n69,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n108,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n43,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n91,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n49,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n96,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n78,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n142,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n98,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n146,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n135,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n29,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n143,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n50,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n140,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n55,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n62,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n58,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n66,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n115,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n51,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n30,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n124,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n73,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n105,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n21,
    KeyNOTWire_0_63
  );


endmodule


