

module Stat_1321_43_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n45,
  n46,
  n276,
  n274,
  n290,
  n291,
  n267,
  n289,
  n300,
  n265,
  n292,
  n249,
  n297,
  n250,
  n259,
  n264,
  n295,
  n252,
  n279,
  n287,
  n266,
  n261,
  n1042,
  n1188,
  n1193,
  n1196,
  n1189,
  n1191,
  n1186,
  n1194,
  n1187,
  n1195,
  n1220,
  n1251,
  n1237,
  n1235,
  n1244,
  n1333,
  n1335,
  n1337,
  n1336,
  n1334,
  n1366,
  n1367,
  n1365,
  n1364,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input n33;
  input n34;
  input n35;
  input n36;
  input n37;
  input n38;
  input n39;
  input n40;
  input n41;
  input n42;
  input n43;
  input n44;
  input n45;
  input n46;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n276;
  output n274;
  output n290;
  output n291;
  output n267;
  output n289;
  output n300;
  output n265;
  output n292;
  output n249;
  output n297;
  output n250;
  output n259;
  output n264;
  output n295;
  output n252;
  output n279;
  output n287;
  output n266;
  output n261;
  output n1042;
  output n1188;
  output n1193;
  output n1196;
  output n1189;
  output n1191;
  output n1186;
  output n1194;
  output n1187;
  output n1195;
  output n1220;
  output n1251;
  output n1237;
  output n1235;
  output n1244;
  output n1333;
  output n1335;
  output n1337;
  output n1336;
  output n1334;
  output n1366;
  output n1367;
  output n1365;
  output n1364;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n251;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n260;
  wire n262;
  wire n263;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n275;
  wire n277;
  wire n278;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n288;
  wire n293;
  wire n294;
  wire n296;
  wire n298;
  wire n299;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1190;
  wire n1192;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1236;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n96,
    n4
  );


  not
  g1
  (
    KeyWire_0_22,
    n44
  );


  not
  g2
  (
    n128,
    n45
  );


  not
  g3
  (
    n163,
    n37
  );


  buf
  g4
  (
    n196,
    n17
  );


  buf
  g5
  (
    KeyWire_0_56,
    n10
  );


  buf
  g6
  (
    n145,
    n42
  );


  not
  g7
  (
    n117,
    n42
  );


  buf
  g8
  (
    n175,
    n39
  );


  buf
  g9
  (
    n106,
    n14
  );


  buf
  g10
  (
    n164,
    n12
  );


  not
  g11
  (
    n72,
    n1
  );


  buf
  g12
  (
    n202,
    n40
  );


  not
  g13
  (
    n168,
    n30
  );


  not
  g14
  (
    n205,
    n46
  );


  buf
  g15
  (
    n148,
    n39
  );


  buf
  g16
  (
    n182,
    n37
  );


  not
  g17
  (
    n221,
    n26
  );


  buf
  g18
  (
    n55,
    n44
  );


  buf
  g19
  (
    n130,
    n41
  );


  buf
  g20
  (
    n170,
    n4
  );


  not
  g21
  (
    n50,
    n38
  );


  buf
  g22
  (
    n185,
    n14
  );


  buf
  g23
  (
    n198,
    n16
  );


  not
  g24
  (
    n71,
    n8
  );


  not
  g25
  (
    n153,
    n30
  );


  not
  g26
  (
    n85,
    n7
  );


  not
  g27
  (
    n216,
    n26
  );


  not
  g28
  (
    n102,
    n43
  );


  not
  g29
  (
    KeyWire_0_58,
    n9
  );


  buf
  g30
  (
    n220,
    n8
  );


  not
  g31
  (
    n162,
    n32
  );


  buf
  g32
  (
    n230,
    n5
  );


  buf
  g33
  (
    n118,
    n29
  );


  buf
  g34
  (
    n215,
    n31
  );


  not
  g35
  (
    n144,
    n45
  );


  buf
  g36
  (
    n94,
    n11
  );


  not
  g37
  (
    n136,
    n27
  );


  not
  g38
  (
    n60,
    n46
  );


  buf
  g39
  (
    n113,
    n23
  );


  buf
  g40
  (
    n222,
    n26
  );


  not
  g41
  (
    n138,
    n27
  );


  not
  g42
  (
    n83,
    n32
  );


  not
  g43
  (
    n169,
    n21
  );


  not
  g44
  (
    n171,
    n42
  );


  not
  g45
  (
    n193,
    n18
  );


  not
  g46
  (
    n149,
    n19
  );


  not
  g47
  (
    n166,
    n37
  );


  not
  g48
  (
    n223,
    n23
  );


  not
  g49
  (
    n165,
    n24
  );


  not
  g50
  (
    n57,
    n37
  );


  buf
  g51
  (
    n156,
    n35
  );


  not
  g52
  (
    n161,
    n6
  );


  buf
  g53
  (
    n172,
    n41
  );


  buf
  g54
  (
    n99,
    n40
  );


  not
  g55
  (
    n188,
    n3
  );


  not
  g56
  (
    n91,
    n12
  );


  not
  g57
  (
    n115,
    n27
  );


  buf
  g58
  (
    n181,
    n46
  );


  buf
  g59
  (
    n135,
    n24
  );


  buf
  g60
  (
    n108,
    n30
  );


  buf
  g61
  (
    n86,
    n20
  );


  buf
  g62
  (
    n200,
    n23
  );


  not
  g63
  (
    n183,
    n29
  );


  not
  g64
  (
    n167,
    n17
  );


  buf
  g65
  (
    n180,
    n19
  );


  not
  g66
  (
    n142,
    n22
  );


  not
  g67
  (
    n189,
    n21
  );


  buf
  g68
  (
    KeyWire_0_7,
    n35
  );


  not
  g69
  (
    n176,
    n25
  );


  buf
  g70
  (
    n93,
    n35
  );


  not
  g71
  (
    n174,
    n7
  );


  buf
  g72
  (
    n81,
    n18
  );


  not
  g73
  (
    n116,
    n3
  );


  not
  g74
  (
    n125,
    n34
  );


  buf
  g75
  (
    n203,
    n21
  );


  not
  g76
  (
    n208,
    n29
  );


  buf
  g77
  (
    n209,
    n24
  );


  buf
  g78
  (
    n173,
    n9
  );


  buf
  g79
  (
    n67,
    n28
  );


  buf
  g80
  (
    n110,
    n31
  );


  buf
  g81
  (
    n224,
    n34
  );


  buf
  g82
  (
    n62,
    n5
  );


  buf
  g83
  (
    n88,
    n18
  );


  buf
  g84
  (
    n132,
    n38
  );


  buf
  g85
  (
    n104,
    n40
  );


  buf
  g86
  (
    n139,
    n11
  );


  buf
  g87
  (
    n73,
    n13
  );


  not
  g88
  (
    n140,
    n2
  );


  buf
  g89
  (
    n141,
    n44
  );


  buf
  g90
  (
    n84,
    n10
  );


  not
  g91
  (
    n58,
    n6
  );


  not
  g92
  (
    n47,
    n12
  );


  not
  g93
  (
    n226,
    n19
  );


  not
  g94
  (
    n54,
    n42
  );


  not
  g95
  (
    n80,
    n40
  );


  buf
  g96
  (
    KeyWire_0_4,
    n31
  );


  not
  g97
  (
    n147,
    n8
  );


  buf
  g98
  (
    n127,
    n20
  );


  buf
  g99
  (
    n112,
    n46
  );


  buf
  g100
  (
    n61,
    n17
  );


  not
  g101
  (
    n69,
    n16
  );


  not
  g102
  (
    n56,
    n2
  );


  buf
  g103
  (
    n160,
    n44
  );


  buf
  g104
  (
    n66,
    n1
  );


  buf
  g105
  (
    n214,
    n15
  );


  not
  g106
  (
    n105,
    n16
  );


  buf
  g107
  (
    n70,
    n6
  );


  buf
  g108
  (
    n119,
    n33
  );


  buf
  g109
  (
    n100,
    n3
  );


  buf
  g110
  (
    n199,
    n10
  );


  buf
  g111
  (
    n122,
    n33
  );


  not
  g112
  (
    n228,
    n1
  );


  not
  g113
  (
    n103,
    n28
  );


  not
  g114
  (
    n129,
    n25
  );


  buf
  g115
  (
    n92,
    n34
  );


  not
  g116
  (
    n146,
    n36
  );


  buf
  g117
  (
    n109,
    n29
  );


  not
  g118
  (
    n89,
    n36
  );


  not
  g119
  (
    n229,
    n25
  );


  not
  g120
  (
    n178,
    n20
  );


  not
  g121
  (
    n78,
    n43
  );


  buf
  g122
  (
    n133,
    n15
  );


  buf
  g123
  (
    n213,
    n26
  );


  not
  g124
  (
    n225,
    n30
  );


  not
  g125
  (
    n211,
    n2
  );


  buf
  g126
  (
    n151,
    n36
  );


  buf
  g127
  (
    n97,
    n7
  );


  not
  g128
  (
    n48,
    n15
  );


  buf
  g129
  (
    n217,
    n36
  );


  not
  g130
  (
    n77,
    n14
  );


  not
  g131
  (
    n159,
    n4
  );


  buf
  g132
  (
    n64,
    n6
  );


  buf
  g133
  (
    n194,
    n8
  );


  not
  g134
  (
    KeyWire_0_45,
    n28
  );


  not
  g135
  (
    n204,
    n45
  );


  not
  g136
  (
    n177,
    n15
  );


  not
  g137
  (
    n131,
    n41
  );


  not
  g138
  (
    n201,
    n14
  );


  not
  g139
  (
    n187,
    n24
  );


  not
  g140
  (
    n158,
    n11
  );


  not
  g141
  (
    n120,
    n31
  );


  buf
  g142
  (
    n68,
    n33
  );


  buf
  g143
  (
    n49,
    n32
  );


  not
  g144
  (
    n210,
    n13
  );


  not
  g145
  (
    KeyWire_0_12,
    n9
  );


  buf
  g146
  (
    n90,
    n34
  );


  not
  g147
  (
    KeyWire_0_11,
    n43
  );


  buf
  g148
  (
    n101,
    n43
  );


  not
  g149
  (
    KeyWire_0_2,
    n9
  );


  not
  g150
  (
    n114,
    n5
  );


  buf
  g151
  (
    n111,
    n38
  );


  not
  g152
  (
    n79,
    n11
  );


  buf
  g153
  (
    n154,
    n5
  );


  buf
  g154
  (
    KeyWire_0_52,
    n22
  );


  buf
  g155
  (
    n206,
    n22
  );


  not
  g156
  (
    n190,
    n18
  );


  not
  g157
  (
    n150,
    n13
  );


  buf
  g158
  (
    n82,
    n4
  );


  buf
  g159
  (
    n124,
    n25
  );


  buf
  g160
  (
    n121,
    n2
  );


  not
  g161
  (
    n134,
    n39
  );


  buf
  g162
  (
    n74,
    n39
  );


  not
  g163
  (
    n143,
    n23
  );


  not
  g164
  (
    n219,
    n3
  );


  buf
  g165
  (
    n87,
    n35
  );


  not
  g166
  (
    n52,
    n22
  );


  not
  g167
  (
    n76,
    n32
  );


  not
  g168
  (
    n227,
    n33
  );


  buf
  g169
  (
    n126,
    n16
  );


  not
  g170
  (
    n197,
    n19
  );


  buf
  g171
  (
    n98,
    n12
  );


  not
  g172
  (
    n63,
    n17
  );


  not
  g173
  (
    n59,
    n10
  );


  not
  g174
  (
    n184,
    n20
  );


  buf
  g175
  (
    n218,
    n41
  );


  not
  g176
  (
    n186,
    n13
  );


  buf
  g177
  (
    n195,
    n27
  );


  not
  g178
  (
    n179,
    n1
  );


  not
  g179
  (
    KeyWire_0_13,
    n21
  );


  buf
  g180
  (
    n207,
    n28
  );


  buf
  g181
  (
    n157,
    n45
  );


  not
  g182
  (
    n152,
    n38
  );


  buf
  g183
  (
    n123,
    n7
  );


  buf
  g184
  (
    n231,
    n47
  );


  buf
  g185
  (
    n232,
    n48
  );


  not
  g186
  (
    n235,
    n47
  );


  buf
  g187
  (
    n234,
    n47
  );


  not
  g188
  (
    n233,
    n47
  );


  buf
  g189
  (
    n247,
    n233
  );


  not
  g190
  (
    n245,
    n234
  );


  not
  g191
  (
    n236,
    n231
  );


  not
  g192
  (
    n244,
    n233
  );


  buf
  g193
  (
    n241,
    n232
  );


  buf
  g194
  (
    n240,
    n231
  );


  not
  g195
  (
    n237,
    n231
  );


  not
  g196
  (
    n246,
    n233
  );


  not
  g197
  (
    n238,
    n232
  );


  buf
  g198
  (
    n243,
    n232
  );


  buf
  g199
  (
    n242,
    n232
  );


  not
  g200
  (
    n248,
    n231
  );


  buf
  g201
  (
    n239,
    n233
  );


  not
  g202
  (
    n282,
    n239
  );


  not
  g203
  (
    n259,
    n243
  );


  buf
  g204
  (
    n291,
    n243
  );


  not
  g205
  (
    n273,
    n247
  );


  buf
  g206
  (
    n289,
    n241
  );


  buf
  g207
  (
    n286,
    n241
  );


  not
  g208
  (
    n297,
    n238
  );


  not
  g209
  (
    n298,
    n238
  );


  not
  g210
  (
    n249,
    n244
  );


  buf
  g211
  (
    n284,
    n248
  );


  not
  g212
  (
    n283,
    n236
  );


  buf
  g213
  (
    n299,
    n242
  );


  buf
  g214
  (
    n280,
    n247
  );


  not
  g215
  (
    n296,
    n238
  );


  buf
  g216
  (
    n292,
    n245
  );


  not
  g217
  (
    KeyWire_0_53,
    n239
  );


  not
  g218
  (
    n253,
    n244
  );


  buf
  g219
  (
    n261,
    n241
  );


  buf
  g220
  (
    KeyWire_0_63,
    n242
  );


  buf
  g221
  (
    n295,
    n240
  );


  not
  g222
  (
    n290,
    n245
  );


  buf
  g223
  (
    KeyWire_0_46,
    n240
  );


  not
  g224
  (
    n260,
    n246
  );


  not
  g225
  (
    n285,
    n248
  );


  not
  g226
  (
    n277,
    n246
  );


  not
  g227
  (
    n274,
    n245
  );


  buf
  g228
  (
    n256,
    n243
  );


  buf
  g229
  (
    n255,
    n248
  );


  buf
  g230
  (
    n252,
    n244
  );


  buf
  g231
  (
    KeyWire_0_32,
    n244
  );


  not
  g232
  (
    n287,
    n248
  );


  buf
  g233
  (
    n276,
    n236
  );


  not
  g234
  (
    n263,
    n241
  );


  buf
  g235
  (
    n258,
    n236
  );


  not
  g236
  (
    n270,
    n240
  );


  not
  g237
  (
    n271,
    n243
  );


  buf
  g238
  (
    n293,
    n246
  );


  buf
  g239
  (
    n267,
    n240
  );


  not
  g240
  (
    n262,
    n237
  );


  buf
  g241
  (
    n279,
    n247
  );


  not
  g242
  (
    n257,
    n242
  );


  buf
  g243
  (
    n251,
    n242
  );


  buf
  g244
  (
    n281,
    n247
  );


  buf
  g245
  (
    n268,
    n237
  );


  buf
  g246
  (
    n250,
    n237
  );


  not
  g247
  (
    n288,
    n236
  );


  buf
  g248
  (
    n300,
    n238
  );


  buf
  g249
  (
    n265,
    n237
  );


  not
  g250
  (
    n269,
    n245
  );


  not
  g251
  (
    n278,
    n239
  );


  not
  g252
  (
    n254,
    n239
  );


  buf
  g253
  (
    n275,
    n246
  );


  not
  g254
  (
    n309,
    n278
  );


  not
  g255
  (
    n310,
    n269
  );


  not
  g256
  (
    n301,
    n272
  );


  buf
  g257
  (
    n307,
    n273
  );


  not
  g258
  (
    n304,
    n277
  );


  not
  g259
  (
    n302,
    n271
  );


  not
  g260
  (
    n305,
    n270
  );


  not
  g261
  (
    n308,
    n274
  );


  not
  g262
  (
    n303,
    n276
  );


  buf
  g263
  (
    n306,
    n275
  );


  xor
  g264
  (
    n322,
    n293,
    n49
  );


  and
  g265
  (
    n314,
    n303,
    n294,
    n48
  );


  nor
  g266
  (
    n321,
    n48,
    n300,
    n283
  );


  xor
  g267
  (
    n323,
    n296,
    n49,
    n290
  );


  xnor
  g268
  (
    n316,
    n302,
    n49,
    n285
  );


  or
  g269
  (
    n312,
    n289,
    n279,
    n287
  );


  or
  g270
  (
    n311,
    n302,
    n299,
    n284
  );


  and
  g271
  (
    n317,
    n282,
    n297,
    n295
  );


  nor
  g272
  (
    n315,
    n303,
    n301
  );


  xor
  g273
  (
    n319,
    n302,
    n280,
    n303
  );


  nand
  g274
  (
    n313,
    n304,
    n288,
    n291,
    n48
  );


  nor
  g275
  (
    n320,
    n302,
    n298,
    n303,
    n301
  );


  or
  g276
  (
    n318,
    n281,
    n292,
    n301,
    n286
  );


  xor
  g277
  (
    n343,
    n60,
    n57,
    n70,
    n315
  );


  nand
  g278
  (
    n336,
    n51,
    n62,
    n54
  );


  xnor
  g279
  (
    n326,
    n50,
    n318,
    n72,
    n78
  );


  xor
  g280
  (
    n331,
    n63,
    n59,
    n62,
    n60
  );


  xnor
  g281
  (
    n332,
    n67,
    n305,
    n78,
    n313
  );


  and
  g282
  (
    n355,
    n67,
    n64,
    n322
  );


  and
  g283
  (
    n333,
    n57,
    n54,
    n312,
    n313
  );


  nand
  g284
  (
    n368,
    n53,
    n75,
    n72,
    n77
  );


  nor
  g285
  (
    n370,
    n59,
    n74,
    n60,
    n66
  );


  nand
  g286
  (
    n360,
    n307,
    n235,
    n52,
    n309
  );


  xor
  g287
  (
    n329,
    n77,
    n307,
    n317,
    n76
  );


  xor
  g288
  (
    n346,
    n310,
    n72,
    n57,
    n78
  );


  or
  g289
  (
    n362,
    n305,
    n76,
    n316,
    n318
  );


  nand
  g290
  (
    n353,
    n59,
    n67,
    n51
  );


  nand
  g291
  (
    n325,
    n62,
    n58,
    n68,
    n63
  );


  nor
  g292
  (
    n327,
    n69,
    n56,
    n314,
    n76
  );


  and
  g293
  (
    n350,
    n70,
    n322,
    n323,
    n234
  );


  or
  g294
  (
    n339,
    n71,
    n304,
    n58,
    n75
  );


  xor
  g295
  (
    n330,
    n320,
    n53,
    n308,
    n312
  );


  xor
  g296
  (
    n365,
    n313,
    n63,
    n75,
    n317
  );


  xnor
  g297
  (
    n352,
    n74,
    n55,
    n321,
    n312
  );


  xnor
  g298
  (
    n345,
    n309,
    n315,
    n57,
    n65
  );


  xor
  g299
  (
    n371,
    n61,
    n52,
    n78,
    n323
  );


  nand
  g300
  (
    n366,
    n66,
    n319,
    n310,
    n308
  );


  and
  g301
  (
    n328,
    n69,
    n64,
    n51,
    n71
  );


  and
  g302
  (
    n364,
    n315,
    n319,
    n314,
    n321
  );


  and
  g303
  (
    n324,
    n320,
    n311,
    n322,
    n323
  );


  xnor
  g304
  (
    n356,
    n61,
    n52,
    n313,
    n306
  );


  xnor
  g305
  (
    n348,
    n318,
    n318,
    n65,
    n70
  );


  xnor
  g306
  (
    n347,
    n50,
    n307,
    n56,
    n69
  );


  and
  g307
  (
    n354,
    n320,
    n319,
    n234,
    n77
  );


  and
  g308
  (
    n334,
    n52,
    n60,
    n56,
    n309
  );


  and
  g309
  (
    n372,
    n51,
    n55,
    n74,
    n316
  );


  and
  g310
  (
    n351,
    n319,
    n312,
    n68
  );


  or
  g311
  (
    n359,
    n64,
    n235,
    n72,
    n317
  );


  nor
  g312
  (
    n342,
    n314,
    n308,
    n73,
    n310
  );


  and
  g313
  (
    KeyWire_0_31,
    n55,
    n53,
    n320,
    n304
  );


  or
  g314
  (
    n363,
    n304,
    n68,
    n311,
    n323
  );


  nand
  g315
  (
    n373,
    n59,
    n306,
    n307,
    n316
  );


  xor
  g316
  (
    n367,
    n73,
    n305,
    n76,
    n235
  );


  or
  g317
  (
    n361,
    n61,
    n314,
    n56,
    n58
  );


  xor
  g318
  (
    n369,
    n58,
    n70,
    n71,
    n316
  );


  xnor
  g319
  (
    n344,
    n53,
    n50,
    n71,
    n321
  );


  nand
  g320
  (
    n357,
    n65,
    n73,
    n235,
    n62
  );


  nand
  g321
  (
    n349,
    n310,
    n50,
    n308,
    n306
  );


  xnor
  g322
  (
    n358,
    n66,
    n322,
    n69,
    n74
  );


  nor
  g323
  (
    n340,
    n75,
    n317,
    n309,
    n73
  );


  nor
  g324
  (
    n335,
    n61,
    n321,
    n315,
    n54
  );


  and
  g325
  (
    KeyWire_0_21,
    n305,
    n234,
    n65,
    n77
  );


  nor
  g326
  (
    n338,
    n66,
    n63,
    n306,
    n55
  );


  buf
  g327
  (
    n484,
    n326
  );


  not
  g328
  (
    n483,
    n358
  );


  not
  g329
  (
    n448,
    n328
  );


  not
  g330
  (
    n381,
    n362
  );


  buf
  g331
  (
    n415,
    n351
  );


  not
  g332
  (
    n470,
    n367
  );


  buf
  g333
  (
    n440,
    n349
  );


  not
  g334
  (
    n431,
    n361
  );


  not
  g335
  (
    n497,
    n342
  );


  buf
  g336
  (
    n408,
    n344
  );


  not
  g337
  (
    n416,
    n344
  );


  not
  g338
  (
    n459,
    n343
  );


  buf
  g339
  (
    n490,
    n338
  );


  not
  g340
  (
    n442,
    n364
  );


  buf
  g341
  (
    n522,
    n352
  );


  not
  g342
  (
    n520,
    n372
  );


  buf
  g343
  (
    n388,
    n366
  );


  not
  g344
  (
    n404,
    n338
  );


  not
  g345
  (
    n413,
    n359
  );


  buf
  g346
  (
    n529,
    n348
  );


  not
  g347
  (
    n461,
    n326
  );


  buf
  g348
  (
    n449,
    n341
  );


  buf
  g349
  (
    n420,
    n368
  );


  buf
  g350
  (
    n469,
    n348
  );


  buf
  g351
  (
    KeyWire_0_3,
    n336
  );


  buf
  g352
  (
    n504,
    n354
  );


  not
  g353
  (
    n494,
    n372
  );


  buf
  g354
  (
    n527,
    n372
  );


  buf
  g355
  (
    n393,
    n341
  );


  not
  g356
  (
    n441,
    n340
  );


  not
  g357
  (
    n414,
    n345
  );


  not
  g358
  (
    n391,
    n349
  );


  not
  g359
  (
    KeyWire_0_57,
    n364
  );


  buf
  g360
  (
    n512,
    n358
  );


  not
  g361
  (
    n386,
    n357
  );


  not
  g362
  (
    n437,
    n369
  );


  not
  g363
  (
    KeyWire_0_8,
    n347
  );


  not
  g364
  (
    n492,
    n347
  );


  buf
  g365
  (
    KeyWire_0_9,
    n360
  );


  buf
  g366
  (
    n516,
    n364
  );


  buf
  g367
  (
    n411,
    n351
  );


  not
  g368
  (
    n400,
    n333
  );


  buf
  g369
  (
    n427,
    n345
  );


  buf
  g370
  (
    n392,
    n367
  );


  not
  g371
  (
    n397,
    n350
  );


  not
  g372
  (
    n433,
    n345
  );


  not
  g373
  (
    n443,
    n370
  );


  buf
  g374
  (
    n456,
    n357
  );


  not
  g375
  (
    n394,
    n334
  );


  not
  g376
  (
    n517,
    n357
  );


  not
  g377
  (
    n488,
    n369
  );


  not
  g378
  (
    n436,
    n337
  );


  buf
  g379
  (
    n478,
    n325
  );


  buf
  g380
  (
    KeyWire_0_37,
    n343
  );


  buf
  g381
  (
    n434,
    n356
  );


  buf
  g382
  (
    n503,
    n365
  );


  not
  g383
  (
    KeyWire_0_36,
    n350
  );


  buf
  g384
  (
    n514,
    n365
  );


  not
  g385
  (
    n521,
    n352
  );


  buf
  g386
  (
    n487,
    n355
  );


  not
  g387
  (
    n515,
    n362
  );


  buf
  g388
  (
    KeyWire_0_61,
    n369
  );


  not
  g389
  (
    n429,
    n330
  );


  not
  g390
  (
    n455,
    n332
  );


  buf
  g391
  (
    n509,
    n346
  );


  buf
  g392
  (
    n482,
    n371
  );


  buf
  g393
  (
    n380,
    n370
  );


  buf
  g394
  (
    n498,
    n342
  );


  buf
  g395
  (
    n382,
    n368
  );


  not
  g396
  (
    n468,
    n340
  );


  buf
  g397
  (
    n472,
    n364
  );


  buf
  g398
  (
    n402,
    n352
  );


  buf
  g399
  (
    n458,
    n331
  );


  not
  g400
  (
    n405,
    n344
  );


  not
  g401
  (
    KeyWire_0_18,
    n332
  );


  not
  g402
  (
    n438,
    n360
  );


  buf
  g403
  (
    n501,
    n353
  );


  not
  g404
  (
    n467,
    n333
  );


  buf
  g405
  (
    n518,
    n338
  );


  buf
  g406
  (
    n447,
    n370
  );


  not
  g407
  (
    n474,
    n325
  );


  buf
  g408
  (
    n486,
    n368
  );


  buf
  g409
  (
    n396,
    n358
  );


  buf
  g410
  (
    n432,
    n342
  );


  not
  g411
  (
    n430,
    n367
  );


  buf
  g412
  (
    n375,
    n346
  );


  not
  g413
  (
    n511,
    n372
  );


  buf
  g414
  (
    n399,
    n373
  );


  buf
  g415
  (
    KeyWire_0_38,
    n348
  );


  buf
  g416
  (
    n505,
    n329
  );


  buf
  g417
  (
    n460,
    n355
  );


  not
  g418
  (
    n463,
    n365
  );


  not
  g419
  (
    n519,
    n347
  );


  not
  g420
  (
    n446,
    n355
  );


  not
  g421
  (
    KeyWire_0_42,
    n363
  );


  not
  g422
  (
    n513,
    n335
  );


  not
  g423
  (
    n489,
    n362
  );


  buf
  g424
  (
    n435,
    n340
  );


  buf
  g425
  (
    n476,
    n361
  );


  not
  g426
  (
    n454,
    n353
  );


  not
  g427
  (
    n473,
    n335
  );


  buf
  g428
  (
    n525,
    n339
  );


  buf
  g429
  (
    n374,
    n356
  );


  not
  g430
  (
    n428,
    n353
  );


  not
  g431
  (
    n477,
    n354
  );


  buf
  g432
  (
    n526,
    n327
  );


  buf
  g433
  (
    n423,
    n371
  );


  not
  g434
  (
    n450,
    n339
  );


  buf
  g435
  (
    n395,
    n370
  );


  not
  g436
  (
    n409,
    n334
  );


  buf
  g437
  (
    n412,
    n349
  );


  buf
  g438
  (
    n376,
    n368
  );


  buf
  g439
  (
    n496,
    n369
  );


  buf
  g440
  (
    n422,
    n357
  );


  not
  g441
  (
    n407,
    n359
  );


  not
  g442
  (
    n510,
    n356
  );


  not
  g443
  (
    n444,
    n352
  );


  not
  g444
  (
    n418,
    n360
  );


  not
  g445
  (
    n424,
    n361
  );


  not
  g446
  (
    n421,
    n329
  );


  buf
  g447
  (
    n499,
    n366
  );


  buf
  g448
  (
    n453,
    n359
  );


  not
  g449
  (
    n528,
    n363
  );


  not
  g450
  (
    n425,
    n359
  );


  not
  g451
  (
    n485,
    n343
  );


  buf
  g452
  (
    n523,
    n331
  );


  not
  g453
  (
    n377,
    n371
  );


  not
  g454
  (
    n481,
    n330
  );


  not
  g455
  (
    n385,
    n362
  );


  buf
  g456
  (
    n475,
    n339
  );


  not
  g457
  (
    n390,
    n337
  );


  buf
  g458
  (
    n379,
    n328
  );


  not
  g459
  (
    n493,
    n365
  );


  buf
  g460
  (
    n508,
    n366
  );


  buf
  g461
  (
    n383,
    n358
  );


  buf
  g462
  (
    n417,
    n361
  );


  not
  g463
  (
    n445,
    n327
  );


  buf
  g464
  (
    n401,
    n373
  );


  not
  g465
  (
    n480,
    n360
  );


  buf
  g466
  (
    n384,
    n356
  );


  buf
  g467
  (
    n451,
    n363
  );


  not
  g468
  (
    n500,
    n336
  );


  not
  g469
  (
    n398,
    n366
  );


  not
  g470
  (
    n506,
    n346
  );


  not
  g471
  (
    n502,
    n355
  );


  buf
  g472
  (
    n457,
    n354
  );


  buf
  g473
  (
    n495,
    n341
  );


  buf
  g474
  (
    n387,
    n373
  );


  not
  g475
  (
    n466,
    n350
  );


  not
  g476
  (
    n410,
    n353
  );


  buf
  g477
  (
    n524,
    n371
  );


  not
  g478
  (
    KeyWire_0_51,
    n354
  );


  not
  g479
  (
    n479,
    n373
  );


  not
  g480
  (
    n471,
    n367
  );


  buf
  g481
  (
    n439,
    n351
  );


  buf
  g482
  (
    n491,
    n363
  );


  buf
  g483
  (
    n828,
    n430
  );


  buf
  g484
  (
    n640,
    n415
  );


  buf
  g485
  (
    n776,
    n379
  );


  buf
  g486
  (
    n861,
    n119
  );


  not
  g487
  (
    n561,
    n147
  );


  not
  g488
  (
    n549,
    n171
  );


  buf
  g489
  (
    n710,
    n505
  );


  buf
  g490
  (
    n718,
    n483
  );


  not
  g491
  (
    KeyWire_0_26,
    n506
  );


  buf
  g492
  (
    n665,
    n450
  );


  buf
  g493
  (
    n684,
    n418
  );


  buf
  g494
  (
    n730,
    n512
  );


  not
  g495
  (
    n742,
    n139
  );


  buf
  g496
  (
    n530,
    n414
  );


  not
  g497
  (
    n754,
    n175
  );


  not
  g498
  (
    n686,
    n380
  );


  not
  g499
  (
    n743,
    n162
  );


  buf
  g500
  (
    n799,
    n487
  );


  not
  g501
  (
    n801,
    n185
  );


  buf
  g502
  (
    n898,
    n96
  );


  buf
  g503
  (
    n591,
    n184
  );


  not
  g504
  (
    n751,
    n212
  );


  buf
  g505
  (
    n723,
    n438
  );


  not
  g506
  (
    n747,
    n94
  );


  not
  g507
  (
    n794,
    n504
  );


  buf
  g508
  (
    n638,
    n428
  );


  buf
  g509
  (
    n866,
    n161
  );


  buf
  g510
  (
    n726,
    n128
  );


  buf
  g511
  (
    n775,
    n86
  );


  not
  g512
  (
    n681,
    n175
  );


  buf
  g513
  (
    n615,
    n500
  );


  not
  g514
  (
    n873,
    n206
  );


  not
  g515
  (
    n760,
    n118
  );


  buf
  g516
  (
    n863,
    n437
  );


  buf
  g517
  (
    n772,
    n412
  );


  buf
  g518
  (
    n598,
    n135
  );


  not
  g519
  (
    n660,
    n445
  );


  buf
  g520
  (
    n902,
    n402
  );


  buf
  g521
  (
    n541,
    n186
  );


  not
  g522
  (
    n679,
    n151
  );


  not
  g523
  (
    n582,
    n117
  );


  not
  g524
  (
    n663,
    n138
  );


  buf
  g525
  (
    n755,
    n478
  );


  buf
  g526
  (
    n689,
    n188
  );


  not
  g527
  (
    n781,
    n492
  );


  buf
  g528
  (
    n609,
    n175
  );


  buf
  g529
  (
    n651,
    n200
  );


  not
  g530
  (
    n559,
    n512
  );


  not
  g531
  (
    n596,
    n151
  );


  buf
  g532
  (
    n672,
    n504
  );


  not
  g533
  (
    n811,
    n472
  );


  buf
  g534
  (
    n589,
    n211
  );


  buf
  g535
  (
    n763,
    n492
  );


  not
  g536
  (
    n741,
    n442
  );


  buf
  g537
  (
    n789,
    n127
  );


  not
  g538
  (
    n536,
    n518
  );


  buf
  g539
  (
    n753,
    n400
  );


  buf
  g540
  (
    KeyWire_0_5,
    n182
  );


  not
  g541
  (
    n578,
    n196
  );


  buf
  g542
  (
    n719,
    n131
  );


  buf
  g543
  (
    n778,
    n374
  );


  not
  g544
  (
    n603,
    n404
  );


  buf
  g545
  (
    n810,
    n475
  );


  not
  g546
  (
    n709,
    n161
  );


  buf
  g547
  (
    KeyWire_0_16,
    n488
  );


  not
  g548
  (
    n800,
    n420
  );


  not
  g549
  (
    n588,
    n107
  );


  buf
  g550
  (
    n901,
    n167
  );


  not
  g551
  (
    n792,
    n217
  );


  not
  g552
  (
    n568,
    n401
  );


  buf
  g553
  (
    n867,
    n92
  );


  buf
  g554
  (
    n724,
    n415
  );


  buf
  g555
  (
    n740,
    n469
  );


  not
  g556
  (
    n882,
    n386
  );


  not
  g557
  (
    n893,
    n463
  );


  not
  g558
  (
    n853,
    n128
  );


  buf
  g559
  (
    n802,
    n502
  );


  not
  g560
  (
    n645,
    n171
  );


  buf
  g561
  (
    n886,
    n486
  );


  buf
  g562
  (
    n734,
    n211
  );


  buf
  g563
  (
    n661,
    n195
  );


  buf
  g564
  (
    n769,
    n496
  );


  not
  g565
  (
    n881,
    n472
  );


  buf
  g566
  (
    n700,
    n156
  );


  not
  g567
  (
    n795,
    n192
  );


  not
  g568
  (
    n666,
    n381
  );


  buf
  g569
  (
    n696,
    n142
  );


  buf
  g570
  (
    n729,
    n81
  );


  buf
  g571
  (
    n818,
    n488
  );


  buf
  g572
  (
    n783,
    n167
  );


  buf
  g573
  (
    n545,
    n143
  );


  not
  g574
  (
    n532,
    n478
  );


  buf
  g575
  (
    n860,
    n459
  );


  not
  g576
  (
    KeyWire_0_47,
    n220
  );


  not
  g577
  (
    n785,
    n443
  );


  not
  g578
  (
    n564,
    n104
  );


  buf
  g579
  (
    n736,
    n402
  );


  buf
  g580
  (
    n604,
    n475
  );


  buf
  g581
  (
    n637,
    n127
  );


  buf
  g582
  (
    n890,
    n95
  );


  buf
  g583
  (
    n648,
    n145
  );


  buf
  g584
  (
    n551,
    n114
  );


  not
  g585
  (
    n558,
    n114
  );


  buf
  g586
  (
    n832,
    n491
  );


  buf
  g587
  (
    n817,
    n202
  );


  buf
  g588
  (
    n626,
    n446
  );


  buf
  g589
  (
    n906,
    n96
  );


  not
  g590
  (
    n885,
    n431
  );


  not
  g591
  (
    n752,
    n203
  );


  not
  g592
  (
    n616,
    n405
  );


  buf
  g593
  (
    n835,
    n84
  );


  not
  g594
  (
    n593,
    n464
  );


  buf
  g595
  (
    n784,
    n90
  );


  not
  g596
  (
    n805,
    n502
  );


  not
  g597
  (
    n877,
    n137
  );


  buf
  g598
  (
    n838,
    n107
  );


  not
  g599
  (
    n874,
    n415
  );


  not
  g600
  (
    n847,
    n487
  );


  not
  g601
  (
    n618,
    n116
  );


  or
  g602
  (
    n848,
    n422,
    n197,
    n214,
    n381
  );


  nor
  g603
  (
    n819,
    n506,
    n161,
    n474,
    n110
  );


  nand
  g604
  (
    n643,
    n456,
    n416,
    n133,
    n439
  );


  xnor
  g605
  (
    n765,
    n164,
    n403,
    n464,
    n446
  );


  xor
  g606
  (
    n745,
    n460,
    n101,
    n517,
    n127
  );


  and
  g607
  (
    n875,
    n405,
    n148,
    n489,
    n377
  );


  nand
  g608
  (
    n825,
    n90,
    n390,
    n479,
    n427
  );


  nor
  g609
  (
    n617,
    n511,
    n461,
    n449,
    n515
  );


  or
  g610
  (
    n655,
    n410,
    n159,
    n467,
    n109
  );


  or
  g611
  (
    n692,
    n200,
    n377,
    n383,
    n473
  );


  nand
  g612
  (
    n738,
    n429,
    n395,
    n408
  );


  xor
  g613
  (
    n701,
    n165,
    n194,
    n136,
    n215
  );


  nor
  g614
  (
    n815,
    n120,
    n439,
    n387,
    n411
  );


  or
  g615
  (
    n713,
    n467,
    n466,
    n505,
    n211
  );


  xnor
  g616
  (
    n693,
    n477,
    n443,
    n498,
    n93
  );


  or
  g617
  (
    n857,
    n465,
    n401,
    n470,
    n217
  );


  xnor
  g618
  (
    n870,
    n500,
    n114,
    n217,
    n453
  );


  nor
  g619
  (
    n687,
    n186,
    n463,
    n508,
    n456
  );


  xnor
  g620
  (
    n607,
    n444,
    n400,
    n216,
    n399
  );


  xnor
  g621
  (
    n581,
    n199,
    n413,
    n106,
    n475
  );


  nor
  g622
  (
    n602,
    n117,
    n120,
    n401,
    n180
  );


  and
  g623
  (
    n829,
    n391,
    n497,
    n520,
    n119
  );


  xor
  g624
  (
    n814,
    n189,
    n174,
    n457,
    n468
  );


  nand
  g625
  (
    n542,
    n195,
    n152,
    n197
  );


  or
  g626
  (
    n806,
    n154,
    n79,
    n219,
    n87
  );


  and
  g627
  (
    n899,
    n499,
    n91,
    n418,
    n102
  );


  nor
  g628
  (
    n858,
    n176,
    n419,
    n509,
    n440
  );


  nor
  g629
  (
    n635,
    n79,
    n132,
    n396,
    n433
  );


  xnor
  g630
  (
    n614,
    n483,
    n85,
    n115,
    n379
  );


  nand
  g631
  (
    KeyWire_0_35,
    n174,
    n89,
    n98,
    n209
  );


  nand
  g632
  (
    n854,
    n130,
    n192,
    n105,
    n399
  );


  or
  g633
  (
    n534,
    n385,
    n94,
    n82,
    n484
  );


  and
  g634
  (
    n649,
    n87,
    n121,
    n414,
    n124
  );


  xnor
  g635
  (
    n749,
    n503,
    n134,
    n190,
    n158
  );


  and
  g636
  (
    n639,
    n85,
    n217,
    n393,
    n183
  );


  xnor
  g637
  (
    n807,
    n133,
    n100,
    n493,
    n194
  );


  nand
  g638
  (
    n694,
    n445,
    n395,
    n443,
    n193
  );


  xnor
  g639
  (
    n565,
    n437,
    n151,
    n160,
    n122
  );


  nor
  g640
  (
    n884,
    n381,
    n158,
    n449,
    n455
  );


  or
  g641
  (
    n865,
    n422,
    n121,
    n106,
    n434
  );


  and
  g642
  (
    n664,
    n93,
    n82,
    n215,
    n111
  );


  xor
  g643
  (
    n699,
    n517,
    n101,
    n200,
    n180
  );


  and
  g644
  (
    n554,
    n452,
    n462,
    n400,
    n441
  );


  xor
  g645
  (
    n657,
    n488,
    n144,
    n494,
    n432
  );


  nand
  g646
  (
    n897,
    n120,
    n193,
    n449,
    n131
  );


  xor
  g647
  (
    n836,
    n384,
    n148,
    n392,
    n509
  );


  xnor
  g648
  (
    n851,
    n196,
    n154,
    n392,
    n482
  );


  xnor
  g649
  (
    n849,
    n205,
    n132,
    n162,
    n434
  );


  xnor
  g650
  (
    n844,
    n500,
    n146,
    n409,
    n136
  );


  or
  g651
  (
    n889,
    n81,
    n513,
    n170,
    n163
  );


  xor
  g652
  (
    n557,
    n434,
    n190,
    n424,
    n415
  );


  and
  g653
  (
    n803,
    n216,
    n396,
    n391,
    n382
  );


  and
  g654
  (
    n711,
    n407,
    n125,
    n100,
    n384
  );


  xor
  g655
  (
    n563,
    n459,
    n169,
    n374,
    n394
  );


  and
  g656
  (
    n872,
    n495,
    n109,
    n169,
    n448
  );


  xnor
  g657
  (
    n725,
    n431,
    n420,
    n168,
    n171
  );


  nor
  g658
  (
    n780,
    n126,
    n89,
    n221,
    n379
  );


  or
  g659
  (
    n620,
    n178,
    n383,
    n141,
    n503
  );


  xor
  g660
  (
    n864,
    n213,
    n450,
    n186,
    n82
  );


  and
  g661
  (
    n566,
    n409,
    n86,
    n188,
    n458
  );


  xnor
  g662
  (
    n606,
    n152,
    n117,
    n208,
    n383
  );


  xor
  g663
  (
    n612,
    n140,
    n145,
    n482,
    n479
  );


  or
  g664
  (
    n695,
    n514,
    n518,
    n417,
    n477
  );


  xnor
  g665
  (
    n883,
    n110,
    n215,
    n124,
    n166
  );


  nand
  g666
  (
    n600,
    n164,
    n489,
    n456,
    n186
  );


  and
  g667
  (
    n677,
    n465,
    n432,
    n482,
    n471
  );


  xnor
  g668
  (
    n721,
    n475,
    n518,
    n180,
    n204
  );


  and
  g669
  (
    n690,
    n155,
    n375,
    n426,
    n450
  );


  xnor
  g670
  (
    n673,
    n210,
    n109,
    n411,
    n468
  );


  nor
  g671
  (
    n631,
    n91,
    n156,
    n130,
    n135
  );


  xnor
  g672
  (
    n702,
    n416,
    n481,
    n153,
    n508
  );


  xnor
  g673
  (
    n624,
    n98,
    n146,
    n183,
    n154
  );


  xor
  g674
  (
    n714,
    n134,
    n382,
    n490,
    n391
  );


  xor
  g675
  (
    n717,
    n519,
    n513,
    n393,
    n451
  );


  xnor
  g676
  (
    n544,
    n391,
    n490,
    n389,
    n476
  );


  or
  g677
  (
    n548,
    n424,
    n98,
    n410,
    n123
  );


  and
  g678
  (
    n669,
    n385,
    n218,
    n135,
    n130
  );


  and
  g679
  (
    n759,
    n406,
    n515,
    n194,
    n436
  );


  nor
  g680
  (
    n868,
    n480,
    n161,
    n177,
    n166
  );


  nand
  g681
  (
    n895,
    n193,
    n153,
    n150,
    n112
  );


  nor
  g682
  (
    n676,
    n503,
    n119,
    n212,
    n423
  );


  xor
  g683
  (
    n748,
    n402,
    n179,
    n419,
    n113
  );


  xnor
  g684
  (
    n623,
    n385,
    n107,
    n397,
    n388
  );


  and
  g685
  (
    n782,
    n92,
    n88,
    n122,
    n507
  );


  xnor
  g686
  (
    n538,
    n183,
    n181,
    n378,
    n460
  );


  or
  g687
  (
    KeyWire_0_0,
    n462,
    n113,
    n474,
    n213
  );


  xnor
  g688
  (
    n770,
    n215,
    n397,
    n138,
    n468
  );


  xnor
  g689
  (
    n727,
    n476,
    n440,
    n195,
    n150
  );


  or
  g690
  (
    n629,
    n516,
    n439,
    n469,
    n494
  );


  and
  g691
  (
    n758,
    n467,
    n389,
    n426,
    n438
  );


  xor
  g692
  (
    n907,
    n392,
    n455,
    n407,
    n493
  );


  xor
  g693
  (
    n722,
    n417,
    n209,
    n213,
    n433
  );


  or
  g694
  (
    n555,
    n478,
    n513,
    n220,
    n471
  );


  nor
  g695
  (
    n580,
    n138,
    n173,
    n149,
    n146
  );


  or
  g696
  (
    n720,
    n214,
    n407,
    n506,
    n87
  );


  xnor
  g697
  (
    n656,
    n388,
    n495,
    n398,
    n487
  );


  xor
  g698
  (
    n553,
    n458,
    n484,
    n510,
    n409
  );


  and
  g699
  (
    KeyWire_0_34,
    n95,
    n193,
    n481,
    n192
  );


  nor
  g700
  (
    n812,
    n169,
    n141,
    n220,
    n410
  );


  or
  g701
  (
    n641,
    n517,
    n205,
    n472,
    n219
  );


  nor
  g702
  (
    n636,
    n405,
    n81,
    n106,
    n375
  );


  nor
  g703
  (
    n539,
    n489,
    n465,
    n156,
    n433
  );


  nand
  g704
  (
    n790,
    n483,
    n87,
    n181,
    n85
  );


  xor
  g705
  (
    n834,
    n480,
    n121,
    n460,
    n376
  );


  nor
  g706
  (
    n826,
    n84,
    n140,
    n388,
    n406
  );


  nor
  g707
  (
    n628,
    n180,
    n152,
    n126,
    n374
  );


  xor
  g708
  (
    n644,
    n497,
    n482,
    n213,
    n80
  );


  and
  g709
  (
    KeyWire_0_50,
    n88,
    n208,
    n145,
    n454
  );


  nor
  g710
  (
    n599,
    n86,
    n220,
    n125,
    n501
  );


  xor
  g711
  (
    n587,
    n473,
    n168,
    n437,
    n444
  );


  nand
  g712
  (
    n590,
    n208,
    n160,
    n492,
    n440
  );


  and
  g713
  (
    KeyWire_0_28,
    n501,
    n381,
    n425,
    n165
  );


  or
  g714
  (
    n552,
    n378,
    n144,
    n506,
    n173
  );


  xnor
  g715
  (
    n843,
    n420,
    n86,
    n387,
    n82
  );


  nor
  g716
  (
    n712,
    n455,
    n444,
    n499,
    n469
  );


  nor
  g717
  (
    n586,
    n426,
    n83,
    n205,
    n404
  );


  xnor
  g718
  (
    n791,
    n485,
    n182,
    n178,
    n438
  );


  xnor
  g719
  (
    KeyWire_0_59,
    n468,
    n103,
    n90,
    n165
  );


  or
  g720
  (
    n859,
    n483,
    n210,
    n105,
    n198
  );


  xnor
  g721
  (
    n771,
    n502,
    n419,
    n462,
    n408
  );


  nand
  g722
  (
    n633,
    n432,
    n80,
    n118,
    n440
  );


  xor
  g723
  (
    n533,
    n396,
    n96,
    n470,
    n176
  );


  and
  g724
  (
    n766,
    n478,
    n177,
    n131,
    n94
  );


  xor
  g725
  (
    n642,
    n182,
    n387,
    n131,
    n486
  );


  nand
  g726
  (
    n674,
    n163,
    n514,
    n204,
    n168
  );


  nand
  g727
  (
    n824,
    n185,
    n168,
    n403,
    n136
  );


  xor
  g728
  (
    n543,
    n157,
    n417,
    n490,
    n122
  );


  and
  g729
  (
    n579,
    n496,
    n120,
    n196,
    n199
  );


  xnor
  g730
  (
    n671,
    n424,
    n516,
    n108,
    n167
  );


  xnor
  g731
  (
    n869,
    n393,
    n423,
    n218,
    n452
  );


  or
  g732
  (
    n797,
    n187,
    n406,
    n155,
    n499
  );


  xnor
  g733
  (
    KeyWire_0_43,
    n141,
    n441,
    n498,
    n394
  );


  or
  g734
  (
    n597,
    n494,
    n406,
    n105,
    n452
  );


  or
  g735
  (
    n779,
    n382,
    n135,
    n111,
    n169
  );


  or
  g736
  (
    n822,
    n432,
    n421,
    n172,
    n414
  );


  nor
  g737
  (
    n878,
    n377,
    n447,
    n104,
    n380
  );


  xor
  g738
  (
    KeyWire_0_24,
    n111,
    n202,
    n99,
    n431
  );


  or
  g739
  (
    n537,
    n450,
    n140,
    n378,
    n497
  );


  xor
  g740
  (
    n896,
    n103,
    n431,
    n384,
    n121
  );


  nor
  g741
  (
    n575,
    n124,
    n476,
    n212,
    n113
  );


  and
  g742
  (
    n856,
    n101,
    n511,
    n218,
    n451
  );


  and
  g743
  (
    n691,
    n185,
    n516,
    n80,
    n83
  );


  nand
  g744
  (
    KeyWire_0_62,
    n394,
    n508,
    n83,
    n153
  );


  xnor
  g745
  (
    n715,
    n505,
    n221,
    n164,
    n141
  );


  nand
  g746
  (
    n728,
    n409,
    n158,
    n488,
    n427
  );


  xor
  g747
  (
    n608,
    n413,
    n162,
    n412,
    n140
  );


  xnor
  g748
  (
    n768,
    n460,
    n197,
    n108,
    n467
  );


  xor
  g749
  (
    KeyWire_0_17,
    n103,
    n451,
    n170,
    n477
  );


  xnor
  g750
  (
    n621,
    n115,
    n96,
    n130,
    n94
  );


  nand
  g751
  (
    n584,
    n181,
    n209,
    n133,
    n212
  );


  nand
  g752
  (
    n592,
    n112,
    n142,
    n486,
    n204
  );


  or
  g753
  (
    n531,
    n174,
    n157,
    n422,
    n485
  );


  nor
  g754
  (
    n837,
    n173,
    n92,
    n485,
    n126
  );


  nor
  g755
  (
    n594,
    n429,
    n412,
    n427,
    n457
  );


  nand
  g756
  (
    n705,
    n159,
    n405,
    n470,
    n480
  );


  xor
  g757
  (
    n688,
    n436,
    n208,
    n149,
    n176
  );


  nand
  g758
  (
    n845,
    n145,
    n456,
    n132,
    n496
  );


  xor
  g759
  (
    n658,
    n519,
    n485,
    n97,
    n89
  );


  or
  g760
  (
    KeyWire_0_44,
    n137,
    n143,
    n179,
    n453
  );


  nor
  g761
  (
    n703,
    n510,
    n102,
    n459,
    n494
  );


  xnor
  g762
  (
    n787,
    n134,
    n473,
    n118,
    n386
  );


  xnor
  g763
  (
    n830,
    n486,
    n435,
    n157,
    n452
  );


  nor
  g764
  (
    KeyWire_0_29,
    n83,
    n125,
    n509,
    n100
  );


  or
  g765
  (
    n892,
    n453,
    n471,
    n481,
    n79
  );


  nand
  g766
  (
    n573,
    n177,
    n100,
    n400,
    n106
  );


  and
  g767
  (
    n683,
    n143,
    n95,
    n461,
    n205
  );


  nand
  g768
  (
    n680,
    n383,
    n155,
    n462,
    n403
  );


  xnor
  g769
  (
    n887,
    n448,
    n204,
    n93,
    n160
  );


  xnor
  g770
  (
    n850,
    n466,
    n177,
    n144,
    n84
  );


  nand
  g771
  (
    n668,
    n481,
    n487,
    n144,
    n200
  );


  and
  g772
  (
    n746,
    n428,
    n93,
    n512,
    n398
  );


  nand
  g773
  (
    n798,
    n517,
    n191,
    n443,
    n195
  );


  nand
  g774
  (
    n796,
    n419,
    n410,
    n401,
    n201
  );


  xnor
  g775
  (
    n562,
    n423,
    n92,
    n498,
    n510
  );


  xnor
  g776
  (
    n583,
    n179,
    n412,
    n209,
    n89
  );


  or
  g777
  (
    n585,
    n509,
    n417,
    n498,
    n99
  );


  and
  g778
  (
    n737,
    n402,
    n515,
    n110,
    n403
  );


  xnor
  g779
  (
    n808,
    n191,
    n414,
    n503,
    n102
  );


  or
  g780
  (
    n627,
    n88,
    n459,
    n182,
    n375
  );


  nor
  g781
  (
    n756,
    n198,
    n464,
    n448,
    n389
  );


  or
  g782
  (
    n716,
    n464,
    n447,
    n408,
    n152
  );


  or
  g783
  (
    n698,
    n110,
    n80,
    n219,
    n123
  );


  nor
  g784
  (
    n571,
    n188,
    n496,
    n118,
    n125
  );


  and
  g785
  (
    n670,
    n184,
    n477,
    n115,
    n423
  );


  nor
  g786
  (
    n630,
    n377,
    n129,
    n396,
    n149
  );


  xnor
  g787
  (
    n820,
    n99,
    n214,
    n418,
    n484
  );


  nor
  g788
  (
    n823,
    n142,
    n134,
    n136,
    n471
  );


  or
  g789
  (
    n833,
    n476,
    n451,
    n495,
    n385
  );


  and
  g790
  (
    n540,
    n207,
    n379,
    n411,
    n192
  );


  nor
  g791
  (
    n622,
    n172,
    n201,
    n207,
    n189
  );


  xor
  g792
  (
    n706,
    n429,
    n413,
    n436,
    n116
  );


  xor
  g793
  (
    n903,
    n490,
    n492,
    n500,
    n399
  );


  or
  g794
  (
    KeyWire_0_14,
    n109,
    n178,
    n470,
    n173
  );


  and
  g795
  (
    n813,
    n408,
    n430,
    n170,
    n203
  );


  nor
  g796
  (
    n905,
    n184,
    n491,
    n439,
    n420
  );


  xnor
  g797
  (
    n739,
    n123,
    n424,
    n159,
    n444
  );


  or
  g798
  (
    n625,
    n473,
    n147,
    n442,
    n421
  );


  xnor
  g799
  (
    n653,
    n398,
    n507,
    n441,
    n91
  );


  or
  g800
  (
    n535,
    n137,
    n176,
    n447,
    n399
  );


  and
  g801
  (
    n574,
    n148,
    n446,
    n495,
    n463
  );


  xor
  g802
  (
    n762,
    n407,
    n139,
    n101,
    n97
  );


  or
  g803
  (
    n577,
    n202,
    n150,
    n129,
    n123
  );


  or
  g804
  (
    n682,
    n175,
    n153,
    n386,
    n198
  );


  xor
  g805
  (
    n732,
    n515,
    n491,
    n448,
    n505
  );


  or
  g806
  (
    n547,
    n128,
    n187,
    n154,
    n501
  );


  nand
  g807
  (
    n731,
    n81,
    n112,
    n453,
    n147
  );


  and
  g808
  (
    n852,
    n97,
    n115,
    n516,
    n519
  );


  xor
  g809
  (
    n809,
    n170,
    n111,
    n139,
    n397
  );


  nor
  g810
  (
    n891,
    n122,
    n218,
    n211,
    n491
  );


  nor
  g811
  (
    n761,
    n469,
    n404,
    n466,
    n457
  );


  xnor
  g812
  (
    n757,
    n421,
    n458,
    n461,
    n150
  );


  nand
  g813
  (
    n654,
    n104,
    n90,
    n416,
    n435
  );


  nand
  g814
  (
    n816,
    n394,
    n374,
    n442,
    n436
  );


  xor
  g815
  (
    KeyWire_0_41,
    n390,
    n428,
    n172,
    n189
  );


  xnor
  g816
  (
    n841,
    n446,
    n493,
    n190,
    n164
  );


  or
  g817
  (
    n707,
    n404,
    n103,
    n206,
    n105
  );


  xnor
  g818
  (
    n572,
    n416,
    n132,
    n196,
    n457
  );


  and
  g819
  (
    n605,
    n151,
    n214,
    n155,
    n216
  );


  nand
  g820
  (
    n777,
    n454,
    n172,
    n88,
    n163
  );


  xor
  g821
  (
    n613,
    n449,
    n380,
    n474,
    n166
  );


  xnor
  g822
  (
    n888,
    n202,
    n185,
    n437,
    n388
  );


  xnor
  g823
  (
    n842,
    n139,
    n519,
    n430,
    n184
  );


  xnor
  g824
  (
    n786,
    n489,
    n501,
    n375,
    n203
  );


  xor
  g825
  (
    n744,
    n434,
    n162,
    n163,
    n376
  );


  and
  g826
  (
    n685,
    n199,
    n157,
    n507,
    n129
  );


  and
  g827
  (
    n619,
    n113,
    n442,
    n474,
    n507
  );


  xnor
  g828
  (
    n894,
    n376,
    n126,
    n149,
    n426
  );


  and
  g829
  (
    n793,
    n108,
    n188,
    n502,
    n201
  );


  xnor
  g830
  (
    n650,
    n147,
    n479,
    n119,
    n518
  );


  xor
  g831
  (
    KeyWire_0_15,
    n421,
    n210,
    n425,
    n454
  );


  and
  g832
  (
    n601,
    n428,
    n191,
    n376,
    n512
  );


  or
  g833
  (
    KeyWire_0_20,
    n189,
    n397,
    n447,
    n85
  );


  and
  g834
  (
    n652,
    n458,
    n418,
    n178,
    n210
  );


  and
  g835
  (
    n567,
    n386,
    n219,
    n466,
    n514
  );


  xnor
  g836
  (
    n846,
    n137,
    n425,
    n393,
    n191
  );


  nor
  g837
  (
    KeyWire_0_39,
    n148,
    n95,
    n84,
    n190
  );


  and
  g838
  (
    n576,
    n187,
    n480,
    n513,
    n143
  );


  xor
  g839
  (
    n839,
    n497,
    n207,
    n99,
    n156
  );


  nor
  g840
  (
    KeyWire_0_60,
    n398,
    n504,
    n510,
    n465
  );


  xnor
  g841
  (
    n904,
    n413,
    n142,
    n472,
    n216
  );


  and
  g842
  (
    n900,
    n107,
    n499,
    n508,
    n427
  );


  nand
  g843
  (
    n667,
    n166,
    n198,
    n146,
    n390
  );


  xnor
  g844
  (
    n556,
    n389,
    n127,
    n117,
    n380
  );


  nand
  g845
  (
    n788,
    n158,
    n114,
    n203,
    n511
  );


  nor
  g846
  (
    n767,
    n445,
    n422,
    n455,
    n201
  );


  nand
  g847
  (
    n876,
    n104,
    n441,
    n484,
    n425
  );


  nor
  g848
  (
    n773,
    n206,
    n181,
    n461,
    n159
  );


  and
  g849
  (
    n862,
    n165,
    n463,
    n116,
    n199
  );


  nor
  g850
  (
    n570,
    n129,
    n138,
    n133,
    n128
  );


  and
  g851
  (
    n647,
    n387,
    n183,
    n411,
    n429
  );


  nand
  g852
  (
    n708,
    n438,
    n167,
    n511,
    n187
  );


  xor
  g853
  (
    n634,
    n206,
    n179,
    n194,
    n504
  );


  or
  g854
  (
    n871,
    n430,
    n79,
    n395,
    n384
  );


  nand
  g855
  (
    n735,
    n91,
    n479,
    n97,
    n160
  );


  nand
  g856
  (
    n697,
    n445,
    n124,
    n435,
    n108
  );


  nand
  g857
  (
    n632,
    n493,
    n98,
    n435,
    n433
  );


  xnor
  g858
  (
    n831,
    n102,
    n207,
    n378,
    n514
  );


  xnor
  g859
  (
    n659,
    n174,
    n171,
    n454,
    n116
  );


  or
  g860
  (
    n546,
    n112,
    n382,
    n392,
    n390
  );


  not
  g861
  (
    n909,
    n531
  );


  nand
  g862
  (
    n908,
    n520,
    n530
  );


  nor
  g863
  (
    n910,
    n532,
    n534,
    n908,
    n533
  );


  buf
  g864
  (
    n912,
    n910
  );


  not
  g865
  (
    KeyWire_0_25,
    n910
  );


  nand
  g866
  (
    n915,
    n538,
    n540
  );


  xor
  g867
  (
    n913,
    n539,
    n912,
    n536,
    n537
  );


  nand
  g868
  (
    n914,
    n912,
    n535,
    n911,
    n541
  );


  xor
  g869
  (
    n919,
    n545,
    n546,
    n915
  );


  nand
  g870
  (
    n920,
    n544,
    n550,
    n913
  );


  xor
  g871
  (
    n917,
    n547,
    n915
  );


  nand
  g872
  (
    n916,
    n548,
    n912,
    n549
  );


  or
  g873
  (
    n918,
    n912,
    n543,
    n914,
    n542
  );


  buf
  g874
  (
    n921,
    n917
  );


  not
  g875
  (
    n922,
    n916
  );


  not
  g876
  (
    n927,
    n917
  );


  buf
  g877
  (
    n925,
    n916
  );


  not
  g878
  (
    n928,
    n917
  );


  not
  g879
  (
    n924,
    n917
  );


  buf
  g880
  (
    n926,
    n916
  );


  not
  g881
  (
    n923,
    n916
  );


  or
  g882
  (
    n929,
    n919,
    n918,
    n523,
    n520
  );


  nor
  g883
  (
    n934,
    n921,
    n521,
    n919
  );


  nand
  g884
  (
    n932,
    n921,
    n523,
    n922
  );


  xnor
  g885
  (
    n936,
    n918,
    n522,
    n521
  );


  xor
  g886
  (
    n935,
    n522,
    n521,
    n918,
    n520
  );


  xor
  g887
  (
    n933,
    n922,
    n920,
    n522
  );


  or
  g888
  (
    n930,
    n922,
    n922,
    n523,
    n919
  );


  nand
  g889
  (
    n931,
    n921,
    n921,
    n521,
    n918
  );


  not
  g890
  (
    n937,
    n923
  );


  and
  g891
  (
    n938,
    n930,
    n929,
    n923
  );


  xnor
  g892
  (
    n940,
    n938,
    n933,
    n937
  );


  nor
  g893
  (
    n941,
    n936,
    n920,
    n938
  );


  nor
  g894
  (
    n943,
    n937,
    n934,
    n938
  );


  xnor
  g895
  (
    n942,
    n935,
    n932,
    n931,
    n930
  );


  xnor
  g896
  (
    n939,
    n932,
    n935,
    n931,
    n936
  );


  buf
  g897
  (
    n952,
    n923
  );


  not
  g898
  (
    n953,
    n939
  );


  buf
  g899
  (
    n960,
    n939
  );


  buf
  g900
  (
    n951,
    n940
  );


  buf
  g901
  (
    n955,
    n943
  );


  buf
  g902
  (
    n962,
    n941
  );


  buf
  g903
  (
    KeyWire_0_19,
    n942
  );


  buf
  g904
  (
    n950,
    n941
  );


  not
  g905
  (
    KeyWire_0_49,
    n941
  );


  buf
  g906
  (
    n947,
    n943
  );


  buf
  g907
  (
    n956,
    n942
  );


  not
  g908
  (
    n958,
    n940
  );


  not
  g909
  (
    n957,
    n940
  );


  not
  g910
  (
    n945,
    n940
  );


  buf
  g911
  (
    n954,
    n943
  );


  buf
  g912
  (
    n948,
    n942
  );


  not
  g913
  (
    n946,
    n941
  );


  buf
  g914
  (
    n944,
    n938
  );


  nand
  g915
  (
    n961,
    n939,
    n943,
    n942
  );


  buf
  g916
  (
    n992,
    n949
  );


  buf
  g917
  (
    n988,
    n947
  );


  not
  g918
  (
    n1000,
    n956
  );


  buf
  g919
  (
    n1011,
    n954
  );


  buf
  g920
  (
    n974,
    n948
  );


  not
  g921
  (
    n989,
    n956
  );


  not
  g922
  (
    n972,
    n953
  );


  buf
  g923
  (
    n985,
    n954
  );


  buf
  g924
  (
    n965,
    n946
  );


  not
  g925
  (
    n997,
    n956
  );


  not
  g926
  (
    n998,
    n953
  );


  not
  g927
  (
    n1009,
    n955
  );


  buf
  g928
  (
    n973,
    n947
  );


  not
  g929
  (
    n995,
    n957
  );


  buf
  g930
  (
    n979,
    n952
  );


  not
  g931
  (
    n1007,
    n944
  );


  not
  g932
  (
    n994,
    n948
  );


  not
  g933
  (
    n999,
    n946
  );


  buf
  g934
  (
    n1013,
    n957
  );


  buf
  g935
  (
    n966,
    n945
  );


  buf
  g936
  (
    KeyWire_0_23,
    n945
  );


  buf
  g937
  (
    n1012,
    n951
  );


  not
  g938
  (
    n1008,
    n944
  );


  buf
  g939
  (
    n971,
    n944
  );


  not
  g940
  (
    n987,
    n947
  );


  not
  g941
  (
    n1004,
    n944
  );


  not
  g942
  (
    n967,
    n945
  );


  buf
  g943
  (
    n990,
    n955
  );


  not
  g944
  (
    n976,
    n952
  );


  not
  g945
  (
    n984,
    n946
  );


  buf
  g946
  (
    n977,
    n948
  );


  buf
  g947
  (
    n986,
    n954
  );


  not
  g948
  (
    n980,
    n950
  );


  buf
  g949
  (
    KeyWire_0_10,
    n952
  );


  buf
  g950
  (
    n1005,
    n955
  );


  not
  g951
  (
    n1014,
    n953
  );


  buf
  g952
  (
    n1002,
    n951
  );


  buf
  g953
  (
    n975,
    n949
  );


  buf
  g954
  (
    n982,
    n946
  );


  buf
  g955
  (
    n991,
    n951
  );


  buf
  g956
  (
    n981,
    n950
  );


  buf
  g957
  (
    n969,
    n945
  );


  buf
  g958
  (
    n996,
    n951
  );


  buf
  g959
  (
    n993,
    n953
  );


  not
  g960
  (
    n964,
    n954
  );


  buf
  g961
  (
    n1001,
    n947
  );


  buf
  g962
  (
    n1010,
    n950
  );


  not
  g963
  (
    n1003,
    n949
  );


  not
  g964
  (
    n1016,
    n956
  );


  not
  g965
  (
    n970,
    n949
  );


  not
  g966
  (
    n963,
    n955
  );


  buf
  g967
  (
    n968,
    n950
  );


  buf
  g968
  (
    n1006,
    n952
  );


  not
  g969
  (
    n978,
    n948
  );


  xnor
  g970
  (
    n1024,
    n965,
    n966,
    n963,
    n961
  );


  nor
  g971
  (
    n1020,
    n962,
    n960,
    n959
  );


  xor
  g972
  (
    n1026,
    n959,
    n965,
    n961
  );


  xor
  g973
  (
    n1022,
    n967,
    n964,
    n960,
    n958
  );


  nor
  g974
  (
    n1021,
    n967,
    n965,
    n966,
    n961
  );


  and
  g975
  (
    n1023,
    n963,
    n964,
    n962
  );


  xor
  g976
  (
    n1019,
    n962,
    n957,
    n966,
    n965
  );


  or
  g977
  (
    n1017,
    n962,
    n963,
    n959,
    n958
  );


  nor
  g978
  (
    n1025,
    n958,
    n964,
    n963,
    n957
  );


  xnor
  g979
  (
    n1018,
    n958,
    n959,
    n966,
    n960
  );


  xor
  g980
  (
    n1030,
    n968,
    n969
  );


  and
  g981
  (
    n1029,
    n969,
    n971,
    n1020
  );


  nor
  g982
  (
    n1032,
    n967,
    n968,
    n970
  );


  or
  g983
  (
    n1028,
    n1018,
    n969,
    n970
  );


  xor
  g984
  (
    n1031,
    n1021,
    n1017,
    n969,
    n970
  );


  nand
  g985
  (
    n1027,
    n967,
    n1019,
    n1020,
    n968
  );


  not
  g986
  (
    n1035,
    n1032
  );


  buf
  g987
  (
    n1036,
    n1029
  );


  buf
  g988
  (
    n1037,
    n1030
  );


  not
  g989
  (
    n1039,
    n1027
  );


  buf
  g990
  (
    n1034,
    n1032
  );


  not
  g991
  (
    n1038,
    n1028
  );


  not
  g992
  (
    KeyWire_0_54,
    n1031
  );


  buf
  g993
  (
    n1033,
    n1031
  );


  nand
  g994
  (
    n1044,
    n972,
    n986,
    n1038,
    n973
  );


  xor
  g995
  (
    n1071,
    n1039,
    n1040,
    n989,
    n987
  );


  nor
  g996
  (
    n1048,
    n988,
    n1035,
    n979
  );


  xor
  g997
  (
    n1054,
    n1039,
    n524,
    n990,
    n984
  );


  nor
  g998
  (
    n1042,
    n983,
    n988,
    n974,
    n1035
  );


  xor
  g999
  (
    n1072,
    n975,
    n992,
    n971,
    n982
  );


  nor
  g1000
  (
    n1052,
    n981,
    n1037,
    n990,
    n1034
  );


  and
  g1001
  (
    n1050,
    n980,
    n977,
    n989,
    n1039
  );


  nor
  g1002
  (
    n1064,
    n1039,
    n984,
    n975
  );


  or
  g1003
  (
    n1059,
    n1037,
    n972,
    n524,
    n976
  );


  or
  g1004
  (
    n1062,
    n1036,
    n987,
    n1033,
    n552
  );


  nor
  g1005
  (
    n1066,
    n993,
    n989,
    n978,
    n981
  );


  and
  g1006
  (
    n1047,
    n991,
    n974,
    n1040,
    n973
  );


  and
  g1007
  (
    n1061,
    n985,
    n977,
    n1034,
    n983
  );


  xor
  g1008
  (
    n1057,
    n980,
    n986,
    n988,
    n1040
  );


  and
  g1009
  (
    n1053,
    n982,
    n984,
    n973,
    n972
  );


  xor
  g1010
  (
    n1041,
    n1035,
    n979,
    n1036,
    n976
  );


  xnor
  g1011
  (
    n1051,
    n975,
    n551,
    n987,
    n985
  );


  xnor
  g1012
  (
    n1056,
    n1038,
    n985,
    n977,
    n980
  );


  and
  g1013
  (
    n1068,
    n524,
    n1038,
    n983,
    n987
  );


  xnor
  g1014
  (
    n1046,
    n981,
    n978,
    n993
  );


  xor
  g1015
  (
    KeyWire_0_33,
    n972,
    n980,
    n1038,
    n553
  );


  and
  g1016
  (
    n1043,
    n524,
    n992,
    n979,
    n982
  );


  xor
  g1017
  (
    n1058,
    n1033,
    n971,
    n983,
    n975
  );


  xor
  g1018
  (
    n1070,
    n981,
    n974,
    n1036,
    n978
  );


  xnor
  g1019
  (
    n1060,
    n986,
    n1033,
    n978
  );


  xor
  g1020
  (
    n1065,
    n990,
    n976,
    n988,
    n982
  );


  and
  g1021
  (
    n1069,
    n1034,
    n1040,
    n973,
    n990
  );


  xor
  g1022
  (
    n1049,
    n976,
    n974,
    n991,
    n992
  );


  xor
  g1023
  (
    n1055,
    n991,
    n1037,
    n985
  );


  or
  g1024
  (
    n1067,
    n989,
    n991,
    n986,
    n1036
  );


  xor
  g1025
  (
    n1045,
    n992,
    n977,
    n979,
    n1034
  );


  xor
  g1026
  (
    n1116,
    n782,
    n1062,
    n603,
    n792
  );


  or
  g1027
  (
    n1113,
    n735,
    n736,
    n1043,
    n619
  );


  nand
  g1028
  (
    n1151,
    n1043,
    n798,
    n738,
    n872
  );


  or
  g1029
  (
    n1171,
    n617,
    n803,
    n645,
    n1046
  );


  or
  g1030
  (
    n1174,
    n1052,
    n689,
    n828,
    n1064
  );


  or
  g1031
  (
    n1079,
    n831,
    n1063,
    n1059,
    n627
  );


  nand
  g1032
  (
    n1078,
    n837,
    n1064,
    n1062,
    n620
  );


  and
  g1033
  (
    n1074,
    n676,
    n585,
    n783,
    n564
  );


  nor
  g1034
  (
    n1177,
    n829,
    n1063,
    n720,
    n723
  );


  nor
  g1035
  (
    n1143,
    n594,
    n838,
    n573,
    n1045
  );


  xor
  g1036
  (
    n1155,
    n725,
    n1049,
    n652,
    n681
  );


  or
  g1037
  (
    n1110,
    n582,
    n849,
    n698,
    n751
  );


  nor
  g1038
  (
    n1130,
    n1041,
    n1067,
    n571,
    n867
  );


  xnor
  g1039
  (
    n1077,
    n561,
    n661,
    n635,
    n687
  );


  and
  g1040
  (
    n1081,
    n823,
    n760,
    n871,
    n593
  );


  xor
  g1041
  (
    n1105,
    n748,
    n1053,
    n852,
    n622
  );


  xor
  g1042
  (
    n1121,
    n606,
    n1042,
    n670,
    n776
  );


  and
  g1043
  (
    n1088,
    n655,
    n664,
    n638,
    n712
  );


  xor
  g1044
  (
    n1163,
    n879,
    n706,
    n686,
    n809
  );


  and
  g1045
  (
    n1172,
    n814,
    n1057,
    n1058,
    n604
  );


  xnor
  g1046
  (
    n1086,
    n1065,
    n568,
    n589,
    n806
  );


  xnor
  g1047
  (
    n1156,
    n768,
    n673,
    n710,
    n636
  );


  nor
  g1048
  (
    n1099,
    n808,
    n767,
    n764,
    n1051
  );


  nor
  g1049
  (
    n1165,
    n1056,
    n844,
    n1049,
    n816
  );


  xor
  g1050
  (
    KeyWire_0_55,
    n759,
    n684,
    n729,
    n833
  );


  or
  g1051
  (
    n1139,
    n1060,
    n878,
    n810,
    n777
  );


  nand
  g1052
  (
    n1176,
    n790,
    n572,
    n1068,
    n818
  );


  xnor
  g1053
  (
    n1109,
    n1049,
    n1060,
    n701,
    n1052
  );


  nand
  g1054
  (
    KeyWire_0_27,
    n774,
    n1051,
    n567,
    n860
  );


  or
  g1055
  (
    n1140,
    n731,
    n1053,
    n804,
    n1052
  );


  and
  g1056
  (
    KeyWire_0_40,
    n682,
    n794,
    n665,
    n1044
  );


  or
  g1057
  (
    n1104,
    n850,
    n574,
    n609,
    n1067
  );


  xor
  g1058
  (
    n1117,
    n854,
    n740,
    n737,
    n1066
  );


  xnor
  g1059
  (
    n1160,
    n826,
    n1056,
    n679,
    n1048
  );


  and
  g1060
  (
    n1087,
    n1057,
    n784,
    n646,
    n575
  );


  or
  g1061
  (
    n1173,
    n709,
    n598,
    n697,
    n1059
  );


  xor
  g1062
  (
    n1136,
    n848,
    n752,
    n868,
    n874
  );


  nand
  g1063
  (
    n1091,
    n749,
    n692,
    n1050,
    n1053
  );


  xor
  g1064
  (
    n1092,
    n1061,
    n1048,
    n576,
    n663
  );


  or
  g1065
  (
    n1094,
    n578,
    n1051,
    n822,
    n649
  );


  or
  g1066
  (
    n1076,
    n728,
    n858,
    n597,
    n1056
  );


  xnor
  g1067
  (
    n1149,
    n626,
    n743,
    n836,
    n866
  );


  and
  g1068
  (
    n1133,
    n1058,
    n869,
    n827,
    n650
  );


  xor
  g1069
  (
    n1178,
    n654,
    n861,
    n842,
    n602
  );


  xnor
  g1070
  (
    n1168,
    n702,
    n713,
    n840,
    n680
  );


  xnor
  g1071
  (
    n1119,
    n770,
    n715,
    n660,
    n586
  );


  xnor
  g1072
  (
    n1102,
    n1057,
    n820,
    n562,
    n755
  );


  and
  g1073
  (
    n1152,
    n1063,
    n704,
    n730,
    n719
  );


  nor
  g1074
  (
    n1073,
    n560,
    n714,
    n667,
    n747
  );


  or
  g1075
  (
    n1125,
    n726,
    n648,
    n781,
    n1067
  );


  xnor
  g1076
  (
    n1107,
    n1066,
    n640,
    n583,
    n1056
  );


  nand
  g1077
  (
    n1162,
    n769,
    n778,
    n685,
    n839
  );


  and
  g1078
  (
    n1122,
    n847,
    n1043,
    n559,
    n1054
  );


  or
  g1079
  (
    n1100,
    n787,
    n1045,
    n811
  );


  nor
  g1080
  (
    n1128,
    n788,
    n853,
    n718,
    n802
  );


  xor
  g1081
  (
    n1082,
    n876,
    n625,
    n555,
    n1047
  );


  nor
  g1082
  (
    n1118,
    n1043,
    n841,
    n717,
    n616
  );


  nor
  g1083
  (
    n1138,
    n789,
    n851,
    n830,
    n780
  );


  xnor
  g1084
  (
    n1153,
    n1046,
    n668,
    n721,
    n1050
  );


  xor
  g1085
  (
    n1083,
    n639,
    n581,
    n815,
    n596
  );


  xor
  g1086
  (
    n1134,
    n800,
    n1055,
    n587,
    n1048
  );


  or
  g1087
  (
    n1158,
    n753,
    n1041,
    n843,
    n677
  );


  nand
  g1088
  (
    n1101,
    n565,
    n584,
    n1060,
    n666
  );


  nor
  g1089
  (
    n1132,
    n672,
    n577,
    n628,
    n1066
  );


  nor
  g1090
  (
    n1142,
    n1065,
    n659,
    n870,
    n1062
  );


  xor
  g1091
  (
    n1169,
    n556,
    n656,
    n845,
    n591
  );


  nor
  g1092
  (
    n1159,
    n631,
    n641,
    n1057,
    n653
  );


  nor
  g1093
  (
    n1120,
    n1063,
    n807,
    n1045,
    n825
  );


  xnor
  g1094
  (
    n1126,
    n855,
    n621,
    n1064,
    n592
  );


  nand
  g1095
  (
    n1144,
    n1064,
    n745,
    n1049,
    n1046
  );


  xnor
  g1096
  (
    n1108,
    n599,
    n727,
    n793,
    n644
  );


  xor
  g1097
  (
    n1111,
    n796,
    n791,
    n595,
    n766
  );


  and
  g1098
  (
    n1181,
    n691,
    n657,
    n824,
    n744
  );


  xor
  g1099
  (
    n1137,
    n590,
    n683,
    n607,
    n856
  );


  xor
  g1100
  (
    n1179,
    n754,
    n612,
    n630,
    n569
  );


  xor
  g1101
  (
    n1103,
    n1044,
    n1055,
    n554,
    n733
  );


  xnor
  g1102
  (
    n1095,
    n711,
    n690,
    n1041,
    n832
  );


  or
  g1103
  (
    n1175,
    n699,
    n1047,
    n865,
    n724
  );


  or
  g1104
  (
    n1147,
    n757,
    n1067,
    n694,
    n674
  );


  xnor
  g1105
  (
    n1075,
    n614,
    n746,
    n863,
    n608
  );


  nand
  g1106
  (
    n1170,
    n615,
    n819,
    n813,
    n1046
  );


  nor
  g1107
  (
    n1123,
    n765,
    n1065,
    n1052,
    n741
  );


  or
  g1108
  (
    n1096,
    n643,
    n675,
    n1051,
    n618
  );


  nor
  g1109
  (
    n1146,
    n763,
    n864,
    n1055,
    n1054
  );


  xor
  g1110
  (
    n1167,
    n605,
    n821,
    n786,
    n1054
  );


  or
  g1111
  (
    n1150,
    n1061,
    n739,
    n875,
    n563
  );


  or
  g1112
  (
    n1157,
    n801,
    n797,
    n1058,
    n756
  );


  nor
  g1113
  (
    n1090,
    n750,
    n1068,
    n812,
    n742
  );


  nand
  g1114
  (
    n1127,
    n880,
    n805,
    n732,
    n634
  );


  and
  g1115
  (
    n1114,
    n611,
    n734,
    n632,
    n846
  );


  or
  g1116
  (
    n1097,
    n1061,
    n637,
    n633,
    n1048
  );


  xor
  g1117
  (
    n1164,
    n773,
    n795,
    n1044,
    n1065
  );


  nor
  g1118
  (
    n1098,
    n613,
    n873,
    n1059,
    n566
  );


  or
  g1119
  (
    n1148,
    n580,
    n669,
    n775,
    n558
  );


  xnor
  g1120
  (
    n1129,
    n817,
    n658,
    n662,
    n1042
  );


  nor
  g1121
  (
    n1154,
    n1044,
    n610,
    n1050
  );


  or
  g1122
  (
    n1161,
    n557,
    n835,
    n623,
    n1062
  );


  nand
  g1123
  (
    n1124,
    n772,
    n708,
    n722,
    n705
  );


  and
  g1124
  (
    n1180,
    n579,
    n834,
    n1042,
    n688
  );


  xnor
  g1125
  (
    n1084,
    n799,
    n1059,
    n857,
    n624
  );


  xnor
  g1126
  (
    n1112,
    n1066,
    n1053,
    n716,
    n629
  );


  or
  g1127
  (
    n1080,
    n877,
    n1054,
    n1061,
    n700
  );


  xor
  g1128
  (
    n1089,
    n1058,
    n1047,
    n771,
    n600
  );


  nand
  g1129
  (
    n1135,
    n785,
    n642,
    n678,
    n1047
  );


  and
  g1130
  (
    n1131,
    n651,
    n703,
    n1055,
    n862
  );


  xnor
  g1131
  (
    n1115,
    n696,
    n1042,
    n758,
    n707
  );


  nor
  g1132
  (
    n1106,
    n570,
    n693,
    n762,
    n779
  );


  nor
  g1133
  (
    n1093,
    n601,
    n671,
    n588,
    n695
  );


  and
  g1134
  (
    n1166,
    n1060,
    n761,
    n647,
    n859
  );


  or
  g1135
  (
    n1182,
    n1073,
    n1074,
    n1075,
    n1076
  );


  not
  g1136
  (
    n1185,
    n1079
  );


  not
  g1137
  (
    n1184,
    n1182
  );


  xor
  g1138
  (
    n1183,
    n1077,
    n1182,
    n1078
  );


  nand
  g1139
  (
    n1186,
    n889,
    n881,
    n883,
    n888
  );


  xnor
  g1140
  (
    n1196,
    n994,
    n1184,
    n898
  );


  xor
  g1141
  (
    n1192,
    n884,
    n1183,
    n525,
    n895
  );


  nor
  g1142
  (
    n1189,
    n885,
    n1080,
    n900,
    n893
  );


  xor
  g1143
  (
    n1194,
    n891,
    n896,
    n1185,
    n899
  );


  and
  g1144
  (
    n1193,
    n892,
    n897,
    n1184,
    n1068
  );


  and
  g1145
  (
    n1190,
    n1069,
    n1183,
    n994,
    n887
  );


  or
  g1146
  (
    n1191,
    n1185,
    n1183,
    n1069,
    n525
  );


  xor
  g1147
  (
    n1187,
    n993,
    n1081,
    n1068,
    n894
  );


  nand
  g1148
  (
    KeyWire_0_48,
    n525,
    n901,
    n1184,
    n1185
  );


  xnor
  g1149
  (
    n1195,
    n886,
    n1183,
    n882,
    n890
  );


  or
  g1150
  (
    n1198,
    n1195,
    n1084
  );


  xnor
  g1151
  (
    n1197,
    n1082,
    n1083,
    n1196
  );


  and
  g1152
  (
    n1204,
    n1101,
    n1102,
    n1197,
    n1198
  );


  and
  g1153
  (
    n1203,
    n1197,
    n1198,
    n1099,
    n1098
  );


  xnor
  g1154
  (
    n1200,
    n1090,
    n1104,
    n1198,
    n1091
  );


  nand
  g1155
  (
    n1199,
    n1105,
    n1198,
    n1095,
    n1086
  );


  xnor
  g1156
  (
    n1202,
    n1093,
    n1097,
    n1087,
    n1092
  );


  and
  g1157
  (
    n1205,
    n1088,
    n1085,
    n1089,
    n1094
  );


  xor
  g1158
  (
    n1201,
    n1096,
    n1197,
    n1103,
    n1100
  );


  and
  g1159
  (
    n1214,
    n909,
    n925,
    n1204
  );


  and
  g1160
  (
    n1211,
    n1199,
    n1106,
    n1111,
    n924
  );


  xor
  g1161
  (
    n1208,
    n1205,
    n908,
    n924
  );


  nor
  g1162
  (
    n1207,
    n1114,
    n924,
    n909,
    n908
  );


  or
  g1163
  (
    n1213,
    n925,
    n1113,
    n1108,
    n1205
  );


  xor
  g1164
  (
    KeyWire_0_1,
    n1185,
    n1109,
    n1112,
    n525
  );


  xnor
  g1165
  (
    KeyWire_0_30,
    n925,
    n1201,
    n909,
    n924
  );


  nand
  g1166
  (
    n1209,
    n1110,
    n1202,
    n1200,
    n923
  );


  xor
  g1167
  (
    n1212,
    n1107,
    n1203,
    n1204,
    n909
  );


  or
  g1168
  (
    n1221,
    n1207,
    n1209,
    n529,
    n1071
  );


  xor
  g1169
  (
    n1224,
    n1071,
    n526,
    n1211,
    n1209
  );


  or
  g1170
  (
    n1218,
    n529,
    n529,
    n527,
    n1206
  );


  xnor
  g1171
  (
    n1216,
    n527,
    n1069,
    n528,
    n1072
  );


  xnor
  g1172
  (
    n1215,
    n527,
    n1069,
    n1208,
    n528
  );


  xnor
  g1173
  (
    n1217,
    n1210,
    n1210,
    n1072,
    n529
  );


  xnor
  g1174
  (
    n1222,
    n1070,
    n1070,
    n526,
    n1072
  );


  nor
  g1175
  (
    n1219,
    n1208,
    n1071,
    n526,
    n1072
  );


  nand
  g1176
  (
    n1223,
    n1207,
    n1070,
    n1071,
    n528
  );


  nor
  g1177
  (
    n1220,
    n526,
    n528,
    n527,
    n1070
  );


  xnor
  g1178
  (
    n1230,
    n1218,
    n1224,
    n1217,
    n1123
  );


  nand
  g1179
  (
    n1228,
    n1139,
    n1129,
    n1137,
    n1116
  );


  xor
  g1180
  (
    n1231,
    n1117,
    n1119,
    n1219,
    n1115
  );


  nand
  g1181
  (
    n1233,
    n1222,
    n1118,
    n1223,
    n1125
  );


  nor
  g1182
  (
    n1225,
    n1127,
    n1122,
    n1131,
    n1136
  );


  and
  g1183
  (
    n1226,
    n1140,
    n1221,
    n1138,
    n1120
  );


  nor
  g1184
  (
    n1227,
    n1133,
    n1220,
    n1126,
    n1121
  );


  or
  g1185
  (
    n1229,
    n1135,
    n1130,
    n1141,
    n1132
  );


  and
  g1186
  (
    n1232,
    n1216,
    n1124,
    n1134,
    n1128
  );


  or
  g1187
  (
    n1251,
    n1229,
    n223,
    n226,
    n222
  );


  xor
  g1188
  (
    n1248,
    n227,
    n225,
    n230,
    n1227
  );


  nand
  g1189
  (
    n1247,
    n222,
    n926,
    n227,
    n1022
  );


  xor
  g1190
  (
    n1239,
    n222,
    n1226,
    n1142,
    n928
  );


  nand
  g1191
  (
    n1245,
    n927,
    n1225,
    n1021,
    n228
  );


  xnor
  g1192
  (
    n1249,
    n229,
    n229,
    n1143,
    n221
  );


  and
  g1193
  (
    n1243,
    n927,
    n229,
    n1228
  );


  nor
  g1194
  (
    n1242,
    n230,
    n224,
    n926,
    n928
  );


  nand
  g1195
  (
    n1238,
    n1227,
    n1229,
    n225,
    n223
  );


  and
  g1196
  (
    KeyWire_0_6,
    n228,
    n223,
    n226
  );


  xnor
  g1197
  (
    n1240,
    n1022,
    n228,
    n1228,
    n1229
  );


  nor
  g1198
  (
    n1250,
    n1229,
    n230,
    n927,
    n1226
  );


  and
  g1199
  (
    n1236,
    n1227,
    n226,
    n227,
    n926
  );


  nor
  g1200
  (
    n1237,
    n1226,
    n926,
    n1228,
    n224
  );


  or
  g1201
  (
    n1241,
    n226,
    n228,
    n227,
    n221
  );


  nor
  g1202
  (
    n1244,
    n1226,
    n927,
    n225,
    n928
  );


  or
  g1203
  (
    n1234,
    n222,
    n224,
    n1225,
    n1228
  );


  or
  g1204
  (
    n1246,
    n230,
    n225,
    n224,
    n1227
  );


  buf
  g1205
  (
    n1257,
    n1230
  );


  buf
  g1206
  (
    n1260,
    n1232
  );


  not
  g1207
  (
    n1258,
    n1244
  );


  not
  g1208
  (
    n1263,
    n1239
  );


  and
  g1209
  (
    n1253,
    n1149,
    n1146,
    n1249,
    n1238
  );


  nor
  g1210
  (
    n1254,
    n1148,
    n1231
  );


  nor
  g1211
  (
    n1259,
    n1247,
    n1151,
    n1245,
    n1147
  );


  xnor
  g1212
  (
    n1252,
    n1230,
    n1150,
    n1246,
    n1233
  );


  nand
  g1213
  (
    n1256,
    n1145,
    n1232,
    n1231,
    n1233
  );


  and
  g1214
  (
    n1261,
    n1242,
    n1240,
    n1233,
    n1232
  );


  and
  g1215
  (
    n1262,
    n1230,
    n1241,
    n1248,
    n1243
  );


  xor
  g1216
  (
    n1255,
    n1230,
    n1232,
    n1233,
    n1144
  );


  nor
  g1217
  (
    n1267,
    n1259,
    n1255,
    n1001,
    n1009
  );


  and
  g1218
  (
    n1265,
    n1014,
    n1016,
    n1255,
    n1214
  );


  xor
  g1219
  (
    n1278,
    n1254,
    n1012,
    n1258,
    n1002
  );


  nand
  g1220
  (
    n1296,
    n1260,
    n1000,
    n1262,
    n997
  );


  nand
  g1221
  (
    n1272,
    n1252,
    n1260,
    n1005
  );


  or
  g1222
  (
    n1274,
    n1011,
    n1015,
    n1213
  );


  xor
  g1223
  (
    n1294,
    n997,
    n1212,
    n1012,
    n998
  );


  nor
  g1224
  (
    n1276,
    n1007,
    n1008,
    n1003,
    n1009
  );


  or
  g1225
  (
    n1280,
    n1251,
    n1007,
    n999,
    n1008
  );


  or
  g1226
  (
    n1277,
    n1006,
    n1001,
    n1261
  );


  xnor
  g1227
  (
    n1264,
    n1013,
    n1012,
    n1015,
    n1258
  );


  nand
  g1228
  (
    n1286,
    n1007,
    n1254,
    n1258,
    n1010
  );


  nand
  g1229
  (
    n1283,
    n1010,
    n1253,
    n1262
  );


  xnor
  g1230
  (
    n1281,
    n1252,
    n1261,
    n1003,
    n1005
  );


  xnor
  g1231
  (
    n1282,
    n999,
    n998,
    n1256,
    n995
  );


  xor
  g1232
  (
    n1269,
    n1214,
    n1260,
    n1254,
    n1002
  );


  nand
  g1233
  (
    n1301,
    n1253,
    n999,
    n904,
    n1013
  );


  xor
  g1234
  (
    n1279,
    n1004,
    n995,
    n999,
    n994
  );


  xnor
  g1235
  (
    n1297,
    n1260,
    n1010,
    n1255,
    n1003
  );


  or
  g1236
  (
    n1300,
    n996,
    n1009,
    n1257,
    n1015
  );


  or
  g1237
  (
    n1290,
    n1213,
    n995,
    n1006,
    n1012
  );


  xor
  g1238
  (
    n1285,
    n1014,
    n1254,
    n906,
    n998
  );


  xnor
  g1239
  (
    n1289,
    n1259,
    n1262,
    n1261
  );


  nor
  g1240
  (
    n1273,
    n1211,
    n1011,
    n997,
    n1250
  );


  xor
  g1241
  (
    n1291,
    n1008,
    n1258,
    n1007,
    n1003
  );


  nor
  g1242
  (
    n1292,
    n1011,
    n1259,
    n996,
    n1256
  );


  and
  g1243
  (
    n1287,
    n1256,
    n1001,
    n907,
    n902
  );


  or
  g1244
  (
    n1288,
    n995,
    n906,
    n1008,
    n1014
  );


  xnor
  g1245
  (
    n1266,
    n1257,
    n1002,
    n994,
    n1004
  );


  or
  g1246
  (
    n1284,
    n1004,
    n1253,
    n905
  );


  and
  g1247
  (
    n1270,
    n907,
    n996,
    n1005,
    n1010
  );


  and
  g1248
  (
    n1299,
    n1257,
    n1212,
    n1013,
    n1252
  );


  xor
  g1249
  (
    n1271,
    n1006,
    n1011,
    n1256,
    n1016
  );


  xnor
  g1250
  (
    n1295,
    n928,
    n997,
    n1014,
    n1252
  );


  nor
  g1251
  (
    n1298,
    n1000,
    n1016,
    n1255,
    n1257
  );


  xor
  g1252
  (
    n1268,
    n1016,
    n1013,
    n1259,
    n1002
  );


  nor
  g1253
  (
    n1293,
    n1006,
    n1009,
    n1000
  );


  nand
  g1254
  (
    n1275,
    n996,
    n903,
    n998,
    n1004
  );


  not
  g1255
  (
    n1313,
    n1264
  );


  buf
  g1256
  (
    n1309,
    n1263
  );


  buf
  g1257
  (
    n1304,
    n1266
  );


  buf
  g1258
  (
    n1307,
    n1275
  );


  buf
  g1259
  (
    n1302,
    n1269
  );


  buf
  g1260
  (
    n1303,
    n1263
  );


  buf
  g1261
  (
    n1312,
    n1273
  );


  buf
  g1262
  (
    n1310,
    n1268
  );


  buf
  g1263
  (
    n1305,
    n1263
  );


  buf
  g1264
  (
    n1306,
    n1271
  );


  or
  g1265
  (
    n1308,
    n1265,
    n1263
  );


  xnor
  g1266
  (
    n1311,
    n1274,
    n1270,
    n1267,
    n1272
  );


  or
  g1267
  (
    n1328,
    n1155,
    n1303,
    n1279,
    n1305
  );


  nor
  g1268
  (
    n1324,
    n1301,
    n1304,
    n1152,
    n1305
  );


  or
  g1269
  (
    n1322,
    n1289,
    n1285,
    n1283,
    n1282
  );


  and
  g1270
  (
    n1327,
    n1299,
    n1301,
    n1300,
    n1281
  );


  nor
  g1271
  (
    n1326,
    n1292,
    n1293,
    n1305,
    n1303
  );


  or
  g1272
  (
    n1318,
    n1157,
    n1298,
    n1304,
    n1286
  );


  xor
  g1273
  (
    n1317,
    n1276,
    n1297,
    n1291,
    n1302
  );


  nor
  g1274
  (
    n1315,
    n1303,
    n1291,
    n1296,
    n1302
  );


  nor
  g1275
  (
    n1325,
    n1299,
    n1298,
    n1294,
    n1278
  );


  xnor
  g1276
  (
    n1319,
    n1294,
    n1284,
    n1277,
    n1288
  );


  nand
  g1277
  (
    n1316,
    n1293,
    n1300,
    n1303,
    n1286
  );


  nand
  g1278
  (
    n1321,
    n1297,
    n1290,
    n1287,
    n1302
  );


  xnor
  g1279
  (
    n1320,
    n1280,
    n1304,
    n1289,
    n1292
  );


  xnor
  g1280
  (
    n1314,
    n1295,
    n1290,
    n1304,
    n1302
  );


  xnor
  g1281
  (
    n1323,
    n1296,
    n1305,
    n1156,
    n1154
  );


  xnor
  g1282
  (
    n1329,
    n1287,
    n1288,
    n1295,
    n1153
  );


  nor
  g1283
  (
    n1336,
    n1306,
    n1310,
    n1308,
    n1314
  );


  and
  g1284
  (
    n1333,
    n1310,
    n1309,
    n1311,
    n1316
  );


  xnor
  g1285
  (
    n1337,
    n1309,
    n1308,
    n1306,
    n1315
  );


  xnor
  g1286
  (
    n1331,
    n1310,
    n1310,
    n1306,
    n1307
  );


  xnor
  g1287
  (
    n1334,
    n1309,
    n1307,
    n1317,
    n1311
  );


  xor
  g1288
  (
    n1335,
    n1308,
    n1316,
    n1314,
    n1311
  );


  xor
  g1289
  (
    n1332,
    n1308,
    n1307,
    n1309
  );


  and
  g1290
  (
    n1330,
    n1306,
    n1311,
    n1315,
    n1317
  );


  buf
  g1291
  (
    n1339,
    n1336
  );


  not
  g1292
  (
    n1338,
    n1335
  );


  xnor
  g1293
  (
    n1340,
    n1177,
    n1339,
    n1169
  );


  nand
  g1294
  (
    n1346,
    n1175,
    n1167,
    n1171,
    n1162
  );


  nor
  g1295
  (
    n1345,
    n1337,
    n1338,
    n1161,
    n1172
  );


  nor
  g1296
  (
    n1347,
    n1165,
    n1180,
    n1339,
    n1158
  );


  and
  g1297
  (
    n1343,
    n1163,
    n1179,
    n1178,
    n1176
  );


  nor
  g1298
  (
    n1342,
    n1159,
    n1164,
    n1173,
    n1338
  );


  or
  g1299
  (
    n1344,
    n1339,
    n1174,
    n1338,
    n1170
  );


  and
  g1300
  (
    n1341,
    n1160,
    n1168,
    n1338,
    n1166
  );


  xnor
  g1301
  (
    n1362,
    n1319,
    n1345,
    n1343,
    n1181
  );


  or
  g1302
  (
    n1351,
    n1341,
    n1342,
    n1312
  );


  nor
  g1303
  (
    n1361,
    n1323,
    n1343,
    n1344,
    n1313
  );


  xnor
  g1304
  (
    n1359,
    n1321,
    n1344,
    n1328,
    n1342
  );


  nor
  g1305
  (
    n1353,
    n1318,
    n1328,
    n1329,
    n1344
  );


  xor
  g1306
  (
    n1348,
    n1026,
    n1327,
    n1347
  );


  nand
  g1307
  (
    n1349,
    n1345,
    n1325,
    n1322
  );


  or
  g1308
  (
    n1352,
    n1024,
    n1025,
    n1329,
    n1324
  );


  and
  g1309
  (
    n1358,
    n1342,
    n1323,
    n1347,
    n1023
  );


  or
  g1310
  (
    n1356,
    n1026,
    n1327,
    n1319,
    n1341
  );


  nor
  g1311
  (
    n1354,
    n1318,
    n1343,
    n1312,
    n1346
  );


  xnor
  g1312
  (
    n1357,
    n1321,
    n1346,
    n1341,
    n1324
  );


  and
  g1313
  (
    n1363,
    n1312,
    n1313,
    n1320,
    n1345
  );


  xnor
  g1314
  (
    n1360,
    n1320,
    n1313,
    n1322,
    n1347
  );


  nor
  g1315
  (
    n1350,
    n1326,
    n1346,
    n1023,
    n1025
  );


  xor
  g1316
  (
    n1355,
    n1340,
    n1024,
    n1313,
    n1326
  );


  or
  g1317
  (
    n1364,
    n1349,
    n1362,
    n1355,
    n1357
  );


  nor
  g1318
  (
    n1365,
    n1360,
    n1351,
    n1350,
    n1352
  );


  xnor
  g1319
  (
    n1366,
    n1358,
    n1363,
    n1356,
    n1354
  );


  or
  g1320
  (
    n1367,
    n1348,
    n1361,
    n1359,
    n1353
  );


  xor
  KeyGate_0_0
  (
    n821,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1206,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n65,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n389,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n107,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n704,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1235,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n137,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n462,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n465,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n1015,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n95,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n192,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n191,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n764,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n678,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n610,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n804,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n378,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n959,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n569,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n341,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n51,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n983,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n879,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n911,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n675,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1145,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n550,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n750,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1210,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n337,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n294,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n1063,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n662,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n560,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n403,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n507,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n452,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n827,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n1085,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n611,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n419,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n774,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n595,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n155,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n264,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n855,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1188,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n949,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n880,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n426,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n212,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n266,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n1040,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n1141,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n75,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n464,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n53,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n646,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n840,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n406,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n733,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n272,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

