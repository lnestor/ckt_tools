// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1654_26_3 written by SynthGen on 2021/06/15 15:04:54
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1654_26_3 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20,
 n1470, n1534, n1536, n1531, n1530, n1533, n1549, n1558,
 n1563, n1559, n1560, n1566, n1550, n1562, n1561, n1565,
 n1551, n1554, n1567, n1553, n1564, n1664, n1673, n1662,
 n1669, n1674, n1667, n1666, n1671, n1672, n1670, n1663,
 n1665, n1668);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20;

output n1470, n1534, n1536, n1531, n1530, n1533, n1549, n1558,
 n1563, n1559, n1560, n1566, n1550, n1562, n1561, n1565,
 n1551, n1554, n1567, n1553, n1564, n1664, n1673, n1662,
 n1669, n1674, n1667, n1666, n1671, n1672, n1670, n1663,
 n1665, n1668;

wire n21, n22, n23, n24, n25, n26, n27, n28,
 n29, n30, n31, n32, n33, n34, n35, n36,
 n37, n38, n39, n40, n41, n42, n43, n44,
 n45, n46, n47, n48, n49, n50, n51, n52,
 n53, n54, n55, n56, n57, n58, n59, n60,
 n61, n62, n63, n64, n65, n66, n67, n68,
 n69, n70, n71, n72, n73, n74, n75, n76,
 n77, n78, n79, n80, n81, n82, n83, n84,
 n85, n86, n87, n88, n89, n90, n91, n92,
 n93, n94, n95, n96, n97, n98, n99, n100,
 n101, n102, n103, n104, n105, n106, n107, n108,
 n109, n110, n111, n112, n113, n114, n115, n116,
 n117, n118, n119, n120, n121, n122, n123, n124,
 n125, n126, n127, n128, n129, n130, n131, n132,
 n133, n134, n135, n136, n137, n138, n139, n140,
 n141, n142, n143, n144, n145, n146, n147, n148,
 n149, n150, n151, n152, n153, n154, n155, n156,
 n157, n158, n159, n160, n161, n162, n163, n164,
 n165, n166, n167, n168, n169, n170, n171, n172,
 n173, n174, n175, n176, n177, n178, n179, n180,
 n181, n182, n183, n184, n185, n186, n187, n188,
 n189, n190, n191, n192, n193, n194, n195, n196,
 n197, n198, n199, n200, n201, n202, n203, n204,
 n205, n206, n207, n208, n209, n210, n211, n212,
 n213, n214, n215, n216, n217, n218, n219, n220,
 n221, n222, n223, n224, n225, n226, n227, n228,
 n229, n230, n231, n232, n233, n234, n235, n236,
 n237, n238, n239, n240, n241, n242, n243, n244,
 n245, n246, n247, n248, n249, n250, n251, n252,
 n253, n254, n255, n256, n257, n258, n259, n260,
 n261, n262, n263, n264, n265, n266, n267, n268,
 n269, n270, n271, n272, n273, n274, n275, n276,
 n277, n278, n279, n280, n281, n282, n283, n284,
 n285, n286, n287, n288, n289, n290, n291, n292,
 n293, n294, n295, n296, n297, n298, n299, n300,
 n301, n302, n303, n304, n305, n306, n307, n308,
 n309, n310, n311, n312, n313, n314, n315, n316,
 n317, n318, n319, n320, n321, n322, n323, n324,
 n325, n326, n327, n328, n329, n330, n331, n332,
 n333, n334, n335, n336, n337, n338, n339, n340,
 n341, n342, n343, n344, n345, n346, n347, n348,
 n349, n350, n351, n352, n353, n354, n355, n356,
 n357, n358, n359, n360, n361, n362, n363, n364,
 n365, n366, n367, n368, n369, n370, n371, n372,
 n373, n374, n375, n376, n377, n378, n379, n380,
 n381, n382, n383, n384, n385, n386, n387, n388,
 n389, n390, n391, n392, n393, n394, n395, n396,
 n397, n398, n399, n400, n401, n402, n403, n404,
 n405, n406, n407, n408, n409, n410, n411, n412,
 n413, n414, n415, n416, n417, n418, n419, n420,
 n421, n422, n423, n424, n425, n426, n427, n428,
 n429, n430, n431, n432, n433, n434, n435, n436,
 n437, n438, n439, n440, n441, n442, n443, n444,
 n445, n446, n447, n448, n449, n450, n451, n452,
 n453, n454, n455, n456, n457, n458, n459, n460,
 n461, n462, n463, n464, n465, n466, n467, n468,
 n469, n470, n471, n472, n473, n474, n475, n476,
 n477, n478, n479, n480, n481, n482, n483, n484,
 n485, n486, n487, n488, n489, n490, n491, n492,
 n493, n494, n495, n496, n497, n498, n499, n500,
 n501, n502, n503, n504, n505, n506, n507, n508,
 n509, n510, n511, n512, n513, n514, n515, n516,
 n517, n518, n519, n520, n521, n522, n523, n524,
 n525, n526, n527, n528, n529, n530, n531, n532,
 n533, n534, n535, n536, n537, n538, n539, n540,
 n541, n542, n543, n544, n545, n546, n547, n548,
 n549, n550, n551, n552, n553, n554, n555, n556,
 n557, n558, n559, n560, n561, n562, n563, n564,
 n565, n566, n567, n568, n569, n570, n571, n572,
 n573, n574, n575, n576, n577, n578, n579, n580,
 n581, n582, n583, n584, n585, n586, n587, n588,
 n589, n590, n591, n592, n593, n594, n595, n596,
 n597, n598, n599, n600, n601, n602, n603, n604,
 n605, n606, n607, n608, n609, n610, n611, n612,
 n613, n614, n615, n616, n617, n618, n619, n620,
 n621, n622, n623, n624, n625, n626, n627, n628,
 n629, n630, n631, n632, n633, n634, n635, n636,
 n637, n638, n639, n640, n641, n642, n643, n644,
 n645, n646, n647, n648, n649, n650, n651, n652,
 n653, n654, n655, n656, n657, n658, n659, n660,
 n661, n662, n663, n664, n665, n666, n667, n668,
 n669, n670, n671, n672, n673, n674, n675, n676,
 n677, n678, n679, n680, n681, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n758, n759, n760, n761, n762, n763, n764,
 n765, n766, n767, n768, n769, n770, n771, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n865, n866, n867, n868,
 n869, n870, n871, n872, n873, n874, n875, n876,
 n877, n878, n879, n880, n881, n882, n883, n884,
 n885, n886, n887, n888, n889, n890, n891, n892,
 n893, n894, n895, n896, n897, n898, n899, n900,
 n901, n902, n903, n904, n905, n906, n907, n908,
 n909, n910, n911, n912, n913, n914, n915, n916,
 n917, n918, n919, n920, n921, n922, n923, n924,
 n925, n926, n927, n928, n929, n930, n931, n932,
 n933, n934, n935, n936, n937, n938, n939, n940,
 n941, n942, n943, n944, n945, n946, n947, n948,
 n949, n950, n951, n952, n953, n954, n955, n956,
 n957, n958, n959, n960, n961, n962, n963, n964,
 n965, n966, n967, n968, n969, n970, n971, n972,
 n973, n974, n975, n976, n977, n978, n979, n980,
 n981, n982, n983, n984, n985, n986, n987, n988,
 n989, n990, n991, n992, n993, n994, n995, n996,
 n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
 n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
 n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
 n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
 n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
 n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
 n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
 n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
 n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
 n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
 n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
 n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
 n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
 n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
 n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
 n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
 n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
 n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
 n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
 n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
 n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
 n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
 n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
 n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
 n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
 n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
 n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
 n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
 n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
 n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
 n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
 n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
 n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
 n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
 n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
 n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
 n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
 n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
 n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
 n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
 n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
 n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
 n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
 n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
 n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
 n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
 n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
 n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
 n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
 n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
 n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
 n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
 n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
 n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
 n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
 n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
 n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
 n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
 n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
 n1469, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
 n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
 n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
 n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
 n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
 n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
 n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
 n1526, n1527, n1528, n1529, n1532, n1535, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1552, n1555, n1556, n1557, n1568, n1569,
 n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
 n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
 n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
 n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
 n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
 n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
 n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
 n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
 n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
 n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
 n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
 n1658, n1659, n1660, n1661;

not  g0 (n43, n8);
not  g1 (n25, n7);
not  g2 (n32, n14);
buf  g3 (n64, n16);
buf  g4 (n28, n11);
buf  g5 (n53, n20);
buf  g6 (n37, n3);
buf  g7 (n87, n6);
not  g8 (n27, n2);
not  g9 (n39, n1);
buf  g10 (n99, n1);
not  g11 (n30, n6);
buf  g12 (n41, n9);
buf  g13 (n55, n9);
not  g14 (n44, n14);
not  g15 (n98, n10);
buf  g16 (n97, n1);
buf  g17 (n89, n6);
buf  g18 (n96, n19);
buf  g19 (n69, n18);
not  g20 (n58, n15);
not  g21 (n50, n7);
buf  g22 (n67, n14);
buf  g23 (n81, n10);
not  g24 (n42, n19);
not  g25 (n76, n4);
buf  g26 (n29, n4);
not  g27 (n49, n16);
not  g28 (n80, n15);
buf  g29 (n66, n4);
not  g30 (n74, n12);
buf  g31 (n68, n10);
buf  g32 (n51, n8);
buf  g33 (n73, n8);
not  g34 (n94, n10);
buf  g35 (n57, n19);
not  g36 (n75, n18);
not  g37 (n95, n1);
buf  g38 (n84, n14);
not  g39 (n93, n3);
not  g40 (n83, n3);
not  g41 (n52, n11);
not  g42 (n72, n2);
not  g43 (n36, n13);
not  g44 (n54, n5);
buf  g45 (n22, n19);
buf  g46 (n40, n7);
buf  g47 (n24, n3);
buf  g48 (n33, n15);
buf  g49 (n35, n18);
not  g50 (n71, n20);
not  g51 (n85, n17);
not  g52 (n21, n6);
buf  g53 (n46, n15);
buf  g54 (n23, n5);
not  g55 (n61, n4);
buf  g56 (n56, n9);
buf  g57 (n38, n17);
buf  g58 (n60, n16);
buf  g59 (n31, n13);
buf  g60 (n88, n13);
not  g61 (n45, n13);
buf  g62 (n70, n2);
not  g63 (n63, n8);
buf  g64 (n47, n9);
buf  g65 (n34, n12);
not  g66 (n59, n16);
not  g67 (n62, n12);
buf  g68 (n78, n11);
buf  g69 (n86, n17);
not  g70 (n26, n7);
buf  g71 (n48, n5);
not  g72 (n92, n20);
not  g73 (n65, n12);
buf  g74 (n91, n2);
buf  g75 (n79, n11);
buf  g76 (n90, n18);
not  g77 (n77, n17);
buf  g78 (n82, n5);
not  g79 (n260, n91);
not  g80 (n365, n29);
buf  g81 (n289, n85);
buf  g82 (n214, n70);
not  g83 (n272, n92);
buf  g84 (n336, n43);
buf  g85 (n182, n80);
not  g86 (n199, n88);
not  g87 (n195, n54);
not  g88 (n279, n61);
not  g89 (n211, n81);
not  g90 (n244, n40);
buf  g91 (n246, n54);
not  g92 (n406, n53);
not  g93 (n187, n91);
buf  g94 (n183, n69);
not  g95 (n150, n63);
buf  g96 (n278, n41);
not  g97 (n296, n94);
not  g98 (n267, n59);
buf  g99 (n340, n55);
not  g100 (n208, n93);
buf  g101 (n287, n27);
buf  g102 (n378, n57);
buf  g103 (n245, n22);
buf  g104 (n130, n29);
not  g105 (n117, n87);
not  g106 (n361, n98);
not  g107 (n128, n65);
buf  g108 (n152, n87);
not  g109 (n352, n91);
buf  g110 (n312, n64);
buf  g111 (n111, n87);
buf  g112 (n141, n74);
not  g113 (n374, n85);
not  g114 (n298, n77);
buf  g115 (n138, n62);
not  g116 (n324, n78);
not  g117 (n209, n40);
not  g118 (n389, n94);
buf  g119 (n355, n46);
not  g120 (n328, n28);
buf  g121 (n103, n72);
buf  g122 (n113, n70);
not  g123 (n385, n63);
not  g124 (n400, n49);
not  g125 (n230, n23);
buf  g126 (n165, n37);
not  g127 (n292, n57);
not  g128 (n250, n67);
not  g129 (n231, n83);
not  g130 (n251, n22);
not  g131 (n380, n92);
buf  g132 (n176, n84);
not  g133 (n159, n59);
buf  g134 (n110, n51);
buf  g135 (n177, n80);
not  g136 (n268, n30);
not  g137 (n301, n89);
not  g138 (n239, n93);
buf  g139 (n102, n56);
not  g140 (n193, n46);
buf  g141 (n313, n31);
buf  g142 (n133, n75);
buf  g143 (n337, n84);
not  g144 (n242, n28);
buf  g145 (n163, n84);
not  g146 (n330, n88);
not  g147 (n135, n29);
not  g148 (n170, n78);
buf  g149 (n363, n56);
buf  g150 (n302, n27);
not  g151 (n282, n59);
not  g152 (n160, n21);
buf  g153 (n373, n29);
buf  g154 (n100, n86);
buf  g155 (n258, n53);
buf  g156 (n276, n36);
not  g157 (n335, n79);
buf  g158 (n377, n61);
not  g159 (n398, n91);
buf  g160 (n136, n62);
buf  g161 (n118, n87);
not  g162 (n202, n39);
not  g163 (n148, n21);
buf  g164 (n137, n41);
buf  g165 (n174, n50);
not  g166 (n140, n85);
buf  g167 (n353, n35);
buf  g168 (n345, n25);
buf  g169 (n234, n76);
not  g170 (n270, n30);
buf  g171 (n179, n43);
not  g172 (n399, n26);
buf  g173 (n391, n49);
not  g174 (n306, n38);
not  g175 (n387, n44);
buf  g176 (n395, n97);
buf  g177 (n325, n83);
not  g178 (n175, n48);
buf  g179 (n134, n26);
buf  g180 (n265, n64);
not  g181 (n178, n88);
buf  g182 (n358, n79);
not  g183 (n382, n66);
buf  g184 (n210, n38);
buf  g185 (n401, n61);
not  g186 (n331, n98);
not  g187 (n295, n36);
not  g188 (n350, n58);
not  g189 (n294, n86);
not  g190 (n359, n21);
buf  g191 (n261, n92);
buf  g192 (n411, n52);
not  g193 (n354, n70);
buf  g194 (n139, n95);
buf  g195 (n161, n32);
not  g196 (n266, n90);
not  g197 (n415, n82);
buf  g198 (n334, n58);
not  g199 (n362, n97);
not  g200 (n200, n66);
buf  g201 (n184, n97);
buf  g202 (n339, n62);
buf  g203 (n315, n75);
buf  g204 (n189, n77);
buf  g205 (n402, n59);
not  g206 (n311, n30);
buf  g207 (n262, n99);
buf  g208 (n121, n39);
not  g209 (n283, n58);
not  g210 (n277, n81);
not  g211 (n226, n45);
buf  g212 (n299, n42);
not  g213 (n357, n73);
buf  g214 (n143, n42);
not  g215 (n147, n47);
not  g216 (n186, n50);
buf  g217 (n132, n96);
buf  g218 (n213, n76);
buf  g219 (n410, n80);
not  g220 (n156, n65);
not  g221 (n249, n95);
not  g222 (n323, n68);
not  g223 (n407, n28);
not  g224 (n225, n27);
not  g225 (n241, n64);
not  g226 (n351, n72);
not  g227 (n369, n52);
not  g228 (n288, n65);
not  g229 (n316, n44);
not  g230 (n180, n32);
buf  g231 (n341, n34);
not  g232 (n169, n34);
not  g233 (n167, n44);
buf  g234 (n371, n45);
not  g235 (n414, n80);
not  g236 (n349, n93);
buf  g237 (n257, n39);
buf  g238 (n218, n51);
buf  g239 (n412, n73);
buf  g240 (n181, n24);
buf  g241 (n392, n37);
not  g242 (n188, n26);
not  g243 (n236, n35);
not  g244 (n219, n48);
not  g245 (n318, n67);
not  g246 (n381, n71);
not  g247 (n396, n66);
buf  g248 (n403, n31);
buf  g249 (n344, n89);
not  g250 (n112, n90);
not  g251 (n115, n79);
not  g252 (n379, n74);
buf  g253 (n168, n33);
not  g254 (n264, n61);
buf  g255 (n271, n60);
not  g256 (n305, n95);
buf  g257 (n123, n31);
buf  g258 (n206, n25);
buf  g259 (n319, n21);
buf  g260 (n122, n51);
buf  g261 (n338, n69);
not  g262 (n185, n23);
not  g263 (n291, n56);
not  g264 (n198, n76);
not  g265 (n375, n92);
buf  g266 (n393, n54);
buf  g267 (n149, n34);
buf  g268 (n274, n47);
buf  g269 (n275, n23);
not  g270 (n314, n94);
buf  g271 (n290, n99);
buf  g272 (n233, n65);
buf  g273 (n409, n35);
buf  g274 (n194, n81);
not  g275 (n269, n77);
buf  g276 (n366, n39);
not  g277 (n346, n74);
not  g278 (n376, n55);
buf  g279 (n397, n72);
not  g280 (n116, n54);
buf  g281 (n191, n32);
buf  g282 (n307, n97);
not  g283 (n173, n89);
buf  g284 (n166, n68);
not  g285 (n197, n31);
not  g286 (n386, n52);
not  g287 (n105, n23);
buf  g288 (n153, n67);
buf  g289 (n235, n99);
not  g290 (n372, n26);
not  g291 (n259, n58);
buf  g292 (n162, n63);
not  g293 (n104, n32);
buf  g294 (n332, n75);
buf  g295 (n300, n37);
buf  g296 (n190, n55);
not  g297 (n320, n98);
not  g298 (n222, n96);
buf  g299 (n106, n68);
buf  g300 (n216, n60);
buf  g301 (n119, n83);
not  g302 (n326, n25);
buf  g303 (n273, n43);
not  g304 (n303, n48);
not  g305 (n405, n82);
buf  g306 (n221, n85);
buf  g307 (n394, n94);
buf  g308 (n281, n47);
buf  g309 (n240, n88);
buf  g310 (n215, n52);
buf  g311 (n343, n22);
buf  g312 (n146, n76);
buf  g313 (n263, n95);
buf  g314 (n347, n98);
not  g315 (n327, n36);
buf  g316 (n109, n99);
buf  g317 (n120, n35);
not  g318 (n203, n74);
not  g319 (n158, n60);
not  g320 (n333, n96);
buf  g321 (n207, n38);
buf  g322 (n293, n49);
buf  g323 (n157, n77);
not  g324 (n204, n34);
not  g325 (n348, n71);
buf  g326 (n224, n90);
buf  g327 (n253, n53);
buf  g328 (n367, n24);
not  g329 (n232, n86);
buf  g330 (n171, n46);
buf  g331 (n309, n84);
not  g332 (n285, n42);
not  g333 (n254, n81);
not  g334 (n172, n50);
not  g335 (n308, n71);
not  g336 (n126, n41);
not  g337 (n256, n49);
not  g338 (n321, n79);
not  g339 (n280, n72);
not  g340 (n124, n24);
buf  g341 (n404, n64);
buf  g342 (n408, n53);
buf  g343 (n322, n83);
not  g344 (n252, n42);
not  g345 (n101, n55);
buf  g346 (n413, n57);
not  g347 (n286, n96);
buf  g348 (n131, n57);
not  g349 (n304, n86);
not  g350 (n384, n62);
buf  g351 (n196, n51);
not  g352 (n155, n45);
buf  g353 (n114, n43);
not  g354 (n227, n75);
buf  g355 (n229, n36);
buf  g356 (n107, n63);
not  g357 (n238, n56);
buf  g358 (n243, n30);
buf  g359 (n247, n46);
buf  g360 (n164, n33);
not  g361 (n329, n40);
buf  g362 (n228, n38);
buf  g363 (n342, n48);
not  g364 (n370, n45);
buf  g365 (n125, n40);
not  g366 (n145, n66);
buf  g367 (n154, n71);
not  g368 (n388, n50);
buf  g369 (n127, n89);
not  g370 (n144, n60);
not  g371 (n364, n78);
buf  g372 (n129, n44);
not  g373 (n223, n70);
not  g374 (n360, n41);
not  g375 (n201, n33);
buf  g376 (n255, n93);
not  g377 (n356, n68);
not  g378 (n237, n73);
not  g379 (n205, n33);
buf  g380 (n212, n25);
buf  g381 (n368, n82);
not  g382 (n297, n73);
not  g383 (n383, n24);
buf  g384 (n151, n37);
buf  g385 (n310, n78);
not  g386 (n217, n67);
not  g387 (n390, n22);
buf  g388 (n192, n90);
buf  g389 (n284, n69);
not  g390 (n317, n82);
not  g391 (n142, n27);
not  g392 (n220, n47);
not  g393 (n248, n69);
not  g394 (n108, n28);
buf  g395 (n493, n117);
not  g396 (n852, n308);
not  g397 (n622, n230);
not  g398 (n535, n112);
buf  g399 (n869, n376);
not  g400 (n486, n338);
not  g401 (n823, n355);
not  g402 (n692, n281);
buf  g403 (n479, n171);
buf  g404 (n540, n382);
buf  g405 (n641, n162);
buf  g406 (n537, n271);
not  g407 (n560, n257);
not  g408 (n846, n394);
not  g409 (n669, n222);
buf  g410 (n1040, n410);
buf  g411 (n538, n108);
buf  g412 (n1027, n104);
not  g413 (n1076, n360);
not  g414 (n853, n310);
buf  g415 (n1047, n317);
not  g416 (n1063, n120);
buf  g417 (n903, n158);
not  g418 (n627, n216);
not  g419 (n619, n154);
buf  g420 (n562, n201);
buf  g421 (n963, n130);
buf  g422 (n713, n339);
buf  g423 (n832, n174);
buf  g424 (n545, n167);
not  g425 (n950, n121);
buf  g426 (n550, n337);
buf  g427 (n883, n106);
buf  g428 (n567, n228);
not  g429 (n1003, n287);
not  g430 (n732, n132);
buf  g431 (n515, n348);
not  g432 (n1000, n173);
buf  g433 (n766, n288);
not  g434 (n1061, n180);
not  g435 (n881, n249);
buf  g436 (n1065, n218);
not  g437 (n584, n105);
buf  g438 (n977, n128);
not  g439 (n518, n190);
not  g440 (n660, n361);
buf  g441 (n855, n166);
not  g442 (n1088, n155);
not  g443 (n575, n279);
buf  g444 (n542, n239);
not  g445 (n1060, n208);
buf  g446 (n837, n153);
not  g447 (n765, n359);
not  g448 (n462, n272);
not  g449 (n635, n312);
not  g450 (n771, n121);
buf  g451 (n815, n218);
not  g452 (n517, n359);
buf  g453 (n565, n392);
not  g454 (n571, n171);
not  g455 (n1008, n189);
not  g456 (n449, n141);
not  g457 (n893, n151);
buf  g458 (n761, n266);
buf  g459 (n1069, n301);
buf  g460 (n556, n160);
not  g461 (n997, n157);
not  g462 (n500, n397);
buf  g463 (n1015, n306);
not  g464 (n657, n197);
not  g465 (n709, n186);
not  g466 (n530, n295);
buf  g467 (n931, n233);
not  g468 (n616, n205);
buf  g469 (n757, n296);
buf  g470 (n933, n131);
not  g471 (n848, n314);
buf  g472 (n778, n371);
not  g473 (n678, n189);
not  g474 (n896, n385);
buf  g475 (n474, n218);
not  g476 (n593, n319);
buf  g477 (n662, n110);
not  g478 (n473, n408);
not  g479 (n510, n379);
buf  g480 (n1037, n203);
not  g481 (n501, n193);
buf  g482 (n947, n310);
not  g483 (n720, n249);
not  g484 (n453, n262);
buf  g485 (n826, n373);
buf  g486 (n649, n347);
not  g487 (n800, n267);
not  g488 (n839, n331);
not  g489 (n441, n293);
buf  g490 (n604, n347);
not  g491 (n569, n102);
buf  g492 (n605, n306);
buf  g493 (n740, n176);
buf  g494 (n751, n187);
buf  g495 (n798, n366);
buf  g496 (n779, n361);
buf  g497 (n435, n118);
not  g498 (n822, n307);
buf  g499 (n930, n277);
not  g500 (n433, n338);
not  g501 (n489, n339);
buf  g502 (n623, n227);
not  g503 (n610, n411);
buf  g504 (n574, n142);
not  g505 (n541, n407);
not  g506 (n863, n283);
buf  g507 (n776, n308);
buf  g508 (n629, n162);
buf  g509 (n816, n353);
buf  g510 (n882, n198);
buf  g511 (n802, n378);
not  g512 (n705, n235);
buf  g513 (n674, n233);
buf  g514 (n667, n268);
not  g515 (n1032, n276);
not  g516 (n892, n185);
not  g517 (n995, n230);
buf  g518 (n745, n344);
not  g519 (n490, n207);
not  g520 (n1064, n104);
buf  g521 (n675, n390);
buf  g522 (n814, n219);
not  g523 (n828, n249);
buf  g524 (n502, n168);
buf  g525 (n680, n150);
buf  g526 (n718, n135);
not  g527 (n1089, n356);
buf  g528 (n946, n332);
buf  g529 (n483, n161);
buf  g530 (n951, n239);
buf  g531 (n639, n215);
buf  g532 (n938, n115);
not  g533 (n744, n149);
not  g534 (n886, n135);
buf  g535 (n561, n406);
not  g536 (n885, n374);
not  g537 (n417, n404);
not  g538 (n470, n404);
buf  g539 (n819, n266);
not  g540 (n711, n188);
buf  g541 (n955, n362);
not  g542 (n691, n283);
buf  g543 (n1021, n345);
buf  g544 (n971, n382);
not  g545 (n643, n381);
not  g546 (n551, n243);
buf  g547 (n958, n184);
buf  g548 (n914, n107);
buf  g549 (n987, n167);
not  g550 (n498, n302);
buf  g551 (n978, n384);
buf  g552 (n791, n378);
buf  g553 (n508, n140);
buf  g554 (n708, n204);
buf  g555 (n636, n114);
not  g556 (n531, n264);
buf  g557 (n877, n273);
not  g558 (n916, n180);
buf  g559 (n965, n107);
buf  g560 (n484, n157);
buf  g561 (n838, n369);
buf  g562 (n717, n337);
buf  g563 (n577, n103);
not  g564 (n595, n154);
not  g565 (n785, n360);
not  g566 (n661, n321);
buf  g567 (n736, n401);
not  g568 (n650, n255);
buf  g569 (n1093, n133);
not  g570 (n786, n191);
buf  g571 (n976, n297);
not  g572 (n465, n243);
buf  g573 (n889, n294);
not  g574 (n644, n347);
buf  g575 (n617, n333);
buf  g576 (n522, n363);
not  g577 (n509, n319);
buf  g578 (n974, n101);
not  g579 (n1012, n333);
buf  g580 (n741, n390);
buf  g581 (n725, n279);
not  g582 (n799, n336);
buf  g583 (n1042, n254);
not  g584 (n422, n215);
not  g585 (n689, n188);
not  g586 (n983, n275);
buf  g587 (n775, n172);
buf  g588 (n790, n365);
buf  g589 (n469, n257);
buf  g590 (n670, n338);
buf  g591 (n1002, n354);
buf  g592 (n867, n402);
buf  g593 (n1084, n297);
not  g594 (n464, n274);
not  g595 (n549, n240);
buf  g596 (n503, n115);
not  g597 (n957, n350);
not  g598 (n857, n307);
buf  g599 (n637, n332);
not  g600 (n555, n252);
buf  g601 (n1070, n177);
buf  g602 (n701, n199);
not  g603 (n972, n176);
not  g604 (n773, n156);
buf  g605 (n439, n325);
not  g606 (n1011, n286);
buf  g607 (n429, n166);
not  g608 (n625, n224);
not  g609 (n872, n329);
buf  g610 (n559, n407);
buf  g611 (n854, n133);
buf  g612 (n457, n169);
not  g613 (n727, n357);
buf  g614 (n1051, n331);
not  g615 (n1086, n410);
not  g616 (n813, n354);
not  g617 (n654, n269);
buf  g618 (n471, n249);
not  g619 (n621, n366);
buf  g620 (n478, n280);
not  g621 (n1041, n366);
buf  g622 (n835, n246);
not  g623 (n640, n268);
not  g624 (n825, n278);
not  g625 (n612, n203);
buf  g626 (n902, n222);
buf  g627 (n472, n102);
not  g628 (n552, n179);
not  g629 (n658, n409);
not  g630 (n671, n252);
not  g631 (n715, n269);
not  g632 (n1050, n364);
not  g633 (n434, n238);
buf  g634 (n873, n290);
buf  g635 (n841, n222);
not  g636 (n884, n178);
not  g637 (n774, n282);
not  g638 (n1025, n350);
not  g639 (n797, n367);
not  g640 (n737, n147);
buf  g641 (n463, n270);
buf  g642 (n891, n167);
buf  g643 (n672, n149);
buf  g644 (n734, n302);
not  g645 (n467, n301);
buf  g646 (n573, n317);
buf  g647 (n1029, n313);
buf  g648 (n770, n358);
buf  g649 (n438, n272);
buf  g650 (n989, n300);
buf  g651 (n926, n302);
buf  g652 (n716, n220);
buf  g653 (n495, n113);
not  g654 (n921, n389);
buf  g655 (n481, n272);
not  g656 (n809, n176);
buf  g657 (n992, n137);
not  g658 (n862, n392);
not  g659 (n521, n226);
buf  g660 (n525, n335);
buf  g661 (n454, n253);
not  g662 (n927, n138);
not  g663 (n609, n139);
not  g664 (n513, n166);
not  g665 (n805, n262);
not  g666 (n468, n124);
buf  g667 (n499, n386);
not  g668 (n714, n111);
buf  g669 (n952, n250);
buf  g670 (n871, n153);
not  g671 (n594, n334);
not  g672 (n1016, n355);
buf  g673 (n919, n402);
buf  g674 (n423, n390);
buf  g675 (n866, n214);
buf  g676 (n733, n177);
not  g677 (n847, n402);
buf  g678 (n696, n395);
not  g679 (n843, n352);
buf  g680 (n1017, n121);
not  g681 (n943, n164);
not  g682 (n557, n201);
buf  g683 (n748, n320);
not  g684 (n730, n223);
not  g685 (n1052, n183);
buf  g686 (n941, n330);
buf  g687 (n937, n346);
not  g688 (n460, n311);
not  g689 (n910, n223);
not  g690 (n586, n110);
not  g691 (n836, n196);
not  g692 (n447, n145);
not  g693 (n758, n382);
buf  g694 (n874, n406);
not  g695 (n880, n100);
not  g696 (n1020, n386);
buf  g697 (n1005, n168);
buf  g698 (n922, n116);
not  g699 (n1031, n300);
buf  g700 (n631, n130);
not  g701 (n702, n360);
buf  g702 (n1087, n205);
not  g703 (n445, n141);
not  g704 (n1091, n297);
buf  g705 (n959, n251);
buf  g706 (n436, n342);
buf  g707 (n578, n281);
buf  g708 (n749, n112);
buf  g709 (n942, n193);
buf  g710 (n682, n144);
buf  g711 (n628, n250);
not  g712 (n817, n104);
not  g713 (n735, n315);
buf  g714 (n606, n352);
not  g715 (n451, n148);
buf  g716 (n788, n179);
buf  g717 (n608, n280);
not  g718 (n583, n290);
buf  g719 (n679, n350);
buf  g720 (n430, n278);
buf  g721 (n1059, n258);
not  g722 (n1053, n252);
buf  g723 (n900, n122);
buf  g724 (n598, n327);
buf  g725 (n861, n230);
buf  g726 (n684, n219);
not  g727 (n1077, n196);
buf  g728 (n683, n217);
buf  g729 (n655, n370);
not  g730 (n476, n200);
not  g731 (n697, n332);
buf  g732 (n928, n228);
buf  g733 (n796, n298);
buf  g734 (n1028, n220);
not  g735 (n1071, n398);
not  g736 (n829, n270);
buf  g737 (n789, n296);
not  g738 (n783, n263);
buf  g739 (n1045, n206);
not  g740 (n563, n264);
not  g741 (n704, n143);
buf  g742 (n827, n255);
not  g743 (n690, n112);
not  g744 (n1030, n358);
buf  g745 (n935, n372);
not  g746 (n426, n377);
buf  g747 (n738, n397);
not  g748 (n721, n343);
buf  g749 (n968, n199);
not  g750 (n1023, n209);
not  g751 (n820, n397);
not  g752 (n964, n235);
not  g753 (n1090, n101);
buf  g754 (n945, n225);
buf  g755 (n1044, n220);
not  g756 (n554, n129);
buf  g757 (n920, n395);
not  g758 (n793, n225);
not  g759 (n419, n411);
not  g760 (n455, n348);
not  g761 (n494, n211);
not  g762 (n859, n254);
not  g763 (n969, n323);
not  g764 (n833, n329);
not  g765 (n808, n318);
not  g766 (n428, n280);
not  g767 (n596, n327);
not  g768 (n897, n225);
buf  g769 (n876, n110);
not  g770 (n1036, n330);
buf  g771 (n523, n240);
not  g772 (n668, n318);
buf  g773 (n899, n396);
buf  g774 (n1068, n202);
buf  g775 (n801, n380);
buf  g776 (n909, n351);
not  g777 (n1022, n284);
not  g778 (n558, n123);
not  g779 (n782, n377);
buf  g780 (n601, n305);
buf  g781 (n504, n213);
not  g782 (n588, n345);
not  g783 (n547, n214);
not  g784 (n985, n324);
buf  g785 (n967, n176);
buf  g786 (n592, n344);
not  g787 (n458, n353);
not  g788 (n611, n223);
buf  g789 (n582, n178);
not  g790 (n524, n181);
buf  g791 (n663, n242);
not  g792 (n587, n400);
buf  g793 (n564, n398);
not  g794 (n1082, n232);
buf  g795 (n750, n169);
buf  g796 (n784, n192);
buf  g797 (n1066, n203);
buf  g798 (n792, n118);
not  g799 (n681, n271);
buf  g800 (n929, n339);
not  g801 (n607, n182);
not  g802 (n570, n274);
buf  g803 (n795, n330);
buf  g804 (n917, n103);
buf  g805 (n477, n134);
buf  g806 (n768, n147);
buf  g807 (n645, n232);
not  g808 (n528, n140);
not  g809 (n634, n361);
buf  g810 (n1024, n208);
not  g811 (n804, n162);
not  g812 (n485, n283);
buf  g813 (n1001, n293);
buf  g814 (n603, n292);
buf  g815 (n999, n159);
not  g816 (n710, n321);
buf  g817 (n807, n177);
not  g818 (n614, n198);
not  g819 (n1014, n292);
not  g820 (n548, n242);
not  g821 (n894, n168);
not  g822 (n440, n345);
not  g823 (n514, n105);
buf  g824 (n580, n231);
not  g825 (n759, n401);
buf  g826 (n949, n213);
not  g827 (n731, n328);
buf  g828 (n907, n287);
buf  g829 (n461, n221);
buf  g830 (n442, n264);
not  g831 (n986, n259);
buf  g832 (n726, n179);
buf  g833 (n653, n163);
buf  g834 (n539, n222);
not  g835 (n676, n398);
buf  g836 (n1079, n232);
buf  g837 (n1010, n144);
buf  g838 (n437, n288);
buf  g839 (n452, n348);
buf  g840 (n1048, n324);
not  g841 (n719, n324);
buf  g842 (n723, n393);
not  g843 (n1018, n293);
not  g844 (n811, n126);
buf  g845 (n888, n276);
not  g846 (n844, n259);
not  g847 (n879, n307);
buf  g848 (n998, n261);
buf  g849 (n1095, n273);
not  g850 (n1072, n388);
not  g851 (n849, n334);
not  g852 (n572, n221);
not  g853 (n700, n157);
buf  g854 (n693, n284);
buf  g855 (n760, n322);
buf  g856 (n1006, n245);
not  g857 (n911, n286);
not  g858 (n685, n235);
buf  g859 (n906, n356);
not  g860 (n975, n244);
not  g861 (n984, n139);
buf  g862 (n664, n165);
buf  g863 (n993, n327);
not  g864 (n901, n185);
buf  g865 (n520, n237);
buf  g866 (n898, n207);
not  g867 (n446, n178);
buf  g868 (n688, n326);
buf  g869 (n443, n242);
not  g870 (n505, n198);
buf  g871 (n990, n217);
buf  g872 (n746, n132);
not  g873 (n450, n136);
buf  g874 (n544, n375);
not  g875 (n1049, n409);
buf  g876 (n772, n146);
not  g877 (n777, n347);
buf  g878 (n1039, n281);
buf  g879 (n742, n247);
not  g880 (n543, n399);
not  g881 (n724, n165);
buf  g882 (n475, n302);
buf  g883 (n1013, n155);
buf  g884 (n491, n147);
nand g885 (n729, n168, n326, n275, n215);
xor  g886 (n673, n163, n304, n120, n307);
or   g887 (n754, n303, n195, n323, n153);
and  g888 (n591, n253, n108, n206, n164);
nor  g889 (n1067, n404, n125, n256, n389);
nor  g890 (n988, n209, n241, n267, n314);
nor  g891 (n1075, n365, n342, n401, n229);
or   g892 (n599, n363, n160, n159, n319);
nand g893 (n632, n193, n383, n122, n370);
nor  g894 (n581, n189, n273, n368, n291);
nand g895 (n568, n212, n119, n224, n234);
nand g896 (n752, n369, n312, n116, n154);
xor  g897 (n648, n161, n247, n275, n112);
nand g898 (n850, n365, n134, n105, n306);
nor  g899 (n824, n391, n268, n108, n145);
nand g900 (n979, n231, n110, n228, n158);
or   g901 (n851, n103, n270, n286, n381);
nor  g902 (n762, n346, n362, n264, n297);
xnor g903 (n703, n172, n184, n200, n229);
or   g904 (n624, n221, n152, n319, n395);
nor  g905 (n940, n333, n299, n239, n367);
and  g906 (n459, n322, n127, n285, n278);
xor  g907 (n764, n318, n387, n300, n269);
and  g908 (n1056, n363, n246, n170, n395);
nand g909 (n576, n246, n149, n189, n388);
xor  g910 (n780, n122, n100, n263, n339);
nor  g911 (n579, n373, n364, n156, n346);
nor  g912 (n821, n375, n228, n312, n141);
xor  g913 (n456, n375, n310, n234, n371);
nand g914 (n618, n273, n393, n378, n127);
nor  g915 (n466, n239, n374, n304, n109);
xnor g916 (n585, n124, n256, n243, n279);
nor  g917 (n496, n174, n216, n128, n194);
nand g918 (n1057, n231, n119, n350, n109);
xnor g919 (n652, n336, n240, n132, n349);
xor  g920 (n512, n378, n290, n383, n137);
nand g921 (n482, n250, n146, n396, n166);
nor  g922 (n646, n340, n215, n270, n337);
nor  g923 (n781, n191, n182, n207, n201);
or   g924 (n1094, n268, n226, n343, n267);
nor  g925 (n534, n410, n318, n380, n316);
xnor g926 (n1046, n123, n208, n101, n233);
nor  g927 (n944, n358, n299, n255, n130);
xnor g928 (n810, n244, n296, n351, n303);
or   g929 (n638, n195, n133, n320, n211);
or   g930 (n966, n285, n341, n241, n186);
xor  g931 (n812, n237, n374, n128, n230);
nand g932 (n982, n186, n322, n352, n140);
and  g933 (n1081, n134, n351, n106, n399);
and  g934 (n506, n111, n271, n368, n387);
and  g935 (n421, n336, n357, n294, n405);
nor  g936 (n424, n245, n195, n183, n288);
xor  g937 (n834, n180, n245, n254, n127);
and  g938 (n739, n102, n400, n334, n372);
and  g939 (n991, n154, n330, n355, n287);
xor  g940 (n1007, n139, n341, n354, n397);
and  g941 (n895, n276, n204, n306, n341);
nor  g942 (n915, n136, n145, n247, n192);
xor  g943 (n529, n136, n327, n372, n216);
xor  g944 (n698, n214, n258, n175, n393);
xnor g945 (n842, n106, n328, n298, n188);
and  g946 (n1019, n388, n305, n261, n258);
or   g947 (n1073, n411, n202, n210, n190);
or   g948 (n659, n384, n146, n364, n401);
xor  g949 (n553, n301, n294, n402, n132);
or   g950 (n1083, n393, n244, n212, n405);
nor  g951 (n864, n342, n179, n240, n357);
xor  g952 (n527, n238, n316, n282, n285);
xnor g953 (n908, n279, n205, n150, n227);
xor  g954 (n923, n192, n337, n100, n145);
and  g955 (n566, n117, n183, n182, n190);
or   g956 (n590, n299, n356, n407, n105);
nand g957 (n647, n410, n271, n235, n288);
xnor g958 (n633, n373, n114, n251, n213);
nor  g959 (n962, n172, n405, n242, n128);
xor  g960 (n981, n380, n371, n150, n258);
nand g961 (n492, n334, n223, n117, n403);
and  g962 (n706, n164, n317, n380, n217);
nor  g963 (n533, n296, n182, n289, n304);
and  g964 (n980, n243, n206, n126, n198);
and  g965 (n970, n248, n260, n109, n409);
xnor g966 (n677, n343, n108, n130, n400);
xnor g967 (n420, n392, n226, n265, n157);
and  g968 (n722, n344, n196, n116, n256);
and  g969 (n953, n150, n202, n129, n116);
and  g970 (n666, n114, n104, n218, n389);
and  g971 (n615, n260, n206, n156, n143);
or   g972 (n642, n191, n229, n117, n344);
xnor g973 (n1055, n390, n404, n269, n282);
or   g974 (n425, n359, n260, n309, n274);
or   g975 (n427, n379, n199, n316, n267);
nand g976 (n416, n142, n248, n287, n398);
nor  g977 (n1054, n305, n324, n379, n360);
xnor g978 (n487, n408, n409, n190, n412);
or   g979 (n630, n277, n113, n341, n177);
xor  g980 (n961, n118, n391, n263, n311);
xnor g981 (n1026, n276, n331, n303, n151);
xnor g982 (n763, n122, n202, n151, n266);
nand g983 (n767, n227, n155, n171);
or   g984 (n1004, n257, n158, n163, n340);
or   g985 (n532, n394, n386, n148, n241);
nand g986 (n831, n173, n335, n367, n139);
nor  g987 (n806, n201, n187, n370, n251);
nand g988 (n695, n253, n216, n109, n353);
nand g989 (n890, n376, n224, n146, n313);
xor  g990 (n497, n188, n135, n326, n408);
nor  g991 (n516, n308, n396, n259, n362);
nand g992 (n860, n349, n362, n265, n165);
and  g993 (n954, n187, n224, n183, n126);
and  g994 (n665, n320, n346, n121, n204);
nor  g995 (n600, n278, n170, n144, n184);
nor  g996 (n444, n376, n385, n261, n260);
or   g997 (n519, n316, n336, n125, n194);
xnor g998 (n913, n187, n251, n291, n184);
or   g999 (n875, n159, n186, n118, n174);
nor  g1000 (n878, n329, n237, n367, n283);
and  g1001 (n830, n354, n138, n194, n257);
xnor g1002 (n769, n329, n291, n227, n290);
nand g1003 (n694, n289, n160, n148, n115);
and  g1004 (n1009, n387, n169, n163, n325);
nand g1005 (n1062, n234, n196, n328, n385);
nand g1006 (n707, n217, n158, n261, n181);
xor  g1007 (n1080, n204, n408, n138, n120);
nor  g1008 (n743, n391, n236, n368, n308);
nor  g1009 (n794, n169, n374, n199, n131);
and  g1010 (n787, n255, n225, n134, n292);
nand g1011 (n994, n294, n246, n315, n247);
nor  g1012 (n418, n205, n309, n262, n256);
or   g1013 (n948, n210, n200, n252, n203);
xnor g1014 (n613, n220, n181, n148, n403);
nor  g1015 (n712, n389, n233, n207, n301);
or   g1016 (n1074, n236, n387, n136, n388);
or   g1017 (n626, n314, n123, n274, n342);
xor  g1018 (n912, n144, n107, n384, n310);
xnor g1019 (n526, n331, n244, n123, n127);
or   g1020 (n546, n323, n263, n358, n111);
xnor g1021 (n747, n221, n355, n277, n159);
and  g1022 (n840, n232, n372, n379, n275);
nand g1023 (n589, n345, n383, n359, n300);
xnor g1024 (n620, n113, n161, n400, n305);
nand g1025 (n699, n303, n371, n125, n385);
or   g1026 (n1035, n119, n381, n133, n200);
xnor g1027 (n1085, n335, n332, n382, n309);
or   g1028 (n868, n280, n394, n124, n162);
or   g1029 (n536, n321, n238, n152, n383);
nand g1030 (n925, n272, n386, n236, n312);
nor  g1031 (n936, n406, n369, n403, n320);
or   g1032 (n728, n211, n175, n185, n356);
nand g1033 (n756, n135, n293, n321, n226);
xor  g1034 (n845, n311, n114, n368, n210);
nor  g1035 (n865, n192, n153, n396, n101);
xor  g1036 (n904, n335, n309, n214, n370);
or   g1037 (n1058, n171, n131, n237, n140);
xor  g1038 (n597, n143, n147, n131, n265);
and  g1039 (n1034, n392, n209, n314, n377);
and  g1040 (n870, n197, n412, n191, n137);
xnor g1041 (n651, n340, n375, n164, n277);
xor  g1042 (n511, n160, n241, n376, n197);
xnor g1043 (n686, n143, n291, n363, n381);
or   g1044 (n755, n403, n254, n317, n315);
and  g1045 (n918, n366, n238, n315, n100);
nor  g1046 (n488, n265, n209, n170, n156);
nand g1047 (n818, n373, n151, n365, n115);
xnor g1048 (n656, n141, n328, n325, n349);
and  g1049 (n1092, n384, n405, n137, n333);
xor  g1050 (n1038, n142, n194, n173, n284);
xnor g1051 (n687, n348, n338, n304, n234);
xnor g1052 (n934, n236, n295, n292, n357);
and  g1053 (n803, n248, n394, n340, n175);
nand g1054 (n924, n170, n213, n298, n391);
xnor g1055 (n432, n407, n323, n142, n211);
xnor g1056 (n858, n361, n289, n250, n311);
or   g1057 (n887, n178, n313, n138, n219);
or   g1058 (n1078, n266, n172, n411, n295);
xnor g1059 (n956, n102, n181, n289, n325);
or   g1060 (n431, n175, n248, n313, n152);
and  g1061 (n602, n167, n212, n180, n173);
xor  g1062 (n932, n152, n103, n298, n284);
or   g1063 (n480, n353, n322, n369, n165);
xor  g1064 (n960, n219, n107, n406, n120);
nor  g1065 (n973, n253, n245, n299, n349);
nand g1066 (n856, n286, n149, n281, n377);
and  g1067 (n1043, n210, n351, n295, n161);
and  g1068 (n448, n185, n282, n119, n352);
xor  g1069 (n939, n259, n262, n106, n129);
nand g1070 (n905, n229, n193, n212, n197);
and  g1071 (n507, n231, n174, n399, n125);
nor  g1072 (n753, n326, n195, n126, n364);
and  g1073 (n1033, n111, n129, n343, n113);
or   g1074 (n996, n124, n285, n208, n399);
nor  g1075 (n1177, n833, n959, n837, n477);
and  g1076 (n1180, n424, n815, n908, n989);
and  g1077 (n1293, n990, n923, n715, n897);
nand g1078 (n1239, n1020, n503, n1019, n526);
nand g1079 (n1237, n588, n757, n444, n705);
xor  g1080 (n1262, n860, n898, n696, n555);
nor  g1081 (n1186, n587, n490, n805, n676);
xor  g1082 (n1148, n493, n1005, n977, n884);
or   g1083 (n1152, n765, n886, n718, n900);
xor  g1084 (n1282, n418, n611, n453, n760);
nand g1085 (n1295, n974, n854, n995, n879);
xnor g1086 (n1104, n693, n915, n785, n709);
xor  g1087 (n1163, n795, n754, n495, n862);
or   g1088 (n1195, n912, n878, n1016, n1010);
xor  g1089 (n1298, n811, n624, n926, n524);
nand g1090 (n1290, n849, n947, n1011, n672);
nand g1091 (n1146, n561, n716, n830, n1012);
xor  g1092 (n1191, n864, n736, n813, n811);
xnor g1093 (n1208, n652, n514, n697, n892);
xnor g1094 (n1244, n924, n547, n663, n872);
nand g1095 (n1100, n1002, n960, n888, n961);
nor  g1096 (n1199, n501, n835, n567, n979);
xor  g1097 (n1225, n846, n870, n893, n954);
or   g1098 (n1212, n464, n835, n536, n685);
or   g1099 (n1171, n434, n623, n549, n844);
nor  g1100 (n1205, n955, n791, n867, n431);
xor  g1101 (n1162, n866, n527, n558, n695);
and  g1102 (n1232, n479, n806, n1015, n752);
xnor g1103 (n1124, n901, n530, n531, n997);
nand g1104 (n1167, n827, n827, n551, n779);
xnor g1105 (n1200, n605, n968, n822, n586);
xor  g1106 (n1139, n904, n903, n731, n564);
or   g1107 (n1276, n810, n1000, n896, n1014);
or   g1108 (n1134, n712, n772, n644, n668);
or   g1109 (n1230, n840, n435, n670, n509);
and  g1110 (n1248, n919, n593, n667, n452);
nand g1111 (n1271, n849, n993, n944, n544);
or   g1112 (n1273, n1002, n470, n480, n797);
and  g1113 (n1172, n884, n912, n956, n619);
xor  g1114 (n1300, n622, n826, n1013, n891);
nand g1115 (n1217, n528, n1006, n627, n789);
or   g1116 (n1275, n688, n897, n936, n513);
and  g1117 (n1175, n699, n1009, n851, n875);
nand g1118 (n1183, n711, n943, n820, n777);
nand g1119 (n1107, n995, n727, n733, n859);
xnor g1120 (n1301, n655, n516, n601, n525);
nor  g1121 (n1112, n887, n1004, n532, n578);
xnor g1122 (n1133, n649, n810, n836, n512);
or   g1123 (n1122, n914, n816, n475, n502);
nor  g1124 (n1283, n953, n831, n936, n994);
and  g1125 (n1220, n1012, n1018, n819, n454);
and  g1126 (n1259, n665, n987, n476, n871);
and  g1127 (n1294, n463, n700, n738, n429);
nand g1128 (n1238, n876, n800, n929, n683);
nor  g1129 (n1222, n633, n691, n519, n496);
nand g1130 (n1243, n883, n848, n878, n847);
xnor g1131 (n1260, n905, n769, n965, n824);
xor  g1132 (n1128, n973, n838, n679, n573);
nand g1133 (n1157, n591, n756, n637, n857);
xnor g1134 (n1234, n981, n858, n554, n799);
xnor g1135 (n1302, n950, n730, n538, n903);
xnor g1136 (n1142, n782, n874, n879, n949);
or   g1137 (n1156, n446, n837, n545, n872);
xor  g1138 (n1106, n673, n550, n540, n658);
xnor g1139 (n1099, n417, n830, n442, n957);
or   g1140 (n1202, n515, n721, n743, n616);
nand g1141 (n1214, n961, n553, n820, n548);
xnor g1142 (n1140, n943, n900, n500, n966);
and  g1143 (n1120, n462, n801, n582, n626);
and  g1144 (n1263, n653, n937, n796, n969);
nand g1145 (n1228, n902, n487, n981, n917);
and  g1146 (n1278, n976, n893, n945, n805);
or   g1147 (n1129, n425, n468, n771, n600);
nor  g1148 (n1303, n648, n986, n560, n542);
xnor g1149 (n1216, n869, n416, n871, n808);
nor  g1150 (n1102, n971, n823, n876, n840);
and  g1151 (n1241, n589, n909, n783, n920);
and  g1152 (n1115, n533, n889, n845, n1018);
nor  g1153 (n1233, n703, n1013, n786, n952);
nand g1154 (n1279, n860, n657, n508, n801);
or   g1155 (n1181, n1017, n486, n931, n948);
xnor g1156 (n1123, n1016, n1007, n774, n674);
or   g1157 (n1226, n535, n759, n858, n971);
xor  g1158 (n1249, n725, n998, n813, n982);
xnor g1159 (n1207, n984, n829, n456, n428);
xnor g1160 (n1126, n852, n877, n421, n773);
xnor g1161 (n1265, n917, n999, n934, n960);
xor  g1162 (n1143, n471, n967, n887, n1017);
xnor g1163 (n1096, n842, n986, n481, n926);
or   g1164 (n1206, n870, n942, n930, n817);
xnor g1165 (n1145, n720, n598, n510, n608);
nor  g1166 (n1229, n973, n584, n809, n1003);
or   g1167 (n1250, n1001, n916, n602, n1000);
and  g1168 (n1198, n859, n972, n808, n865);
nor  g1169 (n1113, n671, n839, n707, n814);
xor  g1170 (n1187, n898, n645, n574, n557);
and  g1171 (n1246, n677, n1011, n939, n822);
xnor g1172 (n1281, n1005, n613, n802, n992);
nand g1173 (n1192, n844, n906, n698, n997);
and  g1174 (n1103, n940, n940, n841, n812);
or   g1175 (n1296, n992, n809, n761, n794);
and  g1176 (n1125, n459, n629, n896, n890);
xor  g1177 (n1215, n942, n856, n862, n621);
or   g1178 (n1190, n883, n933, n911, n855);
and  g1179 (n1201, n974, n978, n951, n990);
nand g1180 (n1299, n599, n594, n964);
or   g1181 (n1224, n581, n632, n1009, n928);
or   g1182 (n1135, n570, n666, n692, n969);
xor  g1183 (n1151, n534, n450, n838, n953);
xor  g1184 (n1149, n770, n821, n993, n1022);
nor  g1185 (n1253, n473, n485, n925, n932);
and  g1186 (n1130, n520, n1021, n766, n963);
xnor g1187 (n1252, n735, n706, n443, n952);
and  g1188 (n1185, n843, n541, n732, n877);
or   g1189 (n1288, n825, n494, n968, n863);
xor  g1190 (n1173, n918, n910, n1019, n714);
or   g1191 (n1197, n1020, n998, n977, n967);
xor  g1192 (n1169, n938, n441, n704, n921);
or   g1193 (n1223, n895, n1008, n634, n803);
xor  g1194 (n1258, n590, n938, n522, n488);
nand g1195 (n1165, n922, n592, n799, n569);
xor  g1196 (n1257, n618, n669, n498, n628);
and  g1197 (n1236, n987, n426, n848, n744);
xnor g1198 (n1178, n861, n643, n740, n975);
and  g1199 (n1154, n976, n690, n962, n664);
and  g1200 (n1179, n853, n946, n420, n915);
or   g1201 (n1155, n749, n853, n991, n562);
xor  g1202 (n1280, n1006, n905, n576, n478);
or   g1203 (n1210, n874, n607, n640, n972);
xor  g1204 (n1164, n894, n460, n928, n828);
xor  g1205 (n1284, n873, n956, n788, n804);
nand g1206 (n1240, n815, n654, n641, n814);
and  g1207 (n1101, n913, n713, n829, n922);
xor  g1208 (n1161, n529, n873, n566, n930);
nand g1209 (n1221, n596, n511, n764, n914);
xnor g1210 (n1108, n919, n689, n962, n851);
nand g1211 (n1098, n1010, n999, n650, n543);
or   g1212 (n1204, n866, n686, n681, n472);
or   g1213 (n1286, n457, n902, n710, n660);
or   g1214 (n1118, n790, n680, n1021, n780);
xnor g1215 (n1136, n556, n638, n728, n614);
or   g1216 (n1297, n985, n904, n889, n982);
xor  g1217 (n1150, n461, n615, n746, n994);
nor  g1218 (n1196, n836, n931, n955, n857);
or   g1219 (n1255, n925, n839, n436, n568);
xnor g1220 (n1261, n895, n751, n817, n1007);
xor  g1221 (n1245, n662, n924, n842, n438);
or   g1222 (n1254, n647, n885, n523, n1014);
nand g1223 (n1272, n646, n719, n989, n970);
xor  g1224 (n1110, n739, n847, n828, n753);
and  g1225 (n1291, n768, n651, n741, n913);
and  g1226 (n1168, n625, n440, n958, n923);
nor  g1227 (n1159, n894, n583, n984, n921);
xnor g1228 (n1242, n947, n824, n745, n901);
or   g1229 (n1184, n841, n948, n899, n957);
or   g1230 (n1137, n950, n832, n946, n927);
and  g1231 (n1269, n419, n437, n776, n506);
or   g1232 (n1116, n787, n775, n832, n941);
and  g1233 (n1218, n1001, n675, n579, n983);
xnor g1234 (n1211, n678, n609, n935, n423);
or   g1235 (n1287, n864, n880, n935, n635);
nand g1236 (n1251, n868, n932, n869, n701);
nor  g1237 (n1114, n445, n563, n929, n639);
xor  g1238 (n1132, n963, n687, n890, n980);
nand g1239 (n1285, n492, n978, n885, n448);
and  g1240 (n1292, n661, n804, n843, n806);
nor  g1241 (n1189, n737, n821, n834, n880);
nand g1242 (n1182, n927, n798, n708, n758);
and  g1243 (n1188, n875, n439, n484, n742);
nor  g1244 (n1176, n449, n734, n970, n939);
and  g1245 (n1235, n620, n816, n907, n818);
xnor g1246 (n1209, n886, n1008, n944, n933);
and  g1247 (n1111, n604, n762, n636, n539);
xor  g1248 (n1147, n537, n659, n474, n722);
xnor g1249 (n1158, n965, n959, n432, n916);
xor  g1250 (n1174, n507, n767, n455, n991);
nand g1251 (n1267, n585, n717, n726, n631);
nor  g1252 (n1247, n482, n863, n447, n800);
xor  g1253 (n1141, n803, n793, n747, n881);
or   g1254 (n1213, n856, n850, n778, n603);
xor  g1255 (n1153, n682, n855, n945, n834);
xor  g1256 (n1160, n575, n497, n781, n466);
xnor g1257 (n1109, n610, n802, n852, n807);
nor  g1258 (n1170, n867, n918, n565, n642);
nand g1259 (n1144, n818, n577, n909, n427);
nor  g1260 (n1264, n630, n724, n694, n910);
xnor g1261 (n1266, n891, n465, n996, n819);
or   g1262 (n1277, n951, n949, n505, n499);
xnor g1263 (n1268, n954, n433, n521, n572);
xnor g1264 (n1105, n1003, n451, n899, n958);
xnor g1265 (n1193, n518, n597, n823, n469);
nand g1266 (n1203, n888, n1015, n784, n807);
xnor g1267 (n1127, n850, n934, n966, n845);
xor  g1268 (n1289, n941, n906, n571, n702);
and  g1269 (n1131, n868, n552, n979, n812);
nor  g1270 (n1194, n988, n729, n606, n792);
xor  g1271 (n1227, n882, n907, n422, n755);
xor  g1272 (n1274, n996, n846, n580, n831);
and  g1273 (n1219, n882, n825, n483, n612);
or   g1274 (n1256, n908, n975, n430, n892);
nand g1275 (n1097, n983, n504, n750, n920);
or   g1276 (n1121, n684, n559, n861, n985);
xor  g1277 (n1231, n491, n1004, n937, n517);
xnor g1278 (n1117, n865, n763, n748, n546);
nand g1279 (n1166, n617, n881, n723, n826);
nand g1280 (n1270, n595, n833, n980, n854);
and  g1281 (n1138, n911, n988, n656, n797);
nor  g1282 (n1119, n467, n798, n489, n458);
not  g1283 (n1315, n1137);
buf  g1284 (n1351, n1099);
buf  g1285 (n1323, n1128);
not  g1286 (n1307, n1102);
buf  g1287 (n1336, n1097);
not  g1288 (n1327, n1111);
not  g1289 (n1331, n1146);
buf  g1290 (n1317, n1143);
not  g1291 (n1353, n1109);
buf  g1292 (n1343, n1124);
not  g1293 (n1326, n1112);
not  g1294 (n1361, n1123);
not  g1295 (n1335, n1100);
not  g1296 (n1352, n1101);
not  g1297 (n1328, n1148);
buf  g1298 (n1350, n1096);
not  g1299 (n1322, n1139);
buf  g1300 (n1334, n1127);
not  g1301 (n1349, n1119);
not  g1302 (n1314, n1142);
buf  g1303 (n1338, n1133);
not  g1304 (n1324, n1120);
buf  g1305 (n1342, n1151);
buf  g1306 (n1337, n1122);
buf  g1307 (n1345, n1132);
not  g1308 (n1341, n1106);
buf  g1309 (n1306, n1110);
not  g1310 (n1357, n1098);
buf  g1311 (n1308, n1136);
buf  g1312 (n1318, n1135);
not  g1313 (n1358, n1104);
not  g1314 (n1356, n1121);
buf  g1315 (n1313, n1113);
not  g1316 (n1333, n1108);
not  g1317 (n1330, n1150);
buf  g1318 (n1360, n1149);
buf  g1319 (n1305, n1117);
not  g1320 (n1340, n1126);
not  g1321 (n1310, n1141);
buf  g1322 (n1354, n1115);
not  g1323 (n1347, n1125);
buf  g1324 (n1319, n1105);
not  g1325 (n1312, n1118);
buf  g1326 (n1332, n1138);
buf  g1327 (n1311, n1147);
buf  g1328 (n1309, n1140);
buf  g1329 (n1344, n1145);
buf  g1330 (n1325, n1153);
not  g1331 (n1355, n1116);
not  g1332 (n1320, n1131);
buf  g1333 (n1339, n1114);
buf  g1334 (n1348, n1144);
buf  g1335 (n1321, n1107);
buf  g1336 (n1346, n1152);
buf  g1337 (n1316, n1129);
not  g1338 (n1304, n1130);
not  g1339 (n1329, n1134);
buf  g1340 (n1359, n1103);
buf  g1341 (n1366, n1305);
buf  g1342 (n1362, n1305);
not  g1343 (n1363, n1307);
or   g1344 (n1365, n1304, n1306);
xor  g1345 (n1364, n1306, n1304, n1308);
buf  g1346 (n1373, n1363);
not  g1347 (n1375, n1364);
buf  g1348 (n1367, n1362);
buf  g1349 (n1374, n1154);
not  g1350 (n1376, n1362);
not  g1351 (n1371, n1156);
buf  g1352 (n1370, n1160);
or   g1353 (n1368, n1159, n1365, n1363);
nand g1354 (n1372, n1157, n1155, n1158, n1366);
nor  g1355 (n1369, n1364, n1366, n1161, n1162);
not  g1356 (n1380, n1367);
not  g1357 (n1377, n1166);
nand g1358 (n1379, n1163, n1368, n1164, n1167);
nor  g1359 (n1378, n1369, n1168, n1165, n1370);
xor  g1360 (n1384, n1191, n1377, n1188, n1186);
xnor g1361 (n1386, n1378, n1204, n1208, n1201);
nor  g1362 (n1394, n1200, n1169, n1183, n1379);
nand g1363 (n1390, n1206, n1176, n1379, n1172);
nand g1364 (n1393, n1213, n1192, n1178, n1210);
xnor g1365 (n1387, n1190, n1185, n1182, n1195);
or   g1366 (n1381, n1181, n1177, n1377, n1379);
xnor g1367 (n1382, n1194, n1378, n1184, n1380);
xnor g1368 (n1392, n1380, n1205, n1170, n1202);
nand g1369 (n1385, n1377, n1211, n1379, n1380);
xor  g1370 (n1388, n1196, n1207, n1378, n1377);
or   g1371 (n1383, n1214, n1209, n1175, n1197);
and  g1372 (n1389, n1212, n1215, n1380, n1193);
nor  g1373 (n1396, n1180, n1171, n1198, n1203);
xor  g1374 (n1395, n1173, n1179, n1174, n1187);
nor  g1375 (n1391, n1378, n1189, n1216, n1199);
nand g1376 (n1399, n1386, n1317, n1313, n1321);
xor  g1377 (n1405, n1323, n1310, n1309, n1311);
nor  g1378 (n1406, n1319, n1315, n1385, n1310);
nand g1379 (n1402, n1224, n1311, n1226, n1324);
nor  g1380 (n1404, n1321, n1314, n1381, n1323);
xnor g1381 (n1403, n1388, n1396, n1384, n1225);
or   g1382 (n1398, n1315, n1394, n1223, n1312);
xor  g1383 (n1400, n1323, n1317, n1382, n1318);
or   g1384 (n1397, n1320, n1391, n1390, n1219);
or   g1385 (n1409, n1221, n1389, n1393, n1309);
nand g1386 (n1411, n1227, n1316, n1322, n1220);
or   g1387 (n1401, n1312, n1395, n1392, n1322);
nor  g1388 (n1408, n1222, n1321, n1217, n1387);
nor  g1389 (n1410, n1319, n1313, n1228, n1322);
nand g1390 (n1407, n1320, n1318, n1383, n1218);
or   g1391 (n1412, n1320, n1324, n1316, n1314);
nor  g1392 (n1430, n1334, n1343, n1353, n1350);
nor  g1393 (n1423, n1400, n1335, n1339, n1399);
xnor g1394 (n1424, n1332, n1336, n1401, n1346);
nand g1395 (n1443, n1338, n1350, n1352, n1343);
nand g1396 (n1439, n1336, n1337, n1346, n1328);
xor  g1397 (n1431, n1325, n1328, n1327, n1347);
xnor g1398 (n1414, n1334, n1326, n1332, n1346);
xnor g1399 (n1428, n1343, n1345, n1326);
nand g1400 (n1435, n1327, n1410, n1334, n1345);
nor  g1401 (n1444, n1351, n1405, n1328, n1353);
or   g1402 (n1426, n1348, n1342, n1404, n1406);
and  g1403 (n1422, n1399, n1340, n1352, n1339);
xnor g1404 (n1413, n1352, n1347, n1338, n1335);
and  g1405 (n1432, n1407, n1348, n1351, n1335);
or   g1406 (n1421, n1406, n1409, n1412, n1344);
xnor g1407 (n1437, n1331, n1327, n1330, n1404);
and  g1408 (n1418, n1412, n1331, n1336, n1326);
xnor g1409 (n1419, n1411, n1340, n1408, n1402);
xnor g1410 (n1440, n1331, n1351, n1400, n1329);
xor  g1411 (n1427, n1398, n1340, n1341, n1402);
and  g1412 (n1442, n1410, n1347, n1403, n1333);
nand g1413 (n1415, n1329, n1329, n1397, n1407);
and  g1414 (n1420, n1401, n1349, n1409, n1397);
or   g1415 (n1429, n1398, n1408, n1325, n1411);
or   g1416 (n1434, n1353, n1350, n1324, n1341);
or   g1417 (n1433, n1342, n1350, n1349, n1337);
xnor g1418 (n1425, n1405, n1333, n1339, n1345);
xnor g1419 (n1436, n1352, n1342, n1347, n1338);
and  g1420 (n1441, n1344, n1351, n1348, n1330);
nor  g1421 (n1416, n1349, n1344, n1337, n1348);
and  g1422 (n1438, n1325, n1341, n1346, n1333);
nand g1423 (n1417, n1349, n1332, n1330, n1403);
buf  g1424 (n1445, n1238);
not  g1425 (n1460, n1428);
buf  g1426 (n1458, n1232);
not  g1427 (n1455, n1426);
buf  g1428 (n1461, n1420);
buf  g1429 (n1452, n1430);
buf  g1430 (n1463, n1229);
buf  g1431 (n1453, n1424);
buf  g1432 (n1462, n1422);
buf  g1433 (n1465, n1235);
buf  g1434 (n1447, n1425);
not  g1435 (n1457, n1428);
buf  g1436 (n1446, n1233);
buf  g1437 (n1467, n1418);
buf  g1438 (n1466, n1427);
buf  g1439 (n1454, n1415);
not  g1440 (n1464, n1234);
not  g1441 (n1449, n1430);
buf  g1442 (n1450, n1426);
buf  g1443 (n1468, n1413);
nand g1444 (n1459, n1417, n1429);
and  g1445 (n1451, n1421, n1419, n1237, n1230);
xor  g1446 (n1456, n1416, n1423, n1427, n1414);
or   g1447 (n1448, n1231, n1431, n1236, n1429);
nand g1448 (n1476, n1374, n1353, n1449, n1241);
nand g1449 (n1480, n1354, n1450, n1445, n1451);
xor  g1450 (n1478, n1376, n1248, n1451, n1239);
nand g1451 (n1469, n1243, n1448, n1246);
or   g1452 (n1473, n1447, n1250, n1355, n1449);
xor  g1453 (n1475, n1244, n1249, n1450, n1447);
nand g1454 (n1477, n1451, n1450, n1446, n1445);
and  g1455 (n1472, n1451, n1447, n1448, n1247);
and  g1456 (n1481, n1373, n1354, n1445);
xnor g1457 (n1474, n1449, n1446, n1372);
or   g1458 (n1471, n1242, n1371, n1354, n1447);
nand g1459 (n1470, n1446, n1445, n1448, n1449);
xnor g1460 (n1479, n1375, n1450, n1245, n1240);
not  g1461 (n1482, n1474);
buf  g1462 (n1483, n1356);
buf  g1463 (n1486, n1355);
not  g1464 (n1484, n1470);
xnor g1465 (n1487, n1472, n1355);
nand g1466 (n1485, n1471, n1355, n1475, n1473);
xnor g1467 (n1490, n1484, n1358, n1482, n1356);
nor  g1468 (n1491, n1483, n1356, n1357);
xor  g1469 (n1488, n1357, n1251, n1486, n1252);
nand g1470 (n1489, n1487, n1357, n1485);
buf  g1471 (n1505, n1491);
not  g1472 (n1499, n1489);
buf  g1473 (n1506, n1444);
xnor g1474 (n1502, n1438, n1024, n1432);
nand g1475 (n1504, n1489, n1488, n1443, n1437);
xor  g1476 (n1492, n1488, n1254, n1437, n1489);
nand g1477 (n1507, n1443, n1491, n1452, n1435);
xor  g1478 (n1495, n1434, n1440, n1436, n1435);
or   g1479 (n1503, n1490, n1024, n1026, n1442);
nand g1480 (n1500, n1434, n1491, n1440, n1439);
and  g1481 (n1496, n1490, n1488, n1438, n1432);
or   g1482 (n1498, n1491, n1433, n1023, n1441);
nand g1483 (n1501, n1489, n1253, n1441, n1444);
and  g1484 (n1494, n1439, n1023, n1436, n1025);
nor  g1485 (n1497, n1433, n1025, n1022, n1442);
or   g1486 (n1493, n1490, n1490, n1431, n1488);
nor  g1487 (n1523, n1462, n1455, n1497, n1495);
nor  g1488 (n1521, n1460, n1462, n1492, n1463);
nand g1489 (n1524, n1458, n1464, n1496, n1493);
xor  g1490 (n1526, n1456, n1456, n1455, n1463);
xnor g1491 (n1511, n1455, n1466, n1261, n1257);
nand g1492 (n1519, n1453, n1493, n1452, n1460);
xor  g1493 (n1512, n1461, n1453, n1457, n1496);
and  g1494 (n1513, n1259, n1461, n1452, n1463);
nor  g1495 (n1518, n1458, n1465, n1494);
xnor g1496 (n1517, n1455, n1461, n1458);
or   g1497 (n1527, n1460, n1454, n1463, n1465);
or   g1498 (n1508, n1453, n1492, n1495, n1494);
xnor g1499 (n1510, n1457, n1461, n1258, n1454);
xnor g1500 (n1522, n1453, n1457, n1256, n1459);
and  g1501 (n1509, n1495, n1462, n1496, n1459);
xnor g1502 (n1525, n1460, n1494, n1260, n1464);
nor  g1503 (n1520, n1495, n1456, n1454);
nor  g1504 (n1515, n1493, n1465, n1459, n1496);
or   g1505 (n1528, n1494, n1452, n1459, n1255);
nor  g1506 (n1516, n1464, n1493, n1492, n1462);
nor  g1507 (n1514, n1456, n1457, n1464, n1492);
xnor g1508 (n1536, n1478, n1481, n1479, n1271);
xnor g1509 (n1533, n1268, n1262, n1467, n1466);
xor  g1510 (n1531, n1468, n1263, n1270, n1477);
nand g1511 (n1534, n1267, n1480, n1468, n1269);
xor  g1512 (n1537, n1509, n1264, n1468, n1508);
or   g1513 (n1529, n1509, n1468, n1467, n1266);
xor  g1514 (n1532, n1466, n1467, n1508);
nand g1515 (n1535, n1508, n1509, n1265, n1510);
xor  g1516 (n1530, n1509, n1466, n1508, n1476);
xnor g1517 (n1539, n1278, n1534, n1535, n1276);
xor  g1518 (n1540, n1537, n1282, n1281, n1274);
nor  g1519 (n1541, n1280, n1275, n1358, n1273);
or   g1520 (n1538, n1279, n1272, n1277, n1536);
buf  g1521 (n1545, n1539);
buf  g1522 (n1547, n1539);
nand g1523 (n1543, n1538, n1358);
not  g1524 (n1546, n1359);
buf  g1525 (n1542, n1538);
and  g1526 (n1544, n1358, n1538);
xnor g1527 (n1553, n1497, n1500, n1507, n1544);
xnor g1528 (n1555, n1545, n1498, n1511, n1510);
xnor g1529 (n1561, n1501, n1499, n1512);
and  g1530 (n1551, n1513, n1502, n1504);
nor  g1531 (n1552, n1543, n1542, n1500, n1545);
xor  g1532 (n1548, n1546, n1505, n1507, n1501);
and  g1533 (n1558, n1502, n1507, n1500);
xnor g1534 (n1556, n1513, n1546, n1543);
nor  g1535 (n1559, n1359, n1511, n1542);
nor  g1536 (n1557, n1497, n1503, n1505);
nor  g1537 (n1554, n1510, n1505, n1499, n1501);
nand g1538 (n1566, n1544, n1542, n1545, n1503);
nand g1539 (n1560, n1502, n1498, n1499, n1512);
nor  g1540 (n1567, n1543, n1513, n1505, n1283);
and  g1541 (n1550, n1500, n1498, n1546);
xnor g1542 (n1562, n1497, n1544, n1504);
xnor g1543 (n1565, n1542, n1503, n1511, n1499);
nor  g1544 (n1549, n1510, n1506, n1546);
xor  g1545 (n1564, n1504, n1513, n1545, n1506);
xor  g1546 (n1563, n1506, n1501, n1504, n1512);
xnor g1547 (n1572, n1284, n1516, n1566);
xnor g1548 (n1569, n1516, n1515, n1564, n1514);
xnor g1549 (n1571, n1285, n1514, n1286, n1515);
xnor g1550 (n1570, n1514, n1515, n1565, n1287);
xnor g1551 (n1568, n1515, n1567, n1563, n1514);
buf  g1552 (n1576, n1572);
buf  g1553 (n1580, n1570);
not  g1554 (n1581, n1518);
xor  g1555 (n1577, n1519, n1517, n1520);
nand g1556 (n1574, n1568, n1518, n1519);
xnor g1557 (n1575, n1519, n1517);
nor  g1558 (n1573, n1520, n1570, n1519);
or   g1559 (n1582, n1568, n1572);
xnor g1560 (n1579, n1571, n1520, n1518);
xor  g1561 (n1583, n1571, n1569, n1516);
nand g1562 (n1578, n1518, n1520, n1517, n1569);
nor  g1563 (n1597, n1028, n1027, n1581, n1578);
xor  g1564 (n1612, n1575, n1521, n1579, n1578);
nor  g1565 (n1592, n1521, n1540, n1541, n1360);
nand g1566 (n1610, n1524, n1027, n1577, n1578);
or   g1567 (n1603, n1576, n1575, n1540, n1577);
and  g1568 (n1607, n1521, n1360, n1525, n1581);
or   g1569 (n1606, n1583, n1291, n1547, n1290);
nand g1570 (n1601, n1576, n1573, n1525, n1579);
and  g1571 (n1590, n1289, n1581, n1580, n1026);
xor  g1572 (n1613, n412, n1524, n1527, n1523);
nor  g1573 (n1605, n1029, n1524, n1539, n1522);
or   g1574 (n1596, n1527, n1541, n1578, n1582);
or   g1575 (n1588, n1360, n1524, n1527, n1541);
xor  g1576 (n1614, n1288, n1361, n1575, n412);
nor  g1577 (n1598, n1302, n1292, n1573, n1522);
nand g1578 (n1602, n1526, n1574, n1028, n1547);
and  g1579 (n1586, n1527, n1579, n1574, n1522);
xnor g1580 (n1593, n1579, n1528, n1541);
xnor g1581 (n1584, n1523, n1574, n1303, n1580);
xnor g1582 (n1589, n1300, n1583, n1540);
nor  g1583 (n1604, n1580, n1526, n1581);
xnor g1584 (n1599, n1297, n1298, n1575, n1526);
and  g1585 (n1609, n1583, n1580, n1301, n1582);
xnor g1586 (n1611, n1577, n1293, n1547, n1029);
and  g1587 (n1600, n1525, n1576, n1296, n1540);
xor  g1588 (n1587, n1523, n1576, n1582, n1299);
or   g1589 (n1594, n1359, n1577, n1582, n1522);
or   g1590 (n1595, n1361, n1574, n1294, n1528);
xor  g1591 (n1608, n1547, n1360, n1528, n1295);
nor  g1592 (n1591, n1525, n1573, n1521, n1361);
or   g1593 (n1585, n1573, n1523, n1361, n1539);
nor  g1594 (n1656, n1044, n1074, n413, n1052);
xor  g1595 (n1648, n1588, n1606, n1038, n1086);
nand g1596 (n1631, n1070, n1051, n1068, n1093);
and  g1597 (n1642, n1050, n1590, n1586, n1064);
xor  g1598 (n1652, n1076, n1054, n1038);
xnor g1599 (n1647, n1056, n1052, n1065, n1040);
and  g1600 (n1644, n415, n1079, n1613, n1082);
nand g1601 (n1657, n1603, n1089, n1609, n1036);
nor  g1602 (n1640, n1058, n1605, n1080, n415);
xor  g1603 (n1635, n1609, n1043, n1057, n1612);
nand g1604 (n1617, n1614, n1604, n1073, n1047);
and  g1605 (n1646, n1055, n1085, n1597, n1090);
or   g1606 (n1658, n1034, n1036, n1077, n1061);
or   g1607 (n1649, n1065, n1600, n1048, n1033);
or   g1608 (n1660, n414, n1040, n1596, n1598);
nor  g1609 (n1616, n1606, n1091, n1611, n1601);
xor  g1610 (n1636, n1614, n1073, n1030, n1044);
nand g1611 (n1653, n1084, n1602, n1033, n1047);
or   g1612 (n1643, n1050, n1049, n1039, n1072);
and  g1613 (n1615, n1037, n1046, n1080, n1089);
and  g1614 (n1626, n1075, n1083, n1603, n414);
nand g1615 (n1638, n1070, n413, n1076, n414);
or   g1616 (n1637, n1030, n1594, n1045, n1081);
nor  g1617 (n1633, n1088, n1083, n1607, n1041);
or   g1618 (n1628, n1031, n1042, n1589, n1037);
nand g1619 (n1629, n1592, n1591, n1593, n1074);
or   g1620 (n1655, n1599, n1071, n1068, n1062);
nand g1621 (n1624, n1094, n1045, n414, n1595);
nand g1622 (n1622, n413, n1046, n1043, n1091);
and  g1623 (n1659, n1049, n1056, n1600, n1092);
xor  g1624 (n1632, n1093, n1067, n1060, n1081);
nor  g1625 (n1634, n1064, n1072, n1090, n1053);
xor  g1626 (n1639, n1039, n1087, n1058, n1063);
and  g1627 (n1627, n1032, n1077, n1088, n1605);
xnor g1628 (n1641, n1610, n1079, n1084, n1055);
or   g1629 (n1623, n1032, n1053, n1601, n1599);
xnor g1630 (n1630, n1041, n1057, n1612, n1082);
nor  g1631 (n1619, n1078, n415, n1608, n1059);
and  g1632 (n1650, n1069, n1066, n1059, n1602);
or   g1633 (n1620, n1604, n1060, n1585, n1063);
xor  g1634 (n1661, n1078, n1608, n415, n1587);
and  g1635 (n1625, n1042, n1048, n413, n1034);
xor  g1636 (n1651, n1071, n1031, n1085, n1061);
nor  g1637 (n1645, n1610, n1051, n1035, n1086);
nor  g1638 (n1618, n1069, n1092, n1067, n1087);
and  g1639 (n1654, n1066, n1613, n1075, n1611);
xor  g1640 (n1621, n1607, n1584, n1062, n1035);
nor  g1641 (n1663, n1654, n1627, n1621, n1624);
or   g1642 (n1667, n1638, n1635, n1628, n1619);
xor  g1643 (n1668, n1637, n1655, n1623, n1094);
nor  g1644 (n1670, n1095, n1641, n1643, n1631);
nand g1645 (n1669, n1646, n1633, n1640, n1653);
nand g1646 (n1666, n1652, n1642, n1648, n1659);
nand g1647 (n1674, n1639, n1657, n1636, n1658);
nor  g1648 (n1665, n20, n1632, n1661, n1647);
xnor g1649 (n1673, n1615, n1630, n1651, n1625);
xnor g1650 (n1671, n1649, n1622, n1645, n1620);
nor  g1651 (n1672, n1661, n1626, n1660, n1656);
xnor g1652 (n1664, n1644, n1617, n1650, n1616);
and  g1653 (n1662, n1629, n1618, n1634, n1095);
endmodule
