

module Stat_1546_16_7
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n1463,
  n1525,
  n1491,
  n1498,
  n1529,
  n1523,
  n1486,
  n1482,
  n1494,
  n1527,
  n1502,
  n1478,
  n1514,
  n1493,
  n1499,
  n1518,
  n1507,
  n1517,
  n1492,
  n1475,
  n1533,
  n1509,
  n1508,
  n1496,
  n1503,
  n1459,
  n1563,
  n1565,
  n1566,
  n1562,
  n1561,
  n1564,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1463;
  output n1525;
  output n1491;
  output n1498;
  output n1529;
  output n1523;
  output n1486;
  output n1482;
  output n1494;
  output n1527;
  output n1502;
  output n1478;
  output n1514;
  output n1493;
  output n1499;
  output n1518;
  output n1507;
  output n1517;
  output n1492;
  output n1475;
  output n1533;
  output n1509;
  output n1508;
  output n1496;
  output n1503;
  output n1459;
  output n1563;
  output n1565;
  output n1566;
  output n1562;
  output n1561;
  output n1564;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1476;
  wire n1477;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1495;
  wire n1497;
  wire n1500;
  wire n1501;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1515;
  wire n1516;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1524;
  wire n1526;
  wire n1528;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n90,
    n6
  );


  not
  g1
  (
    n36,
    n12
  );


  buf
  g2
  (
    n86,
    n12
  );


  not
  g3
  (
    n26,
    n18
  );


  not
  g4
  (
    n80,
    n14
  );


  not
  g5
  (
    n21,
    n4
  );


  buf
  g6
  (
    n66,
    n2
  );


  not
  g7
  (
    n67,
    n19
  );


  not
  g8
  (
    n69,
    n19
  );


  buf
  g9
  (
    n62,
    n19
  );


  not
  g10
  (
    n54,
    n5
  );


  not
  g11
  (
    n61,
    n18
  );


  buf
  g12
  (
    n33,
    n14
  );


  not
  g13
  (
    n79,
    n12
  );


  buf
  g14
  (
    n31,
    n15
  );


  not
  g15
  (
    n45,
    n20
  );


  buf
  g16
  (
    n58,
    n9
  );


  buf
  g17
  (
    n64,
    n7
  );


  buf
  g18
  (
    KeyWire_0_1,
    n7
  );


  buf
  g19
  (
    n73,
    n20
  );


  buf
  g20
  (
    n60,
    n15
  );


  buf
  g21
  (
    n55,
    n3
  );


  not
  g22
  (
    n40,
    n4
  );


  buf
  g23
  (
    n38,
    n17
  );


  buf
  g24
  (
    n50,
    n11
  );


  buf
  g25
  (
    n24,
    n18
  );


  buf
  g26
  (
    n43,
    n2
  );


  not
  g27
  (
    n87,
    n11
  );


  not
  g28
  (
    n84,
    n7
  );


  not
  g29
  (
    n37,
    n12
  );


  buf
  g30
  (
    n100,
    n18
  );


  buf
  g31
  (
    n99,
    n17
  );


  not
  g32
  (
    n30,
    n2
  );


  buf
  g33
  (
    n97,
    n2
  );


  not
  g34
  (
    n49,
    n4
  );


  buf
  g35
  (
    n44,
    n6
  );


  buf
  g36
  (
    n94,
    n20
  );


  not
  g37
  (
    n82,
    n1
  );


  buf
  g38
  (
    n65,
    n10
  );


  buf
  g39
  (
    n93,
    n1
  );


  not
  g40
  (
    n63,
    n11
  );


  not
  g41
  (
    n35,
    n16
  );


  buf
  g42
  (
    n76,
    n13
  );


  buf
  g43
  (
    n32,
    n13
  );


  not
  g44
  (
    n74,
    n8
  );


  buf
  g45
  (
    n28,
    n3
  );


  not
  g46
  (
    n56,
    n17
  );


  buf
  g47
  (
    n34,
    n13
  );


  not
  g48
  (
    n72,
    n20
  );


  buf
  g49
  (
    n78,
    n9
  );


  buf
  g50
  (
    n27,
    n19
  );


  not
  g51
  (
    n91,
    n14
  );


  not
  g52
  (
    n85,
    n7
  );


  not
  g53
  (
    n42,
    n17
  );


  not
  g54
  (
    n71,
    n8
  );


  not
  g55
  (
    n52,
    n8
  );


  not
  g56
  (
    n47,
    n11
  );


  buf
  g57
  (
    n22,
    n4
  );


  not
  g58
  (
    n57,
    n14
  );


  buf
  g59
  (
    n81,
    n16
  );


  not
  g60
  (
    n23,
    n3
  );


  buf
  g61
  (
    n96,
    n9
  );


  buf
  g62
  (
    n92,
    n10
  );


  not
  g63
  (
    n70,
    n13
  );


  buf
  g64
  (
    n25,
    n6
  );


  buf
  g65
  (
    n51,
    n1
  );


  buf
  g66
  (
    n68,
    n5
  );


  not
  g67
  (
    n29,
    n9
  );


  not
  g68
  (
    n48,
    n6
  );


  not
  g69
  (
    n53,
    n3
  );


  buf
  g70
  (
    n98,
    n16
  );


  buf
  g71
  (
    n75,
    n5
  );


  buf
  g72
  (
    n46,
    n10
  );


  buf
  g73
  (
    n83,
    n5
  );


  buf
  g74
  (
    n39,
    n15
  );


  not
  g75
  (
    n89,
    n15
  );


  buf
  g76
  (
    n88,
    n10
  );


  not
  g77
  (
    n77,
    n1
  );


  buf
  g78
  (
    n95,
    n8
  );


  buf
  g79
  (
    n41,
    n16
  );


  buf
  g80
  (
    n317,
    n26
  );


  buf
  g81
  (
    n110,
    n30
  );


  not
  g82
  (
    n320,
    n30
  );


  buf
  g83
  (
    n183,
    n62
  );


  not
  g84
  (
    n177,
    n35
  );


  not
  g85
  (
    n247,
    n65
  );


  buf
  g86
  (
    n234,
    n51
  );


  buf
  g87
  (
    n132,
    n32
  );


  buf
  g88
  (
    n202,
    n51
  );


  not
  g89
  (
    n187,
    n48
  );


  buf
  g90
  (
    n149,
    n21
  );


  not
  g91
  (
    n163,
    n61
  );


  buf
  g92
  (
    n270,
    n68
  );


  buf
  g93
  (
    n190,
    n38
  );


  not
  g94
  (
    n304,
    n47
  );


  not
  g95
  (
    n221,
    n42
  );


  not
  g96
  (
    n273,
    n49
  );


  not
  g97
  (
    n294,
    n34
  );


  buf
  g98
  (
    n167,
    n45
  );


  not
  g99
  (
    n267,
    n70
  );


  buf
  g100
  (
    n271,
    n69
  );


  not
  g101
  (
    n170,
    n53
  );


  not
  g102
  (
    n291,
    n39
  );


  buf
  g103
  (
    n116,
    n61
  );


  buf
  g104
  (
    n251,
    n74
  );


  buf
  g105
  (
    n309,
    n40
  );


  not
  g106
  (
    n269,
    n58
  );


  not
  g107
  (
    n161,
    n50
  );


  buf
  g108
  (
    n101,
    n56
  );


  buf
  g109
  (
    n121,
    n27
  );


  not
  g110
  (
    n112,
    n27
  );


  buf
  g111
  (
    n287,
    n56
  );


  not
  g112
  (
    n254,
    n22
  );


  not
  g113
  (
    n168,
    n44
  );


  not
  g114
  (
    n148,
    n72
  );


  not
  g115
  (
    n272,
    n41
  );


  buf
  g116
  (
    n201,
    n32
  );


  not
  g117
  (
    n244,
    n66
  );


  not
  g118
  (
    n230,
    n45
  );


  buf
  g119
  (
    n240,
    n67
  );


  not
  g120
  (
    n138,
    n29
  );


  not
  g121
  (
    n150,
    n21
  );


  not
  g122
  (
    n140,
    n70
  );


  not
  g123
  (
    n172,
    n47
  );


  not
  g124
  (
    n278,
    n22
  );


  not
  g125
  (
    n152,
    n33
  );


  not
  g126
  (
    n281,
    n46
  );


  buf
  g127
  (
    n204,
    n68
  );


  buf
  g128
  (
    n292,
    n39
  );


  not
  g129
  (
    n319,
    n40
  );


  not
  g130
  (
    n127,
    n31
  );


  buf
  g131
  (
    n295,
    n65
  );


  not
  g132
  (
    n166,
    n49
  );


  not
  g133
  (
    n308,
    n69
  );


  buf
  g134
  (
    n178,
    n65
  );


  buf
  g135
  (
    n155,
    n55
  );


  not
  g136
  (
    n113,
    n59
  );


  buf
  g137
  (
    n164,
    n44
  );


  buf
  g138
  (
    n122,
    n42
  );


  not
  g139
  (
    n257,
    n22
  );


  not
  g140
  (
    n195,
    n34
  );


  not
  g141
  (
    n198,
    n24
  );


  buf
  g142
  (
    n186,
    n71
  );


  not
  g143
  (
    n282,
    n64
  );


  not
  g144
  (
    n139,
    n28
  );


  not
  g145
  (
    n249,
    n24
  );


  buf
  g146
  (
    n252,
    n61
  );


  not
  g147
  (
    n258,
    n55
  );


  not
  g148
  (
    n214,
    n46
  );


  not
  g149
  (
    n297,
    n28
  );


  not
  g150
  (
    n222,
    n59
  );


  buf
  g151
  (
    n275,
    n56
  );


  buf
  g152
  (
    n268,
    n54
  );


  buf
  g153
  (
    n266,
    n25
  );


  not
  g154
  (
    n318,
    n46
  );


  buf
  g155
  (
    n174,
    n25
  );


  not
  g156
  (
    n236,
    n62
  );


  buf
  g157
  (
    n165,
    n72
  );


  buf
  g158
  (
    n211,
    n33
  );


  not
  g159
  (
    n147,
    n56
  );


  not
  g160
  (
    n238,
    n51
  );


  buf
  g161
  (
    n302,
    n71
  );


  buf
  g162
  (
    n115,
    n72
  );


  not
  g163
  (
    n231,
    n57
  );


  not
  g164
  (
    n216,
    n23
  );


  buf
  g165
  (
    n185,
    n66
  );


  not
  g166
  (
    n108,
    n48
  );


  not
  g167
  (
    n248,
    n40
  );


  buf
  g168
  (
    n310,
    n33
  );


  buf
  g169
  (
    n215,
    n54
  );


  not
  g170
  (
    n223,
    n39
  );


  not
  g171
  (
    n137,
    n42
  );


  not
  g172
  (
    n109,
    n24
  );


  buf
  g173
  (
    n158,
    n67
  );


  buf
  g174
  (
    n182,
    n62
  );


  not
  g175
  (
    n134,
    n41
  );


  not
  g176
  (
    n144,
    n68
  );


  not
  g177
  (
    n301,
    n63
  );


  buf
  g178
  (
    n306,
    n54
  );


  not
  g179
  (
    n184,
    n53
  );


  buf
  g180
  (
    n171,
    n55
  );


  not
  g181
  (
    n135,
    n57
  );


  buf
  g182
  (
    n243,
    n29
  );


  buf
  g183
  (
    n225,
    n38
  );


  buf
  g184
  (
    n197,
    n64
  );


  buf
  g185
  (
    n262,
    n43
  );


  buf
  g186
  (
    n298,
    n36
  );


  not
  g187
  (
    n123,
    n73
  );


  not
  g188
  (
    n286,
    n75
  );


  not
  g189
  (
    n189,
    n75
  );


  buf
  g190
  (
    n232,
    n23
  );


  buf
  g191
  (
    n284,
    n75
  );


  buf
  g192
  (
    n207,
    n67
  );


  not
  g193
  (
    n142,
    n60
  );


  not
  g194
  (
    n241,
    n23
  );


  not
  g195
  (
    n194,
    n70
  );


  buf
  g196
  (
    n299,
    n73
  );


  not
  g197
  (
    n176,
    n63
  );


  buf
  g198
  (
    n235,
    n37
  );


  not
  g199
  (
    n255,
    n49
  );


  not
  g200
  (
    n143,
    n44
  );


  not
  g201
  (
    n226,
    n70
  );


  buf
  g202
  (
    n125,
    n64
  );


  buf
  g203
  (
    n120,
    n37
  );


  not
  g204
  (
    n102,
    n31
  );


  not
  g205
  (
    n175,
    n36
  );


  not
  g206
  (
    n229,
    n69
  );


  buf
  g207
  (
    n233,
    n69
  );


  not
  g208
  (
    n114,
    n26
  );


  buf
  g209
  (
    n276,
    n48
  );


  buf
  g210
  (
    n191,
    n49
  );


  buf
  g211
  (
    n316,
    n50
  );


  buf
  g212
  (
    n300,
    n48
  );


  buf
  g213
  (
    n129,
    n57
  );


  buf
  g214
  (
    n307,
    n37
  );


  buf
  g215
  (
    n133,
    n25
  );


  not
  g216
  (
    n131,
    n73
  );


  not
  g217
  (
    n289,
    n72
  );


  buf
  g218
  (
    n192,
    n52
  );


  buf
  g219
  (
    n200,
    n27
  );


  buf
  g220
  (
    KeyWire_0_9,
    n53
  );


  buf
  g221
  (
    n136,
    n68
  );


  buf
  g222
  (
    n224,
    n74
  );


  not
  g223
  (
    n228,
    n35
  );


  buf
  g224
  (
    n103,
    n50
  );


  not
  g225
  (
    n181,
    n47
  );


  not
  g226
  (
    n314,
    n52
  );


  not
  g227
  (
    n218,
    n45
  );


  not
  g228
  (
    n104,
    n52
  );


  buf
  g229
  (
    n303,
    n30
  );


  not
  g230
  (
    n315,
    n59
  );


  buf
  g231
  (
    n203,
    n57
  );


  not
  g232
  (
    n246,
    n73
  );


  not
  g233
  (
    n124,
    n23
  );


  not
  g234
  (
    n146,
    n64
  );


  not
  g235
  (
    n293,
    n28
  );


  not
  g236
  (
    n126,
    n43
  );


  not
  g237
  (
    n154,
    n59
  );


  not
  g238
  (
    n162,
    n71
  );


  buf
  g239
  (
    n217,
    n67
  );


  buf
  g240
  (
    n212,
    n33
  );


  buf
  g241
  (
    n219,
    n40
  );


  buf
  g242
  (
    n209,
    n26
  );


  not
  g243
  (
    n105,
    n71
  );


  not
  g244
  (
    n261,
    n74
  );


  not
  g245
  (
    n242,
    n58
  );


  not
  g246
  (
    n111,
    n32
  );


  buf
  g247
  (
    n106,
    n66
  );


  buf
  g248
  (
    n279,
    n46
  );


  not
  g249
  (
    n199,
    n31
  );


  buf
  g250
  (
    n274,
    n35
  );


  not
  g251
  (
    n296,
    n50
  );


  not
  g252
  (
    n151,
    n74
  );


  not
  g253
  (
    n118,
    n22
  );


  not
  g254
  (
    n265,
    n41
  );


  not
  g255
  (
    n188,
    n42
  );


  buf
  g256
  (
    n169,
    n51
  );


  buf
  g257
  (
    n206,
    n21
  );


  not
  g258
  (
    n312,
    n24
  );


  not
  g259
  (
    n260,
    n65
  );


  buf
  g260
  (
    n205,
    n28
  );


  buf
  g261
  (
    n264,
    n38
  );


  buf
  g262
  (
    n173,
    n27
  );


  buf
  g263
  (
    n157,
    n34
  );


  buf
  g264
  (
    n107,
    n60
  );


  buf
  g265
  (
    n256,
    n60
  );


  not
  g266
  (
    n196,
    n63
  );


  buf
  g267
  (
    n160,
    n38
  );


  buf
  g268
  (
    n253,
    n44
  );


  buf
  g269
  (
    n213,
    n61
  );


  not
  g270
  (
    n227,
    n66
  );


  buf
  g271
  (
    n239,
    n36
  );


  not
  g272
  (
    n263,
    n45
  );


  buf
  g273
  (
    n220,
    n25
  );


  not
  g274
  (
    n277,
    n31
  );


  not
  g275
  (
    n280,
    n58
  );


  not
  g276
  (
    n117,
    n36
  );


  buf
  g277
  (
    n145,
    n29
  );


  buf
  g278
  (
    n130,
    n30
  );


  buf
  g279
  (
    n153,
    n32
  );


  not
  g280
  (
    n290,
    n58
  );


  buf
  g281
  (
    n193,
    n21
  );


  buf
  g282
  (
    n128,
    n39
  );


  buf
  g283
  (
    n179,
    n62
  );


  buf
  g284
  (
    n288,
    n34
  );


  not
  g285
  (
    n159,
    n53
  );


  buf
  g286
  (
    n208,
    n35
  );


  buf
  g287
  (
    n305,
    n52
  );


  not
  g288
  (
    n119,
    n75
  );


  buf
  g289
  (
    n311,
    n55
  );


  buf
  g290
  (
    n156,
    n41
  );


  buf
  g291
  (
    n250,
    n54
  );


  not
  g292
  (
    n283,
    n60
  );


  buf
  g293
  (
    n259,
    n63
  );


  buf
  g294
  (
    n285,
    n43
  );


  buf
  g295
  (
    n245,
    n29
  );


  buf
  g296
  (
    n237,
    n37
  );


  not
  g297
  (
    n180,
    n43
  );


  not
  g298
  (
    n210,
    n47
  );


  buf
  g299
  (
    n313,
    n26
  );


  not
  g300
  (
    n460,
    n222
  );


  buf
  g301
  (
    n406,
    n126
  );


  not
  g302
  (
    n339,
    n173
  );


  not
  g303
  (
    n374,
    n163
  );


  not
  g304
  (
    n356,
    n261
  );


  not
  g305
  (
    n545,
    n179
  );


  buf
  g306
  (
    n376,
    n224
  );


  not
  g307
  (
    n405,
    n237
  );


  not
  g308
  (
    n440,
    n117
  );


  not
  g309
  (
    n365,
    n183
  );


  not
  g310
  (
    n515,
    n271
  );


  not
  g311
  (
    n419,
    n184
  );


  buf
  g312
  (
    n443,
    n174
  );


  not
  g313
  (
    n409,
    n284
  );


  not
  g314
  (
    n527,
    n243
  );


  not
  g315
  (
    n341,
    n121
  );


  buf
  g316
  (
    n422,
    n266
  );


  buf
  g317
  (
    n368,
    n118
  );


  buf
  g318
  (
    n474,
    n102
  );


  buf
  g319
  (
    n383,
    n84
  );


  not
  g320
  (
    n471,
    n238
  );


  buf
  g321
  (
    n458,
    n259
  );


  not
  g322
  (
    n377,
    n215
  );


  not
  g323
  (
    n507,
    n201
  );


  not
  g324
  (
    n476,
    n293
  );


  buf
  g325
  (
    n509,
    n290
  );


  buf
  g326
  (
    n516,
    n153
  );


  not
  g327
  (
    n431,
    n185
  );


  buf
  g328
  (
    n540,
    n195
  );


  buf
  g329
  (
    n353,
    n228
  );


  buf
  g330
  (
    n326,
    n278
  );


  buf
  g331
  (
    n352,
    n143
  );


  buf
  g332
  (
    n434,
    n107
  );


  not
  g333
  (
    n459,
    n263
  );


  not
  g334
  (
    n529,
    n210
  );


  buf
  g335
  (
    n541,
    n76
  );


  not
  g336
  (
    n416,
    n258
  );


  not
  g337
  (
    n512,
    n283
  );


  not
  g338
  (
    n508,
    n247
  );


  not
  g339
  (
    n518,
    n231
  );


  buf
  g340
  (
    n501,
    n249
  );


  buf
  g341
  (
    n487,
    n133
  );


  not
  g342
  (
    n333,
    n214
  );


  not
  g343
  (
    n468,
    n157
  );


  buf
  g344
  (
    n382,
    n138
  );


  buf
  g345
  (
    n534,
    n113
  );


  not
  g346
  (
    KeyWire_0_4,
    n223
  );


  not
  g347
  (
    n371,
    n241
  );


  not
  g348
  (
    n522,
    n274
  );


  not
  g349
  (
    n343,
    n263
  );


  not
  g350
  (
    n400,
    n140
  );


  buf
  g351
  (
    n439,
    n269
  );


  not
  g352
  (
    n362,
    n123
  );


  buf
  g353
  (
    n322,
    n113
  );


  buf
  g354
  (
    n499,
    n229
  );


  not
  g355
  (
    n526,
    n144
  );


  not
  g356
  (
    n415,
    n181
  );


  buf
  g357
  (
    n493,
    n203
  );


  not
  g358
  (
    n513,
    n235
  );


  not
  g359
  (
    n506,
    n260
  );


  not
  g360
  (
    n327,
    n191
  );


  not
  g361
  (
    n480,
    n79
  );


  not
  g362
  (
    n418,
    n172
  );


  buf
  g363
  (
    n449,
    n160
  );


  buf
  g364
  (
    n373,
    n233
  );


  buf
  g365
  (
    n543,
    n130
  );


  buf
  g366
  (
    n492,
    n115
  );


  buf
  g367
  (
    n452,
    n209
  );


  buf
  g368
  (
    n359,
    n242
  );


  not
  g369
  (
    n519,
    n234
  );


  buf
  g370
  (
    n329,
    n256
  );


  buf
  g371
  (
    n425,
    n134
  );


  buf
  g372
  (
    n454,
    n233
  );


  buf
  g373
  (
    n325,
    n125
  );


  buf
  g374
  (
    n496,
    n200
  );


  not
  g375
  (
    n504,
    n298
  );


  buf
  g376
  (
    n494,
    n204
  );


  not
  g377
  (
    n530,
    n248
  );


  not
  g378
  (
    n427,
    n83
  );


  not
  g379
  (
    n336,
    n121
  );


  buf
  g380
  (
    n453,
    n301
  );


  buf
  g381
  (
    n503,
    n146
  );


  not
  g382
  (
    n381,
    n163
  );


  not
  g383
  (
    n348,
    n179
  );


  not
  g384
  (
    n389,
    n83
  );


  buf
  g385
  (
    n472,
    n268
  );


  xor
  g386
  (
    n528,
    n126,
    n114,
    n160,
    n218
  );


  nor
  g387
  (
    n505,
    n300,
    n217,
    n287,
    n144
  );


  or
  g388
  (
    n510,
    n78,
    n290,
    n188,
    n133
  );


  xor
  g389
  (
    n392,
    n199,
    n133,
    n267,
    n106
  );


  xor
  g390
  (
    n364,
    n277,
    n114,
    n128,
    n298
  );


  nor
  g391
  (
    n435,
    n186,
    n135,
    n256,
    n187
  );


  xnor
  g392
  (
    n489,
    n276,
    n109,
    n157,
    n232
  );


  nor
  g393
  (
    n429,
    n270,
    n300,
    n173,
    n76
  );


  xnor
  g394
  (
    n398,
    n164,
    n268,
    n168,
    n244
  );


  nor
  g395
  (
    n369,
    n220,
    n205,
    n166,
    n128
  );


  nand
  g396
  (
    n464,
    n129,
    n299,
    n140,
    n303
  );


  nand
  g397
  (
    n331,
    n103,
    n225,
    n282,
    n297
  );


  and
  g398
  (
    n450,
    n249,
    n127,
    n260,
    n152
  );


  nor
  g399
  (
    n384,
    n136,
    n277,
    n214,
    n302
  );


  and
  g400
  (
    n470,
    n206,
    n119,
    n216,
    n207
  );


  nand
  g401
  (
    n342,
    n169,
    n120,
    n181,
    n165
  );


  or
  g402
  (
    n536,
    n81,
    n268,
    n219,
    n195
  );


  xnor
  g403
  (
    n351,
    n270,
    n81,
    n208,
    n281
  );


  xnor
  g404
  (
    n495,
    n246,
    n131,
    n222,
    n176
  );


  nand
  g405
  (
    n535,
    n147,
    n271,
    n261,
    n186
  );


  and
  g406
  (
    n403,
    n250,
    n151,
    n303,
    n249
  );


  xnor
  g407
  (
    n484,
    n265,
    n186,
    n141,
    n213
  );


  or
  g408
  (
    n532,
    n105,
    n191,
    n187,
    n142
  );


  xnor
  g409
  (
    n511,
    n114,
    n232,
    n178,
    n211
  );


  xor
  g410
  (
    n396,
    n107,
    n83,
    n280,
    n164
  );


  nand
  g411
  (
    n391,
    n208,
    n239,
    n178,
    n250
  );


  and
  g412
  (
    KeyWire_0_11,
    n255,
    n122,
    n252,
    n292
  );


  xnor
  g413
  (
    n481,
    n202,
    n262,
    n240,
    n259
  );


  xnor
  g414
  (
    n433,
    n188,
    n223,
    n226,
    n242
  );


  xnor
  g415
  (
    n525,
    n266,
    n77,
    n119,
    n182
  );


  nand
  g416
  (
    n500,
    n175,
    n161,
    n168,
    n103
  );


  or
  g417
  (
    n537,
    n273,
    n206,
    n181,
    n101
  );


  or
  g418
  (
    n442,
    n279,
    n253,
    n178,
    n290
  );


  xnor
  g419
  (
    n413,
    n251,
    n245,
    n182,
    n104
  );


  nor
  g420
  (
    n401,
    n300,
    n169,
    n301,
    n154
  );


  nand
  g421
  (
    n432,
    n123,
    n199,
    n197
  );


  nand
  g422
  (
    n441,
    n256,
    n198,
    n156,
    n289
  );


  xor
  g423
  (
    n482,
    n156,
    n205,
    n183,
    n157
  );


  xor
  g424
  (
    n363,
    n223,
    n166,
    n211,
    n177
  );


  nand
  g425
  (
    n335,
    n278,
    n279,
    n159,
    n229
  );


  nand
  g426
  (
    n358,
    n167,
    n221,
    n158,
    n185
  );


  and
  g427
  (
    n350,
    n299,
    n155,
    n250,
    n105
  );


  xor
  g428
  (
    n379,
    n215,
    n287,
    n125,
    n255
  );


  and
  g429
  (
    n324,
    n276,
    n255,
    n280,
    n227
  );


  nor
  g430
  (
    n466,
    n248,
    n102,
    n138,
    n153
  );


  xnor
  g431
  (
    n390,
    n130,
    n201,
    n207,
    n239
  );


  nand
  g432
  (
    n447,
    n122,
    n270,
    n110,
    n267
  );


  or
  g433
  (
    n323,
    n231,
    n171,
    n286,
    n122
  );


  nand
  g434
  (
    n349,
    n116,
    n247,
    n280,
    n151
  );


  xor
  g435
  (
    n437,
    n111,
    n190,
    n288,
    n212
  );


  and
  g436
  (
    n491,
    n292,
    n170,
    n293,
    n214
  );


  xor
  g437
  (
    n361,
    n198,
    n182,
    n272,
    n170
  );


  and
  g438
  (
    n355,
    n175,
    n275,
    n172,
    n174
  );


  and
  g439
  (
    n385,
    n200,
    n207,
    n166,
    n108
  );


  xor
  g440
  (
    n370,
    n264,
    n237,
    n297,
    n233
  );


  xor
  g441
  (
    n485,
    n272,
    n171,
    n149,
    n284
  );


  xnor
  g442
  (
    n465,
    n170,
    n202,
    n302,
    n184
  );


  or
  g443
  (
    n539,
    n248,
    n298,
    n148,
    n136
  );


  or
  g444
  (
    n531,
    n262,
    n302,
    n78,
    n116
  );


  nand
  g445
  (
    n520,
    n160,
    n81,
    n176,
    n303
  );


  or
  g446
  (
    n330,
    n210,
    n132,
    n301,
    n111
  );


  xor
  g447
  (
    n546,
    n162,
    n197,
    n154,
    n165
  );


  nor
  g448
  (
    n486,
    n196,
    n299,
    n135,
    n149
  );


  or
  g449
  (
    n430,
    n209,
    n130,
    n200,
    n115
  );


  and
  g450
  (
    n414,
    n269,
    n258,
    n302,
    n267
  );


  xor
  g451
  (
    n372,
    n108,
    n193,
    n163,
    n284
  );


  nand
  g452
  (
    n448,
    n81,
    n209,
    n198,
    n303
  );


  nor
  g453
  (
    n347,
    n286,
    n82,
    n183,
    n254
  );


  xor
  g454
  (
    n490,
    n220,
    n80,
    n116,
    n297
  );


  xor
  g455
  (
    n388,
    n257,
    n192,
    n241,
    n235
  );


  or
  g456
  (
    n475,
    n145,
    n105,
    n172,
    n296
  );


  and
  g457
  (
    n445,
    n266,
    n145,
    n289,
    n298
  );


  xnor
  g458
  (
    n338,
    n126,
    n272,
    n230,
    n228
  );


  nand
  g459
  (
    n340,
    n239,
    n230,
    n154,
    n139
  );


  nand
  g460
  (
    n514,
    n127,
    n82,
    n243,
    n190
  );


  xnor
  g461
  (
    n420,
    n137,
    n104,
    n112,
    n203
  );


  or
  g462
  (
    n438,
    n238,
    n143,
    n106,
    n152
  );


  xnor
  g463
  (
    n542,
    n218,
    n234,
    n80,
    n196
  );


  and
  g464
  (
    n360,
    n190,
    n79,
    n228,
    n222
  );


  or
  g465
  (
    n344,
    n211,
    n79,
    n296,
    n110
  );


  nor
  g466
  (
    n544,
    n164,
    n131,
    n294,
    n144
  );


  xor
  g467
  (
    n473,
    n257,
    n254,
    n106,
    n76
  );


  and
  g468
  (
    n428,
    n136,
    n213,
    n296,
    n253
  );


  nand
  g469
  (
    n497,
    n244,
    n218,
    n247,
    n278
  );


  nor
  g470
  (
    n446,
    n216,
    n243,
    n118,
    n111
  );


  and
  g471
  (
    n479,
    n204,
    n158,
    n225,
    n219
  );


  xnor
  g472
  (
    n457,
    n288,
    n245,
    n224,
    n155
  );


  xor
  g473
  (
    n521,
    n151,
    n155,
    n240,
    n188
  );


  or
  g474
  (
    n467,
    n78,
    n192,
    n179,
    n221
  );


  xnor
  g475
  (
    n517,
    n252,
    n78,
    n156,
    n147
  );


  and
  g476
  (
    n451,
    n177,
    n109,
    n120,
    n221
  );


  xor
  g477
  (
    n334,
    n153,
    n115,
    n206,
    n212
  );


  nor
  g478
  (
    n488,
    n118,
    n124,
    n208,
    n162
  );


  or
  g479
  (
    n523,
    n140,
    n150,
    n142,
    n77
  );


  nor
  g480
  (
    n478,
    n264,
    n251,
    n224,
    n82
  );


  xor
  g481
  (
    n462,
    n236,
    n257,
    n176,
    n273
  );


  nand
  g482
  (
    n444,
    n125,
    n197,
    n132,
    n230
  );


  or
  g483
  (
    n456,
    n137,
    n152,
    n189,
    n205
  );


  or
  g484
  (
    n423,
    n103,
    n139,
    n235,
    n289
  );


  nor
  g485
  (
    n502,
    n263,
    n227,
    n194,
    n301
  );


  xor
  g486
  (
    n533,
    n102,
    n246,
    n137,
    n295
  );


  and
  g487
  (
    KeyWire_0_14,
    n161,
    n80,
    n194,
    n237
  );


  and
  g488
  (
    n436,
    n229,
    n117,
    n134,
    n219
  );


  xnor
  g489
  (
    n463,
    n141,
    n77,
    n225,
    n236
  );


  and
  g490
  (
    n346,
    n107,
    n77,
    n238,
    n261
  );


  xor
  g491
  (
    n387,
    n204,
    n226,
    n80,
    n167
  );


  xnor
  g492
  (
    n332,
    n226,
    n201,
    n149,
    n177
  );


  and
  g493
  (
    n424,
    n244,
    n210,
    n271,
    n104
  );


  or
  g494
  (
    n408,
    n124,
    n134,
    n254,
    n251
  );


  xnor
  g495
  (
    n367,
    n131,
    n110,
    n165,
    n121
  );


  nor
  g496
  (
    n378,
    n277,
    n253,
    n241,
    n203
  );


  nand
  g497
  (
    n461,
    n101,
    n293,
    n196,
    n124
  );


  nand
  g498
  (
    n426,
    n185,
    n232,
    n240,
    n167
  );


  or
  g499
  (
    n407,
    n215,
    n274,
    n297,
    n173
  );


  or
  g500
  (
    n397,
    n252,
    n194,
    n212,
    n216
  );


  nor
  g501
  (
    n386,
    n262,
    n119,
    n132,
    n117
  );


  nor
  g502
  (
    n477,
    n264,
    n150,
    n174,
    n180
  );


  xnor
  g503
  (
    n375,
    n217,
    n286,
    n161,
    n180
  );


  xor
  g504
  (
    n345,
    n287,
    n171,
    n288,
    n193
  );


  xor
  g505
  (
    n321,
    n138,
    n227,
    n79,
    n275
  );


  xnor
  g506
  (
    n394,
    n145,
    n294,
    n282,
    n265
  );


  or
  g507
  (
    n498,
    n213,
    n295,
    n139,
    n283
  );


  xor
  g508
  (
    n547,
    n128,
    n175,
    n195,
    n299
  );


  xnor
  g509
  (
    n395,
    n184,
    n231,
    n112,
    n189
  );


  and
  g510
  (
    n366,
    n234,
    n141,
    n108,
    n291
  );


  or
  g511
  (
    n483,
    n76,
    n142,
    n159,
    n265
  );


  xnor
  g512
  (
    n357,
    n242,
    n84,
    n236,
    n285
  );


  and
  g513
  (
    n337,
    n259,
    n273,
    n295,
    n169
  );


  and
  g514
  (
    n411,
    n101,
    n220,
    n162,
    n292
  );


  nand
  g515
  (
    n399,
    n294,
    n127,
    n202,
    n146
  );


  xnor
  g516
  (
    n538,
    n113,
    n148,
    n275,
    n246
  );


  or
  g517
  (
    n404,
    n109,
    n269,
    n192,
    n187
  );


  xor
  g518
  (
    n417,
    n146,
    n285,
    n291,
    n279
  );


  nor
  g519
  (
    n469,
    n193,
    n191,
    n281,
    n112
  );


  xnor
  g520
  (
    n402,
    n159,
    n150,
    n260,
    n276
  );


  or
  g521
  (
    n412,
    n281,
    n129,
    n283,
    n291
  );


  and
  g522
  (
    n421,
    n245,
    n180,
    n274,
    n300
  );


  and
  g523
  (
    n354,
    n135,
    n148,
    n285,
    n129
  );


  nand
  g524
  (
    n524,
    n147,
    n189,
    n168,
    n120
  );


  xor
  g525
  (
    n393,
    n158,
    n82,
    n282,
    n258
  );


  and
  g526
  (
    n328,
    n83,
    n217,
    n123,
    n143
  );


  not
  g527
  (
    n645,
    n452
  );


  not
  g528
  (
    n611,
    n324
  );


  buf
  g529
  (
    n663,
    n416
  );


  buf
  g530
  (
    n629,
    n448
  );


  buf
  g531
  (
    n615,
    n439
  );


  buf
  g532
  (
    n674,
    n359
  );


  not
  g533
  (
    n596,
    n380
  );


  buf
  g534
  (
    n631,
    n85
  );


  buf
  g535
  (
    n719,
    n388
  );


  not
  g536
  (
    n591,
    n417
  );


  not
  g537
  (
    n580,
    n455
  );


  buf
  g538
  (
    n609,
    n481
  );


  buf
  g539
  (
    n599,
    n94
  );


  buf
  g540
  (
    n640,
    n85
  );


  buf
  g541
  (
    n664,
    n415
  );


  buf
  g542
  (
    n604,
    n100
  );


  buf
  g543
  (
    n630,
    n428
  );


  buf
  g544
  (
    n634,
    n311
  );


  not
  g545
  (
    n561,
    n394
  );


  buf
  g546
  (
    n633,
    n312
  );


  buf
  g547
  (
    n650,
    n98
  );


  not
  g548
  (
    n704,
    n446
  );


  not
  g549
  (
    n742,
    n440
  );


  buf
  g550
  (
    n660,
    n427
  );


  not
  g551
  (
    n684,
    n97
  );


  not
  g552
  (
    n657,
    n382
  );


  not
  g553
  (
    n573,
    n87
  );


  buf
  g554
  (
    n667,
    n511
  );


  buf
  g555
  (
    n593,
    n411
  );


  not
  g556
  (
    n701,
    n392
  );


  not
  g557
  (
    n605,
    n85
  );


  buf
  g558
  (
    n679,
    n307
  );


  buf
  g559
  (
    n705,
    n406
  );


  not
  g560
  (
    n707,
    n404
  );


  buf
  g561
  (
    n736,
    n459
  );


  not
  g562
  (
    n597,
    n316
  );


  not
  g563
  (
    n565,
    n508
  );


  not
  g564
  (
    n623,
    n438
  );


  not
  g565
  (
    n571,
    n515
  );


  buf
  g566
  (
    n672,
    n342
  );


  not
  g567
  (
    n733,
    n376
  );


  buf
  g568
  (
    n618,
    n349
  );


  not
  g569
  (
    n551,
    n365
  );


  buf
  g570
  (
    n602,
    n89
  );


  buf
  g571
  (
    n643,
    n357
  );


  buf
  g572
  (
    n635,
    n305
  );


  buf
  g573
  (
    n713,
    n310
  );


  buf
  g574
  (
    n612,
    n89
  );


  buf
  g575
  (
    n708,
    n477
  );


  not
  g576
  (
    n566,
    n328
  );


  not
  g577
  (
    n686,
    n435
  );


  not
  g578
  (
    n590,
    n307
  );


  not
  g579
  (
    KeyWire_0_5,
    n378
  );


  buf
  g580
  (
    n671,
    n410
  );


  buf
  g581
  (
    n681,
    n308
  );


  not
  g582
  (
    n562,
    n93
  );


  buf
  g583
  (
    n740,
    n315
  );


  buf
  g584
  (
    n584,
    n311
  );


  buf
  g585
  (
    n606,
    n432
  );


  not
  g586
  (
    n550,
    n479
  );


  not
  g587
  (
    n711,
    n387
  );


  not
  g588
  (
    n730,
    n316
  );


  buf
  g589
  (
    n668,
    n311
  );


  not
  g590
  (
    n720,
    n494
  );


  not
  g591
  (
    n636,
    n419
  );


  not
  g592
  (
    n601,
    n96
  );


  buf
  g593
  (
    n626,
    n495
  );


  not
  g594
  (
    n610,
    n91
  );


  not
  g595
  (
    n552,
    n513
  );


  not
  g596
  (
    n715,
    n100
  );


  not
  g597
  (
    n678,
    n466
  );


  not
  g598
  (
    n653,
    n306
  );


  buf
  g599
  (
    n581,
    n84
  );


  buf
  g600
  (
    n718,
    n492
  );


  not
  g601
  (
    n728,
    n85
  );


  not
  g602
  (
    n559,
    n97
  );


  buf
  g603
  (
    n556,
    n354
  );


  buf
  g604
  (
    n680,
    n443
  );


  not
  g605
  (
    n613,
    n506
  );


  buf
  g606
  (
    n706,
    n409
  );


  buf
  g607
  (
    n638,
    n457
  );


  buf
  g608
  (
    n557,
    n95
  );


  buf
  g609
  (
    n568,
    n503
  );


  buf
  g610
  (
    n688,
    n92
  );


  not
  g611
  (
    n710,
    n336
  );


  not
  g612
  (
    n691,
    n96
  );


  buf
  g613
  (
    n689,
    n97
  );


  buf
  g614
  (
    n716,
    n423
  );


  not
  g615
  (
    n553,
    n491
  );


  not
  g616
  (
    n614,
    n488
  );


  not
  g617
  (
    n641,
    n489
  );


  buf
  g618
  (
    n739,
    n86
  );


  not
  g619
  (
    n594,
    n414
  );


  buf
  g620
  (
    n735,
    n306
  );


  buf
  g621
  (
    n575,
    n451
  );


  not
  g622
  (
    n700,
    n335
  );


  not
  g623
  (
    n703,
    n312
  );


  not
  g624
  (
    n697,
    n326
  );


  not
  g625
  (
    n627,
    n313
  );


  not
  g626
  (
    n589,
    n308
  );


  buf
  g627
  (
    n558,
    n361
  );


  buf
  g628
  (
    n620,
    n304
  );


  not
  g629
  (
    n669,
    n444
  );


  buf
  g630
  (
    n628,
    n313
  );


  buf
  g631
  (
    n579,
    n442
  );


  buf
  g632
  (
    n665,
    n486
  );


  not
  g633
  (
    n651,
    n436
  );


  buf
  g634
  (
    n659,
    n454
  );


  buf
  g635
  (
    n731,
    n310
  );


  not
  g636
  (
    n675,
    n314
  );


  not
  g637
  (
    n570,
    n373
  );


  buf
  g638
  (
    n685,
    n329
  );


  buf
  g639
  (
    n572,
    n305
  );


  not
  g640
  (
    n548,
    n356
  );


  buf
  g641
  (
    n624,
    n458
  );


  not
  g642
  (
    n616,
    n421
  );


  buf
  g643
  (
    n673,
    n424
  );


  buf
  g644
  (
    n648,
    n86
  );


  not
  g645
  (
    n586,
    n316
  );


  not
  g646
  (
    n587,
    n429
  );


  not
  g647
  (
    n646,
    n325
  );


  buf
  g648
  (
    n682,
    n447
  );


  not
  g649
  (
    n617,
    n497
  );


  not
  g650
  (
    n658,
    n343
  );


  not
  g651
  (
    n555,
    n398
  );


  not
  g652
  (
    n621,
    n306
  );


  buf
  g653
  (
    n694,
    n433
  );


  buf
  g654
  (
    n737,
    n500
  );


  buf
  g655
  (
    n569,
    n100
  );


  buf
  g656
  (
    n738,
    n482
  );


  buf
  g657
  (
    n709,
    n456
  );


  not
  g658
  (
    n662,
    n305
  );


  not
  g659
  (
    n560,
    n352
  );


  not
  g660
  (
    n693,
    n98
  );


  buf
  g661
  (
    n725,
    n445
  );


  buf
  g662
  (
    n639,
    n345
  );


  buf
  g663
  (
    n600,
    n304
  );


  buf
  g664
  (
    n717,
    n425
  );


  not
  g665
  (
    n702,
    n467
  );


  buf
  g666
  (
    n690,
    n314
  );


  not
  g667
  (
    n695,
    n91
  );


  not
  g668
  (
    n577,
    n93
  );


  buf
  g669
  (
    n696,
    n490
  );


  not
  g670
  (
    n724,
    n311
  );


  not
  g671
  (
    n727,
    n371
  );


  not
  g672
  (
    n699,
    n431
  );


  not
  g673
  (
    n632,
    n512
  );


  not
  g674
  (
    n692,
    n95
  );


  not
  g675
  (
    n676,
    n94
  );


  buf
  g676
  (
    n567,
    n363
  );


  buf
  g677
  (
    n582,
    n89
  );


  not
  g678
  (
    n607,
    n99
  );


  buf
  g679
  (
    n712,
    n348
  );


  not
  g680
  (
    n656,
    n366
  );


  not
  g681
  (
    n732,
    n453
  );


  not
  g682
  (
    n649,
    n322
  );


  and
  g683
  (
    n588,
    n450,
    n313
  );


  xnor
  g684
  (
    n574,
    n333,
    n402,
    n370,
    n496
  );


  nand
  g685
  (
    n592,
    n405,
    n400,
    n386,
    n360
  );


  nand
  g686
  (
    n564,
    n99,
    n86,
    n468,
    n408
  );


  xor
  g687
  (
    n677,
    n501,
    n499,
    n312,
    n384
  );


  xor
  g688
  (
    n647,
    n341,
    n92,
    n337,
    n315
  );


  xnor
  g689
  (
    n734,
    n91,
    n87,
    n389,
    n434
  );


  nor
  g690
  (
    n603,
    n465,
    n310,
    n472,
    n93
  );


  or
  g691
  (
    n655,
    n351,
    n464,
    n347,
    n474
  );


  or
  g692
  (
    n563,
    n355,
    n304,
    n485,
    n407
  );


  xor
  g693
  (
    n578,
    n470,
    n375,
    n330,
    n381
  );


  or
  g694
  (
    n576,
    n92,
    n98,
    n484,
    n397
  );


  nand
  g695
  (
    n654,
    n88,
    n314,
    n476,
    n430
  );


  xnor
  g696
  (
    n585,
    n475,
    n95,
    n327,
    n372
  );


  and
  g697
  (
    n595,
    n514,
    n391,
    n364,
    n502
  );


  nand
  g698
  (
    n683,
    n305,
    n307,
    n96,
    n340
  );


  xnor
  g699
  (
    n554,
    n353,
    n88,
    n437,
    n498
  );


  xor
  g700
  (
    n625,
    n505,
    n480,
    n312,
    n393
  );


  xnor
  g701
  (
    n642,
    n493,
    n91,
    n509,
    n516
  );


  nor
  g702
  (
    n652,
    n99,
    n88,
    n403,
    n315
  );


  or
  g703
  (
    n743,
    n469,
    n358,
    n462,
    n308
  );


  xor
  g704
  (
    n661,
    n390,
    n441,
    n315,
    n420
  );


  nand
  g705
  (
    n666,
    n323,
    n321,
    n399,
    n395
  );


  nand
  g706
  (
    n687,
    n86,
    n473,
    n385,
    n309
  );


  xor
  g707
  (
    n729,
    n461,
    n426,
    n487,
    n344
  );


  xnor
  g708
  (
    n723,
    n379,
    n94,
    n84,
    n362
  );


  and
  g709
  (
    n549,
    n346,
    n368,
    n510,
    n307
  );


  nor
  g710
  (
    n637,
    n483,
    n309,
    n316,
    n313
  );


  nor
  g711
  (
    n622,
    n89,
    n90,
    n504,
    n93
  );


  nand
  g712
  (
    n698,
    n88,
    n87,
    n460,
    n422
  );


  xor
  g713
  (
    n714,
    n95,
    n90,
    n507,
    n367
  );


  xnor
  g714
  (
    n608,
    n369,
    n478,
    n308,
    n374
  );


  xnor
  g715
  (
    n726,
    n98,
    n304,
    n306,
    n413
  );


  and
  g716
  (
    n741,
    n92,
    n383,
    n309,
    n471
  );


  nand
  g717
  (
    n619,
    n96,
    n401,
    n314,
    n310
  );


  nand
  g718
  (
    n721,
    n90,
    n334,
    n331,
    n396
  );


  nor
  g719
  (
    n670,
    n94,
    n100,
    n97,
    n377
  );


  nand
  g720
  (
    n583,
    n412,
    n99,
    n87,
    n350
  );


  nand
  g721
  (
    n644,
    n418,
    n338,
    n309,
    n332
  );


  or
  g722
  (
    n722,
    n463,
    n90,
    n449,
    n339
  );


  or
  g723
  (
    n744,
    n548,
    n317
  );


  xnor
  g724
  (
    n746,
    n528,
    n523,
    n526,
    n517
  );


  or
  g725
  (
    n747,
    n518,
    n521,
    n524,
    n527
  );


  xnor
  g726
  (
    n745,
    n520,
    n744
  );


  xnor
  g727
  (
    n748,
    n744,
    n522,
    n519,
    n525
  );


  nor
  g728
  (
    n750,
    n572,
    n748,
    n747,
    n577
  );


  nor
  g729
  (
    n754,
    n550,
    n573,
    n563,
    n556
  );


  nor
  g730
  (
    n753,
    n746,
    n564,
    n748,
    n566
  );


  or
  g731
  (
    n758,
    n568,
    n561,
    n558,
    n578
  );


  nor
  g732
  (
    n752,
    n554,
    n557,
    n747,
    n574
  );


  nand
  g733
  (
    n756,
    n745,
    n551,
    n746,
    n553
  );


  or
  g734
  (
    n755,
    n549,
    n747,
    n565,
    n559
  );


  nand
  g735
  (
    n757,
    n560,
    n562,
    n555,
    n746
  );


  or
  g736
  (
    n751,
    n567,
    n552,
    n570,
    n748
  );


  xnor
  g737
  (
    n749,
    n575,
    n576,
    n571,
    n569
  );


  not
  g738
  (
    n782,
    n755
  );


  not
  g739
  (
    n768,
    n753
  );


  not
  g740
  (
    n776,
    n756
  );


  buf
  g741
  (
    n766,
    n754
  );


  buf
  g742
  (
    n770,
    n751
  );


  not
  g743
  (
    n771,
    n758
  );


  not
  g744
  (
    n777,
    n752
  );


  not
  g745
  (
    n772,
    n758
  );


  not
  g746
  (
    n778,
    n756
  );


  buf
  g747
  (
    n759,
    n755
  );


  not
  g748
  (
    n761,
    n749
  );


  buf
  g749
  (
    n781,
    n758
  );


  not
  g750
  (
    n783,
    n751
  );


  not
  g751
  (
    n767,
    n753
  );


  not
  g752
  (
    n775,
    n757
  );


  not
  g753
  (
    n780,
    n754
  );


  buf
  g754
  (
    n773,
    n754
  );


  not
  g755
  (
    n763,
    n752
  );


  not
  g756
  (
    n762,
    n756
  );


  not
  g757
  (
    n764,
    n750
  );


  buf
  g758
  (
    n769,
    n755
  );


  buf
  g759
  (
    n784,
    n753
  );


  not
  g760
  (
    KeyWire_0_15,
    n751
  );


  not
  g761
  (
    n760,
    n752
  );


  not
  g762
  (
    n779,
    n757
  );


  buf
  g763
  (
    n774,
    n757
  );


  buf
  g764
  (
    n812,
    n777
  );


  not
  g765
  (
    n824,
    n760
  );


  buf
  g766
  (
    n877,
    n768
  );


  not
  g767
  (
    n788,
    n781
  );


  buf
  g768
  (
    n855,
    n765
  );


  buf
  g769
  (
    n836,
    n778
  );


  buf
  g770
  (
    n800,
    n759
  );


  not
  g771
  (
    n882,
    n759
  );


  not
  g772
  (
    n846,
    n771
  );


  buf
  g773
  (
    n806,
    n782
  );


  not
  g774
  (
    n814,
    n762
  );


  not
  g775
  (
    n833,
    n774
  );


  not
  g776
  (
    n880,
    n769
  );


  not
  g777
  (
    n826,
    n780
  );


  buf
  g778
  (
    n818,
    n766
  );


  not
  g779
  (
    n799,
    n783
  );


  not
  g780
  (
    n866,
    n762
  );


  not
  g781
  (
    n858,
    n764
  );


  buf
  g782
  (
    n862,
    n775
  );


  buf
  g783
  (
    n870,
    n766
  );


  not
  g784
  (
    KeyWire_0_10,
    n768
  );


  not
  g785
  (
    n813,
    n774
  );


  not
  g786
  (
    n817,
    n776
  );


  buf
  g787
  (
    n840,
    n773
  );


  buf
  g788
  (
    n848,
    n781
  );


  not
  g789
  (
    n825,
    n781
  );


  buf
  g790
  (
    n881,
    n771
  );


  not
  g791
  (
    n793,
    n783
  );


  buf
  g792
  (
    n875,
    n781
  );


  not
  g793
  (
    n790,
    n780
  );


  not
  g794
  (
    n802,
    n772
  );


  not
  g795
  (
    n809,
    n766
  );


  buf
  g796
  (
    n831,
    n769
  );


  not
  g797
  (
    n786,
    n771
  );


  buf
  g798
  (
    n837,
    n771
  );


  buf
  g799
  (
    n865,
    n763
  );


  buf
  g800
  (
    n873,
    n770
  );


  not
  g801
  (
    n829,
    n768
  );


  buf
  g802
  (
    n798,
    n761
  );


  not
  g803
  (
    n816,
    n779
  );


  buf
  g804
  (
    n797,
    n783
  );


  not
  g805
  (
    n871,
    n775
  );


  buf
  g806
  (
    n839,
    n767
  );


  not
  g807
  (
    n808,
    n767
  );


  not
  g808
  (
    n860,
    n772
  );


  not
  g809
  (
    n803,
    n780
  );


  not
  g810
  (
    n787,
    n764
  );


  buf
  g811
  (
    n847,
    n780
  );


  not
  g812
  (
    n796,
    n772
  );


  not
  g813
  (
    n819,
    n778
  );


  buf
  g814
  (
    n820,
    n778
  );


  buf
  g815
  (
    n864,
    n763
  );


  not
  g816
  (
    n856,
    n770
  );


  not
  g817
  (
    n867,
    n773
  );


  buf
  g818
  (
    n854,
    n779
  );


  buf
  g819
  (
    n879,
    n759
  );


  buf
  g820
  (
    n876,
    n777
  );


  buf
  g821
  (
    n834,
    n773
  );


  buf
  g822
  (
    n841,
    n759
  );


  not
  g823
  (
    n807,
    n777
  );


  not
  g824
  (
    n811,
    n775
  );


  buf
  g825
  (
    n835,
    n776
  );


  buf
  g826
  (
    n853,
    n782
  );


  buf
  g827
  (
    n850,
    n762
  );


  buf
  g828
  (
    n838,
    n782
  );


  buf
  g829
  (
    n844,
    n768
  );


  buf
  g830
  (
    n789,
    n764
  );


  buf
  g831
  (
    n863,
    n777
  );


  buf
  g832
  (
    n851,
    n767
  );


  buf
  g833
  (
    n842,
    n762
  );


  not
  g834
  (
    n792,
    n763
  );


  buf
  g835
  (
    n795,
    n776
  );


  not
  g836
  (
    n815,
    n782
  );


  not
  g837
  (
    n843,
    n765
  );


  not
  g838
  (
    n801,
    n770
  );


  not
  g839
  (
    n883,
    n761
  );


  not
  g840
  (
    n852,
    n764
  );


  buf
  g841
  (
    n884,
    n769
  );


  not
  g842
  (
    n823,
    n766
  );


  not
  g843
  (
    n861,
    n776
  );


  buf
  g844
  (
    n878,
    n765
  );


  not
  g845
  (
    n805,
    n783
  );


  buf
  g846
  (
    n869,
    n779
  );


  not
  g847
  (
    n832,
    n765
  );


  not
  g848
  (
    n785,
    n775
  );


  buf
  g849
  (
    n859,
    n773
  );


  not
  g850
  (
    n794,
    n774
  );


  buf
  g851
  (
    n791,
    n760
  );


  buf
  g852
  (
    n821,
    n760
  );


  not
  g853
  (
    n845,
    n770
  );


  not
  g854
  (
    n810,
    n763
  );


  not
  g855
  (
    n822,
    n778
  );


  buf
  g856
  (
    n827,
    n772
  );


  not
  g857
  (
    n874,
    n769
  );


  buf
  g858
  (
    n868,
    n761
  );


  buf
  g859
  (
    n857,
    n779
  );


  not
  g860
  (
    n849,
    n760
  );


  not
  g861
  (
    n830,
    n767
  );


  buf
  g862
  (
    n872,
    n761
  );


  buf
  g863
  (
    n828,
    n774
  );


  buf
  g864
  (
    n913,
    n635
  );


  buf
  g865
  (
    n927,
    n733
  );


  not
  g866
  (
    n915,
    n851
  );


  buf
  g867
  (
    n1039,
    n864
  );


  buf
  g868
  (
    n1018,
    n861
  );


  buf
  g869
  (
    n1035,
    n809
  );


  buf
  g870
  (
    n1154,
    n820
  );


  buf
  g871
  (
    n980,
    n730
  );


  not
  g872
  (
    n1032,
    n821
  );


  not
  g873
  (
    n1082,
    n792
  );


  not
  g874
  (
    n1074,
    n863
  );


  not
  g875
  (
    n1093,
    n855
  );


  buf
  g876
  (
    KeyWire_0_2,
    n738
  );


  not
  g877
  (
    n1157,
    n801
  );


  not
  g878
  (
    n897,
    n809
  );


  buf
  g879
  (
    n1110,
    n664
  );


  not
  g880
  (
    n933,
    n811
  );


  buf
  g881
  (
    n1105,
    n698
  );


  not
  g882
  (
    n986,
    n863
  );


  not
  g883
  (
    n1048,
    n858
  );


  not
  g884
  (
    n941,
    n819
  );


  buf
  g885
  (
    n999,
    n737
  );


  buf
  g886
  (
    n968,
    n840
  );


  buf
  g887
  (
    n1175,
    n849
  );


  buf
  g888
  (
    n902,
    n827
  );


  buf
  g889
  (
    n1111,
    n677
  );


  not
  g890
  (
    n1191,
    n854
  );


  buf
  g891
  (
    n997,
    n815
  );


  buf
  g892
  (
    n1083,
    n692
  );


  buf
  g893
  (
    n960,
    n796
  );


  not
  g894
  (
    n992,
    n822
  );


  buf
  g895
  (
    n994,
    n690
  );


  buf
  g896
  (
    n905,
    n785
  );


  not
  g897
  (
    n910,
    n825
  );


  not
  g898
  (
    n1084,
    n856
  );


  buf
  g899
  (
    n936,
    n863
  );


  not
  g900
  (
    n985,
    n718
  );


  not
  g901
  (
    n1180,
    n803
  );


  buf
  g902
  (
    n956,
    n658
  );


  buf
  g903
  (
    n885,
    n843
  );


  not
  g904
  (
    n945,
    n688
  );


  not
  g905
  (
    n1041,
    n829
  );


  buf
  g906
  (
    n906,
    n597
  );


  not
  g907
  (
    n1079,
    n828
  );


  not
  g908
  (
    n1062,
    n611
  );


  buf
  g909
  (
    n1134,
    n828
  );


  not
  g910
  (
    n955,
    n691
  );


  buf
  g911
  (
    n1028,
    n599
  );


  buf
  g912
  (
    n1000,
    n835
  );


  not
  g913
  (
    n1203,
    n729
  );


  buf
  g914
  (
    n1137,
    n711
  );


  buf
  g915
  (
    n1046,
    n603
  );


  buf
  g916
  (
    n916,
    n847
  );


  buf
  g917
  (
    n1081,
    n824
  );


  not
  g918
  (
    n969,
    n813
  );


  not
  g919
  (
    n888,
    n634
  );


  buf
  g920
  (
    n1104,
    n721
  );


  not
  g921
  (
    n944,
    n801
  );


  not
  g922
  (
    n1050,
    n802
  );


  buf
  g923
  (
    n1068,
    n797
  );


  not
  g924
  (
    n1135,
    n742
  );


  buf
  g925
  (
    n967,
    n789
  );


  not
  g926
  (
    n1099,
    n829
  );


  not
  g927
  (
    n958,
    n795
  );


  not
  g928
  (
    n935,
    n815
  );


  buf
  g929
  (
    n1113,
    n840
  );


  not
  g930
  (
    n1179,
    n789
  );


  buf
  g931
  (
    n1070,
    n596
  );


  buf
  g932
  (
    n1063,
    n855
  );


  buf
  g933
  (
    n975,
    n709
  );


  not
  g934
  (
    n1114,
    n808
  );


  not
  g935
  (
    n1036,
    n706
  );


  buf
  g936
  (
    n1017,
    n838
  );


  buf
  g937
  (
    n1056,
    n666
  );


  buf
  g938
  (
    n1077,
    n612
  );


  not
  g939
  (
    n1078,
    n805
  );


  not
  g940
  (
    n1069,
    n717
  );


  not
  g941
  (
    n962,
    n799
  );


  not
  g942
  (
    n1166,
    n845
  );


  not
  g943
  (
    n922,
    n680
  );


  buf
  g944
  (
    n1176,
    n819
  );


  buf
  g945
  (
    n1181,
    n852
  );


  not
  g946
  (
    n921,
    n623
  );


  buf
  g947
  (
    n928,
    n843
  );


  not
  g948
  (
    n1119,
    n615
  );


  buf
  g949
  (
    n1043,
    n788
  );


  buf
  g950
  (
    n1075,
    n839
  );


  buf
  g951
  (
    n1015,
    n810
  );


  buf
  g952
  (
    n1193,
    n794
  );


  not
  g953
  (
    n891,
    n859
  );


  buf
  g954
  (
    n946,
    n839
  );


  not
  g955
  (
    n1141,
    n636
  );


  buf
  g956
  (
    n1100,
    n823
  );


  buf
  g957
  (
    n1138,
    n805
  );


  buf
  g958
  (
    n887,
    n860
  );


  not
  g959
  (
    n1040,
    n791
  );


  buf
  g960
  (
    n1072,
    n837
  );


  not
  g961
  (
    n1092,
    n847
  );


  buf
  g962
  (
    n965,
    n724
  );


  not
  g963
  (
    n886,
    n788
  );


  not
  g964
  (
    KeyWire_0_6,
    n581
  );


  not
  g965
  (
    n981,
    n857
  );


  buf
  g966
  (
    n1001,
    n786
  );


  not
  g967
  (
    n1156,
    n619
  );


  not
  g968
  (
    n1080,
    n719
  );


  buf
  g969
  (
    n1065,
    n826
  );


  buf
  g970
  (
    n924,
    n847
  );


  not
  g971
  (
    n943,
    n618
  );


  not
  g972
  (
    n996,
    n827
  );


  not
  g973
  (
    n1085,
    n841
  );


  buf
  g974
  (
    n1064,
    n837
  );


  not
  g975
  (
    n1186,
    n804
  );


  not
  g976
  (
    n959,
    n813
  );


  buf
  g977
  (
    n1169,
    n734
  );


  not
  g978
  (
    n972,
    n814
  );


  not
  g979
  (
    n1006,
    n731
  );


  not
  g980
  (
    n1044,
    n630
  );


  buf
  g981
  (
    n939,
    n732
  );


  not
  g982
  (
    n1031,
    n830
  );


  not
  g983
  (
    n1025,
    n687
  );


  not
  g984
  (
    n973,
    n696
  );


  buf
  g985
  (
    n953,
    n656
  );


  xnor
  g986
  (
    n1117,
    n796,
    n742
  );


  xor
  g987
  (
    n1132,
    n793,
    n836
  );


  or
  g988
  (
    n1027,
    n685,
    n644
  );


  nand
  g989
  (
    n1158,
    n854,
    n848
  );


  or
  g990
  (
    n1020,
    n791,
    n731
  );


  xor
  g991
  (
    n1182,
    n732,
    n849
  );


  nand
  g992
  (
    n1188,
    n591,
    n812
  );


  or
  g993
  (
    n1033,
    n674,
    n663
  );


  nor
  g994
  (
    n1047,
    n818,
    n785
  );


  xnor
  g995
  (
    n993,
    n735,
    n846
  );


  xnor
  g996
  (
    n966,
    n856,
    n815
  );


  nand
  g997
  (
    n1002,
    n741,
    n614
  );


  xnor
  g998
  (
    n923,
    n828,
    n833
  );


  xor
  g999
  (
    n952,
    n793,
    n800
  );


  nor
  g1000
  (
    n1071,
    n832,
    n824
  );


  nor
  g1001
  (
    n1194,
    n829,
    n700
  );


  xnor
  g1002
  (
    n1124,
    n835,
    n786
  );


  xor
  g1003
  (
    n909,
    n844,
    n831
  );


  and
  g1004
  (
    n1143,
    n795,
    n842
  );


  xnor
  g1005
  (
    n1202,
    n857,
    n836
  );


  xnor
  g1006
  (
    n1121,
    n832,
    n647
  );


  xor
  g1007
  (
    n964,
    n851,
    n651
  );


  or
  g1008
  (
    n1059,
    n739,
    n816
  );


  buf
  g1009
  (
    n1103,
    n787
  );


  xor
  g1010
  (
    n950,
    n843,
    n616
  );


  or
  g1011
  (
    n1171,
    n794,
    n733
  );


  nand
  g1012
  (
    n1115,
    n725,
    n852
  );


  and
  g1013
  (
    n977,
    n862,
    n683
  );


  and
  g1014
  (
    n1190,
    n586,
    n530
  );


  nor
  g1015
  (
    n934,
    n825,
    n788
  );


  nand
  g1016
  (
    n930,
    n791,
    n678
  );


  nand
  g1017
  (
    n988,
    n673,
    n822
  );


  nor
  g1018
  (
    n1004,
    n637,
    n830
  );


  nand
  g1019
  (
    n1096,
    n842,
    n811
  );


  nand
  g1020
  (
    n991,
    n810,
    n856
  );


  xnor
  g1021
  (
    n1162,
    n798,
    n844
  );


  nand
  g1022
  (
    n1153,
    n828,
    n845
  );


  and
  g1023
  (
    n948,
    n833,
    n799
  );


  xnor
  g1024
  (
    n1197,
    n794,
    n592
  );


  nand
  g1025
  (
    n1185,
    n854,
    n845
  );


  nor
  g1026
  (
    n1090,
    n857,
    n662
  );


  xnor
  g1027
  (
    n1026,
    n807,
    n801
  );


  xnor
  g1028
  (
    n1189,
    n583,
    n813
  );


  xnor
  g1029
  (
    n925,
    n860,
    n731
  );


  xor
  g1030
  (
    n1016,
    n858,
    n808
  );


  or
  g1031
  (
    n983,
    n531,
    n642
  );


  or
  g1032
  (
    n907,
    n851,
    n667
  );


  nand
  g1033
  (
    n1142,
    n855,
    n832
  );


  nor
  g1034
  (
    n1178,
    n864,
    n829
  );


  nor
  g1035
  (
    n1195,
    n805,
    n861
  );


  or
  g1036
  (
    n1184,
    n806,
    n802
  );


  xnor
  g1037
  (
    n1150,
    n860,
    n812
  );


  or
  g1038
  (
    n937,
    n584,
    n638
  );


  and
  g1039
  (
    n917,
    n736,
    n633
  );


  xnor
  g1040
  (
    n1010,
    n580,
    n827
  );


  nand
  g1041
  (
    n1003,
    n625,
    n804
  );


  nor
  g1042
  (
    n1055,
    n834,
    n846
  );


  nand
  g1043
  (
    n990,
    n679,
    n617
  );


  xnor
  g1044
  (
    n1107,
    n807,
    n852
  );


  and
  g1045
  (
    n1042,
    n601,
    n834
  );


  nor
  g1046
  (
    n1024,
    n854,
    n799
  );


  nor
  g1047
  (
    n1172,
    n851,
    n815
  );


  nand
  g1048
  (
    n1076,
    n837,
    n650
  );


  xnor
  g1049
  (
    n1147,
    n847,
    n813
  );


  or
  g1050
  (
    n1136,
    n787,
    n786
  );


  xor
  g1051
  (
    n1174,
    n801,
    n802
  );


  and
  g1052
  (
    n1089,
    n826,
    n831
  );


  nand
  g1053
  (
    n1061,
    n839,
    n669
  );


  xnor
  g1054
  (
    n1097,
    n697,
    n714
  );


  xor
  g1055
  (
    n1161,
    n846,
    n838
  );


  nand
  g1056
  (
    n898,
    n627,
    n814
  );


  xnor
  g1057
  (
    n1034,
    n823,
    n631
  );


  nand
  g1058
  (
    n987,
    n824,
    n806
  );


  nand
  g1059
  (
    n1022,
    n689,
    n792
  );


  nand
  g1060
  (
    n931,
    n864,
    n708
  );


  or
  g1061
  (
    n963,
    n817,
    n598
  );


  and
  g1062
  (
    n1102,
    n585,
    n661
  );


  and
  g1063
  (
    n1094,
    n742,
    n798
  );


  or
  g1064
  (
    n1123,
    n713,
    n808
  );


  and
  g1065
  (
    n1170,
    n837,
    n582
  );


  or
  g1066
  (
    n1200,
    n842,
    n701
  );


  nand
  g1067
  (
    n1122,
    n643,
    n622
  );


  xor
  g1068
  (
    n1101,
    n820,
    n646
  );


  nor
  g1069
  (
    n1149,
    n695,
    n785
  );


  nor
  g1070
  (
    n1155,
    n738,
    n741
  );


  xor
  g1071
  (
    n1152,
    n818,
    n607
  );


  and
  g1072
  (
    n1045,
    n826,
    n588
  );


  or
  g1073
  (
    n1037,
    n862,
    n818
  );


  xnor
  g1074
  (
    n1183,
    n848,
    n816
  );


  nand
  g1075
  (
    n1198,
    n860,
    n729
  );


  xnor
  g1076
  (
    n1066,
    n838,
    n859
  );


  nor
  g1077
  (
    n1125,
    n817,
    n814
  );


  and
  g1078
  (
    n961,
    n670,
    n608
  );


  xnor
  g1079
  (
    n912,
    n858,
    n831
  );


  and
  g1080
  (
    n1086,
    n807,
    n733
  );


  and
  g1081
  (
    KeyWire_0_13,
    n739,
    n628
  );


  or
  g1082
  (
    n1073,
    n735,
    n729
  );


  nor
  g1083
  (
    n1007,
    n800,
    n833
  );


  xnor
  g1084
  (
    n1173,
    n740,
    n676
  );


  xnor
  g1085
  (
    n1112,
    n848,
    n827
  );


  nand
  g1086
  (
    n1029,
    n693,
    n672
  );


  nor
  g1087
  (
    n976,
    n841,
    n853
  );


  and
  g1088
  (
    n1011,
    n817,
    n639
  );


  or
  g1089
  (
    n1019,
    n812,
    n853
  );


  xnor
  g1090
  (
    n1030,
    n791,
    n675
  );


  xnor
  g1091
  (
    n1098,
    n822,
    n816
  );


  nor
  g1092
  (
    n957,
    n727,
    n800
  );


  xnor
  g1093
  (
    n938,
    n853,
    n787
  );


  nand
  g1094
  (
    n949,
    n788,
    n738
  );


  nand
  g1095
  (
    n1140,
    n648,
    n823
  );


  nor
  g1096
  (
    n1005,
    n832,
    n654
  );


  xnor
  g1097
  (
    n1196,
    n862,
    n640
  );


  xor
  g1098
  (
    n893,
    n793,
    n657
  );


  and
  g1099
  (
    n932,
    n716,
    n850
  );


  nand
  g1100
  (
    n911,
    n792,
    n825
  );


  nand
  g1101
  (
    n995,
    n819,
    n807
  );


  xor
  g1102
  (
    n1187,
    n532,
    n736
  );


  and
  g1103
  (
    n1160,
    n850,
    n734
  );


  nor
  g1104
  (
    n998,
    n798,
    n800
  );


  and
  g1105
  (
    n1058,
    n715,
    n712
  );


  nor
  g1106
  (
    n942,
    n653,
    n681
  );


  xnor
  g1107
  (
    n894,
    n668,
    n789
  );


  nand
  g1108
  (
    n892,
    n795,
    n812
  );


  and
  g1109
  (
    n904,
    n684,
    n579
  );


  and
  g1110
  (
    n954,
    n795,
    n853
  );


  and
  g1111
  (
    n889,
    n810,
    n835
  );


  or
  g1112
  (
    n908,
    n797,
    n809
  );


  and
  g1113
  (
    n1106,
    n844,
    n621
  );


  and
  g1114
  (
    n1139,
    n734,
    n641
  );


  and
  g1115
  (
    n929,
    n590,
    n722
  );


  and
  g1116
  (
    n1116,
    n822,
    n741
  );


  xnor
  g1117
  (
    n1151,
    n613,
    n737
  );


  nor
  g1118
  (
    n974,
    n694,
    n740
  );


  or
  g1119
  (
    n1053,
    n834,
    n814
  );


  xor
  g1120
  (
    n895,
    n852,
    n833
  );


  xnor
  g1121
  (
    n984,
    n859,
    n726
  );


  xor
  g1122
  (
    n926,
    n816,
    n834
  );


  or
  g1123
  (
    n1051,
    n803,
    n849
  );


  nor
  g1124
  (
    n1057,
    n686,
    n863
  );


  and
  g1125
  (
    n918,
    n728,
    n624
  );


  nor
  g1126
  (
    n1087,
    n820,
    n841
  );


  xor
  g1127
  (
    n1126,
    n793,
    n804
  );


  xor
  g1128
  (
    n914,
    n823,
    n794
  );


  nand
  g1129
  (
    n1133,
    n705,
    n682
  );


  and
  g1130
  (
    n1008,
    n802,
    n790
  );


  or
  g1131
  (
    n1091,
    n626,
    n858
  );


  and
  g1132
  (
    n1128,
    n606,
    n737
  );


  or
  g1133
  (
    n951,
    n723,
    n595
  );


  and
  g1134
  (
    n896,
    n806,
    n820
  );


  buf
  g1135
  (
    n1067,
    n821
  );


  and
  g1136
  (
    n940,
    n826,
    n817
  );


  xnor
  g1137
  (
    n903,
    n649,
    n710
  );


  xor
  g1138
  (
    n1127,
    n609,
    n655
  );


  nand
  g1139
  (
    KeyWire_0_8,
    n805,
    n804
  );


  nor
  g1140
  (
    n1192,
    n605,
    n797
  );


  nand
  g1141
  (
    n890,
    n840,
    n660
  );


  and
  g1142
  (
    n1012,
    n819,
    n789
  );


  and
  g1143
  (
    n1130,
    n841,
    n671
  );


  nand
  g1144
  (
    n1120,
    n629,
    n849
  );


  nand
  g1145
  (
    n1146,
    n587,
    n856
  );


  nor
  g1146
  (
    n1088,
    n796,
    n809
  );


  nand
  g1147
  (
    n1199,
    n790,
    n620
  );


  nand
  g1148
  (
    n920,
    n529,
    n730
  );


  xor
  g1149
  (
    n1052,
    n740,
    n848
  );


  nor
  g1150
  (
    n1131,
    n836,
    n811
  );


  xnor
  g1151
  (
    n1049,
    n799,
    n846
  );


  xnor
  g1152
  (
    n1009,
    n600,
    n593
  );


  xor
  g1153
  (
    n1164,
    n702,
    n707
  );


  xor
  g1154
  (
    n978,
    n803,
    n659
  );


  xor
  g1155
  (
    n1168,
    n861,
    n843
  );


  nor
  g1156
  (
    n1013,
    n803,
    n821
  );


  or
  g1157
  (
    n1129,
    n861,
    n830
  );


  xnor
  g1158
  (
    n1054,
    n703,
    n792
  );


  or
  g1159
  (
    n1038,
    n844,
    n862
  );


  xor
  g1160
  (
    n1118,
    n796,
    n632
  );


  nor
  g1161
  (
    n1144,
    n604,
    n811
  );


  or
  g1162
  (
    n1148,
    n699,
    n840
  );


  nand
  g1163
  (
    n1167,
    n652,
    n735
  );


  nor
  g1164
  (
    n1165,
    n730,
    n835
  );


  xnor
  g1165
  (
    n1095,
    n786,
    n790
  );


  nand
  g1166
  (
    n900,
    n842,
    n857
  );


  nand
  g1167
  (
    n901,
    n830,
    n798
  );


  or
  g1168
  (
    n1109,
    n790,
    n797
  );


  or
  g1169
  (
    n1145,
    n855,
    n732
  );


  xnor
  g1170
  (
    n1021,
    n824,
    n836
  );


  and
  g1171
  (
    n1023,
    n859,
    n736
  );


  nand
  g1172
  (
    n1108,
    n825,
    n850
  );


  xor
  g1173
  (
    n979,
    n845,
    n831
  );


  nand
  g1174
  (
    n1159,
    n665,
    n594
  );


  xor
  g1175
  (
    n919,
    n704,
    n810
  );


  and
  g1176
  (
    n1060,
    n589,
    n602
  );


  nor
  g1177
  (
    n899,
    n808,
    n806
  );


  xnor
  g1178
  (
    n947,
    n818,
    n743
  );


  xor
  g1179
  (
    n989,
    n720,
    n839
  );


  xor
  g1180
  (
    n1201,
    n610,
    n838
  );


  or
  g1181
  (
    n982,
    n645,
    n850
  );


  nand
  g1182
  (
    n1163,
    n739,
    n785
  );


  or
  g1183
  (
    n1316,
    n892,
    n1005,
    n977,
    n1077
  );


  xnor
  g1184
  (
    n1450,
    n942,
    n1124,
    n939,
    n1095
  );


  and
  g1185
  (
    n1214,
    n1167,
    n986,
    n1054,
    n1156
  );


  and
  g1186
  (
    n1287,
    n1054,
    n1109,
    n960,
    n943
  );


  nor
  g1187
  (
    n1357,
    n1175,
    n1039,
    n985,
    n1144
  );


  and
  g1188
  (
    n1205,
    n978,
    n1145,
    n962,
    n1104
  );


  or
  g1189
  (
    n1431,
    n1018,
    n1017,
    n1047,
    n1118
  );


  xor
  g1190
  (
    n1406,
    n1162,
    n890,
    n1048,
    n894
  );


  nor
  g1191
  (
    n1266,
    n537,
    n1112,
    n1053
  );


  xnor
  g1192
  (
    n1427,
    n1114,
    n1086,
    n927,
    n971
  );


  and
  g1193
  (
    n1363,
    n1050,
    n1020,
    n866,
    n980
  );


  xnor
  g1194
  (
    n1428,
    n1016,
    n1076,
    n1156,
    n1055
  );


  or
  g1195
  (
    n1283,
    n1037,
    n1188,
    n1104,
    n931
  );


  nand
  g1196
  (
    n1423,
    n995,
    n903,
    n1109,
    n1171
  );


  nand
  g1197
  (
    n1255,
    n1149,
    n1135,
    n1035,
    n1151
  );


  or
  g1198
  (
    n1442,
    n962,
    n1128,
    n1096,
    n1178
  );


  xnor
  g1199
  (
    n1319,
    n915,
    n937,
    n910,
    n1155
  );


  and
  g1200
  (
    n1347,
    n1119,
    n1144,
    n943,
    n941
  );


  nor
  g1201
  (
    n1365,
    n945,
    n989,
    n1142,
    n905
  );


  xor
  g1202
  (
    n1400,
    n971,
    n1140,
    n1089,
    n1057
  );


  and
  g1203
  (
    n1208,
    n1011,
    n1022,
    n1045,
    n1082
  );


  nor
  g1204
  (
    n1223,
    n1113,
    n1078,
    n905,
    n1014
  );


  xnor
  g1205
  (
    n1366,
    n1083,
    n951,
    n957,
    n1019
  );


  nand
  g1206
  (
    n1437,
    n1013,
    n1169,
    n546,
    n981
  );


  xnor
  g1207
  (
    n1349,
    n1115,
    n1027,
    n1106,
    n1075
  );


  nand
  g1208
  (
    n1443,
    n1150,
    n1033,
    n940,
    n1184
  );


  xnor
  g1209
  (
    n1305,
    n1170,
    n967,
    n968,
    n1021
  );


  and
  g1210
  (
    n1254,
    n949,
    n1142,
    n907,
    n1199
  );


  or
  g1211
  (
    n1271,
    n1068,
    n1065,
    n1060,
    n1159
  );


  nor
  g1212
  (
    KeyWire_0_7,
    n1100,
    n948,
    n1201,
    n1032
  );


  and
  g1213
  (
    n1438,
    n983,
    n1085,
    n998,
    n934
  );


  xnor
  g1214
  (
    n1394,
    n1009,
    n1121,
    n541,
    n1074
  );


  or
  g1215
  (
    n1293,
    n1111,
    n1193,
    n1058,
    n1047
  );


  nor
  g1216
  (
    n1215,
    n1182,
    n892,
    n961,
    n867
  );


  nor
  g1217
  (
    n1265,
    n1062,
    n1038,
    n1184,
    n1019
  );


  and
  g1218
  (
    n1294,
    n938,
    n916,
    n1130,
    n1021
  );


  xnor
  g1219
  (
    n1327,
    n1189,
    n973,
    n982,
    n909
  );


  nor
  g1220
  (
    n1419,
    n1080,
    n1138,
    n995,
    n1098
  );


  and
  g1221
  (
    n1219,
    n902,
    n975,
    n1050,
    n1087
  );


  nand
  g1222
  (
    n1310,
    n1160,
    n933,
    n1153,
    n978
  );


  xor
  g1223
  (
    n1247,
    n1071,
    n1147,
    n1183,
    n982
  );


  nand
  g1224
  (
    n1441,
    n1192,
    n1191,
    n960,
    n900
  );


  and
  g1225
  (
    n1226,
    n940,
    n1082,
    n1002,
    n1042
  );


  nor
  g1226
  (
    n1430,
    n1191,
    n1108,
    n926,
    n1060
  );


  nor
  g1227
  (
    n1352,
    n1070,
    n1196,
    n1129,
    n952
  );


  xor
  g1228
  (
    n1401,
    n1167,
    n923,
    n931,
    n1124
  );


  nor
  g1229
  (
    n1417,
    n1146,
    n913,
    n535,
    n944
  );


  xnor
  g1230
  (
    n1248,
    n1189,
    n1103,
    n898,
    n940
  );


  xor
  g1231
  (
    n1222,
    n908,
    n1193,
    n1034,
    n1042
  );


  nand
  g1232
  (
    n1342,
    n1093,
    n926,
    n865,
    n543
  );


  nor
  g1233
  (
    n1403,
    n961,
    n937,
    n1127,
    n902
  );


  xnor
  g1234
  (
    n1295,
    n904,
    n924,
    n1023,
    n1151
  );


  xnor
  g1235
  (
    n1416,
    n1049,
    n1083,
    n1097,
    n963
  );


  nor
  g1236
  (
    n1371,
    n886,
    n935,
    n534,
    n987
  );


  xor
  g1237
  (
    n1377,
    n1193,
    n1136,
    n953,
    n1012
  );


  xor
  g1238
  (
    n1360,
    n1164,
    n984,
    n1179,
    n1161
  );


  or
  g1239
  (
    n1367,
    n1016,
    n1186,
    n1015,
    n999
  );


  nand
  g1240
  (
    n1324,
    n1068,
    n1190,
    n895,
    n901
  );


  or
  g1241
  (
    n1429,
    n955,
    n1067,
    n1074,
    n1022
  );


  nor
  g1242
  (
    n1236,
    n1063,
    n1131,
    n885,
    n911
  );


  and
  g1243
  (
    n1315,
    n1176,
    n1073,
    n317,
    n1072
  );


  xor
  g1244
  (
    n1333,
    n1086,
    n1153,
    n1188,
    n1176
  );


  nand
  g1245
  (
    n1420,
    n987,
    n983,
    n999,
    n969
  );


  xnor
  g1246
  (
    n1243,
    n1198,
    n1004,
    n1056,
    n1188
  );


  xor
  g1247
  (
    n1321,
    n1199,
    n1196,
    n885,
    n784
  );


  and
  g1248
  (
    n1313,
    n890,
    n1113,
    n1081,
    n1173
  );


  and
  g1249
  (
    n1433,
    n960,
    n1158,
    n954,
    n1186
  );


  nor
  g1250
  (
    n1256,
    n1099,
    n536,
    n1125,
    n914
  );


  and
  g1251
  (
    n1372,
    n991,
    n1037,
    n1087,
    n958
  );


  nor
  g1252
  (
    n1232,
    n1084,
    n943,
    n1151,
    n1130
  );


  xor
  g1253
  (
    n1206,
    n533,
    n864,
    n900,
    n1041
  );


  nand
  g1254
  (
    n1239,
    n1121,
    n866,
    n976,
    n1001
  );


  nor
  g1255
  (
    n1241,
    n952,
    n1090,
    n917,
    n1034
  );


  nor
  g1256
  (
    n1339,
    n1036,
    n954,
    n1168,
    n1126
  );


  xnor
  g1257
  (
    n1369,
    n973,
    n903,
    n1180
  );


  and
  g1258
  (
    n1233,
    n1128,
    n1070,
    n1142,
    n1016
  );


  xor
  g1259
  (
    n1355,
    n1000,
    n1181,
    n1066,
    n994
  );


  nand
  g1260
  (
    n1252,
    n969,
    n969,
    n318,
    n1025
  );


  xnor
  g1261
  (
    n1302,
    n545,
    n1174,
    n980,
    n1073
  );


  or
  g1262
  (
    n1399,
    n986,
    n1103,
    n1185,
    n1097
  );


  and
  g1263
  (
    n1453,
    n893,
    n1113,
    n1169,
    n891
  );


  and
  g1264
  (
    n1273,
    n909,
    n950,
    n1127,
    n917
  );


  and
  g1265
  (
    n1303,
    n1030,
    n1080,
    n1126,
    n920
  );


  or
  g1266
  (
    n1370,
    n1198,
    n1035,
    n922,
    n1170
  );


  and
  g1267
  (
    n1413,
    n1105,
    n1131,
    n901,
    n978
  );


  or
  g1268
  (
    n1411,
    n1189,
    n1052,
    n1171,
    n1071
  );


  nor
  g1269
  (
    n1238,
    n991,
    n947,
    n1193,
    n938
  );


  xor
  g1270
  (
    n1314,
    n932,
    n938,
    n892,
    n318
  );


  nor
  g1271
  (
    n1362,
    n1194,
    n1119,
    n1019,
    n1200
  );


  and
  g1272
  (
    n1277,
    n1154,
    n934,
    n1096,
    n1145
  );


  nand
  g1273
  (
    n1359,
    n1079,
    n996,
    n930,
    n894
  );


  and
  g1274
  (
    n1312,
    n975,
    n975,
    n1143,
    n1089
  );


  xnor
  g1275
  (
    n1436,
    n993,
    n318,
    n1160,
    n867
  );


  nor
  g1276
  (
    n1358,
    n539,
    n977,
    n1165,
    n1136
  );


  nand
  g1277
  (
    n1336,
    n921,
    n1005,
    n1043,
    n895
  );


  nor
  g1278
  (
    n1398,
    n1107,
    n1036,
    n1202,
    n909
  );


  xnor
  g1279
  (
    n1282,
    n979,
    n946,
    n1057,
    n1163
  );


  xnor
  g1280
  (
    n1424,
    n1200,
    n951,
    n1175,
    n1187
  );


  xnor
  g1281
  (
    n1404,
    n1067,
    n1134,
    n1052,
    n961
  );


  xor
  g1282
  (
    n1261,
    n1164,
    n930,
    n956,
    n925
  );


  xor
  g1283
  (
    n1383,
    n1069,
    n915,
    n1163,
    n1143
  );


  xnor
  g1284
  (
    n1304,
    n948,
    n1011,
    n1010,
    n1040
  );


  xor
  g1285
  (
    n1422,
    n1044,
    n1075,
    n1099,
    n956
  );


  nand
  g1286
  (
    n1325,
    n1111,
    n1095,
    n1088,
    n1002
  );


  nor
  g1287
  (
    n1229,
    n988,
    n886,
    n1140,
    n1121
  );


  nor
  g1288
  (
    n1446,
    n979,
    n985,
    n993,
    n1078
  );


  xor
  g1289
  (
    n1439,
    n1083,
    n950,
    n1060,
    n999
  );


  or
  g1290
  (
    n1393,
    n867,
    n1129,
    n1017,
    n939
  );


  xor
  g1291
  (
    n1328,
    n1015,
    n887,
    n1065,
    n968
  );


  or
  g1292
  (
    n1410,
    n972,
    n1026,
    n1154,
    n1007
  );


  nor
  g1293
  (
    n1402,
    n1041,
    n922,
    n933,
    n1061
  );


  xnor
  g1294
  (
    n1204,
    n544,
    n1030,
    n1129,
    n1058
  );


  or
  g1295
  (
    n1418,
    n913,
    n926,
    n988,
    n1156
  );


  xor
  g1296
  (
    n1386,
    n1102,
    n1197,
    n1020,
    n317
  );


  or
  g1297
  (
    n1257,
    n1175,
    n1183,
    n963,
    n981
  );


  xor
  g1298
  (
    n1290,
    n1130,
    n1029,
    n970,
    n889
  );


  xnor
  g1299
  (
    n1220,
    n887,
    n1051,
    n1150,
    n1161
  );


  xnor
  g1300
  (
    n1384,
    n1085,
    n1177,
    n1123,
    n1153
  );


  nor
  g1301
  (
    n1381,
    n1123,
    n1147,
    n918,
    n1199
  );


  or
  g1302
  (
    n1311,
    n1073,
    n990,
    n1046
  );


  nand
  g1303
  (
    n1298,
    n910,
    n1079,
    n1088
  );


  nor
  g1304
  (
    n1249,
    n965,
    n936,
    n1008,
    n984
  );


  xnor
  g1305
  (
    n1269,
    n1122,
    n1014,
    n1006,
    n1103
  );


  nor
  g1306
  (
    n1289,
    n1149,
    n1051,
    n928,
    n1057
  );


  xnor
  g1307
  (
    n1322,
    n985,
    n1003,
    n1123,
    n1132
  );


  nor
  g1308
  (
    n1234,
    n1139,
    n910,
    n1064,
    n1116
  );


  nor
  g1309
  (
    n1380,
    n1023,
    n1100,
    n924,
    n1091
  );


  nand
  g1310
  (
    n1262,
    n984,
    n917,
    n923,
    n929
  );


  xor
  g1311
  (
    n1331,
    n1004,
    n1035,
    n784,
    n1032
  );


  or
  g1312
  (
    n1391,
    n904,
    n1111,
    n1183,
    n1046
  );


  and
  g1313
  (
    n1407,
    n1114,
    n1061,
    n1069,
    n1009
  );


  xor
  g1314
  (
    n1280,
    n1195,
    n970,
    n866,
    n1106
  );


  nand
  g1315
  (
    n1267,
    n991,
    n1098,
    n1169,
    n1199
  );


  nand
  g1316
  (
    n1337,
    n994,
    n1145,
    n1104,
    n1001
  );


  xor
  g1317
  (
    n1409,
    n1181,
    n1105,
    n896,
    n1085
  );


  or
  g1318
  (
    n1452,
    n921,
    n930,
    n1010,
    n1006
  );


  nor
  g1319
  (
    n1382,
    n1038,
    n1100,
    n1012,
    n1196
  );


  xnor
  g1320
  (
    n1346,
    n1157,
    n911,
    n1171,
    n1091
  );


  xor
  g1321
  (
    n1445,
    n992,
    n867,
    n997,
    n1013
  );


  or
  g1322
  (
    n1387,
    n895,
    n1118,
    n1036,
    n1165
  );


  nand
  g1323
  (
    n1350,
    n888,
    n1058,
    n1042,
    n986
  );


  and
  g1324
  (
    n1218,
    n929,
    n866,
    n1056,
    n1168
  );


  and
  g1325
  (
    n1224,
    n914,
    n1115,
    n939,
    n865
  );


  xor
  g1326
  (
    n1318,
    n1184,
    n1030,
    n966,
    n1094
  );


  nand
  g1327
  (
    n1434,
    n1051,
    n1059,
    n1007,
    n941
  );


  xnor
  g1328
  (
    n1211,
    n1192,
    n1026,
    n888,
    n1055
  );


  nor
  g1329
  (
    n1270,
    n1063,
    n1032,
    n1052,
    n907
  );


  nand
  g1330
  (
    n1213,
    n1024,
    n996,
    n1077,
    n989
  );


  nand
  g1331
  (
    n1374,
    n1062,
    n913,
    n1102,
    n1201
  );


  nand
  g1332
  (
    n1291,
    n1141,
    n1003,
    n1028,
    n967
  );


  xnor
  g1333
  (
    n1345,
    n919,
    n1202,
    n992,
    n1172
  );


  nand
  g1334
  (
    n1397,
    n1096,
    n1004,
    n988,
    n1141
  );


  xor
  g1335
  (
    n1415,
    n1161,
    n1068,
    n1080,
    n1143
  );


  or
  g1336
  (
    n1225,
    n911,
    n1010,
    n1037,
    n1093
  );


  nor
  g1337
  (
    n1242,
    n1196,
    n1078,
    n950,
    n1191
  );


  nor
  g1338
  (
    n1356,
    n959,
    n1163,
    n1162,
    n1170
  );


  xnor
  g1339
  (
    n1296,
    n891,
    n977,
    n1089,
    n1031
  );


  and
  g1340
  (
    n1454,
    n901,
    n1155,
    n889,
    n1131
  );


  xor
  g1341
  (
    n1405,
    n1133,
    n1065,
    n894,
    n1102
  );


  nor
  g1342
  (
    n1344,
    n896,
    n953,
    n885,
    n1202
  );


  xnor
  g1343
  (
    n1448,
    n1197,
    n1075,
    n1117,
    n1008
  );


  xnor
  g1344
  (
    n1260,
    n1134,
    n915,
    n1031,
    n932
  );


  nor
  g1345
  (
    n1447,
    n1061,
    n1027,
    n1007,
    n1048
  );


  nor
  g1346
  (
    n1329,
    n1108,
    n1072,
    n1200,
    n1110
  );


  or
  g1347
  (
    n1368,
    n1012,
    n1194,
    n1088,
    n1053
  );


  xor
  g1348
  (
    n1272,
    n1137,
    n865,
    n1027,
    n1015
  );


  and
  g1349
  (
    n1292,
    n1172,
    n1122,
    n1039,
    n920
  );


  and
  g1350
  (
    n1279,
    n966,
    n900,
    n972,
    n904
  );


  nand
  g1351
  (
    n1392,
    n1201,
    n1140,
    n1187,
    n944
  );


  and
  g1352
  (
    n1309,
    n1147,
    n1092,
    n1044,
    n1148
  );


  nand
  g1353
  (
    n1245,
    n908,
    n1045,
    n1198,
    n1025
  );


  or
  g1354
  (
    n1246,
    n931,
    n1077,
    n1041,
    n1101
  );


  nand
  g1355
  (
    n1408,
    n1059,
    n1076,
    n918,
    n996
  );


  xor
  g1356
  (
    n1301,
    n1137,
    n997,
    n919,
    n1136
  );


  xor
  g1357
  (
    n1351,
    n891,
    n924,
    n1064,
    n932
  );


  xnor
  g1358
  (
    n1230,
    n1185,
    n1126,
    n1107,
    n1064
  );


  nand
  g1359
  (
    n1396,
    n1101,
    n887,
    n1168,
    n925
  );


  nand
  g1360
  (
    n1412,
    n1022,
    n1135,
    n914,
    n1190
  );


  and
  g1361
  (
    n1251,
    n946,
    n1092,
    n1086,
    n1028
  );


  nor
  g1362
  (
    n1212,
    n1141,
    n902,
    n1198,
    n927
  );


  xnor
  g1363
  (
    n1209,
    n890,
    n1014,
    n982,
    n1040
  );


  nor
  g1364
  (
    n1281,
    n1005,
    n962,
    n1062,
    n1092
  );


  xor
  g1365
  (
    n1231,
    n1197,
    n1047,
    n1195,
    n956
  );


  nor
  g1366
  (
    n1263,
    n987,
    n1098,
    n905,
    n912
  );


  nand
  g1367
  (
    n1285,
    n1187,
    n920,
    n1024,
    n1133
  );


  nand
  g1368
  (
    n1250,
    n1002,
    n1185,
    n1106,
    n1097
  );


  xor
  g1369
  (
    n1395,
    n1018,
    n1134,
    n1120,
    n1001
  );


  xnor
  g1370
  (
    n1300,
    n916,
    n1117,
    n1090,
    n983
  );


  or
  g1371
  (
    n1343,
    n997,
    n1178,
    n957,
    n897
  );


  xor
  g1372
  (
    n1237,
    n1152,
    n921,
    n865,
    n937
  );


  nand
  g1373
  (
    n1414,
    n1081,
    n995,
    n964,
    n1177
  );


  or
  g1374
  (
    n1216,
    n1173,
    n1031,
    n929,
    n1093
  );


  nand
  g1375
  (
    n1455,
    n1094,
    n1066,
    n540,
    n1013
  );


  xnor
  g1376
  (
    n1320,
    n970,
    n1190,
    n1197
  );


  xor
  g1377
  (
    n1354,
    n907,
    n1139,
    n1091,
    n1101
  );


  and
  g1378
  (
    n1364,
    n949,
    n1050,
    n992,
    n1081
  );


  xnor
  g1379
  (
    n1449,
    n893,
    n936,
    n966,
    n1155
  );


  and
  g1380
  (
    n1276,
    n974,
    n1046,
    n928
  );


  xnor
  g1381
  (
    n1335,
    n1072,
    n918,
    n954,
    n317
  );


  xor
  g1382
  (
    n1299,
    n919,
    n1148,
    n1011,
    n1152
  );


  and
  g1383
  (
    n1228,
    n906,
    n1162,
    n967,
    n965
  );


  nand
  g1384
  (
    n1244,
    n994,
    n973,
    n945,
    n972
  );


  or
  g1385
  (
    n1306,
    n1000,
    n319,
    n1180,
    n1165
  );


  or
  g1386
  (
    n1385,
    n1024,
    n922,
    n981,
    n1033
  );


  nor
  g1387
  (
    n1286,
    n1176,
    n1132,
    n1201,
    n955
  );


  and
  g1388
  (
    n1284,
    n993,
    n946,
    n949,
    n1115
  );


  or
  g1389
  (
    n1264,
    n1159,
    n1074,
    n1138,
    n1167
  );


  xnor
  g1390
  (
    n1390,
    n944,
    n989,
    n964,
    n953
  );


  nand
  g1391
  (
    n1258,
    n1084,
    n1090,
    n1038,
    n1116
  );


  xnor
  g1392
  (
    n1334,
    n898,
    n1095,
    n968,
    n1182
  );


  xnor
  g1393
  (
    n1361,
    n1125,
    n1116,
    n936,
    n979
  );


  nor
  g1394
  (
    n1210,
    n1044,
    n1008,
    n980,
    n1146
  );


  xor
  g1395
  (
    n1317,
    n897,
    n974,
    n941,
    n959
  );


  xnor
  g1396
  (
    n1217,
    n1181,
    n1023,
    n1118,
    n1040
  );


  or
  g1397
  (
    n1451,
    n1017,
    n942,
    n1187,
    n1067
  );


  nor
  g1398
  (
    n1432,
    n963,
    n1109,
    n1174,
    n1146
  );


  nor
  g1399
  (
    n1375,
    n898,
    n1133,
    n1076,
    n1082
  );


  xor
  g1400
  (
    n1221,
    n964,
    n1087,
    n1160,
    n976
  );


  and
  g1401
  (
    n1340,
    n1195,
    n1182,
    n923,
    n1071
  );


  xor
  g1402
  (
    n1373,
    n1158,
    n1020,
    n1192,
    n908
  );


  or
  g1403
  (
    n1235,
    n899,
    n1159,
    n1148,
    n1194
  );


  nand
  g1404
  (
    n1338,
    n1105,
    n1000,
    n1164,
    n1070
  );


  or
  g1405
  (
    n1288,
    n1189,
    n886,
    n1139,
    n1003
  );


  xor
  g1406
  (
    n1341,
    n925,
    n935,
    n906,
    n1026
  );


  xor
  g1407
  (
    n1268,
    n958,
    n1033,
    n1124,
    n998
  );


  or
  g1408
  (
    n1253,
    n1173,
    n916,
    n945,
    n1117
  );


  xnor
  g1409
  (
    n1227,
    n965,
    n542,
    n912,
    n1149
  );


  xor
  g1410
  (
    n1444,
    n976,
    n1120,
    n1192,
    n974
  );


  or
  g1411
  (
    n1421,
    n889,
    n1049,
    n1006,
    n1045
  );


  or
  g1412
  (
    n1207,
    n1158,
    n1157,
    n1112,
    n957
  );


  or
  g1413
  (
    n1297,
    n1180,
    n1157,
    n927,
    n899
  );


  and
  g1414
  (
    n1240,
    n1144,
    n998,
    n955,
    n933
  );


  nand
  g1415
  (
    n1308,
    n899,
    n1191,
    n1110,
    n896
  );


  and
  g1416
  (
    n1440,
    n959,
    n318,
    n1029,
    n1066
  );


  nor
  g1417
  (
    n1348,
    n1029,
    n784,
    n1055,
    n1054
  );


  nand
  g1418
  (
    n1326,
    n935,
    n1069,
    n1174,
    n538
  );


  nor
  g1419
  (
    KeyWire_0_12,
    n951,
    n1009,
    n1048,
    n1049
  );


  nand
  g1420
  (
    n1353,
    n1059,
    n1154,
    n1120,
    n1152
  );


  xor
  g1421
  (
    n1425,
    n1132,
    n1128,
    n1084,
    n1056
  );


  nor
  g1422
  (
    n1274,
    n897,
    n1018,
    n1122,
    n1135
  );


  or
  g1423
  (
    n1323,
    n1177,
    n1112,
    n1166,
    n1172
  );


  xnor
  g1424
  (
    n1376,
    n1099,
    n1179,
    n1021,
    n1119
  );


  xnor
  g1425
  (
    n1275,
    n971,
    n1188,
    n1138,
    n1043
  );


  or
  g1426
  (
    n1330,
    n1028,
    n947,
    n906,
    n1186
  );


  or
  g1427
  (
    n1435,
    n990,
    n952,
    n1166,
    n1127
  );


  and
  g1428
  (
    n1278,
    n942,
    n1195,
    n1107,
    n958
  );


  xnor
  g1429
  (
    n1388,
    n1108,
    n1166,
    n784,
    n1110
  );


  xnor
  g1430
  (
    n1379,
    n934,
    n1125,
    n1094,
    n1200
  );


  or
  g1431
  (
    n1307,
    n1043,
    n1178,
    n1194,
    n888
  );


  or
  g1432
  (
    n1378,
    n1025,
    n912,
    n1034,
    n1150
  );


  and
  g1433
  (
    n1259,
    n1039,
    n947,
    n1063,
    n893
  );


  and
  g1434
  (
    n1332,
    n948,
    n1114,
    n1137,
    n1179
  );


  and
  g1435
  (
    n1490,
    n874,
    n1333,
    n1252,
    n1389
  );


  or
  g1436
  (
    n1491,
    n1368,
    n1272,
    n1214,
    n1381
  );


  and
  g1437
  (
    n1506,
    n1255,
    n1344,
    n1445,
    n1356
  );


  nor
  g1438
  (
    n1468,
    n1406,
    n1265,
    n1401,
    n1335
  );


  and
  g1439
  (
    n1505,
    n1339,
    n879,
    n1232,
    n1338
  );


  nor
  g1440
  (
    n1525,
    n1247,
    n1436,
    n1443,
    n882
  );


  nor
  g1441
  (
    n1476,
    n870,
    n874,
    n1439,
    n1395
  );


  and
  g1442
  (
    n1530,
    n1270,
    n1345,
    n1405,
    n1329
  );


  nand
  g1443
  (
    n1519,
    n1256,
    n1334,
    n1298,
    n1316
  );


  and
  g1444
  (
    n1517,
    n1322,
    n1274,
    n1262,
    n1300
  );


  and
  g1445
  (
    n1469,
    n1371,
    n1303,
    n1390,
    n878
  );


  and
  g1446
  (
    n1477,
    n1435,
    n1281,
    n1350,
    n1205
  );


  xnor
  g1447
  (
    n1532,
    n1319,
    n1400,
    n883,
    n884
  );


  nor
  g1448
  (
    n1486,
    n1427,
    n1293,
    n884,
    n1432
  );


  nor
  g1449
  (
    KeyWire_0_3,
    n875,
    n1245,
    n1299,
    n1424
  );


  xnor
  g1450
  (
    n1484,
    n1292,
    n1328,
    n880,
    n1301
  );


  xor
  g1451
  (
    n1461,
    n1446,
    n1348,
    n1433,
    n1280
  );


  or
  g1452
  (
    n1531,
    n1275,
    n1239,
    n1407,
    n1285
  );


  or
  g1453
  (
    n1528,
    n1236,
    n877,
    n881,
    n872
  );


  xnor
  g1454
  (
    n1466,
    n1217,
    n872,
    n876,
    n1209
  );


  xnor
  g1455
  (
    n1485,
    n1307,
    n1417,
    n879,
    n1314
  );


  or
  g1456
  (
    n1503,
    n1414,
    n1398,
    n1244,
    n1373
  );


  nor
  g1457
  (
    n1533,
    n1277,
    n1206,
    n1404,
    n1393
  );


  or
  g1458
  (
    n1499,
    n1367,
    n1355,
    n1224,
    n870
  );


  nor
  g1459
  (
    n1480,
    n1421,
    n1331,
    n880,
    n883
  );


  xnor
  g1460
  (
    n1475,
    n1219,
    n1380,
    n1359,
    n1324
  );


  xor
  g1461
  (
    n1498,
    n873,
    n877,
    n1394,
    n1366
  );


  xor
  g1462
  (
    n1523,
    n1410,
    n1431,
    n1341,
    n1212
  );


  nor
  g1463
  (
    n1459,
    n1235,
    n1411,
    n881,
    n1408
  );


  nor
  g1464
  (
    n1464,
    n870,
    n1415,
    n1440,
    n1305
  );


  xor
  g1465
  (
    n1512,
    n1388,
    n871,
    n1309,
    n1254
  );


  and
  g1466
  (
    n1487,
    n868,
    n884,
    n1250,
    n883
  );


  xor
  g1467
  (
    n1467,
    n1267,
    n1430,
    n879,
    n1418
  );


  or
  g1468
  (
    n1500,
    n1297,
    n1276,
    n1361,
    n1286
  );


  nand
  g1469
  (
    n1479,
    n875,
    n873,
    n1241,
    n1231
  );


  xnor
  g1470
  (
    n1510,
    n1357,
    n1447,
    n1279,
    n878
  );


  or
  g1471
  (
    n1513,
    n1258,
    n1249,
    n877,
    n872
  );


  nand
  g1472
  (
    n1527,
    n1396,
    n1336,
    n1374,
    n1317
  );


  xor
  g1473
  (
    n1516,
    n872,
    n1240,
    n1383,
    n1321
  );


  and
  g1474
  (
    n1495,
    n1438,
    n1437,
    n1386,
    n873
  );


  and
  g1475
  (
    n1470,
    n874,
    n871,
    n877,
    n1378
  );


  and
  g1476
  (
    n1481,
    n1320,
    n1211,
    n1234,
    n882
  );


  or
  g1477
  (
    n1508,
    n1312,
    n1372,
    n1210,
    n1248
  );


  xor
  g1478
  (
    n1511,
    n1229,
    n1364,
    n1428,
    n1340
  );


  xnor
  g1479
  (
    n1493,
    n1327,
    n871,
    n1360,
    n868
  );


  or
  g1480
  (
    n1473,
    n1352,
    n869,
    n1422,
    n1294
  );


  nand
  g1481
  (
    n1465,
    n1330,
    n1419,
    n1441,
    n880
  );


  nand
  g1482
  (
    n1496,
    n1243,
    n1337,
    n1295,
    n1399
  );


  xnor
  g1483
  (
    n1524,
    n1376,
    n874,
    n1226,
    n1308
  );


  nand
  g1484
  (
    n1494,
    n1259,
    n1444,
    n1332,
    n1261
  );


  or
  g1485
  (
    n1501,
    n878,
    n1375,
    n1402,
    n1273
  );


  xor
  g1486
  (
    n1521,
    n1213,
    n1278,
    n1425,
    n880
  );


  or
  g1487
  (
    n1489,
    n1325,
    n1379,
    n1369,
    n869
  );


  xor
  g1488
  (
    n1460,
    n1343,
    n1288,
    n1271,
    n1310
  );


  xor
  g1489
  (
    n1483,
    n875,
    n1208,
    n1223,
    n1326
  );


  or
  g1490
  (
    n1514,
    n1423,
    n1429,
    n1260,
    n1304
  );


  and
  g1491
  (
    n1504,
    n1426,
    n1221,
    n1238,
    n1323
  );


  nor
  g1492
  (
    n1488,
    n1370,
    n881,
    n1387,
    n873
  );


  nand
  g1493
  (
    n1462,
    n884,
    n1349,
    n1403,
    n876
  );


  nand
  g1494
  (
    n1458,
    n1434,
    n870,
    n1230,
    n1358
  );


  and
  g1495
  (
    n1507,
    n1220,
    n881,
    n1242,
    n1266
  );


  nor
  g1496
  (
    n1522,
    n1420,
    n1233,
    n1346,
    n1204
  );


  xnor
  g1497
  (
    n1520,
    n1397,
    n1354,
    n1313,
    n1264
  );


  nor
  g1498
  (
    n1492,
    n883,
    n1385,
    n1215,
    n1382
  );


  or
  g1499
  (
    n1518,
    n1287,
    n1257,
    n1225,
    n1228
  );


  or
  g1500
  (
    n1526,
    n869,
    n1284,
    n876,
    n879
  );


  xnor
  g1501
  (
    n1478,
    n1353,
    n875,
    n1384,
    n1302
  );


  xor
  g1502
  (
    n1529,
    n1311,
    n1318,
    n1296,
    n1269
  );


  nand
  g1503
  (
    n1457,
    n1347,
    n1216,
    n1253,
    n871
  );


  nand
  g1504
  (
    n1509,
    n1291,
    n878,
    n882,
    n1282
  );


  or
  g1505
  (
    n1471,
    n1283,
    n1412,
    n1289,
    n1315
  );


  xnor
  g1506
  (
    n1456,
    n1207,
    n1237,
    n1218,
    n1351
  );


  xor
  g1507
  (
    n1474,
    n1413,
    n876,
    n882,
    n1391
  );


  nand
  g1508
  (
    n1482,
    n869,
    n1365,
    n1263,
    n1377
  );


  xnor
  g1509
  (
    n1472,
    n868,
    n1227,
    n1222,
    n1342
  );


  xnor
  g1510
  (
    n1502,
    n1246,
    n1290,
    n1363,
    n1268
  );


  xnor
  g1511
  (
    n1515,
    n1442,
    n1392,
    n1416,
    n1409
  );


  nand
  g1512
  (
    n1497,
    n1251,
    n868,
    n1306,
    n1362
  );


  xnor
  g1513
  (
    n1534,
    n1482,
    n1203
  );


  nand
  g1514
  (
    n1535,
    n1202,
    n1483,
    n1203
  );


  buf
  g1515
  (
    n1540,
    n1534
  );


  not
  g1516
  (
    n1538,
    n1451
  );


  xor
  g1517
  (
    n1536,
    n1449,
    n1535
  );


  or
  g1518
  (
    n1537,
    n1448,
    n1452
  );


  or
  g1519
  (
    n1539,
    n1535,
    n1450,
    n1534
  );


  or
  g1520
  (
    n1551,
    n320,
    n1514,
    n1493,
    n1521
  );


  xnor
  g1521
  (
    n1548,
    n1524,
    n1537,
    n1453,
    n1497
  );


  and
  g1522
  (
    n1556,
    n1496,
    n1502,
    n1494,
    n1539
  );


  xor
  g1523
  (
    n1547,
    n1501,
    n1510,
    n1512,
    n1499
  );


  and
  g1524
  (
    n1554,
    n1511,
    n1536,
    n1489
  );


  xor
  g1525
  (
    n1555,
    n1532,
    n1537,
    n1506
  );


  or
  g1526
  (
    n1553,
    n1538,
    n1495,
    n1523,
    n1519
  );


  nor
  g1527
  (
    n1552,
    n1503,
    n1539,
    n1540,
    n320
  );


  xnor
  g1528
  (
    n1559,
    n1486,
    n743,
    n1513,
    n1531
  );


  or
  g1529
  (
    n1558,
    n1539,
    n319,
    n320,
    n1538
  );


  nand
  g1530
  (
    n1549,
    n1536,
    n1518,
    n1508,
    n320
  );


  or
  g1531
  (
    n1560,
    n1498,
    n1526,
    n1500,
    n1540
  );


  or
  g1532
  (
    n1543,
    n1484,
    n1515,
    n1529,
    n743
  );


  or
  g1533
  (
    KeyWire_0_0,
    n1505,
    n319,
    n1485,
    n1522
  );


  nor
  g1534
  (
    n1546,
    n1540,
    n1487,
    n1538,
    n1539
  );


  xnor
  g1535
  (
    n1541,
    n1540,
    n1516,
    n1492,
    n1504
  );


  and
  g1536
  (
    n1545,
    n319,
    n1490,
    n1533,
    n1525
  );


  and
  g1537
  (
    n1544,
    n1517,
    n1520,
    n1536,
    n1537
  );


  nand
  g1538
  (
    n1550,
    n1538,
    n1507,
    n1530,
    n1527
  );


  xnor
  g1539
  (
    n1542,
    n1528,
    n1488,
    n1509,
    n1491
  );


  and
  g1540
  (
    n1564,
    n1546,
    n1548,
    n1558,
    n1554
  );


  nand
  g1541
  (
    n1563,
    n1541,
    n1557,
    n1556,
    n547
  );


  xor
  g1542
  (
    n1561,
    n1454,
    n1543,
    n1535,
    n1547
  );


  xnor
  g1543
  (
    n1566,
    n1559,
    n1455,
    n1545,
    n1549
  );


  xor
  g1544
  (
    n1562,
    n1552,
    n1555,
    n1553,
    n1544
  );


  and
  g1545
  (
    n1565,
    n1560,
    n1542,
    n1551,
    n1550
  );


  xnor
  KeyGate_0_0
  (
    n1557,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n59,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n970,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1463,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n455,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n598,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1177,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1426,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n971,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n141,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n804,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n410,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1389,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1014,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n380,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n765,
    KeyNOTWire_0_15
  );


endmodule

