// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1321_43_4 written by SynthGen on 2021/06/15 15:04:52
module Stat_1321_43_4( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46,
 n276, n274, n290, n291, n267, n289, n300, n265,
 n292, n249, n297, n250, n259, n264, n295, n252,
 n279, n287, n266, n261, n1042, n1188, n1193, n1196,
 n1189, n1191, n1186, n1194, n1187, n1195, n1220, n1251,
 n1237, n1235, n1244, n1333, n1335, n1337, n1336, n1334,
 n1366, n1367, n1365, n1364);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46;

output n276, n274, n290, n291, n267, n289, n300, n265,
 n292, n249, n297, n250, n259, n264, n295, n252,
 n279, n287, n266, n261, n1042, n1188, n1193, n1196,
 n1189, n1191, n1186, n1194, n1187, n1195, n1220, n1251,
 n1237, n1235, n1244, n1333, n1335, n1337, n1336, n1334,
 n1366, n1367, n1365, n1364;

wire n47, n48, n49, n50, n51, n52, n53, n54,
 n55, n56, n57, n58, n59, n60, n61, n62,
 n63, n64, n65, n66, n67, n68, n69, n70,
 n71, n72, n73, n74, n75, n76, n77, n78,
 n79, n80, n81, n82, n83, n84, n85, n86,
 n87, n88, n89, n90, n91, n92, n93, n94,
 n95, n96, n97, n98, n99, n100, n101, n102,
 n103, n104, n105, n106, n107, n108, n109, n110,
 n111, n112, n113, n114, n115, n116, n117, n118,
 n119, n120, n121, n122, n123, n124, n125, n126,
 n127, n128, n129, n130, n131, n132, n133, n134,
 n135, n136, n137, n138, n139, n140, n141, n142,
 n143, n144, n145, n146, n147, n148, n149, n150,
 n151, n152, n153, n154, n155, n156, n157, n158,
 n159, n160, n161, n162, n163, n164, n165, n166,
 n167, n168, n169, n170, n171, n172, n173, n174,
 n175, n176, n177, n178, n179, n180, n181, n182,
 n183, n184, n185, n186, n187, n188, n189, n190,
 n191, n192, n193, n194, n195, n196, n197, n198,
 n199, n200, n201, n202, n203, n204, n205, n206,
 n207, n208, n209, n210, n211, n212, n213, n214,
 n215, n216, n217, n218, n219, n220, n221, n222,
 n223, n224, n225, n226, n227, n228, n229, n230,
 n231, n232, n233, n234, n235, n236, n237, n238,
 n239, n240, n241, n242, n243, n244, n245, n246,
 n247, n248, n251, n253, n254, n255, n256, n257,
 n258, n260, n262, n263, n268, n269, n270, n271,
 n272, n273, n275, n277, n278, n280, n281, n282,
 n283, n284, n285, n286, n288, n293, n294, n296,
 n298, n299, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n487, n488, n489, n490,
 n491, n492, n493, n494, n495, n496, n497, n498,
 n499, n500, n501, n502, n503, n504, n505, n506,
 n507, n508, n509, n510, n511, n512, n513, n514,
 n515, n516, n517, n518, n519, n520, n521, n522,
 n523, n524, n525, n526, n527, n528, n529, n530,
 n531, n532, n533, n534, n535, n536, n537, n538,
 n539, n540, n541, n542, n543, n544, n545, n546,
 n547, n548, n549, n550, n551, n552, n553, n554,
 n555, n556, n557, n558, n559, n560, n561, n562,
 n563, n564, n565, n566, n567, n568, n569, n570,
 n571, n572, n573, n574, n575, n576, n577, n578,
 n579, n580, n581, n582, n583, n584, n585, n586,
 n587, n588, n589, n590, n591, n592, n593, n594,
 n595, n596, n597, n598, n599, n600, n601, n602,
 n603, n604, n605, n606, n607, n608, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n660, n661, n662, n663, n664, n665, n666,
 n667, n668, n669, n670, n671, n672, n673, n674,
 n675, n676, n677, n678, n679, n680, n681, n682,
 n683, n684, n685, n686, n687, n688, n689, n690,
 n691, n692, n693, n694, n695, n696, n697, n698,
 n699, n700, n701, n702, n703, n704, n705, n706,
 n707, n708, n709, n710, n711, n712, n713, n714,
 n715, n716, n717, n718, n719, n720, n721, n722,
 n723, n724, n725, n726, n727, n728, n729, n730,
 n731, n732, n733, n734, n735, n736, n737, n738,
 n739, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1043,
 n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
 n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
 n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
 n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
 n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
 n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
 n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
 n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
 n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
 n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
 n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
 n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
 n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
 n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
 n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
 n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
 n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
 n1180, n1181, n1182, n1183, n1184, n1185, n1190, n1192,
 n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
 n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
 n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1221,
 n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
 n1230, n1231, n1232, n1233, n1234, n1236, n1238, n1239,
 n1240, n1241, n1242, n1243, n1245, n1246, n1247, n1248,
 n1249, n1250, n1252, n1253, n1254, n1255, n1256, n1257,
 n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
 n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
 n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
 n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
 n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
 n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
 n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
 n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
 n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
 n1330, n1331, n1332, n1338, n1339, n1340, n1341, n1342,
 n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
 n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
 n1359, n1360, n1361, n1362, n1363;

not  g0 (n96, n4);
not  g1 (n51, n44);
not  g2 (n128, n45);
not  g3 (n163, n37);
buf  g4 (n196, n17);
buf  g5 (n75, n10);
buf  g6 (n145, n42);
not  g7 (n117, n42);
buf  g8 (n175, n39);
buf  g9 (n106, n14);
buf  g10 (n164, n12);
not  g11 (n72, n1);
buf  g12 (n202, n40);
not  g13 (n168, n30);
not  g14 (n205, n46);
buf  g15 (n148, n39);
buf  g16 (n182, n37);
not  g17 (n221, n26);
buf  g18 (n55, n44);
buf  g19 (n130, n41);
buf  g20 (n170, n4);
not  g21 (n50, n38);
buf  g22 (n185, n14);
buf  g23 (n198, n16);
not  g24 (n71, n8);
not  g25 (n153, n30);
not  g26 (n85, n7);
not  g27 (n216, n26);
not  g28 (n102, n43);
not  g29 (n53, n9);
buf  g30 (n220, n8);
not  g31 (n162, n32);
buf  g32 (n230, n5);
buf  g33 (n118, n29);
buf  g34 (n215, n31);
not  g35 (n144, n45);
buf  g36 (n94, n11);
not  g37 (n136, n27);
not  g38 (n60, n46);
buf  g39 (n113, n23);
buf  g40 (n222, n26);
not  g41 (n138, n27);
not  g42 (n83, n32);
not  g43 (n169, n21);
not  g44 (n171, n42);
not  g45 (n193, n18);
not  g46 (n149, n19);
not  g47 (n166, n37);
not  g48 (n223, n23);
not  g49 (n165, n24);
not  g50 (n57, n37);
buf  g51 (n156, n35);
not  g52 (n161, n6);
buf  g53 (n172, n41);
buf  g54 (n99, n40);
not  g55 (n188, n3);
not  g56 (n91, n12);
not  g57 (n115, n27);
buf  g58 (n181, n46);
buf  g59 (n135, n24);
buf  g60 (n108, n30);
buf  g61 (n86, n20);
buf  g62 (n200, n23);
not  g63 (n183, n29);
not  g64 (n167, n17);
buf  g65 (n180, n19);
not  g66 (n142, n22);
not  g67 (n189, n21);
buf  g68 (n137, n35);
not  g69 (n176, n25);
buf  g70 (n93, n35);
not  g71 (n174, n7);
buf  g72 (n81, n18);
not  g73 (n116, n3);
not  g74 (n125, n34);
buf  g75 (n203, n21);
not  g76 (n208, n29);
buf  g77 (n209, n24);
buf  g78 (n173, n9);
buf  g79 (n67, n28);
buf  g80 (n110, n31);
buf  g81 (n224, n34);
buf  g82 (n62, n5);
buf  g83 (n88, n18);
buf  g84 (n132, n38);
buf  g85 (n104, n40);
buf  g86 (n139, n11);
buf  g87 (n73, n13);
not  g88 (n140, n2);
buf  g89 (n141, n44);
buf  g90 (n84, n10);
not  g91 (n58, n6);
not  g92 (n47, n12);
not  g93 (n226, n19);
not  g94 (n54, n42);
not  g95 (n80, n40);
buf  g96 (n107, n31);
not  g97 (n147, n8);
buf  g98 (n127, n20);
buf  g99 (n112, n46);
buf  g100 (n61, n17);
not  g101 (n69, n16);
not  g102 (n56, n2);
buf  g103 (n160, n44);
buf  g104 (n66, n1);
buf  g105 (n214, n15);
not  g106 (n105, n16);
buf  g107 (n70, n6);
buf  g108 (n119, n33);
buf  g109 (n100, n3);
buf  g110 (n199, n10);
buf  g111 (n122, n33);
not  g112 (n228, n1);
not  g113 (n103, n28);
not  g114 (n129, n25);
buf  g115 (n92, n34);
not  g116 (n146, n36);
buf  g117 (n109, n29);
not  g118 (n89, n36);
not  g119 (n229, n25);
not  g120 (n178, n20);
not  g121 (n78, n43);
buf  g122 (n133, n15);
buf  g123 (n213, n26);
not  g124 (n225, n30);
not  g125 (n211, n2);
buf  g126 (n151, n36);
buf  g127 (n97, n7);
not  g128 (n48, n15);
buf  g129 (n217, n36);
not  g130 (n77, n14);
not  g131 (n159, n4);
buf  g132 (n64, n6);
buf  g133 (n194, n8);
not  g134 (n155, n28);
not  g135 (n204, n45);
not  g136 (n177, n15);
not  g137 (n131, n41);
not  g138 (n201, n14);
not  g139 (n187, n24);
not  g140 (n158, n11);
not  g141 (n120, n31);
buf  g142 (n68, n33);
buf  g143 (n49, n32);
not  g144 (n210, n13);
not  g145 (n192, n9);
buf  g146 (n90, n34);
not  g147 (n95, n43);
buf  g148 (n101, n43);
not  g149 (n65, n9);
not  g150 (n114, n5);
buf  g151 (n111, n38);
not  g152 (n79, n11);
buf  g153 (n154, n5);
buf  g154 (n212, n22);
buf  g155 (n206, n22);
not  g156 (n190, n18);
not  g157 (n150, n13);
buf  g158 (n82, n4);
buf  g159 (n124, n25);
buf  g160 (n121, n2);
not  g161 (n134, n39);
buf  g162 (n74, n39);
not  g163 (n143, n23);
not  g164 (n219, n3);
buf  g165 (n87, n35);
not  g166 (n52, n22);
not  g167 (n76, n32);
not  g168 (n227, n33);
buf  g169 (n126, n16);
not  g170 (n197, n19);
buf  g171 (n98, n12);
not  g172 (n63, n17);
not  g173 (n59, n10);
not  g174 (n184, n20);
buf  g175 (n218, n41);
not  g176 (n186, n13);
buf  g177 (n195, n27);
not  g178 (n179, n1);
not  g179 (n191, n21);
buf  g180 (n207, n28);
buf  g181 (n157, n45);
not  g182 (n152, n38);
buf  g183 (n123, n7);
buf  g184 (n231, n47);
buf  g185 (n232, n48);
not  g186 (n235, n47);
buf  g187 (n234, n47);
not  g188 (n233, n47);
buf  g189 (n247, n233);
not  g190 (n245, n234);
not  g191 (n236, n231);
not  g192 (n244, n233);
buf  g193 (n241, n232);
buf  g194 (n240, n231);
not  g195 (n237, n231);
not  g196 (n246, n233);
not  g197 (n238, n232);
buf  g198 (n243, n232);
buf  g199 (n242, n232);
not  g200 (n248, n231);
buf  g201 (n239, n233);
not  g202 (n282, n239);
not  g203 (n259, n243);
buf  g204 (n291, n243);
not  g205 (n273, n247);
buf  g206 (n289, n241);
buf  g207 (n286, n241);
not  g208 (n297, n238);
not  g209 (n298, n238);
not  g210 (n249, n244);
buf  g211 (n284, n248);
not  g212 (n283, n236);
buf  g213 (n299, n242);
buf  g214 (n280, n247);
not  g215 (n296, n238);
buf  g216 (n292, n245);
not  g217 (n266, n239);
not  g218 (n253, n244);
buf  g219 (n261, n241);
buf  g220 (n272, n242);
buf  g221 (n295, n240);
not  g222 (n290, n245);
buf  g223 (n264, n240);
not  g224 (n260, n246);
not  g225 (n285, n248);
not  g226 (n277, n246);
not  g227 (n274, n245);
buf  g228 (n256, n243);
buf  g229 (n255, n248);
buf  g230 (n252, n244);
buf  g231 (n294, n244);
not  g232 (n287, n248);
buf  g233 (n276, n236);
not  g234 (n263, n241);
buf  g235 (n258, n236);
not  g236 (n270, n240);
not  g237 (n271, n243);
buf  g238 (n293, n246);
buf  g239 (n267, n240);
not  g240 (n262, n237);
buf  g241 (n279, n247);
not  g242 (n257, n242);
buf  g243 (n251, n242);
buf  g244 (n281, n247);
buf  g245 (n268, n237);
buf  g246 (n250, n237);
not  g247 (n288, n236);
buf  g248 (n300, n238);
buf  g249 (n265, n237);
not  g250 (n269, n245);
not  g251 (n278, n239);
not  g252 (n254, n239);
buf  g253 (n275, n246);
not  g254 (n309, n278);
not  g255 (n310, n269);
not  g256 (n301, n272);
buf  g257 (n307, n273);
not  g258 (n304, n277);
not  g259 (n302, n271);
not  g260 (n305, n270);
not  g261 (n308, n274);
not  g262 (n303, n276);
buf  g263 (n306, n275);
xor  g264 (n322, n293, n49);
and  g265 (n314, n303, n294, n48);
nor  g266 (n321, n48, n300, n283);
xor  g267 (n323, n296, n49, n290);
xnor g268 (n316, n302, n49, n285);
or   g269 (n312, n289, n279, n287);
or   g270 (n311, n302, n299, n284);
and  g271 (n317, n282, n297, n295);
nor  g272 (n315, n303, n301);
xor  g273 (n319, n302, n280, n303);
nand g274 (n313, n304, n288, n291, n48);
nor  g275 (n320, n302, n298, n303, n301);
or   g276 (n318, n281, n292, n301, n286);
xor  g277 (n343, n60, n57, n70, n315);
nand g278 (n336, n51, n62, n54);
xnor g279 (n326, n50, n318, n72, n78);
xor  g280 (n331, n63, n59, n62, n60);
xnor g281 (n332, n67, n305, n78, n313);
and  g282 (n355, n67, n64, n322);
and  g283 (n333, n57, n54, n312, n313);
nand g284 (n368, n53, n75, n72, n77);
nor  g285 (n370, n59, n74, n60, n66);
nand g286 (n360, n307, n235, n52, n309);
xor  g287 (n329, n77, n307, n317, n76);
xor  g288 (n346, n310, n72, n57, n78);
or   g289 (n362, n305, n76, n316, n318);
nand g290 (n353, n59, n67, n51);
nand g291 (n325, n62, n58, n68, n63);
nor  g292 (n327, n69, n56, n314, n76);
and  g293 (n350, n70, n322, n323, n234);
or   g294 (n339, n71, n304, n58, n75);
xor  g295 (n330, n320, n53, n308, n312);
xor  g296 (n365, n313, n63, n75, n317);
xnor g297 (n352, n74, n55, n321, n312);
xnor g298 (n345, n309, n315, n57, n65);
xor  g299 (n371, n61, n52, n78, n323);
nand g300 (n366, n66, n319, n310, n308);
and  g301 (n328, n69, n64, n51, n71);
and  g302 (n364, n315, n319, n314, n321);
and  g303 (n324, n320, n311, n322, n323);
xnor g304 (n356, n61, n52, n313, n306);
xnor g305 (n348, n318, n318, n65, n70);
xnor g306 (n347, n50, n307, n56, n69);
and  g307 (n354, n320, n319, n234, n77);
and  g308 (n334, n52, n60, n56, n309);
and  g309 (n372, n51, n55, n74, n316);
and  g310 (n351, n319, n312, n68);
or   g311 (n359, n64, n235, n72, n317);
nor  g312 (n342, n314, n308, n73, n310);
and  g313 (n337, n55, n53, n320, n304);
or   g314 (n363, n304, n68, n311, n323);
nand g315 (n373, n59, n306, n307, n316);
xor  g316 (n367, n73, n305, n76, n235);
or   g317 (n361, n61, n314, n56, n58);
xor  g318 (n369, n58, n70, n71, n316);
xnor g319 (n344, n53, n50, n71, n321);
nand g320 (n357, n65, n73, n235, n62);
nand g321 (n349, n310, n50, n308, n306);
xnor g322 (n358, n66, n322, n69, n74);
nor  g323 (n340, n75, n317, n309, n73);
nor  g324 (n335, n61, n321, n315, n54);
and  g325 (n341, n305, n234, n65, n77);
nor  g326 (n338, n66, n63, n306, n55);
buf  g327 (n484, n326);
not  g328 (n483, n358);
not  g329 (n448, n328);
not  g330 (n381, n362);
buf  g331 (n415, n351);
not  g332 (n470, n367);
buf  g333 (n440, n349);
not  g334 (n431, n361);
not  g335 (n497, n342);
buf  g336 (n408, n344);
not  g337 (n416, n344);
not  g338 (n459, n343);
buf  g339 (n490, n338);
not  g340 (n442, n364);
buf  g341 (n522, n352);
not  g342 (n520, n372);
buf  g343 (n388, n366);
not  g344 (n404, n338);
not  g345 (n413, n359);
buf  g346 (n529, n348);
not  g347 (n461, n326);
buf  g348 (n449, n341);
buf  g349 (n420, n368);
buf  g350 (n469, n348);
buf  g351 (n389, n336);
buf  g352 (n504, n354);
not  g353 (n494, n372);
buf  g354 (n527, n372);
buf  g355 (n393, n341);
not  g356 (n441, n340);
not  g357 (n414, n345);
not  g358 (n391, n349);
not  g359 (n464, n364);
buf  g360 (n512, n358);
not  g361 (n386, n357);
not  g362 (n437, n369);
not  g363 (n462, n347);
not  g364 (n492, n347);
buf  g365 (n465, n360);
buf  g366 (n516, n364);
buf  g367 (n411, n351);
not  g368 (n400, n333);
buf  g369 (n427, n345);
buf  g370 (n392, n367);
not  g371 (n397, n350);
not  g372 (n433, n345);
not  g373 (n443, n370);
buf  g374 (n456, n357);
not  g375 (n394, n334);
not  g376 (n517, n357);
not  g377 (n488, n369);
not  g378 (n436, n337);
buf  g379 (n478, n325);
buf  g380 (n507, n343);
buf  g381 (n434, n356);
buf  g382 (n503, n365);
not  g383 (n403, n350);
buf  g384 (n514, n365);
not  g385 (n521, n352);
buf  g386 (n487, n355);
not  g387 (n515, n362);
buf  g388 (n406, n369);
not  g389 (n429, n330);
not  g390 (n455, n332);
buf  g391 (n509, n346);
buf  g392 (n482, n371);
buf  g393 (n380, n370);
buf  g394 (n498, n342);
buf  g395 (n382, n368);
not  g396 (n468, n340);
buf  g397 (n472, n364);
buf  g398 (n402, n352);
buf  g399 (n458, n331);
not  g400 (n405, n344);
not  g401 (n378, n332);
not  g402 (n438, n360);
buf  g403 (n501, n353);
not  g404 (n467, n333);
buf  g405 (n518, n338);
buf  g406 (n447, n370);
not  g407 (n474, n325);
buf  g408 (n486, n368);
buf  g409 (n396, n358);
buf  g410 (n432, n342);
not  g411 (n430, n367);
buf  g412 (n375, n346);
not  g413 (n511, n372);
buf  g414 (n399, n373);
buf  g415 (n452, n348);
buf  g416 (n505, n329);
buf  g417 (n460, n355);
not  g418 (n463, n365);
not  g419 (n519, n347);
not  g420 (n446, n355);
not  g421 (n419, n363);
not  g422 (n513, n335);
not  g423 (n489, n362);
buf  g424 (n435, n340);
buf  g425 (n476, n361);
not  g426 (n454, n353);
not  g427 (n473, n335);
buf  g428 (n525, n339);
buf  g429 (n374, n356);
not  g430 (n428, n353);
not  g431 (n477, n354);
buf  g432 (n526, n327);
buf  g433 (n423, n371);
not  g434 (n450, n339);
buf  g435 (n395, n370);
not  g436 (n409, n334);
buf  g437 (n412, n349);
buf  g438 (n376, n368);
buf  g439 (n496, n369);
buf  g440 (n422, n357);
not  g441 (n407, n359);
not  g442 (n510, n356);
not  g443 (n444, n352);
not  g444 (n418, n360);
not  g445 (n424, n361);
not  g446 (n421, n329);
buf  g447 (n499, n366);
buf  g448 (n453, n359);
not  g449 (n528, n363);
not  g450 (n425, n359);
not  g451 (n485, n343);
buf  g452 (n523, n331);
not  g453 (n377, n371);
not  g454 (n481, n330);
not  g455 (n385, n362);
buf  g456 (n475, n339);
not  g457 (n390, n337);
buf  g458 (n379, n328);
not  g459 (n493, n365);
buf  g460 (n508, n366);
buf  g461 (n383, n358);
buf  g462 (n417, n361);
not  g463 (n445, n327);
buf  g464 (n401, n373);
not  g465 (n480, n360);
buf  g466 (n384, n356);
buf  g467 (n451, n363);
not  g468 (n500, n336);
not  g469 (n398, n366);
not  g470 (n506, n346);
not  g471 (n502, n355);
buf  g472 (n457, n354);
buf  g473 (n495, n341);
buf  g474 (n387, n373);
not  g475 (n466, n350);
not  g476 (n410, n353);
buf  g477 (n524, n371);
not  g478 (n426, n354);
not  g479 (n479, n373);
not  g480 (n471, n367);
buf  g481 (n439, n351);
buf  g482 (n491, n363);
buf  g483 (n828, n430);
buf  g484 (n640, n415);
buf  g485 (n776, n379);
buf  g486 (n861, n119);
not  g487 (n561, n147);
not  g488 (n549, n171);
buf  g489 (n710, n505);
buf  g490 (n718, n483);
not  g491 (n675, n506);
buf  g492 (n665, n450);
buf  g493 (n684, n418);
buf  g494 (n730, n512);
not  g495 (n742, n139);
buf  g496 (n530, n414);
not  g497 (n754, n175);
not  g498 (n686, n380);
not  g499 (n743, n162);
buf  g500 (n799, n487);
not  g501 (n801, n185);
buf  g502 (n898, n96);
buf  g503 (n591, n184);
not  g504 (n751, n212);
buf  g505 (n723, n438);
not  g506 (n747, n94);
not  g507 (n794, n504);
buf  g508 (n638, n428);
buf  g509 (n866, n161);
buf  g510 (n726, n128);
buf  g511 (n775, n86);
not  g512 (n681, n175);
buf  g513 (n615, n500);
not  g514 (n873, n206);
not  g515 (n760, n118);
buf  g516 (n863, n437);
buf  g517 (n772, n412);
buf  g518 (n598, n135);
not  g519 (n660, n445);
buf  g520 (n902, n402);
buf  g521 (n541, n186);
not  g522 (n679, n151);
not  g523 (n582, n117);
not  g524 (n663, n138);
buf  g525 (n755, n478);
buf  g526 (n689, n188);
not  g527 (n781, n492);
buf  g528 (n609, n175);
buf  g529 (n651, n200);
not  g530 (n559, n512);
not  g531 (n596, n151);
buf  g532 (n672, n504);
not  g533 (n811, n472);
buf  g534 (n589, n211);
buf  g535 (n763, n492);
not  g536 (n741, n442);
buf  g537 (n789, n127);
not  g538 (n536, n518);
buf  g539 (n753, n400);
buf  g540 (n704, n182);
not  g541 (n578, n196);
buf  g542 (n719, n131);
buf  g543 (n778, n374);
not  g544 (n603, n404);
buf  g545 (n810, n475);
not  g546 (n709, n161);
buf  g547 (n610, n488);
not  g548 (n800, n420);
not  g549 (n588, n107);
buf  g550 (n901, n167);
not  g551 (n792, n217);
not  g552 (n568, n401);
buf  g553 (n867, n92);
buf  g554 (n724, n415);
buf  g555 (n740, n469);
not  g556 (n882, n386);
not  g557 (n893, n463);
not  g558 (n853, n128);
buf  g559 (n802, n502);
not  g560 (n645, n171);
buf  g561 (n886, n486);
buf  g562 (n734, n211);
buf  g563 (n661, n195);
buf  g564 (n769, n496);
not  g565 (n881, n472);
buf  g566 (n700, n156);
not  g567 (n795, n192);
not  g568 (n666, n381);
buf  g569 (n696, n142);
buf  g570 (n729, n81);
buf  g571 (n818, n488);
buf  g572 (n783, n167);
buf  g573 (n545, n143);
not  g574 (n532, n478);
buf  g575 (n860, n459);
not  g576 (n855, n220);
not  g577 (n785, n443);
not  g578 (n564, n104);
buf  g579 (n736, n402);
buf  g580 (n604, n475);
buf  g581 (n637, n127);
buf  g582 (n890, n95);
buf  g583 (n648, n145);
buf  g584 (n551, n114);
not  g585 (n558, n114);
buf  g586 (n832, n491);
buf  g587 (n817, n202);
buf  g588 (n626, n446);
buf  g589 (n906, n96);
not  g590 (n885, n431);
not  g591 (n752, n203);
not  g592 (n616, n405);
buf  g593 (n835, n84);
not  g594 (n593, n464);
buf  g595 (n784, n90);
not  g596 (n805, n502);
not  g597 (n877, n137);
buf  g598 (n838, n107);
not  g599 (n874, n415);
not  g600 (n847, n487);
not  g601 (n618, n116);
or   g602 (n848, n422, n197, n214, n381);
nor  g603 (n819, n506, n161, n474, n110);
nand g604 (n643, n456, n416, n133, n439);
xnor g605 (n765, n164, n403, n464, n446);
xor  g606 (n745, n460, n101, n517, n127);
and  g607 (n875, n405, n148, n489, n377);
nand g608 (n825, n90, n390, n479, n427);
nor  g609 (n617, n511, n461, n449, n515);
or   g610 (n655, n410, n159, n467, n109);
or   g611 (n692, n200, n377, n383, n473);
nand g612 (n738, n429, n395, n408);
xor  g613 (n701, n165, n194, n136, n215);
nor  g614 (n815, n120, n439, n387, n411);
or   g615 (n713, n467, n466, n505, n211);
xnor g616 (n693, n477, n443, n498, n93);
or   g617 (n857, n465, n401, n470, n217);
xnor g618 (n870, n500, n114, n217, n453);
nor  g619 (n687, n186, n463, n508, n456);
xnor g620 (n607, n444, n400, n216, n399);
xnor g621 (n581, n199, n413, n106, n475);
nor  g622 (n602, n117, n120, n401, n180);
and  g623 (n829, n391, n497, n520, n119);
xor  g624 (n814, n189, n174, n457, n468);
nand g625 (n542, n195, n152, n197);
or   g626 (n806, n154, n79, n219, n87);
and  g627 (n899, n499, n91, n418, n102);
nor  g628 (n858, n176, n419, n509, n440);
nor  g629 (n635, n79, n132, n396, n433);
xnor g630 (n614, n483, n85, n115, n379);
nand g631 (n560, n174, n89, n98, n209);
nand g632 (n854, n130, n192, n105, n399);
or   g633 (n534, n385, n94, n82, n484);
and  g634 (n649, n87, n121, n414, n124);
xnor g635 (n749, n503, n134, n190, n158);
and  g636 (n639, n85, n217, n393, n183);
xnor g637 (n807, n133, n100, n493, n194);
nand g638 (n694, n445, n395, n443, n193);
xnor g639 (n565, n437, n151, n160, n122);
nor  g640 (n884, n381, n158, n449, n455);
or   g641 (n865, n422, n121, n106, n434);
and  g642 (n664, n93, n82, n215, n111);
xor  g643 (n699, n517, n101, n200, n180);
and  g644 (n554, n452, n462, n400, n441);
xor  g645 (n657, n488, n144, n494, n432);
nand g646 (n897, n120, n193, n449, n131);
xor  g647 (n836, n384, n148, n392, n509);
xnor g648 (n851, n196, n154, n392, n482);
xnor g649 (n849, n205, n132, n162, n434);
xnor g650 (n844, n500, n146, n409, n136);
or   g651 (n889, n81, n513, n170, n163);
xor  g652 (n557, n434, n190, n424, n415);
and  g653 (n803, n216, n396, n391, n382);
and  g654 (n711, n407, n125, n100, n384);
xor  g655 (n563, n459, n169, n374, n394);
and  g656 (n872, n495, n109, n169, n448);
xnor g657 (n725, n431, n420, n168, n171);
nor  g658 (n780, n126, n89, n221, n379);
or   g659 (n620, n178, n383, n141, n503);
xor  g660 (n864, n213, n450, n186, n82);
and  g661 (n566, n409, n86, n188, n458);
xnor g662 (n606, n152, n117, n208, n383);
xor  g663 (n612, n140, n145, n482, n479);
or   g664 (n695, n514, n518, n417, n477);
xnor g665 (n883, n110, n215, n124, n166);
nand g666 (n600, n164, n489, n456, n186);
and  g667 (n677, n465, n432, n482, n471);
xnor g668 (n721, n475, n518, n180, n204);
and  g669 (n690, n155, n375, n426, n450);
xnor g670 (n673, n210, n109, n411, n468);
nor  g671 (n631, n91, n156, n130, n135);
xnor g672 (n702, n416, n481, n153, n508);
xnor g673 (n624, n98, n146, n183, n154);
xor  g674 (n714, n134, n382, n490, n391);
xor  g675 (n717, n519, n513, n393, n451);
xnor g676 (n544, n391, n490, n389, n476);
or   g677 (n548, n424, n98, n410, n123);
and  g678 (n669, n385, n218, n135, n130);
and  g679 (n759, n406, n515, n194, n436);
nor  g680 (n868, n480, n161, n177, n166);
nand g681 (n895, n193, n153, n150, n112);
nor  g682 (n676, n503, n119, n212, n423);
xor  g683 (n748, n402, n179, n419, n113);
xnor g684 (n623, n385, n107, n397, n388);
and  g685 (n782, n92, n88, n122, n507);
xnor g686 (n538, n183, n181, n378, n460);
or   g687 (n821, n462, n113, n474, n213);
xnor g688 (n770, n215, n397, n138, n468);
xnor g689 (n727, n476, n440, n195, n150);
or   g690 (n629, n516, n439, n469, n494);
and  g691 (n758, n467, n389, n426, n438);
xor  g692 (n907, n392, n455, n407, n493);
xor  g693 (n722, n417, n209, n213, n433);
or   g694 (n555, n478, n513, n220, n471);
nor  g695 (n580, n138, n173, n149, n146);
or   g696 (n720, n214, n407, n506, n87);
xnor g697 (n656, n388, n495, n398, n487);
xor  g698 (n553, n458, n484, n510, n409);
and  g699 (n662, n95, n193, n481, n192);
nor  g700 (n812, n169, n141, n220, n410);
or   g701 (n641, n517, n205, n472, n219);
nor  g702 (n636, n405, n81, n106, n375);
nor  g703 (n539, n489, n465, n156, n433);
nand g704 (n790, n483, n87, n181, n85);
xor  g705 (n834, n480, n121, n460, n376);
nor  g706 (n826, n84, n140, n388, n406);
nor  g707 (n628, n180, n152, n126, n374);
xor  g708 (n644, n497, n482, n213, n80);
and  g709 (n880, n88, n208, n145, n454);
nor  g710 (n599, n86, n220, n125, n501);
xor  g711 (n587, n473, n168, n437, n444);
nand g712 (n590, n208, n160, n492, n440);
and  g713 (n550, n501, n381, n425, n165);
or   g714 (n552, n378, n144, n506, n173);
xnor g715 (n843, n420, n86, n387, n82);
nor  g716 (n712, n455, n444, n499, n469);
nor  g717 (n586, n426, n83, n205, n404);
xnor g718 (n791, n485, n182, n178, n438);
xnor g719 (n646, n468, n103, n90, n165);
or   g720 (n859, n483, n210, n105, n198);
xnor g721 (n771, n502, n419, n462, n408);
nand g722 (n633, n432, n80, n118, n440);
xor  g723 (n533, n396, n96, n470, n176);
and  g724 (n766, n478, n177, n131, n94);
xor  g725 (n642, n182, n387, n131, n486);
nand g726 (n674, n163, n514, n204, n168);
nand g727 (n824, n185, n168, n403, n136);
xor  g728 (n543, n157, n417, n490, n122);
and  g729 (n579, n496, n120, n196, n199);
xnor g730 (n671, n424, n516, n108, n167);
xnor g731 (n869, n393, n423, n218, n452);
or   g732 (n797, n187, n406, n155, n499);
xnor g733 (n774, n141, n441, n498, n394);
or   g734 (n597, n494, n406, n105, n452);
or   g735 (n779, n382, n135, n111, n169);
or   g736 (n822, n432, n421, n172, n414);
nor  g737 (n878, n377, n447, n104, n380);
xor  g738 (n879, n111, n202, n99, n431);
or   g739 (n537, n450, n140, n378, n497);
xor  g740 (n896, n103, n431, n384, n121);
nor  g741 (n575, n124, n476, n212, n113);
and  g742 (n856, n101, n511, n218, n451);
and  g743 (n691, n185, n516, n80, n83);
nand g744 (n733, n394, n508, n83, n153);
xnor g745 (n715, n505, n221, n164, n141);
nand g746 (n728, n409, n158, n488, n427);
xor  g747 (n608, n413, n162, n412, n140);
xnor g748 (n768, n460, n197, n108, n467);
xor  g749 (n804, n103, n451, n170, n477);
xnor g750 (n621, n115, n96, n130, n94);
nand g751 (n584, n181, n209, n133, n212);
nand g752 (n592, n112, n142, n486, n204);
or   g753 (n531, n174, n157, n422, n485);
nor  g754 (n837, n173, n92, n485, n126);
nor  g755 (n594, n429, n412, n427, n457);
nand g756 (n705, n159, n405, n470, n480);
xor  g757 (n688, n436, n208, n149, n176);
nand g758 (n845, n145, n456, n132, n496);
xor  g759 (n658, n519, n485, n97, n89);
or   g760 (n595, n137, n143, n179, n453);
nor  g761 (n703, n510, n102, n459, n494);
xnor g762 (n787, n134, n473, n118, n386);
xnor g763 (n830, n486, n435, n157, n452);
nor  g764 (n750, n83, n125, n509, n100);
or   g765 (n892, n453, n471, n481, n79);
nand g766 (n573, n177, n100, n400, n106);
and  g767 (n683, n143, n95, n461, n205);
nand g768 (n680, n383, n155, n462, n403);
xnor g769 (n887, n448, n204, n93, n160);
xnor g770 (n850, n466, n177, n144, n84);
nand g771 (n668, n481, n487, n144, n200);
and  g772 (n746, n428, n93, n512, n398);
nand g773 (n798, n517, n191, n443, n195);
nand g774 (n796, n419, n410, n401, n201);
xnor g775 (n562, n423, n92, n498, n510);
xnor g776 (n583, n179, n412, n209, n89);
or   g777 (n585, n509, n417, n498, n99);
and  g778 (n737, n402, n515, n110, n403);
xnor g779 (n808, n191, n414, n503, n102);
or   g780 (n627, n88, n459, n182, n375);
nor  g781 (n756, n198, n464, n448, n389);
or   g782 (n716, n464, n447, n408, n152);
or   g783 (n698, n110, n80, n219, n123);
nor  g784 (n571, n188, n496, n118, n125);
and  g785 (n670, n184, n477, n115, n423);
nor  g786 (n630, n377, n129, n396, n149);
xnor g787 (n820, n99, n214, n418, n484);
nor  g788 (n823, n142, n134, n136, n471);
or   g789 (n833, n476, n451, n495, n385);
and  g790 (n540, n207, n379, n411, n192);
nor  g791 (n622, n172, n201, n207, n189);
xor  g792 (n706, n429, n413, n436, n116);
xor  g793 (n903, n490, n492, n500, n399);
or   g794 (n764, n109, n178, n470, n173);
and  g795 (n813, n408, n430, n170, n203);
nor  g796 (n905, n184, n491, n439, n420);
xnor g797 (n739, n123, n424, n159, n444);
or   g798 (n625, n473, n147, n442, n421);
xnor g799 (n653, n398, n507, n441, n91);
or   g800 (n535, n137, n176, n447, n399);
and  g801 (n574, n148, n446, n495, n463);
xor  g802 (n762, n407, n139, n101, n97);
or   g803 (n577, n202, n150, n129, n123);
or   g804 (n682, n175, n153, n386, n198);
xor  g805 (n732, n515, n491, n448, n505);
or   g806 (n547, n128, n187, n154, n501);
nand g807 (n731, n81, n112, n453, n147);
and  g808 (n852, n97, n115, n516, n519);
xor  g809 (n809, n170, n111, n139, n397);
nor  g810 (n891, n122, n218, n211, n491);
nor  g811 (n761, n469, n404, n466, n457);
xnor g812 (n757, n421, n458, n461, n150);
nand g813 (n654, n104, n90, n416, n435);
nand g814 (n816, n394, n374, n442, n436);
xor  g815 (n611, n390, n428, n172, n189);
xnor g816 (n841, n446, n493, n190, n164);
or   g817 (n707, n404, n103, n206, n105);
xnor g818 (n572, n416, n132, n196, n457);
and  g819 (n605, n151, n214, n155, n216);
nand g820 (n777, n454, n172, n88, n163);
xor  g821 (n613, n449, n380, n474, n166);
xnor g822 (n888, n202, n185, n437, n388);
xnor g823 (n842, n139, n519, n430, n184);
xnor g824 (n786, n489, n501, n375, n203);
xor  g825 (n744, n434, n162, n163, n376);
and  g826 (n685, n199, n157, n507, n129);
and  g827 (n619, n113, n442, n474, n507);
xnor g828 (n894, n376, n126, n149, n426);
and  g829 (n793, n108, n188, n502, n201);
xnor g830 (n650, n147, n479, n119, n518);
xor  g831 (n678, n421, n210, n425, n454);
and  g832 (n601, n428, n191, n376, n512);
or   g833 (n569, n189, n397, n447, n85);
and  g834 (n652, n458, n418, n178, n210);
and  g835 (n567, n386, n219, n466, n514);
xnor g836 (n846, n137, n425, n393, n191);
nor  g837 (n827, n148, n95, n84, n190);
and  g838 (n576, n187, n480, n513, n143);
xor  g839 (n839, n497, n207, n99, n156);
nor  g840 (n840, n398, n504, n510, n465);
xnor g841 (n904, n413, n142, n472, n216);
and  g842 (n900, n107, n499, n508, n427);
nand g843 (n667, n166, n198, n146, n390);
xnor g844 (n556, n389, n127, n117, n380);
nand g845 (n788, n158, n114, n203, n511);
nor  g846 (n767, n445, n422, n455, n201);
nand g847 (n876, n104, n441, n484, n425);
nor  g848 (n773, n206, n181, n461, n159);
and  g849 (n862, n165, n463, n116, n199);
nor  g850 (n570, n129, n138, n133, n128);
and  g851 (n647, n387, n183, n411, n429);
nand g852 (n708, n438, n167, n511, n187);
xor  g853 (n634, n206, n179, n194, n504);
or   g854 (n871, n430, n79, n395, n384);
nand g855 (n735, n91, n479, n97, n160);
nand g856 (n697, n445, n124, n435, n108);
nand g857 (n632, n493, n98, n435, n433);
xnor g858 (n831, n102, n207, n378, n514);
xnor g859 (n659, n174, n171, n454, n116);
or   g860 (n546, n112, n382, n392, n390);
not  g861 (n909, n531);
nand g862 (n908, n520, n530);
nor  g863 (n910, n532, n534, n908, n533);
buf  g864 (n912, n910);
not  g865 (n911, n910);
nand g866 (n915, n538, n540);
xor  g867 (n913, n539, n912, n536, n537);
nand g868 (n914, n912, n535, n911, n541);
xor  g869 (n919, n545, n546, n915);
nand g870 (n920, n544, n550, n913);
xor  g871 (n917, n547, n915);
nand g872 (n916, n548, n912, n549);
or   g873 (n918, n912, n543, n914, n542);
buf  g874 (n921, n917);
not  g875 (n922, n916);
not  g876 (n927, n917);
buf  g877 (n925, n916);
not  g878 (n928, n917);
not  g879 (n924, n917);
buf  g880 (n926, n916);
not  g881 (n923, n916);
or   g882 (n929, n919, n918, n523, n520);
nor  g883 (n934, n921, n521, n919);
nand g884 (n932, n921, n523, n922);
xnor g885 (n936, n918, n522, n521);
xor  g886 (n935, n522, n521, n918, n520);
xor  g887 (n933, n922, n920, n522);
or   g888 (n930, n922, n922, n523, n919);
nand g889 (n931, n921, n921, n521, n918);
not  g890 (n937, n923);
and  g891 (n938, n930, n929, n923);
xnor g892 (n940, n938, n933, n937);
nor  g893 (n941, n936, n920, n938);
nor  g894 (n943, n937, n934, n938);
xnor g895 (n942, n935, n932, n931, n930);
xnor g896 (n939, n932, n935, n931, n936);
buf  g897 (n952, n923);
not  g898 (n953, n939);
buf  g899 (n960, n939);
buf  g900 (n951, n940);
buf  g901 (n955, n943);
buf  g902 (n962, n941);
buf  g903 (n959, n942);
buf  g904 (n950, n941);
not  g905 (n949, n941);
buf  g906 (n947, n943);
buf  g907 (n956, n942);
not  g908 (n958, n940);
not  g909 (n957, n940);
not  g910 (n945, n940);
buf  g911 (n954, n943);
buf  g912 (n948, n942);
not  g913 (n946, n941);
buf  g914 (n944, n938);
nand g915 (n961, n939, n943, n942);
buf  g916 (n992, n949);
buf  g917 (n988, n947);
not  g918 (n1000, n956);
buf  g919 (n1011, n954);
buf  g920 (n974, n948);
not  g921 (n989, n956);
not  g922 (n972, n953);
buf  g923 (n985, n954);
buf  g924 (n965, n946);
not  g925 (n997, n956);
not  g926 (n998, n953);
not  g927 (n1009, n955);
buf  g928 (n973, n947);
not  g929 (n995, n957);
buf  g930 (n979, n952);
not  g931 (n1007, n944);
not  g932 (n994, n948);
not  g933 (n999, n946);
buf  g934 (n1013, n957);
buf  g935 (n966, n945);
buf  g936 (n983, n945);
buf  g937 (n1012, n951);
not  g938 (n1008, n944);
buf  g939 (n971, n944);
not  g940 (n987, n947);
not  g941 (n1004, n944);
not  g942 (n967, n945);
buf  g943 (n990, n955);
not  g944 (n976, n952);
not  g945 (n984, n946);
buf  g946 (n977, n948);
buf  g947 (n986, n954);
not  g948 (n980, n950);
buf  g949 (n1015, n952);
buf  g950 (n1005, n955);
not  g951 (n1014, n953);
buf  g952 (n1002, n951);
buf  g953 (n975, n949);
buf  g954 (n982, n946);
buf  g955 (n991, n951);
buf  g956 (n981, n950);
buf  g957 (n969, n945);
buf  g958 (n996, n951);
buf  g959 (n993, n953);
not  g960 (n964, n954);
buf  g961 (n1001, n947);
buf  g962 (n1010, n950);
not  g963 (n1003, n949);
not  g964 (n1016, n956);
not  g965 (n970, n949);
not  g966 (n963, n955);
buf  g967 (n968, n950);
buf  g968 (n1006, n952);
not  g969 (n978, n948);
xnor g970 (n1024, n965, n966, n963, n961);
nor  g971 (n1020, n962, n960, n959);
xor  g972 (n1026, n959, n965, n961);
xor  g973 (n1022, n967, n964, n960, n958);
nor  g974 (n1021, n967, n965, n966, n961);
and  g975 (n1023, n963, n964, n962);
xor  g976 (n1019, n962, n957, n966, n965);
or   g977 (n1017, n962, n963, n959, n958);
nor  g978 (n1025, n958, n964, n963, n957);
xnor g979 (n1018, n958, n959, n966, n960);
xor  g980 (n1030, n968, n969);
and  g981 (n1029, n969, n971, n1020);
nor  g982 (n1032, n967, n968, n970);
or   g983 (n1028, n1018, n969, n970);
xor  g984 (n1031, n1021, n1017, n969, n970);
nand g985 (n1027, n967, n1019, n1020, n968);
not  g986 (n1035, n1032);
buf  g987 (n1036, n1029);
buf  g988 (n1037, n1030);
not  g989 (n1039, n1027);
buf  g990 (n1034, n1032);
not  g991 (n1038, n1028);
not  g992 (n1040, n1031);
buf  g993 (n1033, n1031);
nand g994 (n1044, n972, n986, n1038, n973);
xor  g995 (n1071, n1039, n1040, n989, n987);
nor  g996 (n1048, n988, n1035, n979);
xor  g997 (n1054, n1039, n524, n990, n984);
nor  g998 (n1042, n983, n988, n974, n1035);
xor  g999 (n1072, n975, n992, n971, n982);
nor  g1000 (n1052, n981, n1037, n990, n1034);
and  g1001 (n1050, n980, n977, n989, n1039);
nor  g1002 (n1064, n1039, n984, n975);
or   g1003 (n1059, n1037, n972, n524, n976);
or   g1004 (n1062, n1036, n987, n1033, n552);
nor  g1005 (n1066, n993, n989, n978, n981);
and  g1006 (n1047, n991, n974, n1040, n973);
and  g1007 (n1061, n985, n977, n1034, n983);
xor  g1008 (n1057, n980, n986, n988, n1040);
and  g1009 (n1053, n982, n984, n973, n972);
xor  g1010 (n1041, n1035, n979, n1036, n976);
xnor g1011 (n1051, n975, n551, n987, n985);
xnor g1012 (n1056, n1038, n985, n977, n980);
and  g1013 (n1068, n524, n1038, n983, n987);
xnor g1014 (n1046, n981, n978, n993);
xor  g1015 (n1063, n972, n980, n1038, n553);
and  g1016 (n1043, n524, n992, n979, n982);
xor  g1017 (n1058, n1033, n971, n983, n975);
xor  g1018 (n1070, n981, n974, n1036, n978);
xnor g1019 (n1060, n986, n1033, n978);
xor  g1020 (n1065, n990, n976, n988, n982);
and  g1021 (n1069, n1034, n1040, n973, n990);
xor  g1022 (n1049, n976, n974, n991, n992);
xor  g1023 (n1055, n991, n1037, n985);
or   g1024 (n1067, n989, n991, n986, n1036);
xor  g1025 (n1045, n992, n977, n979, n1034);
xor  g1026 (n1116, n782, n1062, n603, n792);
or   g1027 (n1113, n735, n736, n1043, n619);
nand g1028 (n1151, n1043, n798, n738, n872);
or   g1029 (n1171, n617, n803, n645, n1046);
or   g1030 (n1174, n1052, n689, n828, n1064);
or   g1031 (n1079, n831, n1063, n1059, n627);
nand g1032 (n1078, n837, n1064, n1062, n620);
and  g1033 (n1074, n676, n585, n783, n564);
nor  g1034 (n1177, n829, n1063, n720, n723);
nor  g1035 (n1143, n594, n838, n573, n1045);
xor  g1036 (n1155, n725, n1049, n652, n681);
or   g1037 (n1110, n582, n849, n698, n751);
nor  g1038 (n1130, n1041, n1067, n571, n867);
xnor g1039 (n1077, n561, n661, n635, n687);
and  g1040 (n1081, n823, n760, n871, n593);
xor  g1041 (n1105, n748, n1053, n852, n622);
xor  g1042 (n1121, n606, n1042, n670, n776);
and  g1043 (n1088, n655, n664, n638, n712);
xor  g1044 (n1163, n879, n706, n686, n809);
and  g1045 (n1172, n814, n1057, n1058, n604);
xnor g1046 (n1086, n1065, n568, n589, n806);
xnor g1047 (n1156, n768, n673, n710, n636);
nor  g1048 (n1099, n808, n767, n764, n1051);
nor  g1049 (n1165, n1056, n844, n1049, n816);
xor  g1050 (n1141, n759, n684, n729, n833);
or   g1051 (n1139, n1060, n878, n810, n777);
nand g1052 (n1176, n790, n572, n1068, n818);
xnor g1053 (n1109, n1049, n1060, n701, n1052);
nand g1054 (n1145, n774, n1051, n567, n860);
or   g1055 (n1140, n731, n1053, n804, n1052);
and  g1056 (n1085, n682, n794, n665, n1044);
or   g1057 (n1104, n850, n574, n609, n1067);
xor  g1058 (n1117, n854, n740, n737, n1066);
xnor g1059 (n1160, n826, n1056, n679, n1048);
and  g1060 (n1087, n1057, n784, n646, n575);
or   g1061 (n1173, n709, n598, n697, n1059);
xor  g1062 (n1136, n848, n752, n868, n874);
nand g1063 (n1091, n749, n692, n1050, n1053);
xor  g1064 (n1092, n1061, n1048, n576, n663);
or   g1065 (n1094, n578, n1051, n822, n649);
or   g1066 (n1076, n728, n858, n597, n1056);
xnor g1067 (n1149, n626, n743, n836, n866);
and  g1068 (n1133, n1058, n869, n827, n650);
xor  g1069 (n1178, n654, n861, n842, n602);
xnor g1070 (n1168, n702, n713, n840, n680);
xnor g1071 (n1119, n770, n715, n660, n586);
xnor g1072 (n1102, n1057, n820, n562, n755);
and  g1073 (n1152, n1063, n704, n730, n719);
nor  g1074 (n1073, n560, n714, n667, n747);
or   g1075 (n1125, n726, n648, n781, n1067);
xnor g1076 (n1107, n1066, n640, n583, n1056);
nand g1077 (n1162, n769, n778, n685, n839);
and  g1078 (n1122, n847, n1043, n559, n1054);
or   g1079 (n1100, n787, n1045, n811);
nor  g1080 (n1128, n788, n853, n718, n802);
xor  g1081 (n1082, n876, n625, n555, n1047);
nor  g1082 (n1118, n1043, n841, n717, n616);
nor  g1083 (n1138, n789, n851, n830, n780);
xnor g1084 (n1153, n1046, n668, n721, n1050);
xor  g1085 (n1083, n639, n581, n815, n596);
xor  g1086 (n1134, n800, n1055, n587, n1048);
or   g1087 (n1158, n753, n1041, n843, n677);
nand g1088 (n1101, n565, n584, n1060, n666);
nor  g1089 (n1132, n672, n577, n628, n1066);
nor  g1090 (n1142, n1065, n659, n870, n1062);
xor  g1091 (n1169, n556, n656, n845, n591);
nor  g1092 (n1159, n631, n641, n1057, n653);
nor  g1093 (n1120, n1063, n807, n1045, n825);
xnor g1094 (n1126, n855, n621, n1064, n592);
nand g1095 (n1144, n1064, n745, n1049, n1046);
xnor g1096 (n1108, n599, n727, n793, n644);
xor  g1097 (n1111, n796, n791, n595, n766);
and  g1098 (n1181, n691, n657, n824, n744);
xor  g1099 (n1137, n590, n683, n607, n856);
xor  g1100 (n1179, n754, n612, n630, n569);
xor  g1101 (n1103, n1044, n1055, n554, n733);
xnor g1102 (n1095, n711, n690, n1041, n832);
or   g1103 (n1175, n699, n1047, n865, n724);
or   g1104 (n1147, n757, n1067, n694, n674);
xnor g1105 (n1075, n614, n746, n863, n608);
nand g1106 (n1170, n615, n819, n813, n1046);
nor  g1107 (n1123, n765, n1065, n1052, n741);
or   g1108 (n1096, n643, n675, n1051, n618);
nor  g1109 (n1146, n763, n864, n1055, n1054);
xor  g1110 (n1167, n605, n821, n786, n1054);
or   g1111 (n1150, n1061, n739, n875, n563);
or   g1112 (n1157, n801, n797, n1058, n756);
nor  g1113 (n1090, n750, n1068, n812, n742);
nand g1114 (n1127, n880, n805, n732, n634);
and  g1115 (n1114, n611, n734, n632, n846);
or   g1116 (n1097, n1061, n637, n633, n1048);
xor  g1117 (n1164, n773, n795, n1044, n1065);
nor  g1118 (n1098, n613, n873, n1059, n566);
or   g1119 (n1148, n580, n669, n775, n558);
xnor g1120 (n1129, n817, n658, n662, n1042);
nor  g1121 (n1154, n1044, n610, n1050);
or   g1122 (n1161, n557, n835, n623, n1062);
nand g1123 (n1124, n772, n708, n722, n705);
and  g1124 (n1180, n579, n834, n1042, n688);
xnor g1125 (n1084, n799, n1059, n857, n624);
xnor g1126 (n1112, n1066, n1053, n716, n629);
or   g1127 (n1080, n877, n1054, n1061, n700);
xor  g1128 (n1089, n1058, n1047, n771, n600);
nand g1129 (n1135, n785, n642, n678, n1047);
and  g1130 (n1131, n651, n703, n1055, n862);
xnor g1131 (n1115, n696, n1042, n758, n707);
nor  g1132 (n1106, n570, n693, n762, n779);
nor  g1133 (n1093, n601, n671, n588, n695);
and  g1134 (n1166, n1060, n761, n647, n859);
or   g1135 (n1182, n1073, n1074, n1075, n1076);
not  g1136 (n1185, n1079);
not  g1137 (n1184, n1182);
xor  g1138 (n1183, n1077, n1182, n1078);
nand g1139 (n1186, n889, n881, n883, n888);
xnor g1140 (n1196, n994, n1184, n898);
xor  g1141 (n1192, n884, n1183, n525, n895);
nor  g1142 (n1189, n885, n1080, n900, n893);
xor  g1143 (n1194, n891, n896, n1185, n899);
and  g1144 (n1193, n892, n897, n1184, n1068);
and  g1145 (n1190, n1069, n1183, n994, n887);
or   g1146 (n1191, n1185, n1183, n1069, n525);
xor  g1147 (n1187, n993, n1081, n1068, n894);
nand g1148 (n1188, n525, n901, n1184, n1185);
xnor g1149 (n1195, n886, n1183, n882, n890);
or   g1150 (n1198, n1195, n1084);
xnor g1151 (n1197, n1082, n1083, n1196);
and  g1152 (n1204, n1101, n1102, n1197, n1198);
and  g1153 (n1203, n1197, n1198, n1099, n1098);
xnor g1154 (n1200, n1090, n1104, n1198, n1091);
nand g1155 (n1199, n1105, n1198, n1095, n1086);
xnor g1156 (n1202, n1093, n1097, n1087, n1092);
and  g1157 (n1205, n1088, n1085, n1089, n1094);
xor  g1158 (n1201, n1096, n1197, n1103, n1100);
and  g1159 (n1214, n909, n925, n1204);
and  g1160 (n1211, n1199, n1106, n1111, n924);
xor  g1161 (n1208, n1205, n908, n924);
nor  g1162 (n1207, n1114, n924, n909, n908);
or   g1163 (n1213, n925, n1113, n1108, n1205);
xor  g1164 (n1206, n1185, n1109, n1112, n525);
xnor g1165 (n1210, n925, n1201, n909, n924);
nand g1166 (n1209, n1110, n1202, n1200, n923);
xor  g1167 (n1212, n1107, n1203, n1204, n909);
or   g1168 (n1221, n1207, n1209, n529, n1071);
xor  g1169 (n1224, n1071, n526, n1211, n1209);
or   g1170 (n1218, n529, n529, n527, n1206);
xnor g1171 (n1216, n527, n1069, n528, n1072);
xnor g1172 (n1215, n527, n1069, n1208, n528);
xnor g1173 (n1217, n1210, n1210, n1072, n529);
xnor g1174 (n1222, n1070, n1070, n526, n1072);
nor  g1175 (n1219, n1208, n1071, n526, n1072);
nand g1176 (n1223, n1207, n1070, n1071, n528);
nor  g1177 (n1220, n526, n528, n527, n1070);
xnor g1178 (n1230, n1218, n1224, n1217, n1123);
nand g1179 (n1228, n1139, n1129, n1137, n1116);
xor  g1180 (n1231, n1117, n1119, n1219, n1115);
nand g1181 (n1233, n1222, n1118, n1223, n1125);
nor  g1182 (n1225, n1127, n1122, n1131, n1136);
and  g1183 (n1226, n1140, n1221, n1138, n1120);
nor  g1184 (n1227, n1133, n1220, n1126, n1121);
or   g1185 (n1229, n1135, n1130, n1141, n1132);
and  g1186 (n1232, n1216, n1124, n1134, n1128);
or   g1187 (n1251, n1229, n223, n226, n222);
xor  g1188 (n1248, n227, n225, n230, n1227);
nand g1189 (n1247, n222, n926, n227, n1022);
xor  g1190 (n1239, n222, n1226, n1142, n928);
nand g1191 (n1245, n927, n1225, n1021, n228);
xnor g1192 (n1249, n229, n229, n1143, n221);
and  g1193 (n1243, n927, n229, n1228);
nor  g1194 (n1242, n230, n224, n926, n928);
nand g1195 (n1238, n1227, n1229, n225, n223);
and  g1196 (n1235, n228, n223, n226);
xnor g1197 (n1240, n1022, n228, n1228, n1229);
nor  g1198 (n1250, n1229, n230, n927, n1226);
and  g1199 (n1236, n1227, n226, n227, n926);
nor  g1200 (n1237, n1226, n926, n1228, n224);
or   g1201 (n1241, n226, n228, n227, n221);
nor  g1202 (n1244, n1226, n927, n225, n928);
or   g1203 (n1234, n222, n224, n1225, n1228);
or   g1204 (n1246, n230, n225, n224, n1227);
buf  g1205 (n1257, n1230);
buf  g1206 (n1260, n1232);
not  g1207 (n1258, n1244);
not  g1208 (n1263, n1239);
and  g1209 (n1253, n1149, n1146, n1249, n1238);
nor  g1210 (n1254, n1148, n1231);
nor  g1211 (n1259, n1247, n1151, n1245, n1147);
xnor g1212 (n1252, n1230, n1150, n1246, n1233);
nand g1213 (n1256, n1145, n1232, n1231, n1233);
and  g1214 (n1261, n1242, n1240, n1233, n1232);
and  g1215 (n1262, n1230, n1241, n1248, n1243);
xor  g1216 (n1255, n1230, n1232, n1233, n1144);
nor  g1217 (n1267, n1259, n1255, n1001, n1009);
and  g1218 (n1265, n1014, n1016, n1255, n1214);
xor  g1219 (n1278, n1254, n1012, n1258, n1002);
nand g1220 (n1296, n1260, n1000, n1262, n997);
nand g1221 (n1272, n1252, n1260, n1005);
or   g1222 (n1274, n1011, n1015, n1213);
xor  g1223 (n1294, n997, n1212, n1012, n998);
nor  g1224 (n1276, n1007, n1008, n1003, n1009);
or   g1225 (n1280, n1251, n1007, n999, n1008);
or   g1226 (n1277, n1006, n1001, n1261);
xnor g1227 (n1264, n1013, n1012, n1015, n1258);
nand g1228 (n1286, n1007, n1254, n1258, n1010);
nand g1229 (n1283, n1010, n1253, n1262);
xnor g1230 (n1281, n1252, n1261, n1003, n1005);
xnor g1231 (n1282, n999, n998, n1256, n995);
xor  g1232 (n1269, n1214, n1260, n1254, n1002);
nand g1233 (n1301, n1253, n999, n904, n1013);
xor  g1234 (n1279, n1004, n995, n999, n994);
xnor g1235 (n1297, n1260, n1010, n1255, n1003);
or   g1236 (n1300, n996, n1009, n1257, n1015);
or   g1237 (n1290, n1213, n995, n1006, n1012);
xor  g1238 (n1285, n1014, n1254, n906, n998);
xnor g1239 (n1289, n1259, n1262, n1261);
nor  g1240 (n1273, n1211, n1011, n997, n1250);
xor  g1241 (n1291, n1008, n1258, n1007, n1003);
nor  g1242 (n1292, n1011, n1259, n996, n1256);
and  g1243 (n1287, n1256, n1001, n907, n902);
or   g1244 (n1288, n995, n906, n1008, n1014);
xnor g1245 (n1266, n1257, n1002, n994, n1004);
or   g1246 (n1284, n1004, n1253, n905);
and  g1247 (n1270, n907, n996, n1005, n1010);
and  g1248 (n1299, n1257, n1212, n1013, n1252);
xor  g1249 (n1271, n1006, n1011, n1256, n1016);
xnor g1250 (n1295, n928, n997, n1014, n1252);
nor  g1251 (n1298, n1000, n1016, n1255, n1257);
xor  g1252 (n1268, n1016, n1013, n1259, n1002);
nor  g1253 (n1293, n1006, n1009, n1000);
nand g1254 (n1275, n996, n903, n998, n1004);
not  g1255 (n1313, n1264);
buf  g1256 (n1309, n1263);
buf  g1257 (n1304, n1266);
buf  g1258 (n1307, n1275);
buf  g1259 (n1302, n1269);
buf  g1260 (n1303, n1263);
buf  g1261 (n1312, n1273);
buf  g1262 (n1310, n1268);
buf  g1263 (n1305, n1263);
buf  g1264 (n1306, n1271);
or   g1265 (n1308, n1265, n1263);
xnor g1266 (n1311, n1274, n1270, n1267, n1272);
or   g1267 (n1328, n1155, n1303, n1279, n1305);
nor  g1268 (n1324, n1301, n1304, n1152, n1305);
or   g1269 (n1322, n1289, n1285, n1283, n1282);
and  g1270 (n1327, n1299, n1301, n1300, n1281);
nor  g1271 (n1326, n1292, n1293, n1305, n1303);
or   g1272 (n1318, n1157, n1298, n1304, n1286);
xor  g1273 (n1317, n1276, n1297, n1291, n1302);
nor  g1274 (n1315, n1303, n1291, n1296, n1302);
nor  g1275 (n1325, n1299, n1298, n1294, n1278);
xnor g1276 (n1319, n1294, n1284, n1277, n1288);
nand g1277 (n1316, n1293, n1300, n1303, n1286);
nand g1278 (n1321, n1297, n1290, n1287, n1302);
xnor g1279 (n1320, n1280, n1304, n1289, n1292);
xnor g1280 (n1314, n1295, n1290, n1304, n1302);
xnor g1281 (n1323, n1296, n1305, n1156, n1154);
xnor g1282 (n1329, n1287, n1288, n1295, n1153);
nor  g1283 (n1336, n1306, n1310, n1308, n1314);
and  g1284 (n1333, n1310, n1309, n1311, n1316);
xnor g1285 (n1337, n1309, n1308, n1306, n1315);
xnor g1286 (n1331, n1310, n1310, n1306, n1307);
xnor g1287 (n1334, n1309, n1307, n1317, n1311);
xor  g1288 (n1335, n1308, n1316, n1314, n1311);
xor  g1289 (n1332, n1308, n1307, n1309);
and  g1290 (n1330, n1306, n1311, n1315, n1317);
buf  g1291 (n1339, n1336);
not  g1292 (n1338, n1335);
xnor g1293 (n1340, n1177, n1339, n1169);
nand g1294 (n1346, n1175, n1167, n1171, n1162);
nor  g1295 (n1345, n1337, n1338, n1161, n1172);
nor  g1296 (n1347, n1165, n1180, n1339, n1158);
and  g1297 (n1343, n1163, n1179, n1178, n1176);
nor  g1298 (n1342, n1159, n1164, n1173, n1338);
or   g1299 (n1344, n1339, n1174, n1338, n1170);
and  g1300 (n1341, n1160, n1168, n1338, n1166);
xnor g1301 (n1362, n1319, n1345, n1343, n1181);
or   g1302 (n1351, n1341, n1342, n1312);
nor  g1303 (n1361, n1323, n1343, n1344, n1313);
xnor g1304 (n1359, n1321, n1344, n1328, n1342);
nor  g1305 (n1353, n1318, n1328, n1329, n1344);
xor  g1306 (n1348, n1026, n1327, n1347);
nand g1307 (n1349, n1345, n1325, n1322);
or   g1308 (n1352, n1024, n1025, n1329, n1324);
and  g1309 (n1358, n1342, n1323, n1347, n1023);
or   g1310 (n1356, n1026, n1327, n1319, n1341);
nor  g1311 (n1354, n1318, n1343, n1312, n1346);
xnor g1312 (n1357, n1321, n1346, n1341, n1324);
and  g1313 (n1363, n1312, n1313, n1320, n1345);
xnor g1314 (n1360, n1320, n1313, n1322, n1347);
nor  g1315 (n1350, n1326, n1346, n1023, n1025);
xor  g1316 (n1355, n1340, n1024, n1313, n1326);
or   g1317 (n1364, n1349, n1362, n1355, n1357);
nor  g1318 (n1365, n1360, n1351, n1350, n1352);
xnor g1319 (n1366, n1358, n1363, n1356, n1354);
or   g1320 (n1367, n1348, n1361, n1359, n1353);
endmodule
