

module Stat_100_58
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n108,
  n113,
  n110,
  n105,
  n128,
  n129,
  n131,
  n107,
  n122,
  n118,
  n115,
  n127,
  n130,
  n121,
  n102,
  n103,
  n106,
  n132,
  n124,
  n104,
  n125,
  n119,
  n123,
  n116,
  n117,
  n120,
  n109,
  n126,
  n101,
  n114,
  n111,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n112;
  output n108;
  output n113;
  output n110;
  output n105;
  output n128;
  output n129;
  output n131;
  output n107;
  output n122;
  output n118;
  output n115;
  output n127;
  output n130;
  output n121;
  output n102;
  output n103;
  output n106;
  output n132;
  output n124;
  output n104;
  output n125;
  output n119;
  output n123;
  output n116;
  output n117;
  output n120;
  output n109;
  output n126;
  output n101;
  output n114;
  output n111;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    KeyWire_0_60,
    n17
  );


  not
  g1
  (
    KeyWire_0_62,
    n16
  );


  buf
  g2
  (
    KeyWire_0_11,
    n13
  );


  not
  g3
  (
    n45,
    n13
  );


  buf
  g4
  (
    KeyWire_0_38,
    n10
  );


  not
  g5
  (
    KeyWire_0_5,
    n12
  );


  not
  g6
  (
    KeyWire_0_30,
    n16
  );


  buf
  g7
  (
    KeyWire_0_12,
    n9
  );


  not
  g8
  (
    KeyWire_0_39,
    n15
  );


  buf
  g9
  (
    KeyWire_0_3,
    n17
  );


  buf
  g10
  (
    n61,
    n14
  );


  buf
  g11
  (
    KeyWire_0_32,
    n18
  );


  buf
  g12
  (
    KeyWire_0_10,
    n1
  );


  not
  g13
  (
    n40,
    n14
  );


  buf
  g14
  (
    n72,
    n18
  );


  not
  g15
  (
    n43,
    n5
  );


  buf
  g16
  (
    n55,
    n19
  );


  not
  g17
  (
    KeyWire_0_58,
    n17
  );


  not
  g18
  (
    KeyWire_0_46,
    n11
  );


  not
  g19
  (
    KeyWire_0_61,
    n16
  );


  buf
  g20
  (
    KeyWire_0_55,
    n9
  );


  not
  g21
  (
    n62,
    n11
  );


  not
  g22
  (
    n41,
    n8
  );


  not
  g23
  (
    KeyWire_0_2,
    n11
  );


  buf
  g24
  (
    n39,
    n4
  );


  buf
  g25
  (
    n35,
    n12
  );


  not
  g26
  (
    KeyWire_0_6,
    n3
  );


  not
  g27
  (
    n36,
    n12
  );


  buf
  g28
  (
    KeyWire_0_15,
    n19
  );


  buf
  g29
  (
    KeyWire_0_16,
    n6
  );


  buf
  g30
  (
    n68,
    n9
  );


  not
  g31
  (
    KeyWire_0_20,
    n13
  );


  buf
  g32
  (
    KeyWire_0_18,
    n18
  );


  buf
  g33
  (
    KeyWire_0_63,
    n2
  );


  buf
  g34
  (
    n33,
    n7
  );


  not
  g35
  (
    n64,
    n15
  );


  buf
  g36
  (
    n59,
    n15
  );


  not
  g37
  (
    KeyWire_0_44,
    n10
  );


  buf
  g38
  (
    n54,
    n14
  );


  buf
  g39
  (
    KeyWire_0_33,
    n10
  );


  buf
  g40
  (
    KeyWire_0_48,
    n37
  );


  buf
  g41
  (
    KeyWire_0_19,
    n40
  );


  buf
  g42
  (
    n80,
    n38
  );


  buf
  g43
  (
    KeyWire_0_51,
    n34
  );


  not
  g44
  (
    KeyWire_0_27,
    n36
  );


  buf
  g45
  (
    n74,
    n40
  );


  not
  g46
  (
    n79,
    n35
  );


  nor
  g47
  (
    KeyWire_0_42,
    n33,
    n39,
    n40
  );


  buf
  g48
  (
    KeyWire_0_7,
    n73
  );


  not
  g49
  (
    KeyWire_0_1,
    n75
  );


  not
  g50
  (
    KeyWire_0_56,
    n74
  );


  not
  g51
  (
    KeyWire_0_8,
    n77
  );


  not
  g52
  (
    KeyWire_0_23,
    n76
  );


  nand
  g53
  (
    n96,
    n22,
    n80,
    n81,
    n27
  );


  and
  g54
  (
    n98,
    n32,
    n21,
    n84
  );


  xnor
  g55
  (
    n91,
    n24,
    n78,
    n27,
    n20
  );


  xnor
  g56
  (
    n99,
    n30,
    n85,
    n32
  );


  nand
  g57
  (
    n88,
    n19,
    n25,
    n84,
    n24
  );


  nor
  g58
  (
    KeyWire_0_25,
    n22,
    n84,
    n32,
    n21
  );


  xnor
  g59
  (
    KeyWire_0_22,
    n85,
    n29,
    n23,
    n82
  );


  xor
  g60
  (
    KeyWire_0_37,
    n80,
    n83,
    n31,
    n81
  );


  xor
  g61
  (
    KeyWire_0_50,
    n82,
    n31,
    n27
  );


  xor
  g62
  (
    n86,
    n22,
    n25,
    n83,
    n26
  );


  nand
  g63
  (
    n87,
    n30,
    n30,
    n25,
    n20
  );


  and
  g64
  (
    KeyWire_0_49,
    n23,
    n26,
    n83,
    n82
  );


  and
  g65
  (
    n90,
    n20,
    n79,
    n28,
    n29
  );


  nor
  g66
  (
    n95,
    n23,
    n26,
    n29,
    n24
  );


  or
  g67
  (
    KeyWire_0_35,
    n81,
    n28,
    n80
  );


  nor
  g68
  (
    n121,
    n44,
    n65,
    n56,
    n63
  );


  and
  g69
  (
    KeyWire_0_41,
    n59,
    n52,
    n45,
    n72
  );


  xor
  g70
  (
    KeyWire_0_40,
    n67,
    n62,
    n86,
    n98
  );


  and
  g71
  (
    n123,
    n49,
    n59,
    n65,
    n55
  );


  or
  g72
  (
    n109,
    n93,
    n69,
    n96
  );


  nand
  g73
  (
    KeyWire_0_34,
    n54,
    n70,
    n92,
    n58
  );


  xor
  g74
  (
    KeyWire_0_24,
    n69,
    n43,
    n94,
    n62
  );


  and
  g75
  (
    n125,
    n95,
    n61,
    n93,
    n42
  );


  xor
  g76
  (
    KeyWire_0_21,
    n53,
    n59,
    n60,
    n54
  );


  or
  g77
  (
    KeyWire_0_45,
    n94,
    n51,
    n64,
    n66
  );


  nand
  g78
  (
    n124,
    n46,
    n57,
    n92,
    n47
  );


  xnor
  g79
  (
    KeyWire_0_9,
    n93,
    n72,
    n98,
    n71
  );


  or
  g80
  (
    KeyWire_0_14,
    n56,
    n97,
    n50,
    n64
  );


  nor
  g81
  (
    KeyWire_0_43,
    n42,
    n55,
    n53,
    n63
  );


  and
  g82
  (
    KeyWire_0_17,
    n52,
    n100,
    n97,
    n91
  );


  nor
  g83
  (
    n114,
    n99,
    n94,
    n100,
    n57
  );


  nor
  g84
  (
    n110,
    n98,
    n45,
    n69,
    n61
  );


  or
  g85
  (
    KeyWire_0_59,
    n95,
    n70,
    n87,
    n68
  );


  xor
  g86
  (
    KeyWire_0_4,
    n50,
    n49,
    n43,
    n71
  );


  and
  g87
  (
    KeyWire_0_31,
    n48,
    n56,
    n67,
    n51
  );


  or
  g88
  (
    KeyWire_0_0,
    n61,
    n41,
    n90,
    n70
  );


  xnor
  g89
  (
    KeyWire_0_28,
    n48,
    n62,
    n64,
    n57
  );


  and
  g90
  (
    KeyWire_0_52,
    n50,
    n51,
    n44,
    n41
  );


  xor
  g91
  (
    KeyWire_0_54,
    n45,
    n66,
    n49,
    n99
  );


  nand
  g92
  (
    KeyWire_0_13,
    n60,
    n52,
    n42,
    n97
  );


  nand
  g93
  (
    KeyWire_0_26,
    n96,
    n68,
    n65,
    n63
  );


  and
  g94
  (
    KeyWire_0_47,
    n71,
    n67,
    n89,
    n53
  );


  nor
  g95
  (
    KeyWire_0_36,
    n66,
    n72,
    n55,
    n100
  );


  or
  g96
  (
    n117,
    n46,
    n68,
    n43,
    n47
  );


  or
  g97
  (
    KeyWire_0_57,
    n58,
    n41,
    n95,
    n54
  );


  nand
  g98
  (
    KeyWire_0_53,
    n44,
    n88,
    n58,
    n60
  );


  nor
  g99
  (
    KeyWire_0_29,
    n48,
    n99,
    n47,
    n46
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n131,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n84,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n56,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n42,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n111,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n49,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n38,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n82,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n85,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n119,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n71,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n70,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n58,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n105,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n107,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n34,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n57,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n116,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n69,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n76,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n37,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n129,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n100,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n81,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n106,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n97,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n115,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n75,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n118,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n103,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n67,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n104,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n50,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n60,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n132,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n92,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n128,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n93,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n66,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n46,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n126,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n108,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n73,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n122,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n51,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n130,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n52,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n112,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n77,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n89,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n94,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n78,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n113,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n127,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n120,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n47,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n83,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n101,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n48,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n102,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n63,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n65,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n53,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n44,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

