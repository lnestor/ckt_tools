

module Stat_725_1628
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n655,
  n652,
  n667,
  n666,
  n662,
  n669,
  n653,
  n665,
  n661,
  n651,
  n736,
  n740,
  n737,
  n742,
  n743,
  n738,
  n741,
  n739,
  n746,
  n744,
  n745,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n655;
  output n652;
  output n667;
  output n666;
  output n662;
  output n669;
  output n653;
  output n665;
  output n661;
  output n651;
  output n736;
  output n740;
  output n737;
  output n742;
  output n743;
  output n738;
  output n741;
  output n739;
  output n746;
  output n744;
  output n745;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n654;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n663;
  wire n664;
  wire n668;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n83,
    n15
  );


  buf
  g1
  (
    KeyWire_0_6,
    n1
  );


  buf
  g2
  (
    n88,
    n9
  );


  not
  g3
  (
    n61,
    n11
  );


  not
  g4
  (
    n73,
    n1
  );


  buf
  g5
  (
    n27,
    n16
  );


  buf
  g6
  (
    KeyWire_0_19,
    n10
  );


  not
  g7
  (
    n23,
    n7
  );


  buf
  g8
  (
    n69,
    n9
  );


  not
  g9
  (
    n95,
    n3
  );


  not
  g10
  (
    n25,
    n2
  );


  not
  g11
  (
    n22,
    n8
  );


  not
  g12
  (
    n29,
    n11
  );


  buf
  g13
  (
    n91,
    n15
  );


  buf
  g14
  (
    n85,
    n19
  );


  buf
  g15
  (
    n47,
    n6
  );


  buf
  g16
  (
    n32,
    n8
  );


  not
  g17
  (
    n39,
    n13
  );


  not
  g18
  (
    n36,
    n11
  );


  not
  g19
  (
    n89,
    n19
  );


  not
  g20
  (
    n78,
    n8
  );


  not
  g21
  (
    n55,
    n19
  );


  buf
  g22
  (
    n60,
    n13
  );


  buf
  g23
  (
    n41,
    n18
  );


  buf
  g24
  (
    n96,
    n5
  );


  buf
  g25
  (
    n70,
    n10
  );


  buf
  g26
  (
    n72,
    n7
  );


  not
  g27
  (
    n24,
    n12
  );


  buf
  g28
  (
    n86,
    n4
  );


  buf
  g29
  (
    n74,
    n14
  );


  buf
  g30
  (
    n75,
    n12
  );


  not
  g31
  (
    n77,
    n6
  );


  buf
  g32
  (
    n57,
    n10
  );


  not
  g33
  (
    n43,
    n11
  );


  buf
  g34
  (
    n71,
    n15
  );


  buf
  g35
  (
    n54,
    n10
  );


  buf
  g36
  (
    n53,
    n7
  );


  buf
  g37
  (
    n48,
    n5
  );


  not
  g38
  (
    n44,
    n1
  );


  buf
  g39
  (
    n40,
    n17
  );


  buf
  g40
  (
    n58,
    n4
  );


  buf
  g41
  (
    n67,
    n2
  );


  buf
  g42
  (
    n63,
    n9
  );


  buf
  g43
  (
    n81,
    n17
  );


  not
  g44
  (
    n82,
    n14
  );


  buf
  g45
  (
    n76,
    n2
  );


  not
  g46
  (
    n90,
    n12
  );


  buf
  g47
  (
    n34,
    n6
  );


  not
  g48
  (
    n26,
    n17
  );


  not
  g49
  (
    n31,
    n15
  );


  buf
  g50
  (
    n84,
    n18
  );


  not
  g51
  (
    n62,
    n14
  );


  not
  g52
  (
    n51,
    n16
  );


  buf
  g53
  (
    n94,
    n13
  );


  not
  g54
  (
    n56,
    n5
  );


  buf
  g55
  (
    n59,
    n8
  );


  buf
  g56
  (
    n79,
    n12
  );


  not
  g57
  (
    n80,
    n3
  );


  buf
  g58
  (
    n35,
    n13
  );


  buf
  g59
  (
    n52,
    n18
  );


  not
  g60
  (
    n92,
    n4
  );


  not
  g61
  (
    n50,
    n16
  );


  not
  g62
  (
    n65,
    n3
  );


  not
  g63
  (
    n87,
    n6
  );


  not
  g64
  (
    n37,
    n4
  );


  not
  g65
  (
    n49,
    n17
  );


  not
  g66
  (
    n30,
    n9
  );


  not
  g67
  (
    n45,
    n14
  );


  buf
  g68
  (
    n66,
    n2
  );


  buf
  g69
  (
    n93,
    n18
  );


  buf
  g70
  (
    n38,
    n1
  );


  buf
  g71
  (
    n68,
    n3
  );


  not
  g72
  (
    n42,
    n7
  );


  buf
  g73
  (
    n64,
    n16
  );


  buf
  g74
  (
    n46,
    n5
  );


  not
  g75
  (
    n314,
    n34
  );


  buf
  g76
  (
    n174,
    n54
  );


  buf
  g77
  (
    n225,
    n62
  );


  buf
  g78
  (
    n210,
    n76
  );


  buf
  g79
  (
    n132,
    n73
  );


  not
  g80
  (
    n187,
    n50
  );


  buf
  g81
  (
    n195,
    n89
  );


  buf
  g82
  (
    n276,
    n76
  );


  not
  g83
  (
    n136,
    n58
  );


  not
  g84
  (
    n113,
    n80
  );


  not
  g85
  (
    n162,
    n27
  );


  not
  g86
  (
    n232,
    n85
  );


  buf
  g87
  (
    n266,
    n29
  );


  buf
  g88
  (
    n101,
    n45
  );


  not
  g89
  (
    n285,
    n28
  );


  buf
  g90
  (
    n161,
    n88
  );


  buf
  g91
  (
    n298,
    n38
  );


  buf
  g92
  (
    n323,
    n27
  );


  buf
  g93
  (
    n197,
    n28
  );


  buf
  g94
  (
    n228,
    n70
  );


  not
  g95
  (
    n190,
    n30
  );


  not
  g96
  (
    n185,
    n80
  );


  buf
  g97
  (
    n203,
    n47
  );


  buf
  g98
  (
    n299,
    n77
  );


  not
  g99
  (
    n194,
    n34
  );


  buf
  g100
  (
    n319,
    n79
  );


  buf
  g101
  (
    n175,
    n56
  );


  not
  g102
  (
    n144,
    n43
  );


  not
  g103
  (
    n109,
    n44
  );


  not
  g104
  (
    n155,
    n55
  );


  buf
  g105
  (
    n215,
    n54
  );


  not
  g106
  (
    n333,
    n36
  );


  buf
  g107
  (
    n240,
    n51
  );


  not
  g108
  (
    n116,
    n82
  );


  buf
  g109
  (
    n158,
    n82
  );


  not
  g110
  (
    n335,
    n47
  );


  not
  g111
  (
    n224,
    n25
  );


  buf
  g112
  (
    n238,
    n86
  );


  not
  g113
  (
    n310,
    n83
  );


  buf
  g114
  (
    n153,
    n32
  );


  not
  g115
  (
    n184,
    n59
  );


  buf
  g116
  (
    n246,
    n78
  );


  buf
  g117
  (
    n294,
    n31
  );


  not
  g118
  (
    n181,
    n41
  );


  not
  g119
  (
    n111,
    n54
  );


  not
  g120
  (
    n98,
    n29
  );


  not
  g121
  (
    n103,
    n75
  );


  buf
  g122
  (
    n318,
    n36
  );


  not
  g123
  (
    n202,
    n74
  );


  buf
  g124
  (
    n163,
    n69
  );


  not
  g125
  (
    n325,
    n83
  );


  buf
  g126
  (
    n239,
    n52
  );


  buf
  g127
  (
    n313,
    n55
  );


  not
  g128
  (
    n262,
    n76
  );


  buf
  g129
  (
    n105,
    n84
  );


  buf
  g130
  (
    n265,
    n65
  );


  buf
  g131
  (
    n193,
    n29
  );


  not
  g132
  (
    n229,
    n81
  );


  not
  g133
  (
    n307,
    n31
  );


  not
  g134
  (
    n251,
    n35
  );


  not
  g135
  (
    KeyWire_0_11,
    n88
  );


  not
  g136
  (
    n221,
    n61
  );


  not
  g137
  (
    n334,
    n68
  );


  buf
  g138
  (
    n283,
    n66
  );


  not
  g139
  (
    n315,
    n74
  );


  buf
  g140
  (
    n237,
    n40
  );


  buf
  g141
  (
    n308,
    n64
  );


  not
  g142
  (
    n254,
    n74
  );


  buf
  g143
  (
    n128,
    n43
  );


  buf
  g144
  (
    n167,
    n67
  );


  not
  g145
  (
    KeyWire_0_23,
    n56
  );


  buf
  g146
  (
    n118,
    n61
  );


  not
  g147
  (
    n189,
    n37
  );


  not
  g148
  (
    n258,
    n57
  );


  buf
  g149
  (
    n231,
    n57
  );


  buf
  g150
  (
    n134,
    n87
  );


  not
  g151
  (
    n164,
    n28
  );


  buf
  g152
  (
    n279,
    n67
  );


  buf
  g153
  (
    n226,
    n48
  );


  not
  g154
  (
    n133,
    n22
  );


  buf
  g155
  (
    n168,
    n37
  );


  buf
  g156
  (
    KeyWire_0_14,
    n24
  );


  buf
  g157
  (
    n198,
    n75
  );


  not
  g158
  (
    n119,
    n44
  );


  not
  g159
  (
    n250,
    n84
  );


  not
  g160
  (
    n110,
    n56
  );


  not
  g161
  (
    n192,
    n69
  );


  buf
  g162
  (
    n263,
    n70
  );


  not
  g163
  (
    n150,
    n62
  );


  buf
  g164
  (
    n270,
    n41
  );


  buf
  g165
  (
    n145,
    n72
  );


  buf
  g166
  (
    n141,
    n72
  );


  buf
  g167
  (
    n274,
    n46
  );


  buf
  g168
  (
    n146,
    n50
  );


  not
  g169
  (
    n303,
    n59
  );


  not
  g170
  (
    n324,
    n63
  );


  buf
  g171
  (
    n252,
    n71
  );


  not
  g172
  (
    KeyWire_0_16,
    n57
  );


  buf
  g173
  (
    n205,
    n31
  );


  buf
  g174
  (
    n234,
    n69
  );


  not
  g175
  (
    n320,
    n60
  );


  not
  g176
  (
    n242,
    n41
  );


  not
  g177
  (
    n269,
    n30
  );


  not
  g178
  (
    n166,
    n64
  );


  buf
  g179
  (
    n121,
    n65
  );


  not
  g180
  (
    n165,
    n87
  );


  buf
  g181
  (
    n117,
    n86
  );


  not
  g182
  (
    n309,
    n63
  );


  buf
  g183
  (
    n329,
    n26
  );


  buf
  g184
  (
    n212,
    n38
  );


  buf
  g185
  (
    n209,
    n71
  );


  buf
  g186
  (
    n100,
    n23
  );


  not
  g187
  (
    n312,
    n58
  );


  buf
  g188
  (
    n247,
    n57
  );


  not
  g189
  (
    n173,
    n47
  );


  buf
  g190
  (
    n301,
    n51
  );


  buf
  g191
  (
    n260,
    n52
  );


  not
  g192
  (
    n122,
    n79
  );


  buf
  g193
  (
    n152,
    n50
  );


  buf
  g194
  (
    n326,
    n68
  );


  buf
  g195
  (
    n142,
    n43
  );


  not
  g196
  (
    n330,
    n73
  );


  not
  g197
  (
    n104,
    n39
  );


  not
  g198
  (
    n275,
    n58
  );


  buf
  g199
  (
    n256,
    n50
  );


  not
  g200
  (
    n139,
    n49
  );


  not
  g201
  (
    n183,
    n84
  );


  buf
  g202
  (
    n179,
    n29
  );


  buf
  g203
  (
    n293,
    n61
  );


  not
  g204
  (
    n147,
    n34
  );


  not
  g205
  (
    n340,
    n67
  );


  not
  g206
  (
    n255,
    n30
  );


  buf
  g207
  (
    n259,
    n53
  );


  not
  g208
  (
    n126,
    n39
  );


  buf
  g209
  (
    n223,
    n43
  );


  not
  g210
  (
    n108,
    n79
  );


  not
  g211
  (
    n114,
    n35
  );


  not
  g212
  (
    n268,
    n49
  );


  buf
  g213
  (
    KeyWire_0_18,
    n35
  );


  buf
  g214
  (
    n339,
    n47
  );


  not
  g215
  (
    n159,
    n38
  );


  buf
  g216
  (
    n273,
    n80
  );


  not
  g217
  (
    n154,
    n60
  );


  not
  g218
  (
    n218,
    n87
  );


  not
  g219
  (
    KeyWire_0_27,
    n42
  );


  buf
  g220
  (
    n213,
    n83
  );


  not
  g221
  (
    n135,
    n26
  );


  buf
  g222
  (
    n115,
    n77
  );


  buf
  g223
  (
    n148,
    n89
  );


  buf
  g224
  (
    n287,
    n30
  );


  buf
  g225
  (
    n151,
    n71
  );


  buf
  g226
  (
    n180,
    n64
  );


  not
  g227
  (
    n149,
    n66
  );


  buf
  g228
  (
    n337,
    n41
  );


  not
  g229
  (
    n143,
    n75
  );


  not
  g230
  (
    n284,
    n81
  );


  buf
  g231
  (
    n176,
    n34
  );


  buf
  g232
  (
    n156,
    n82
  );


  not
  g233
  (
    n343,
    n64
  );


  not
  g234
  (
    n131,
    n51
  );


  not
  g235
  (
    n206,
    n65
  );


  buf
  g236
  (
    n169,
    n66
  );


  not
  g237
  (
    n196,
    n75
  );


  buf
  g238
  (
    n140,
    n25
  );


  buf
  g239
  (
    n130,
    n89
  );


  not
  g240
  (
    n177,
    n48
  );


  buf
  g241
  (
    n278,
    n81
  );


  buf
  g242
  (
    n137,
    n73
  );


  not
  g243
  (
    n248,
    n87
  );


  buf
  g244
  (
    n305,
    n74
  );


  buf
  g245
  (
    n297,
    n36
  );


  not
  g246
  (
    n342,
    n83
  );


  buf
  g247
  (
    n97,
    n82
  );


  not
  g248
  (
    n188,
    n76
  );


  not
  g249
  (
    n244,
    n56
  );


  not
  g250
  (
    n295,
    n42
  );


  not
  g251
  (
    n316,
    n45
  );


  not
  g252
  (
    n331,
    n88
  );


  buf
  g253
  (
    n200,
    n52
  );


  not
  g254
  (
    n160,
    n69
  );


  buf
  g255
  (
    n280,
    n23
  );


  buf
  g256
  (
    n272,
    n49
  );


  not
  g257
  (
    n328,
    n77
  );


  not
  g258
  (
    n300,
    n86
  );


  buf
  g259
  (
    n220,
    n46
  );


  not
  g260
  (
    n230,
    n31
  );


  buf
  g261
  (
    n282,
    n85
  );


  not
  g262
  (
    n171,
    n37
  );


  not
  g263
  (
    n204,
    n45
  );


  not
  g264
  (
    n292,
    n33
  );


  buf
  g265
  (
    n107,
    n48
  );


  not
  g266
  (
    n243,
    n60
  );


  buf
  g267
  (
    n214,
    n52
  );


  not
  g268
  (
    n302,
    n62
  );


  not
  g269
  (
    n341,
    n89
  );


  buf
  g270
  (
    n261,
    n85
  );


  not
  g271
  (
    n127,
    n62
  );


  not
  g272
  (
    n112,
    n55
  );


  not
  g273
  (
    n306,
    n72
  );


  buf
  g274
  (
    n102,
    n53
  );


  not
  g275
  (
    n120,
    n33
  );


  not
  g276
  (
    n201,
    n48
  );


  buf
  g277
  (
    n321,
    n58
  );


  buf
  g278
  (
    n277,
    n70
  );


  buf
  g279
  (
    n235,
    n65
  );


  buf
  g280
  (
    n327,
    n53
  );


  buf
  g281
  (
    n317,
    n68
  );


  not
  g282
  (
    n216,
    n40
  );


  buf
  g283
  (
    n172,
    n39
  );


  buf
  g284
  (
    KeyWire_0_26,
    n70
  );


  not
  g285
  (
    n191,
    n63
  );


  not
  g286
  (
    KeyWire_0_31,
    n44
  );


  not
  g287
  (
    n99,
    n37
  );


  buf
  g288
  (
    n322,
    n85
  );


  not
  g289
  (
    n182,
    n78
  );


  not
  g290
  (
    n124,
    n35
  );


  not
  g291
  (
    n222,
    n28
  );


  not
  g292
  (
    n288,
    n24
  );


  not
  g293
  (
    n249,
    n60
  );


  not
  g294
  (
    n253,
    n88
  );


  buf
  g295
  (
    n336,
    n46
  );


  not
  g296
  (
    n227,
    n33
  );


  buf
  g297
  (
    n286,
    n81
  );


  not
  g298
  (
    n233,
    n45
  );


  not
  g299
  (
    n123,
    n78
  );


  not
  g300
  (
    n311,
    n38
  );


  buf
  g301
  (
    n106,
    n72
  );


  not
  g302
  (
    n291,
    n84
  );


  buf
  g303
  (
    n217,
    n63
  );


  not
  g304
  (
    n219,
    n55
  );


  not
  g305
  (
    n271,
    n44
  );


  buf
  g306
  (
    n186,
    n54
  );


  not
  g307
  (
    n267,
    n59
  );


  buf
  g308
  (
    n199,
    n46
  );


  not
  g309
  (
    n170,
    n33
  );


  buf
  g310
  (
    n264,
    n61
  );


  buf
  g311
  (
    n129,
    n32
  );


  buf
  g312
  (
    n208,
    n22
  );


  buf
  g313
  (
    n290,
    n73
  );


  not
  g314
  (
    n207,
    n67
  );


  not
  g315
  (
    n338,
    n79
  );


  buf
  g316
  (
    n304,
    n78
  );


  not
  g317
  (
    n257,
    n77
  );


  buf
  g318
  (
    n211,
    n86
  );


  xor
  g319
  (
    n138,
    n66,
    n59,
    n51,
    n40
  );


  nor
  g320
  (
    n241,
    n68,
    n71,
    n80,
    n42
  );


  nand
  g321
  (
    n332,
    n49,
    n42,
    n40,
    n32
  );


  xnor
  g322
  (
    n296,
    n32,
    n53,
    n36,
    n39
  );


  nor
  g323
  (
    n398,
    n148,
    n220,
    n289,
    n173
  );


  nor
  g324
  (
    n349,
    n237,
    n157,
    n281,
    n211
  );


  xor
  g325
  (
    n387,
    n215,
    n20,
    n194,
    n231
  );


  nand
  g326
  (
    n361,
    n299,
    n306,
    n122,
    n201
  );


  nor
  g327
  (
    n393,
    n310,
    n171,
    n240,
    n169
  );


  or
  g328
  (
    n382,
    n307,
    n185,
    n142,
    n241
  );


  or
  g329
  (
    n375,
    n101,
    n236,
    n188,
    n219
  );


  nand
  g330
  (
    n372,
    n164,
    n167,
    n116,
    n223
  );


  nand
  g331
  (
    n383,
    n277,
    n229,
    n301,
    n121
  );


  nand
  g332
  (
    n359,
    n295,
    n276,
    n257,
    n153
  );


  or
  g333
  (
    n391,
    n292,
    n120,
    n177,
    n224
  );


  and
  g334
  (
    n351,
    n287,
    n114,
    n228,
    n245
  );


  xnor
  g335
  (
    n370,
    n19,
    n104,
    n181,
    n258
  );


  nand
  g336
  (
    n397,
    n172,
    n217,
    n238,
    n191
  );


  xnor
  g337
  (
    n380,
    n165,
    n105,
    n242,
    n274
  );


  nand
  g338
  (
    n368,
    n260,
    n108,
    n226,
    n133
  );


  and
  g339
  (
    n388,
    n145,
    n197,
    n192,
    n244
  );


  xor
  g340
  (
    n399,
    n221,
    n235,
    n267,
    n204
  );


  nand
  g341
  (
    n350,
    n202,
    n168,
    n162,
    n302
  );


  nor
  g342
  (
    n371,
    n175,
    n268,
    n225,
    n273
  );


  nand
  g343
  (
    n377,
    n113,
    n152,
    n198,
    n271
  );


  nand
  g344
  (
    n374,
    n111,
    n283,
    n186,
    n174
  );


  or
  g345
  (
    n355,
    n20,
    n208,
    n146,
    n115
  );


  or
  g346
  (
    n354,
    n130,
    n117,
    n139,
    n239
  );


  or
  g347
  (
    n353,
    n259,
    n147,
    n161,
    n183
  );


  or
  g348
  (
    n348,
    n97,
    n288,
    n230,
    n280
  );


  or
  g349
  (
    n386,
    n232,
    n207,
    n166,
    n286
  );


  xor
  g350
  (
    n362,
    n284,
    n123,
    n218,
    n250
  );


  nand
  g351
  (
    n392,
    n137,
    n243,
    n227,
    n21
  );


  or
  g352
  (
    n345,
    n265,
    n159,
    n189,
    n216
  );


  nor
  g353
  (
    n395,
    n107,
    n135,
    n21,
    n170
  );


  nor
  g354
  (
    n363,
    n253,
    n300,
    n119,
    n297
  );


  nand
  g355
  (
    n352,
    n263,
    n141,
    n213,
    n149
  );


  xor
  g356
  (
    n385,
    n180,
    n196,
    n247,
    n200
  );


  nand
  g357
  (
    n347,
    n126,
    n210,
    n151,
    n282
  );


  or
  g358
  (
    n390,
    n234,
    n291,
    n251,
    n193
  );


  or
  g359
  (
    n389,
    n311,
    n304,
    n278,
    n285
  );


  xnor
  g360
  (
    n369,
    n182,
    n118,
    n270,
    n296
  );


  xnor
  g361
  (
    n364,
    n261,
    n233,
    n248,
    n127
  );


  and
  g362
  (
    n360,
    n294,
    n195,
    n184,
    n214
  );


  nand
  g363
  (
    n384,
    n102,
    n178,
    n99,
    n179
  );


  and
  g364
  (
    n358,
    n144,
    n190,
    n138,
    n106
  );


  or
  g365
  (
    n378,
    n110,
    n103,
    n112,
    n212
  );


  nand
  g366
  (
    n365,
    n209,
    n21,
    n269,
    n132
  );


  xor
  g367
  (
    n367,
    n303,
    n205,
    n131,
    n21
  );


  and
  g368
  (
    n394,
    n155,
    n143,
    n279,
    n203
  );


  and
  g369
  (
    n376,
    n252,
    n124,
    n187,
    n128
  );


  or
  g370
  (
    n381,
    n199,
    n98,
    n256,
    n255
  );


  and
  g371
  (
    n373,
    n298,
    n266,
    n129,
    n160
  );


  or
  g372
  (
    n379,
    n254,
    n20,
    n308,
    n305
  );


  xor
  g373
  (
    n396,
    n154,
    n264,
    n158,
    n100
  );


  nor
  g374
  (
    n366,
    n206,
    n262,
    n150,
    n125
  );


  or
  g375
  (
    n400,
    n272,
    n249,
    n109,
    n290
  );


  nor
  g376
  (
    n346,
    n275,
    n140,
    n176,
    n20
  );


  nor
  g377
  (
    n357,
    n293,
    n134,
    n222,
    n163
  );


  and
  g378
  (
    n356,
    n156,
    n136,
    n309,
    n246
  );


  buf
  g379
  (
    n404,
    n372
  );


  buf
  g380
  (
    n403,
    n360
  );


  not
  g381
  (
    n406,
    n350
  );


  buf
  g382
  (
    KeyWire_0_13,
    n363
  );


  not
  g383
  (
    n405,
    n357
  );


  not
  g384
  (
    n415,
    n349
  );


  buf
  g385
  (
    n401,
    n347
  );


  buf
  g386
  (
    n408,
    n90
  );


  buf
  g387
  (
    n417,
    n355
  );


  buf
  g388
  (
    n409,
    n354
  );


  buf
  g389
  (
    n412,
    n345
  );


  buf
  g390
  (
    n410,
    n367
  );


  xor
  g391
  (
    n413,
    n348,
    n362,
    n358,
    n365
  );


  xor
  g392
  (
    n411,
    n90,
    n90,
    n353,
    n359
  );


  xor
  g393
  (
    n407,
    n370,
    n366,
    n352,
    n361
  );


  nor
  g394
  (
    n414,
    n346,
    n368,
    n90,
    n351
  );


  xor
  g395
  (
    n402,
    n371,
    n369,
    n356,
    n364
  );


  not
  g396
  (
    n430,
    n318
  );


  not
  g397
  (
    n429,
    n93
  );


  or
  g398
  (
    n424,
    n324,
    n91
  );


  and
  g399
  (
    n420,
    n92,
    n401,
    n414,
    n410
  );


  nor
  g400
  (
    n422,
    n321,
    n404,
    n406,
    n91
  );


  or
  g401
  (
    n428,
    n92,
    n325,
    n327,
    n93
  );


  nand
  g402
  (
    n419,
    n94,
    n416,
    n412,
    n314
  );


  nand
  g403
  (
    n421,
    n409,
    n402,
    n91,
    n94
  );


  or
  g404
  (
    n427,
    n96,
    n320,
    n403,
    n95
  );


  nor
  g405
  (
    n426,
    n91,
    n319,
    n405,
    n93
  );


  xnor
  g406
  (
    n423,
    n323,
    n92,
    n95,
    n313
  );


  xnor
  g407
  (
    n418,
    n92,
    n315,
    n93,
    n408
  );


  nor
  g408
  (
    n431,
    n411,
    n94,
    n415,
    n326
  );


  and
  g409
  (
    n433,
    n95,
    n407,
    n96
  );


  or
  g410
  (
    n432,
    n413,
    n317,
    n322,
    n316
  );


  xor
  g411
  (
    n425,
    n94,
    n95,
    n96,
    n312
  );


  not
  g412
  (
    n489,
    n426
  );


  buf
  g413
  (
    n485,
    n423
  );


  buf
  g414
  (
    n475,
    n422
  );


  buf
  g415
  (
    n477,
    n430
  );


  buf
  g416
  (
    n470,
    n431
  );


  buf
  g417
  (
    n480,
    n422
  );


  buf
  g418
  (
    n454,
    n374
  );


  not
  g419
  (
    n436,
    n427
  );


  not
  g420
  (
    n441,
    n423
  );


  not
  g421
  (
    n478,
    n419
  );


  buf
  g422
  (
    n490,
    n427
  );


  buf
  g423
  (
    n450,
    n420
  );


  buf
  g424
  (
    n443,
    n419
  );


  not
  g425
  (
    n474,
    n421
  );


  not
  g426
  (
    n471,
    n429
  );


  buf
  g427
  (
    n469,
    n418
  );


  buf
  g428
  (
    n465,
    n425
  );


  buf
  g429
  (
    n444,
    n420
  );


  not
  g430
  (
    n440,
    n425
  );


  not
  g431
  (
    n484,
    n418
  );


  buf
  g432
  (
    n488,
    n424
  );


  buf
  g433
  (
    n479,
    n421
  );


  buf
  g434
  (
    n461,
    n418
  );


  buf
  g435
  (
    n456,
    n420
  );


  buf
  g436
  (
    n448,
    n376
  );


  not
  g437
  (
    n437,
    n426
  );


  buf
  g438
  (
    n439,
    n426
  );


  not
  g439
  (
    n468,
    n422
  );


  buf
  g440
  (
    KeyWire_0_2,
    n429
  );


  buf
  g441
  (
    n457,
    n424
  );


  buf
  g442
  (
    n449,
    n378
  );


  buf
  g443
  (
    n452,
    n377
  );


  buf
  g444
  (
    n473,
    n431
  );


  buf
  g445
  (
    n486,
    n428
  );


  not
  g446
  (
    n434,
    n431
  );


  buf
  g447
  (
    n438,
    n428
  );


  buf
  g448
  (
    n451,
    n430
  );


  buf
  g449
  (
    n482,
    n424
  );


  not
  g450
  (
    n472,
    n431
  );


  buf
  g451
  (
    n447,
    n430
  );


  buf
  g452
  (
    n435,
    n421
  );


  buf
  g453
  (
    n442,
    n422
  );


  not
  g454
  (
    n464,
    n429
  );


  not
  g455
  (
    n467,
    n432
  );


  buf
  g456
  (
    n476,
    n430
  );


  not
  g457
  (
    n462,
    n373
  );


  not
  g458
  (
    n453,
    n425
  );


  buf
  g459
  (
    n455,
    n424
  );


  not
  g460
  (
    n445,
    n421
  );


  buf
  g461
  (
    n466,
    n420
  );


  not
  g462
  (
    n459,
    n427
  );


  not
  g463
  (
    n458,
    n375
  );


  not
  g464
  (
    n487,
    n428
  );


  and
  g465
  (
    KeyWire_0_7,
    n423,
    n425
  );


  or
  g466
  (
    n481,
    n427,
    n419
  );


  nor
  g467
  (
    n446,
    n428,
    n429
  );


  or
  g468
  (
    n483,
    n426,
    n418,
    n423,
    n419
  );


  not
  g469
  (
    n513,
    n436
  );


  buf
  g470
  (
    n511,
    n434
  );


  buf
  g471
  (
    n509,
    n440
  );


  buf
  g472
  (
    n514,
    n438
  );


  buf
  g473
  (
    n517,
    n437
  );


  not
  g474
  (
    n499,
    n437
  );


  not
  g475
  (
    n494,
    n439
  );


  buf
  g476
  (
    n498,
    n438
  );


  not
  g477
  (
    n510,
    n381
  );


  buf
  g478
  (
    n502,
    n439
  );


  not
  g479
  (
    n497,
    n435
  );


  not
  g480
  (
    n506,
    n441
  );


  buf
  g481
  (
    n508,
    n382
  );


  buf
  g482
  (
    n515,
    n439
  );


  buf
  g483
  (
    n500,
    n436
  );


  not
  g484
  (
    n491,
    n434
  );


  not
  g485
  (
    n493,
    n380
  );


  buf
  g486
  (
    n504,
    n435
  );


  buf
  g487
  (
    n512,
    n383
  );


  buf
  g488
  (
    n505,
    n438
  );


  not
  g489
  (
    n503,
    n441
  );


  not
  g490
  (
    n495,
    n440
  );


  not
  g491
  (
    n492,
    n439
  );


  not
  g492
  (
    KeyWire_0_24,
    n437
  );


  not
  g493
  (
    n516,
    n436
  );


  nor
  g494
  (
    n496,
    n436,
    n440
  );


  xnor
  g495
  (
    n507,
    n437,
    n441,
    n438,
    n379
  );


  buf
  g496
  (
    n519,
    n495
  );


  buf
  g497
  (
    n525,
    n493
  );


  buf
  g498
  (
    n532,
    n492
  );


  buf
  g499
  (
    n526,
    n492
  );


  not
  g500
  (
    n531,
    n494
  );


  buf
  g501
  (
    n528,
    n495
  );


  buf
  g502
  (
    n520,
    n494
  );


  buf
  g503
  (
    n521,
    n417
  );


  not
  g504
  (
    n529,
    n495
  );


  buf
  g505
  (
    n523,
    n494
  );


  not
  g506
  (
    n518,
    n492
  );


  buf
  g507
  (
    n522,
    n493
  );


  not
  g508
  (
    n533,
    n491
  );


  buf
  g509
  (
    n524,
    n491
  );


  buf
  g510
  (
    n527,
    n492
  );


  buf
  g511
  (
    KeyWire_0_3,
    n493
  );


  or
  g512
  (
    n530,
    n494,
    n493
  );


  or
  g513
  (
    n544,
    n531,
    n433,
    n451
  );


  nand
  g514
  (
    n551,
    n453,
    n445,
    n529
  );


  or
  g515
  (
    n541,
    n443,
    n432,
    n523,
    n518
  );


  or
  g516
  (
    n539,
    n433,
    n443,
    n445,
    n446
  );


  and
  g517
  (
    n547,
    n520,
    n445,
    n528,
    n443
  );


  and
  g518
  (
    n535,
    n446,
    n450,
    n447,
    n525
  );


  xor
  g519
  (
    n549,
    n447,
    n452,
    n433,
    n441
  );


  nor
  g520
  (
    n538,
    n526,
    n450,
    n449,
    n442
  );


  nor
  g521
  (
    n546,
    n524,
    n442,
    n533,
    n453
  );


  and
  g522
  (
    n542,
    n450,
    n447,
    n446,
    n522
  );


  xnor
  g523
  (
    KeyWire_0_12,
    n527,
    n446,
    n534,
    n449
  );


  nor
  g524
  (
    n550,
    n448,
    n442,
    n452,
    n444
  );


  xnor
  g525
  (
    n548,
    n444,
    n534,
    n451,
    n452
  );


  nand
  g526
  (
    KeyWire_0_0,
    n443,
    n444,
    n448,
    n452
  );


  nand
  g527
  (
    n537,
    n449,
    n521,
    n432,
    n448
  );


  nand
  g528
  (
    n543,
    n442,
    n532,
    n444,
    n451
  );


  xnor
  g529
  (
    n545,
    n432,
    n448,
    n530,
    n453
  );


  or
  g530
  (
    n540,
    n450,
    n519,
    n449,
    n447
  );


  xnor
  g531
  (
    n563,
    n461,
    n465,
    n502,
    n547
  );


  and
  g532
  (
    n564,
    n547,
    n501,
    n476,
    n488
  );


  xor
  g533
  (
    n583,
    n474,
    n498,
    n487,
    n536
  );


  xnor
  g534
  (
    n606,
    n539,
    n471,
    n470,
    n466
  );


  nor
  g535
  (
    n562,
    n501,
    n550,
    n467,
    n500
  );


  and
  g536
  (
    n565,
    n542,
    n470,
    n549,
    n468
  );


  and
  g537
  (
    n582,
    n501,
    n488,
    n480,
    n546
  );


  or
  g538
  (
    n610,
    n458,
    n495,
    n487,
    n546
  );


  or
  g539
  (
    n574,
    n501,
    n540,
    n542,
    n502
  );


  nor
  g540
  (
    n560,
    n540,
    n481,
    n461,
    n545
  );


  and
  g541
  (
    KeyWire_0_21,
    n476,
    n477,
    n463,
    n458
  );


  nand
  g542
  (
    n601,
    n478,
    n543,
    n467,
    n474
  );


  or
  g543
  (
    n586,
    n486,
    n459,
    n535,
    n476
  );


  and
  g544
  (
    n557,
    n482,
    n460,
    n475,
    n465
  );


  nand
  g545
  (
    KeyWire_0_29,
    n458,
    n483,
    n478
  );


  nor
  g546
  (
    n608,
    n459,
    n503,
    n486,
    n499
  );


  nand
  g547
  (
    n568,
    n504,
    n475,
    n482,
    n544
  );


  nand
  g548
  (
    n592,
    n474,
    n546,
    n548,
    n455
  );


  nand
  g549
  (
    n587,
    n469,
    n473,
    n455,
    n483
  );


  and
  g550
  (
    n578,
    n488,
    n473,
    n543,
    n468
  );


  or
  g551
  (
    n599,
    n477,
    n484,
    n462,
    n453
  );


  nor
  g552
  (
    n554,
    n464,
    n485,
    n470,
    n478
  );


  nand
  g553
  (
    n593,
    n502,
    n471,
    n485,
    n538
  );


  nand
  g554
  (
    n604,
    n504,
    n462,
    n479,
    n457
  );


  nor
  g555
  (
    n588,
    n539,
    n541,
    n547,
    n468
  );


  and
  g556
  (
    n584,
    n504,
    n549,
    n539,
    n497
  );


  or
  g557
  (
    n571,
    n484,
    n464,
    n465,
    n474
  );


  or
  g558
  (
    n556,
    n497,
    n500,
    n460,
    n498
  );


  nand
  g559
  (
    n573,
    n503,
    n460,
    n481,
    n470
  );


  xnor
  g560
  (
    n569,
    n466,
    n484,
    n487,
    n467
  );


  and
  g561
  (
    KeyWire_0_30,
    n542,
    n469,
    n496
  );


  xnor
  g562
  (
    n600,
    n460,
    n455,
    n486,
    n483
  );


  nand
  g563
  (
    n579,
    n500,
    n543,
    n537,
    n497
  );


  nor
  g564
  (
    n581,
    n454,
    n538,
    n477,
    n482
  );


  nor
  g565
  (
    n555,
    n536,
    n548,
    n462,
    n472
  );


  nor
  g566
  (
    n570,
    n472,
    n546,
    n503,
    n457
  );


  or
  g567
  (
    n566,
    n463,
    n475,
    n464,
    n476
  );


  xor
  g568
  (
    n580,
    n504,
    n544,
    n542,
    n467
  );


  and
  g569
  (
    KeyWire_0_9,
    n539,
    n502,
    n536,
    n484
  );


  and
  g570
  (
    n596,
    n549,
    n479,
    n463,
    n544
  );


  or
  g571
  (
    n597,
    n548,
    n547,
    n540,
    n535
  );


  nand
  g572
  (
    n577,
    n498,
    n454,
    n545,
    n536
  );


  xnor
  g573
  (
    KeyWire_0_10,
    n541,
    n544,
    n497,
    n475
  );


  and
  g574
  (
    n567,
    n537,
    n471,
    n480,
    n473
  );


  and
  g575
  (
    n595,
    n463,
    n454,
    n496,
    n538
  );


  nor
  g576
  (
    n576,
    n454,
    n498,
    n485,
    n469
  );


  or
  g577
  (
    n559,
    n549,
    n479,
    n466,
    n500
  );


  and
  g578
  (
    n591,
    n459,
    n464,
    n481,
    n456
  );


  nand
  g579
  (
    n609,
    n543,
    n461,
    n499,
    n473
  );


  xnor
  g580
  (
    n598,
    n537,
    n459,
    n457,
    n541
  );


  xnor
  g581
  (
    n611,
    n545,
    n538,
    n481,
    n456
  );


  xor
  g582
  (
    n561,
    n478,
    n485,
    n462,
    n461
  );


  nand
  g583
  (
    n553,
    n472,
    n487,
    n496,
    n471
  );


  xnor
  g584
  (
    n585,
    n457,
    n480,
    n458,
    n472
  );


  nand
  g585
  (
    n572,
    n486,
    n456,
    n503,
    n465
  );


  and
  g586
  (
    n607,
    n466,
    n499,
    n456,
    n540
  );


  xnor
  g587
  (
    n558,
    n480,
    n455,
    n468,
    n499
  );


  nor
  g588
  (
    n589,
    n479,
    n545,
    n541,
    n548
  );


  xor
  g589
  (
    n603,
    n477,
    n537,
    n469,
    n482
  );


  buf
  g590
  (
    KeyWire_0_25,
    n505
  );


  buf
  g591
  (
    n617,
    n507
  );


  buf
  g592
  (
    n614,
    n557
  );


  not
  g593
  (
    n621,
    n556
  );


  not
  g594
  (
    n613,
    n507
  );


  not
  g595
  (
    n618,
    n554
  );


  buf
  g596
  (
    n623,
    n507
  );


  not
  g597
  (
    n619,
    n507
  );


  or
  g598
  (
    n612,
    n558,
    n506,
    n557,
    n505
  );


  or
  g599
  (
    n622,
    n555,
    n506,
    n559,
    n505
  );


  xor
  g600
  (
    n615,
    n553,
    n555,
    n559,
    n506
  );


  xor
  g601
  (
    n620,
    n556,
    n505,
    n558,
    n506
  );


  not
  g602
  (
    n647,
    n392
  );


  buf
  g603
  (
    n639,
    n620
  );


  not
  g604
  (
    n643,
    n619
  );


  not
  g605
  (
    n633,
    n384
  );


  not
  g606
  (
    n644,
    n616
  );


  buf
  g607
  (
    n626,
    n389
  );


  buf
  g608
  (
    n641,
    n612
  );


  not
  g609
  (
    n632,
    n612
  );


  not
  g610
  (
    n645,
    n614
  );


  not
  g611
  (
    n629,
    n617
  );


  not
  g612
  (
    n637,
    n621
  );


  not
  g613
  (
    n630,
    n621
  );


  buf
  g614
  (
    n638,
    n618
  );


  buf
  g615
  (
    n634,
    n621
  );


  not
  g616
  (
    n631,
    n391
  );


  not
  g617
  (
    n627,
    n615
  );


  buf
  g618
  (
    n642,
    n622
  );


  buf
  g619
  (
    n624,
    n613
  );


  not
  g620
  (
    n640,
    n388
  );


  buf
  g621
  (
    n625,
    n620
  );


  nor
  g622
  (
    n635,
    n613,
    n622
  );


  xnor
  g623
  (
    n628,
    n386,
    n616,
    n385,
    n393
  );


  xnor
  g624
  (
    n636,
    n387,
    n615,
    n617,
    n618
  );


  nor
  g625
  (
    n646,
    n614,
    n619,
    n621,
    n390
  );


  nand
  g626
  (
    n665,
    n625,
    n552,
    n561,
    n572
  );


  xnor
  g627
  (
    n669,
    n508,
    n581,
    n580,
    n509
  );


  and
  g628
  (
    n664,
    n509,
    n566,
    n395,
    n574
  );


  nor
  g629
  (
    n663,
    n626,
    n577,
    n576,
    n624
  );


  nor
  g630
  (
    n648,
    n510,
    n508,
    n551,
    n627
  );


  xor
  g631
  (
    n672,
    n394,
    n564,
    n561,
    n584
  );


  nand
  g632
  (
    n666,
    n625,
    n550,
    n576,
    n509
  );


  xnor
  g633
  (
    n670,
    n396,
    n579,
    n624,
    n573
  );


  nor
  g634
  (
    KeyWire_0_20,
    n628,
    n629,
    n568,
    n574
  );


  xnor
  g635
  (
    n660,
    n583,
    n562,
    n552,
    n575
  );


  or
  g636
  (
    n651,
    n585,
    n585,
    n575,
    n577
  );


  nor
  g637
  (
    n655,
    n582,
    n398,
    n560,
    n584
  );


  nor
  g638
  (
    n654,
    n509,
    n400,
    n569,
    n571
  );


  and
  g639
  (
    n661,
    n579,
    n628,
    n567,
    n510
  );


  xor
  g640
  (
    n652,
    n626,
    n563,
    n551,
    n630
  );


  nor
  g641
  (
    n673,
    n629,
    n580,
    n627,
    n624
  );


  or
  g642
  (
    n650,
    n550,
    n508,
    n628
  );


  xnor
  g643
  (
    n668,
    n582,
    n565,
    n572,
    n573
  );


  xor
  g644
  (
    n671,
    n551,
    n628,
    n586,
    n630
  );


  xnor
  g645
  (
    n656,
    n570,
    n578,
    n624,
    n625
  );


  nor
  g646
  (
    n658,
    n552,
    n578,
    n563,
    n550
  );


  or
  g647
  (
    n649,
    n560,
    n629,
    n569,
    n551
  );


  nor
  g648
  (
    n653,
    n571,
    n566,
    n565,
    n562
  );


  nand
  g649
  (
    n657,
    n625,
    n568,
    n570,
    n626
  );


  and
  g650
  (
    n667,
    n629,
    n567,
    n564,
    n397
  );


  nand
  g651
  (
    n662,
    n627,
    n399,
    n581,
    n552
  );


  xnor
  g652
  (
    n674,
    n583,
    n627,
    n626,
    n630
  );


  xnor
  g653
  (
    n689,
    n596,
    n659,
    n605,
    n660
  );


  or
  g654
  (
    n680,
    n662,
    n602,
    n586,
    n665
  );


  xor
  g655
  (
    n682,
    n610,
    n611,
    n600,
    n668
  );


  or
  g656
  (
    KeyWire_0_15,
    n664,
    n599,
    n593
  );


  xor
  g657
  (
    n684,
    n606,
    n597,
    n666,
    n607
  );


  or
  g658
  (
    n686,
    n667,
    n598,
    n673,
    n591
  );


  xnor
  g659
  (
    n685,
    n594,
    n588,
    n605
  );


  xor
  g660
  (
    n690,
    n604,
    n597,
    n601,
    n606
  );


  or
  g661
  (
    n691,
    n590,
    n604,
    n589,
    n603
  );


  nor
  g662
  (
    n681,
    n661,
    n599,
    n595,
    n670
  );


  nand
  g663
  (
    n679,
    n601,
    n663,
    n609,
    n600
  );


  and
  g664
  (
    n676,
    n592,
    n592,
    n669,
    n589
  );


  and
  g665
  (
    n675,
    n610,
    n591,
    n658,
    n608
  );


  xnor
  g666
  (
    n687,
    n608,
    n671,
    n603,
    n611
  );


  nor
  g667
  (
    n678,
    n609,
    n595,
    n587,
    n596
  );


  nand
  g668
  (
    n683,
    n607,
    n590,
    n594,
    n598
  );


  xor
  g669
  (
    n688,
    n602,
    n674,
    n587,
    n672
  );


  xnor
  g670
  (
    n735,
    n515,
    n690,
    n513,
    n639
  );


  xor
  g671
  (
    n719,
    n489,
    n512,
    n635,
    n647
  );


  or
  g672
  (
    KeyWire_0_1,
    n642,
    n687,
    n646,
    n637
  );


  and
  g673
  (
    n714,
    n513,
    n513,
    n636,
    n640
  );


  and
  g674
  (
    n726,
    n682,
    n514,
    n642,
    n340
  );


  xnor
  g675
  (
    n696,
    n640,
    n635,
    n623,
    n684
  );


  or
  g676
  (
    n708,
    n644,
    n515,
    n339,
    n334
  );


  xnor
  g677
  (
    n724,
    n490,
    n676,
    n516,
    n517
  );


  xor
  g678
  (
    n698,
    n329,
    n634,
    n623,
    n690
  );


  xor
  g679
  (
    n718,
    n517,
    n643,
    n641,
    n489
  );


  nor
  g680
  (
    n720,
    n622,
    n515,
    n335,
    n642
  );


  nor
  g681
  (
    n722,
    n512,
    n488,
    n631,
    n647
  );


  nand
  g682
  (
    n715,
    n632,
    n511,
    n644,
    n678
  );


  xor
  g683
  (
    n702,
    n639,
    n640,
    n685,
    n510
  );


  and
  g684
  (
    n734,
    n637,
    n639,
    n678,
    n644
  );


  xnor
  g685
  (
    n699,
    n643,
    n514,
    n684,
    n631
  );


  nand
  g686
  (
    n700,
    n646,
    n676,
    n517,
    n644
  );


  and
  g687
  (
    KeyWire_0_28,
    n689,
    n510,
    n682,
    n685
  );


  nor
  g688
  (
    n733,
    n635,
    n641,
    n638,
    n684
  );


  xor
  g689
  (
    n710,
    n681,
    n634,
    n632,
    n511
  );


  xor
  g690
  (
    n711,
    n633,
    n638,
    n516,
    n689
  );


  and
  g691
  (
    n707,
    n630,
    n638,
    n433,
    n343
  );


  xor
  g692
  (
    n727,
    n342,
    n336,
    n513,
    n681
  );


  and
  g693
  (
    n709,
    n632,
    n647,
    n634,
    n511
  );


  and
  g694
  (
    n695,
    n636,
    n633,
    n689,
    n517
  );


  xor
  g695
  (
    KeyWire_0_17,
    n512,
    n642,
    n687,
    n688
  );


  xnor
  g696
  (
    n701,
    n637,
    n631,
    n632,
    n677
  );


  or
  g697
  (
    n697,
    n641,
    n688,
    n634,
    n344
  );


  nand
  g698
  (
    n713,
    n685,
    n489,
    n516,
    n643
  );


  nand
  g699
  (
    n693,
    n639,
    n490,
    n675,
    n686
  );


  and
  g700
  (
    n716,
    n679,
    n635,
    n688,
    n330
  );


  and
  g701
  (
    n731,
    n623,
    n691,
    n328
  );


  xor
  g702
  (
    n705,
    n514,
    n633,
    n677,
    n643
  );


  nor
  g703
  (
    KeyWire_0_22,
    n337,
    n646,
    n333,
    n641
  );


  xnor
  g704
  (
    n704,
    n647,
    n515,
    n638,
    n623
  );


  nand
  g705
  (
    n706,
    n516,
    n691,
    n512,
    n511
  );


  and
  g706
  (
    n721,
    n686,
    n640,
    n680,
    n675
  );


  and
  g707
  (
    n729,
    n646,
    n680,
    n686,
    n683
  );


  or
  g708
  (
    KeyWire_0_5,
    n679,
    n490,
    n338,
    n622
  );


  xor
  g709
  (
    n703,
    n636,
    n690,
    n489,
    n645
  );


  nor
  g710
  (
    n728,
    n633,
    n645,
    n687,
    n341
  );


  xnor
  g711
  (
    n692,
    n490,
    n631,
    n682,
    n683
  );


  and
  g712
  (
    n723,
    n637,
    n332,
    n636,
    n683
  );


  or
  g713
  (
    n725,
    n331,
    n645,
    n514
  );


  nor
  g714
  (
    KeyWire_0_8,
    n693,
    n696,
    n692,
    n695
  );


  and
  g715
  (
    n739,
    n721,
    n723,
    n701,
    n709
  );


  nand
  g716
  (
    n738,
    n694,
    n727,
    n726,
    n699
  );


  nand
  g717
  (
    n745,
    n735,
    n730,
    n710,
    n717
  );


  xor
  g718
  (
    n740,
    n698,
    n702,
    n706,
    n713
  );


  nor
  g719
  (
    n746,
    n719,
    n708,
    n724,
    n700
  );


  xor
  g720
  (
    n741,
    n729,
    n722,
    n716,
    n715
  );


  xor
  g721
  (
    n742,
    n733,
    n703,
    n705,
    n720
  );


  nor
  g722
  (
    n736,
    n728,
    n732,
    n711,
    n734
  );


  xor
  g723
  (
    n737,
    n697,
    n707,
    n718,
    n712
  );


  and
  g724
  (
    KeyWire_0_4,
    n725,
    n714,
    n731,
    n704
  );


  xor
  KeyGate_0_0
  (
    n536,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n732,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n463,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n534,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n743,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n730,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n33,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n460,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n744,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n602,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n590,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n236,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n552,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n416,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n178,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n677,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n289,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n694,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n245,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n28,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n659,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n575,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n717,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n281,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n501,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n616,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n157,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n125,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n712,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n594,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n605,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n344,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

