

module Stat_2000_301
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1518,
  n1517,
  n1533,
  n2029,
  n2025,
  n2020,
  n2010,
  n2031,
  n2008,
  n2028,
  n2012,
  n2027,
  n2022,
  n2030,
  n2006,
  n2024,
  n2032,
  n2018,
  n2009,
  n2021,
  n2016,
  n2013,
  n2023,
  n2005,
  n2026,
  n2014,
  n2011,
  n2017,
  n2004,
  n2019,
  n2007,
  n2015,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1518;
  output n1517;
  output n1533;
  output n2029;
  output n2025;
  output n2020;
  output n2010;
  output n2031;
  output n2008;
  output n2028;
  output n2012;
  output n2027;
  output n2022;
  output n2030;
  output n2006;
  output n2024;
  output n2032;
  output n2018;
  output n2009;
  output n2021;
  output n2016;
  output n2013;
  output n2023;
  output n2005;
  output n2026;
  output n2014;
  output n2011;
  output n2017;
  output n2004;
  output n2019;
  output n2007;
  output n2015;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;

  not
  g0
  (
    n40,
    n13
  );


  buf
  g1
  (
    n93,
    n21
  );


  buf
  g2
  (
    n83,
    n29
  );


  not
  g3
  (
    n149,
    n8
  );


  not
  g4
  (
    n72,
    n19
  );


  buf
  g5
  (
    n122,
    n31
  );


  not
  g6
  (
    n45,
    n18
  );


  buf
  g7
  (
    n53,
    n23
  );


  not
  g8
  (
    n73,
    n7
  );


  not
  g9
  (
    n139,
    n25
  );


  not
  g10
  (
    n92,
    n32
  );


  buf
  g11
  (
    n87,
    n32
  );


  not
  g12
  (
    n39,
    n11
  );


  not
  g13
  (
    n127,
    n24
  );


  buf
  g14
  (
    n42,
    n11
  );


  buf
  g15
  (
    n134,
    n11
  );


  not
  g16
  (
    n84,
    n15
  );


  not
  g17
  (
    n154,
    n5
  );


  not
  g18
  (
    n75,
    n16
  );


  buf
  g19
  (
    n68,
    n30
  );


  not
  g20
  (
    n88,
    n25
  );


  buf
  g21
  (
    n47,
    n24
  );


  buf
  g22
  (
    n150,
    n12
  );


  not
  g23
  (
    n77,
    n27
  );


  not
  g24
  (
    n36,
    n14
  );


  not
  g25
  (
    n111,
    n3
  );


  buf
  g26
  (
    n58,
    n26
  );


  buf
  g27
  (
    n34,
    n28
  );


  not
  g28
  (
    n144,
    n10
  );


  buf
  g29
  (
    n74,
    n8
  );


  not
  g30
  (
    n104,
    n9
  );


  not
  g31
  (
    n56,
    n2
  );


  not
  g32
  (
    n138,
    n17
  );


  buf
  g33
  (
    n69,
    n6
  );


  not
  g34
  (
    n119,
    n12
  );


  not
  g35
  (
    n136,
    n11
  );


  not
  g36
  (
    n98,
    n31
  );


  not
  g37
  (
    n86,
    n18
  );


  not
  g38
  (
    n35,
    n7
  );


  buf
  g39
  (
    n116,
    n10
  );


  not
  g40
  (
    n153,
    n25
  );


  not
  g41
  (
    n157,
    n21
  );


  buf
  g42
  (
    n85,
    n31
  );


  buf
  g43
  (
    n79,
    n14
  );


  not
  g44
  (
    n33,
    n22
  );


  not
  g45
  (
    n102,
    n28
  );


  not
  g46
  (
    n126,
    n17
  );


  buf
  g47
  (
    n94,
    n27
  );


  buf
  g48
  (
    n140,
    n23
  );


  not
  g49
  (
    n62,
    n3
  );


  not
  g50
  (
    n135,
    n4
  );


  not
  g51
  (
    n55,
    n29
  );


  not
  g52
  (
    n115,
    n18
  );


  buf
  g53
  (
    n108,
    n30
  );


  buf
  g54
  (
    n142,
    n18
  );


  not
  g55
  (
    n123,
    n10
  );


  buf
  g56
  (
    n160,
    n15
  );


  not
  g57
  (
    n89,
    n5
  );


  not
  g58
  (
    n107,
    n26
  );


  not
  g59
  (
    n82,
    n6
  );


  not
  g60
  (
    n132,
    n22
  );


  not
  g61
  (
    n103,
    n2
  );


  not
  g62
  (
    n110,
    n29
  );


  buf
  g63
  (
    n51,
    n14
  );


  buf
  g64
  (
    n120,
    n5
  );


  not
  g65
  (
    n67,
    n20
  );


  buf
  g66
  (
    n97,
    n2
  );


  buf
  g67
  (
    n151,
    n10
  );


  not
  g68
  (
    n60,
    n1
  );


  buf
  g69
  (
    n129,
    n13
  );


  buf
  g70
  (
    n146,
    n7
  );


  buf
  g71
  (
    n99,
    n4
  );


  not
  g72
  (
    n143,
    n6
  );


  buf
  g73
  (
    n91,
    n16
  );


  not
  g74
  (
    n137,
    n27
  );


  not
  g75
  (
    n59,
    n15
  );


  buf
  g76
  (
    n121,
    n5
  );


  not
  g77
  (
    n96,
    n21
  );


  not
  g78
  (
    n61,
    n17
  );


  buf
  g79
  (
    n95,
    n23
  );


  not
  g80
  (
    n57,
    n16
  );


  buf
  g81
  (
    n156,
    n13
  );


  buf
  g82
  (
    n113,
    n26
  );


  buf
  g83
  (
    n125,
    n16
  );


  not
  g84
  (
    n90,
    n25
  );


  not
  g85
  (
    n128,
    n9
  );


  not
  g86
  (
    n152,
    n22
  );


  not
  g87
  (
    n105,
    n19
  );


  buf
  g88
  (
    n41,
    n13
  );


  not
  g89
  (
    n112,
    n23
  );


  buf
  g90
  (
    n117,
    n4
  );


  buf
  g91
  (
    n78,
    n1
  );


  not
  g92
  (
    n106,
    n6
  );


  not
  g93
  (
    n48,
    n28
  );


  not
  g94
  (
    n141,
    n31
  );


  buf
  g95
  (
    n64,
    n2
  );


  not
  g96
  (
    n46,
    n9
  );


  buf
  g97
  (
    n148,
    n1
  );


  buf
  g98
  (
    n101,
    n3
  );


  buf
  g99
  (
    n37,
    n20
  );


  not
  g100
  (
    n65,
    n19
  );


  not
  g101
  (
    n70,
    n7
  );


  not
  g102
  (
    n80,
    n19
  );


  not
  g103
  (
    n50,
    n24
  );


  buf
  g104
  (
    n44,
    n12
  );


  not
  g105
  (
    n118,
    n30
  );


  not
  g106
  (
    n38,
    n24
  );


  not
  g107
  (
    n158,
    n32
  );


  not
  g108
  (
    n71,
    n12
  );


  not
  g109
  (
    n155,
    n26
  );


  buf
  g110
  (
    n130,
    n20
  );


  buf
  g111
  (
    n81,
    n9
  );


  buf
  g112
  (
    n159,
    n4
  );


  buf
  g113
  (
    n43,
    n14
  );


  buf
  g114
  (
    n54,
    n21
  );


  buf
  g115
  (
    n114,
    n1
  );


  not
  g116
  (
    n49,
    n28
  );


  buf
  g117
  (
    n145,
    n17
  );


  buf
  g118
  (
    n124,
    n20
  );


  not
  g119
  (
    n66,
    n22
  );


  not
  g120
  (
    n52,
    n29
  );


  not
  g121
  (
    n147,
    n8
  );


  not
  g122
  (
    n109,
    n30
  );


  not
  g123
  (
    n133,
    n8
  );


  not
  g124
  (
    n76,
    n3
  );


  not
  g125
  (
    n63,
    n15
  );


  not
  g126
  (
    n131,
    n27
  );


  not
  g127
  (
    n100,
    n32
  );


  buf
  g128
  (
    n511,
    n105
  );


  buf
  g129
  (
    n210,
    n47
  );


  buf
  g130
  (
    n394,
    n41
  );


  buf
  g131
  (
    n520,
    n150
  );


  not
  g132
  (
    n221,
    n65
  );


  not
  g133
  (
    n164,
    n124
  );


  buf
  g134
  (
    n633,
    n89
  );


  not
  g135
  (
    n576,
    n78
  );


  buf
  g136
  (
    n339,
    n114
  );


  buf
  g137
  (
    n577,
    n57
  );


  not
  g138
  (
    n224,
    n138
  );


  not
  g139
  (
    n215,
    n72
  );


  buf
  g140
  (
    n338,
    n66
  );


  not
  g141
  (
    n165,
    n60
  );


  buf
  g142
  (
    n312,
    n116
  );


  not
  g143
  (
    n575,
    n145
  );


  buf
  g144
  (
    n260,
    n100
  );


  not
  g145
  (
    n631,
    n149
  );


  buf
  g146
  (
    n421,
    n97
  );


  not
  g147
  (
    n168,
    n134
  );


  not
  g148
  (
    n516,
    n69
  );


  not
  g149
  (
    n550,
    n124
  );


  buf
  g150
  (
    n632,
    n128
  );


  buf
  g151
  (
    n569,
    n73
  );


  not
  g152
  (
    n202,
    n66
  );


  buf
  g153
  (
    n341,
    n38
  );


  not
  g154
  (
    n375,
    n81
  );


  buf
  g155
  (
    n494,
    n76
  );


  buf
  g156
  (
    n248,
    n130
  );


  buf
  g157
  (
    n386,
    n142
  );


  buf
  g158
  (
    n234,
    n84
  );


  buf
  g159
  (
    n324,
    n136
  );


  not
  g160
  (
    n560,
    n117
  );


  not
  g161
  (
    n602,
    n146
  );


  buf
  g162
  (
    n601,
    n109
  );


  buf
  g163
  (
    n505,
    n99
  );


  not
  g164
  (
    n189,
    n45
  );


  not
  g165
  (
    n423,
    n124
  );


  not
  g166
  (
    n586,
    n144
  );


  buf
  g167
  (
    n497,
    n129
  );


  buf
  g168
  (
    n597,
    n97
  );


  not
  g169
  (
    n486,
    n75
  );


  not
  g170
  (
    n384,
    n107
  );


  buf
  g171
  (
    n469,
    n152
  );


  not
  g172
  (
    n618,
    n52
  );


  buf
  g173
  (
    n351,
    n121
  );


  not
  g174
  (
    n363,
    n142
  );


  not
  g175
  (
    n651,
    n153
  );


  not
  g176
  (
    n193,
    n115
  );


  buf
  g177
  (
    n639,
    n141
  );


  not
  g178
  (
    n211,
    n98
  );


  buf
  g179
  (
    n462,
    n46
  );


  not
  g180
  (
    KeyWire_0_7,
    n37
  );


  not
  g181
  (
    n173,
    n42
  );


  buf
  g182
  (
    n258,
    n42
  );


  buf
  g183
  (
    n171,
    n105
  );


  not
  g184
  (
    n656,
    n116
  );


  buf
  g185
  (
    n416,
    n91
  );


  not
  g186
  (
    n245,
    n33
  );


  buf
  g187
  (
    n181,
    n128
  );


  not
  g188
  (
    n251,
    n82
  );


  not
  g189
  (
    n587,
    n63
  );


  buf
  g190
  (
    n540,
    n122
  );


  buf
  g191
  (
    n395,
    n111
  );


  buf
  g192
  (
    n390,
    n149
  );


  not
  g193
  (
    n368,
    n86
  );


  not
  g194
  (
    n412,
    n82
  );


  buf
  g195
  (
    n238,
    n160
  );


  not
  g196
  (
    n428,
    n152
  );


  not
  g197
  (
    n549,
    n48
  );


  buf
  g198
  (
    n242,
    n119
  );


  not
  g199
  (
    n222,
    n99
  );


  not
  g200
  (
    n317,
    n103
  );


  buf
  g201
  (
    n273,
    n43
  );


  buf
  g202
  (
    n272,
    n129
  );


  buf
  g203
  (
    n647,
    n127
  );


  buf
  g204
  (
    n567,
    n37
  );


  not
  g205
  (
    n483,
    n36
  );


  buf
  g206
  (
    n356,
    n88
  );


  buf
  g207
  (
    n225,
    n85
  );


  not
  g208
  (
    n182,
    n78
  );


  buf
  g209
  (
    n452,
    n126
  );


  buf
  g210
  (
    n485,
    n155
  );


  not
  g211
  (
    n546,
    n86
  );


  buf
  g212
  (
    n169,
    n123
  );


  buf
  g213
  (
    n366,
    n34
  );


  not
  g214
  (
    n642,
    n98
  );


  not
  g215
  (
    n187,
    n41
  );


  buf
  g216
  (
    n596,
    n49
  );


  not
  g217
  (
    n345,
    n148
  );


  not
  g218
  (
    n545,
    n74
  );


  not
  g219
  (
    n233,
    n158
  );


  not
  g220
  (
    n209,
    n54
  );


  not
  g221
  (
    n568,
    n159
  );


  not
  g222
  (
    n410,
    n57
  );


  buf
  g223
  (
    n574,
    n144
  );


  buf
  g224
  (
    n229,
    n106
  );


  not
  g225
  (
    n327,
    n47
  );


  buf
  g226
  (
    n179,
    n76
  );


  buf
  g227
  (
    n319,
    n146
  );


  buf
  g228
  (
    n203,
    n72
  );


  buf
  g229
  (
    n277,
    n121
  );


  buf
  g230
  (
    n358,
    n90
  );


  not
  g231
  (
    n623,
    n79
  );


  buf
  g232
  (
    n406,
    n140
  );


  not
  g233
  (
    n611,
    n143
  );


  buf
  g234
  (
    n279,
    n81
  );


  buf
  g235
  (
    n268,
    n126
  );


  not
  g236
  (
    n479,
    n88
  );


  buf
  g237
  (
    n243,
    n106
  );


  buf
  g238
  (
    n544,
    n125
  );


  buf
  g239
  (
    n393,
    n80
  );


  not
  g240
  (
    n638,
    n56
  );


  buf
  g241
  (
    n609,
    n61
  );


  not
  g242
  (
    n409,
    n113
  );


  buf
  g243
  (
    n400,
    n41
  );


  buf
  g244
  (
    n493,
    n87
  );


  not
  g245
  (
    n509,
    n59
  );


  not
  g246
  (
    n401,
    n71
  );


  buf
  g247
  (
    n612,
    n38
  );


  buf
  g248
  (
    n561,
    n45
  );


  buf
  g249
  (
    n335,
    n150
  );


  not
  g250
  (
    n413,
    n64
  );


  buf
  g251
  (
    n392,
    n58
  );


  buf
  g252
  (
    n526,
    n66
  );


  buf
  g253
  (
    n298,
    n121
  );


  buf
  g254
  (
    n269,
    n68
  );


  not
  g255
  (
    n630,
    n88
  );


  not
  g256
  (
    n590,
    n100
  );


  not
  g257
  (
    n192,
    n127
  );


  buf
  g258
  (
    n304,
    n123
  );


  not
  g259
  (
    n226,
    n110
  );


  not
  g260
  (
    n257,
    n50
  );


  buf
  g261
  (
    n278,
    n55
  );


  not
  g262
  (
    n201,
    n113
  );


  not
  g263
  (
    n517,
    n48
  );


  not
  g264
  (
    n283,
    n140
  );


  buf
  g265
  (
    n239,
    n80
  );


  not
  g266
  (
    n220,
    n118
  );


  not
  g267
  (
    n660,
    n128
  );


  not
  g268
  (
    n266,
    n93
  );


  buf
  g269
  (
    n364,
    n87
  );


  buf
  g270
  (
    n637,
    n149
  );


  buf
  g271
  (
    n309,
    n37
  );


  buf
  g272
  (
    n478,
    n39
  );


  not
  g273
  (
    n342,
    n83
  );


  buf
  g274
  (
    n161,
    n79
  );


  not
  g275
  (
    n482,
    n101
  );


  buf
  g276
  (
    n628,
    n93
  );


  not
  g277
  (
    n391,
    n113
  );


  buf
  g278
  (
    n565,
    n153
  );


  not
  g279
  (
    n538,
    n69
  );


  buf
  g280
  (
    n223,
    n112
  );


  buf
  g281
  (
    n326,
    n133
  );


  not
  g282
  (
    n383,
    n75
  );


  buf
  g283
  (
    n484,
    n39
  );


  not
  g284
  (
    n252,
    n139
  );


  buf
  g285
  (
    n417,
    n48
  );


  buf
  g286
  (
    n519,
    n117
  );


  not
  g287
  (
    n175,
    n61
  );


  not
  g288
  (
    n167,
    n53
  );


  not
  g289
  (
    n343,
    n108
  );


  not
  g290
  (
    n284,
    n70
  );


  buf
  g291
  (
    n186,
    n40
  );


  buf
  g292
  (
    n573,
    n135
  );


  not
  g293
  (
    n231,
    n147
  );


  not
  g294
  (
    n206,
    n100
  );


  not
  g295
  (
    n228,
    n102
  );


  buf
  g296
  (
    n473,
    n156
  );


  not
  g297
  (
    n426,
    n152
  );


  buf
  g298
  (
    n359,
    n156
  );


  not
  g299
  (
    n434,
    n82
  );


  buf
  g300
  (
    n604,
    n94
  );


  buf
  g301
  (
    n330,
    n36
  );


  not
  g302
  (
    n552,
    n66
  );


  buf
  g303
  (
    n463,
    n96
  );


  not
  g304
  (
    n293,
    n131
  );


  not
  g305
  (
    n634,
    n125
  );


  not
  g306
  (
    n619,
    n130
  );


  buf
  g307
  (
    n643,
    n136
  );


  buf
  g308
  (
    n502,
    n158
  );


  not
  g309
  (
    n177,
    n92
  );


  not
  g310
  (
    n652,
    n115
  );


  buf
  g311
  (
    n296,
    n44
  );


  buf
  g312
  (
    n444,
    n86
  );


  not
  g313
  (
    n608,
    n60
  );


  buf
  g314
  (
    n297,
    n138
  );


  buf
  g315
  (
    n461,
    n96
  );


  buf
  g316
  (
    n584,
    n94
  );


  not
  g317
  (
    n344,
    n59
  );


  not
  g318
  (
    n610,
    n45
  );


  buf
  g319
  (
    n666,
    n131
  );


  not
  g320
  (
    n476,
    n146
  );


  buf
  g321
  (
    n453,
    n136
  );


  buf
  g322
  (
    n492,
    n152
  );


  not
  g323
  (
    n616,
    n155
  );


  buf
  g324
  (
    n571,
    n39
  );


  not
  g325
  (
    n454,
    n98
  );


  not
  g326
  (
    n564,
    n89
  );


  not
  g327
  (
    n337,
    n116
  );


  buf
  g328
  (
    n289,
    n93
  );


  not
  g329
  (
    n340,
    n125
  );


  buf
  g330
  (
    n503,
    n157
  );


  buf
  g331
  (
    n440,
    n131
  );


  not
  g332
  (
    n262,
    n40
  );


  not
  g333
  (
    n558,
    n62
  );


  not
  g334
  (
    n504,
    n133
  );


  not
  g335
  (
    n166,
    n74
  );


  not
  g336
  (
    n606,
    n39
  );


  not
  g337
  (
    n163,
    n64
  );


  not
  g338
  (
    n559,
    n79
  );


  buf
  g339
  (
    n301,
    n52
  );


  not
  g340
  (
    n362,
    n43
  );


  not
  g341
  (
    n305,
    n124
  );


  not
  g342
  (
    n599,
    n44
  );


  not
  g343
  (
    n236,
    n76
  );


  buf
  g344
  (
    n665,
    n34
  );


  buf
  g345
  (
    n667,
    n59
  );


  buf
  g346
  (
    n672,
    n42
  );


  buf
  g347
  (
    n589,
    n61
  );


  buf
  g348
  (
    n240,
    n65
  );


  buf
  g349
  (
    n331,
    n48
  );


  not
  g350
  (
    n350,
    n64
  );


  not
  g351
  (
    n532,
    n111
  );


  buf
  g352
  (
    n582,
    n38
  );


  buf
  g353
  (
    n622,
    n93
  );


  buf
  g354
  (
    n276,
    n62
  );


  not
  g355
  (
    n663,
    n145
  );


  not
  g356
  (
    n365,
    n73
  );


  buf
  g357
  (
    n661,
    n103
  );


  buf
  g358
  (
    n255,
    n141
  );


  buf
  g359
  (
    n649,
    n55
  );


  buf
  g360
  (
    n199,
    n125
  );


  not
  g361
  (
    n624,
    n104
  );


  not
  g362
  (
    n464,
    n150
  );


  buf
  g363
  (
    n196,
    n145
  );


  buf
  g364
  (
    n399,
    n126
  );


  buf
  g365
  (
    n183,
    n135
  );


  buf
  g366
  (
    n653,
    n123
  );


  not
  g367
  (
    n377,
    n36
  );


  not
  g368
  (
    n581,
    n78
  );


  buf
  g369
  (
    n264,
    n35
  );


  not
  g370
  (
    n360,
    n108
  );


  not
  g371
  (
    n515,
    n95
  );


  not
  g372
  (
    n411,
    n52
  );


  buf
  g373
  (
    n455,
    n108
  );


  not
  g374
  (
    n443,
    n102
  );


  buf
  g375
  (
    n398,
    n84
  );


  not
  g376
  (
    n379,
    n135
  );


  not
  g377
  (
    n306,
    n133
  );


  not
  g378
  (
    n372,
    n64
  );


  buf
  g379
  (
    n354,
    n49
  );


  buf
  g380
  (
    n184,
    n77
  );


  not
  g381
  (
    n525,
    n103
  );


  not
  g382
  (
    n274,
    n88
  );


  not
  g383
  (
    n530,
    n111
  );


  not
  g384
  (
    n570,
    n49
  );


  not
  g385
  (
    n408,
    n122
  );


  buf
  g386
  (
    n265,
    n55
  );


  buf
  g387
  (
    n563,
    n70
  );


  not
  g388
  (
    n430,
    n138
  );


  buf
  g389
  (
    n427,
    n107
  );


  not
  g390
  (
    n246,
    n153
  );


  not
  g391
  (
    n562,
    n65
  );


  not
  g392
  (
    n466,
    n107
  );


  buf
  g393
  (
    n543,
    n117
  );


  not
  g394
  (
    n437,
    n130
  );


  not
  g395
  (
    n635,
    n41
  );


  not
  g396
  (
    n446,
    n109
  );


  buf
  g397
  (
    n664,
    n37
  );


  buf
  g398
  (
    n244,
    n35
  );


  not
  g399
  (
    n347,
    n147
  );


  not
  g400
  (
    n669,
    n67
  );


  not
  g401
  (
    n627,
    n81
  );


  not
  g402
  (
    n321,
    n72
  );


  buf
  g403
  (
    n621,
    n127
  );


  buf
  g404
  (
    n172,
    n103
  );


  buf
  g405
  (
    n442,
    n65
  );


  buf
  g406
  (
    n275,
    n157
  );


  not
  g407
  (
    n548,
    n50
  );


  not
  g408
  (
    n227,
    n54
  );


  buf
  g409
  (
    n620,
    n78
  );


  buf
  g410
  (
    n551,
    n135
  );


  not
  g411
  (
    n303,
    n151
  );


  not
  g412
  (
    n217,
    n140
  );


  not
  g413
  (
    n374,
    n33
  );


  not
  g414
  (
    n299,
    n120
  );


  not
  g415
  (
    n605,
    n63
  );


  buf
  g416
  (
    n369,
    n50
  );


  buf
  g417
  (
    n332,
    n62
  );


  buf
  g418
  (
    n650,
    n156
  );


  buf
  g419
  (
    n470,
    n122
  );


  buf
  g420
  (
    n598,
    n100
  );


  not
  g421
  (
    n388,
    n34
  );


  not
  g422
  (
    n370,
    n81
  );


  not
  g423
  (
    n316,
    n95
  );


  buf
  g424
  (
    n495,
    n159
  );


  buf
  g425
  (
    n381,
    n95
  );


  not
  g426
  (
    n445,
    n97
  );


  buf
  g427
  (
    n522,
    n58
  );


  not
  g428
  (
    n518,
    n115
  );


  not
  g429
  (
    n194,
    n118
  );


  not
  g430
  (
    n180,
    n160
  );


  not
  g431
  (
    n636,
    n80
  );


  buf
  g432
  (
    n472,
    n59
  );


  not
  g433
  (
    n198,
    n54
  );


  not
  g434
  (
    n349,
    n102
  );


  buf
  g435
  (
    n389,
    n57
  );


  buf
  g436
  (
    n310,
    n110
  );


  not
  g437
  (
    n378,
    n102
  );


  buf
  g438
  (
    n448,
    n76
  );


  not
  g439
  (
    n555,
    n94
  );


  not
  g440
  (
    n547,
    n154
  );


  not
  g441
  (
    n415,
    n106
  );


  not
  g442
  (
    n190,
    n49
  );


  not
  g443
  (
    n241,
    n43
  );


  buf
  g444
  (
    n314,
    n33
  );


  buf
  g445
  (
    n407,
    n85
  );


  not
  g446
  (
    n467,
    n77
  );


  not
  g447
  (
    n556,
    n154
  );


  buf
  g448
  (
    n441,
    n61
  );


  buf
  g449
  (
    n281,
    n114
  );


  buf
  g450
  (
    n334,
    n91
  );


  not
  g451
  (
    n254,
    n84
  );


  not
  g452
  (
    n641,
    n143
  );


  not
  g453
  (
    n625,
    n153
  );


  not
  g454
  (
    n496,
    n44
  );


  not
  g455
  (
    n539,
    n150
  );


  buf
  g456
  (
    n487,
    n85
  );


  buf
  g457
  (
    n237,
    n95
  );


  not
  g458
  (
    n500,
    n33
  );


  not
  g459
  (
    n583,
    n87
  );


  not
  g460
  (
    n655,
    n40
  );


  not
  g461
  (
    n480,
    n101
  );


  buf
  g462
  (
    n593,
    n77
  );


  not
  g463
  (
    n535,
    n131
  );


  buf
  g464
  (
    n528,
    n158
  );


  buf
  g465
  (
    n458,
    n36
  );


  buf
  g466
  (
    n536,
    n122
  );


  not
  g467
  (
    n396,
    n132
  );


  buf
  g468
  (
    n670,
    n129
  );


  not
  g469
  (
    n318,
    n84
  );


  buf
  g470
  (
    n585,
    n99
  );


  not
  g471
  (
    n253,
    n155
  );


  not
  g472
  (
    n195,
    n101
  );


  buf
  g473
  (
    n214,
    n90
  );


  buf
  g474
  (
    n307,
    n62
  );


  buf
  g475
  (
    n527,
    n57
  );


  buf
  g476
  (
    n501,
    n53
  );


  buf
  g477
  (
    n270,
    n82
  );


  buf
  g478
  (
    n449,
    n101
  );


  buf
  g479
  (
    n475,
    n58
  );


  not
  g480
  (
    n617,
    n109
  );


  not
  g481
  (
    n197,
    n155
  );


  buf
  g482
  (
    n510,
    n116
  );


  buf
  g483
  (
    n592,
    n151
  );


  buf
  g484
  (
    n422,
    n132
  );


  buf
  g485
  (
    n591,
    n160
  );


  buf
  g486
  (
    n282,
    n83
  );


  buf
  g487
  (
    n603,
    n151
  );


  not
  g488
  (
    n292,
    n112
  );


  buf
  g489
  (
    n300,
    n47
  );


  not
  g490
  (
    n185,
    n104
  );


  not
  g491
  (
    n208,
    n104
  );


  buf
  g492
  (
    n424,
    n99
  );


  not
  g493
  (
    n235,
    n96
  );


  buf
  g494
  (
    n512,
    n110
  );


  buf
  g495
  (
    n523,
    n77
  );


  buf
  g496
  (
    n267,
    n159
  );


  buf
  g497
  (
    n419,
    n106
  );


  buf
  g498
  (
    n614,
    n120
  );


  buf
  g499
  (
    n213,
    n140
  );


  buf
  g500
  (
    n320,
    n51
  );


  not
  g501
  (
    n451,
    n114
  );


  not
  g502
  (
    n465,
    n113
  );


  not
  g503
  (
    n323,
    n115
  );


  buf
  g504
  (
    n348,
    n46
  );


  not
  g505
  (
    n205,
    n128
  );


  buf
  g506
  (
    n600,
    n68
  );


  not
  g507
  (
    n325,
    n44
  );


  not
  g508
  (
    n506,
    n142
  );


  not
  g509
  (
    n477,
    n96
  );


  not
  g510
  (
    n657,
    n120
  );


  buf
  g511
  (
    n488,
    n136
  );


  buf
  g512
  (
    n554,
    n67
  );


  buf
  g513
  (
    n380,
    n85
  );


  not
  g514
  (
    n219,
    n141
  );


  buf
  g515
  (
    n645,
    n92
  );


  buf
  g516
  (
    n191,
    n138
  );


  not
  g517
  (
    n468,
    n147
  );


  not
  g518
  (
    n207,
    n132
  );


  buf
  g519
  (
    n459,
    n79
  );


  not
  g520
  (
    n566,
    n56
  );


  not
  g521
  (
    n481,
    n154
  );


  not
  g522
  (
    n382,
    n43
  );


  not
  g523
  (
    n200,
    n137
  );


  buf
  g524
  (
    n615,
    n119
  );


  not
  g525
  (
    n346,
    n118
  );


  buf
  g526
  (
    n230,
    n83
  );


  buf
  g527
  (
    n232,
    n110
  );


  not
  g528
  (
    n658,
    n120
  );


  buf
  g529
  (
    n668,
    n108
  );


  not
  g530
  (
    n218,
    n139
  );


  buf
  g531
  (
    n367,
    n111
  );


  buf
  g532
  (
    n439,
    n92
  );


  not
  g533
  (
    n287,
    n35
  );


  buf
  g534
  (
    n402,
    n119
  );


  buf
  g535
  (
    n263,
    n52
  );


  buf
  g536
  (
    n286,
    n134
  );


  buf
  g537
  (
    n285,
    n149
  );


  not
  g538
  (
    n542,
    n127
  );


  buf
  g539
  (
    n537,
    n86
  );


  buf
  g540
  (
    n435,
    n73
  );


  buf
  g541
  (
    n438,
    n75
  );


  buf
  g542
  (
    n403,
    n141
  );


  buf
  g543
  (
    n302,
    n71
  );


  buf
  g544
  (
    n534,
    n132
  );


  buf
  g545
  (
    n216,
    n75
  );


  buf
  g546
  (
    n397,
    n156
  );


  buf
  g547
  (
    n414,
    n54
  );


  buf
  g548
  (
    n328,
    n105
  );


  buf
  g549
  (
    n271,
    n139
  );


  buf
  g550
  (
    n170,
    n112
  );


  not
  g551
  (
    n259,
    n90
  );


  buf
  g552
  (
    n256,
    n134
  );


  not
  g553
  (
    n294,
    n46
  );


  not
  g554
  (
    n640,
    n143
  );


  not
  g555
  (
    n489,
    n134
  );


  buf
  g556
  (
    n204,
    n90
  );


  buf
  g557
  (
    n429,
    n71
  );


  buf
  g558
  (
    n247,
    n51
  );


  not
  g559
  (
    n572,
    n89
  );


  not
  g560
  (
    n514,
    n137
  );


  buf
  g561
  (
    n280,
    n60
  );


  buf
  g562
  (
    n595,
    n146
  );


  not
  g563
  (
    n376,
    n118
  );


  buf
  g564
  (
    n553,
    n91
  );


  buf
  g565
  (
    n662,
    n87
  );


  not
  g566
  (
    n594,
    n148
  );


  not
  g567
  (
    n471,
    n105
  );


  buf
  g568
  (
    n521,
    n157
  );


  not
  g569
  (
    n433,
    n89
  );


  buf
  g570
  (
    n371,
    n70
  );


  not
  g571
  (
    n578,
    n55
  );


  buf
  g572
  (
    n654,
    n158
  );


  buf
  g573
  (
    n250,
    n104
  );


  buf
  g574
  (
    n420,
    n139
  );


  not
  g575
  (
    n533,
    n72
  );


  not
  g576
  (
    n405,
    n50
  );


  not
  g577
  (
    n557,
    n35
  );


  not
  g578
  (
    n507,
    n68
  );


  not
  g579
  (
    n425,
    n71
  );


  not
  g580
  (
    n490,
    n63
  );


  buf
  g581
  (
    n513,
    n42
  );


  not
  g582
  (
    n322,
    n129
  );


  not
  g583
  (
    n648,
    n56
  );


  buf
  g584
  (
    n646,
    n114
  );


  buf
  g585
  (
    n531,
    n51
  );


  not
  g586
  (
    n404,
    n69
  );


  buf
  g587
  (
    n671,
    n144
  );


  buf
  g588
  (
    n541,
    n83
  );


  not
  g589
  (
    n431,
    n73
  );


  buf
  g590
  (
    n291,
    n46
  );


  not
  g591
  (
    n607,
    n69
  );


  buf
  g592
  (
    KeyWire_0_6,
    n80
  );


  not
  g593
  (
    n588,
    n40
  );


  not
  g594
  (
    n353,
    n154
  );


  not
  g595
  (
    n311,
    n112
  );


  buf
  g596
  (
    n212,
    n68
  );


  buf
  g597
  (
    n333,
    n67
  );


  not
  g598
  (
    n176,
    n97
  );


  not
  g599
  (
    n290,
    n53
  );


  not
  g600
  (
    n474,
    n51
  );


  not
  g601
  (
    n357,
    n91
  );


  not
  g602
  (
    n460,
    n92
  );


  not
  g603
  (
    n288,
    n117
  );


  not
  g604
  (
    n456,
    n142
  );


  not
  g605
  (
    n373,
    n45
  );


  buf
  g606
  (
    n313,
    n126
  );


  not
  g607
  (
    n315,
    n137
  );


  not
  g608
  (
    n450,
    n159
  );


  buf
  g609
  (
    n336,
    n123
  );


  buf
  g610
  (
    n457,
    n133
  );


  not
  g611
  (
    n436,
    n34
  );


  buf
  g612
  (
    n174,
    n143
  );


  buf
  g613
  (
    n629,
    n47
  );


  buf
  g614
  (
    n644,
    n38
  );


  buf
  g615
  (
    n579,
    n58
  );


  not
  g616
  (
    n613,
    n145
  );


  not
  g617
  (
    n361,
    n60
  );


  not
  g618
  (
    n261,
    n160
  );


  buf
  g619
  (
    n162,
    n98
  );


  buf
  g620
  (
    n580,
    n63
  );


  buf
  g621
  (
    n498,
    n74
  );


  not
  g622
  (
    n355,
    n119
  );


  not
  g623
  (
    n508,
    n137
  );


  buf
  g624
  (
    n249,
    n147
  );


  not
  g625
  (
    n418,
    n130
  );


  buf
  g626
  (
    n659,
    n67
  );


  not
  g627
  (
    n352,
    n148
  );


  not
  g628
  (
    n499,
    n74
  );


  buf
  g629
  (
    n295,
    n157
  );


  buf
  g630
  (
    n447,
    n94
  );


  buf
  g631
  (
    n524,
    n151
  );


  not
  g632
  (
    n308,
    n144
  );


  not
  g633
  (
    n387,
    n148
  );


  not
  g634
  (
    n626,
    n109
  );


  buf
  g635
  (
    n178,
    n70
  );


  buf
  g636
  (
    n529,
    n107
  );


  not
  g637
  (
    n385,
    n121
  );


  not
  g638
  (
    n491,
    n56
  );


  buf
  g639
  (
    n432,
    n53
  );


  nand
  g640
  (
    n695,
    n397,
    n518,
    n426,
    n668
  );


  and
  g641
  (
    n1066,
    n331,
    n231,
    n435,
    n629
  );


  xnor
  g642
  (
    n777,
    n198,
    n655,
    n639,
    n621
  );


  and
  g643
  (
    n778,
    n576,
    n422,
    n233,
    n183
  );


  xor
  g644
  (
    n995,
    n662,
    n645,
    n171,
    n297
  );


  nand
  g645
  (
    n1121,
    n465,
    n351,
    n325,
    n355
  );


  and
  g646
  (
    n979,
    n347,
    n554,
    n444,
    n252
  );


  xor
  g647
  (
    n742,
    n620,
    n428,
    n484,
    n575
  );


  xor
  g648
  (
    n679,
    n356,
    n608,
    n387,
    n571
  );


  nand
  g649
  (
    n826,
    n498,
    n478,
    n602,
    n212
  );


  nor
  g650
  (
    n911,
    n524,
    n544,
    n355,
    n395
  );


  or
  g651
  (
    n868,
    n275,
    n381,
    n436,
    n604
  );


  nor
  g652
  (
    n1007,
    n444,
    n316,
    n261,
    n204
  );


  xnor
  g653
  (
    n1045,
    n480,
    n300,
    n605,
    n630
  );


  nand
  g654
  (
    n1146,
    n575,
    n457,
    n251,
    n553
  );


  or
  g655
  (
    n727,
    n278,
    n665,
    n190,
    n549
  );


  and
  g656
  (
    n1052,
    n495,
    n256,
    n552,
    n493
  );


  and
  g657
  (
    n1006,
    n201,
    n410,
    n350,
    n525
  );


  xnor
  g658
  (
    n1009,
    n191,
    n381,
    n580,
    n211
  );


  xor
  g659
  (
    n1119,
    n176,
    n477,
    n333,
    n256
  );


  xor
  g660
  (
    n717,
    n417,
    n358,
    n479,
    n596
  );


  xnor
  g661
  (
    n1161,
    n265,
    n416,
    n590,
    n496
  );


  nand
  g662
  (
    n903,
    n643,
    n659,
    n258,
    n450
  );


  xnor
  g663
  (
    n1054,
    n412,
    n494,
    n491,
    n177
  );


  xor
  g664
  (
    n1053,
    n573,
    n494,
    n589,
    n331
  );


  nor
  g665
  (
    n1152,
    n338,
    n471,
    n506
  );


  nand
  g666
  (
    n867,
    n269,
    n472,
    n516,
    n356
  );


  and
  g667
  (
    n1100,
    n200,
    n447,
    n585,
    n455
  );


  xor
  g668
  (
    n1117,
    n260,
    n554,
    n656,
    n346
  );


  xnor
  g669
  (
    n988,
    n432,
    n416,
    n407,
    n300
  );


  and
  g670
  (
    n896,
    n468,
    n469,
    n470,
    n345
  );


  nand
  g671
  (
    n949,
    n567,
    n472,
    n238,
    n549
  );


  and
  g672
  (
    n714,
    n450,
    n436,
    n578,
    n236
  );


  xor
  g673
  (
    n1167,
    n378,
    n611,
    n250,
    n565
  );


  xnor
  g674
  (
    n1068,
    n545,
    n164,
    n450,
    n182
  );


  xnor
  g675
  (
    n977,
    n364,
    n605,
    n543,
    n621
  );


  xnor
  g676
  (
    n1180,
    n575,
    n186,
    n667,
    n480
  );


  nand
  g677
  (
    n786,
    n397,
    n172,
    n349,
    n304
  );


  and
  g678
  (
    n1005,
    n454,
    n270,
    n443,
    n595
  );


  xnor
  g679
  (
    n997,
    n322,
    n492,
    n458,
    n486
  );


  xor
  g680
  (
    n1129,
    n510,
    n349,
    n548,
    n402
  );


  nand
  g681
  (
    n893,
    n617,
    n194,
    n546,
    n332
  );


  nand
  g682
  (
    n722,
    n361,
    n213,
    n339,
    n262
  );


  nor
  g683
  (
    n836,
    n276,
    n499,
    n628,
    n342
  );


  nor
  g684
  (
    n890,
    n305,
    n465,
    n164,
    n601
  );


  or
  g685
  (
    n673,
    n569,
    n531,
    n178,
    n233
  );


  or
  g686
  (
    n992,
    n642,
    n462,
    n165,
    n339
  );


  nand
  g687
  (
    n734,
    n451,
    n622,
    n543,
    n578
  );


  or
  g688
  (
    n1091,
    n470,
    n593,
    n216,
    n498
  );


  or
  g689
  (
    n966,
    n551,
    n600,
    n294,
    n412
  );


  or
  g690
  (
    n1151,
    n555,
    n294,
    n420,
    n379
  );


  xnor
  g691
  (
    n1039,
    n359,
    n484,
    n537,
    n659
  );


  or
  g692
  (
    n1124,
    n288,
    n570,
    n383,
    n429
  );


  nor
  g693
  (
    n685,
    n263,
    n534,
    n303,
    n569
  );


  and
  g694
  (
    n955,
    n318,
    n413,
    n489,
    n380
  );


  or
  g695
  (
    n989,
    n191,
    n648,
    n595,
    n219
  );


  or
  g696
  (
    n923,
    n490,
    n409,
    n451,
    n477
  );


  or
  g697
  (
    n1042,
    n432,
    n389,
    n204,
    n227
  );


  nand
  g698
  (
    n858,
    n265,
    n603,
    n565,
    n248
  );


  xor
  g699
  (
    n969,
    n418,
    n622,
    n660,
    n296
  );


  xnor
  g700
  (
    n716,
    n257,
    n234,
    n432,
    n291
  );


  or
  g701
  (
    n880,
    n258,
    n162,
    n271,
    n603
  );


  nand
  g702
  (
    n701,
    n409,
    n566,
    n551,
    n405
  );


  and
  g703
  (
    n1174,
    n416,
    n325,
    n601,
    n339
  );


  xnor
  g704
  (
    n985,
    n360,
    n444,
    n533,
    n542
  );


  or
  g705
  (
    KeyWire_0_15,
    n321,
    n240,
    n179,
    n613
  );


  or
  g706
  (
    n747,
    n611,
    n415,
    n502,
    n404
  );


  xnor
  g707
  (
    n1093,
    n364,
    n267,
    n457,
    n613
  );


  and
  g708
  (
    n1128,
    n618,
    n194,
    n469,
    n432
  );


  nand
  g709
  (
    n1157,
    n525,
    n579,
    n334,
    n578
  );


  nand
  g710
  (
    n774,
    n524,
    n522,
    n558,
    n466
  );


  nand
  g711
  (
    n807,
    n207,
    n476,
    n399,
    n170
  );


  or
  g712
  (
    n901,
    n427,
    n661,
    n509,
    n277
  );


  and
  g713
  (
    n1130,
    n447,
    n667,
    n414,
    n616
  );


  nand
  g714
  (
    n864,
    n319,
    n590,
    n548,
    n564
  );


  nor
  g715
  (
    n1025,
    n601,
    n299,
    n391,
    n576
  );


  nor
  g716
  (
    n1024,
    n165,
    n184,
    n248,
    n252
  );


  xor
  g717
  (
    n908,
    n586,
    n533,
    n582,
    n296
  );


  xnor
  g718
  (
    n682,
    n611,
    n622,
    n405,
    n557
  );


  and
  g719
  (
    n1164,
    n257,
    n402,
    n417,
    n306
  );


  xor
  g720
  (
    n756,
    n255,
    n588,
    n281,
    n309
  );


  xor
  g721
  (
    n741,
    n480,
    n367,
    n473,
    n422
  );


  nor
  g722
  (
    n1016,
    n510,
    n415,
    n624,
    n301
  );


  xnor
  g723
  (
    n761,
    n298,
    n441,
    n494,
    n547
  );


  and
  g724
  (
    n1044,
    n219,
    n328,
    n214,
    n199
  );


  nor
  g725
  (
    n866,
    n414,
    n172,
    n250,
    n427
  );


  nor
  g726
  (
    n1060,
    n396,
    n373,
    n323,
    n421
  );


  nand
  g727
  (
    n793,
    n443,
    n236,
    n251,
    n313
  );


  nand
  g728
  (
    n764,
    n506,
    n337,
    n517,
    n361
  );


  xnor
  g729
  (
    n721,
    n530,
    n641,
    n564,
    n492
  );


  and
  g730
  (
    n849,
    n232,
    n599,
    n475,
    n662
  );


  nand
  g731
  (
    n1020,
    n651,
    n285,
    n348,
    n618
  );


  xnor
  g732
  (
    n1163,
    n585,
    n338,
    n527,
    n330
  );


  or
  g733
  (
    n938,
    n281,
    n612,
    n249,
    n561
  );


  xor
  g734
  (
    n1059,
    n375,
    n188,
    n410,
    n222
  );


  or
  g735
  (
    n863,
    n195,
    n567,
    n248,
    n302
  );


  and
  g736
  (
    n677,
    n247,
    n394,
    n218
  );


  nor
  g737
  (
    n1023,
    n368,
    n538,
    n589,
    n280
  );


  nor
  g738
  (
    n841,
    n457,
    n557,
    n363,
    n621
  );


  or
  g739
  (
    n944,
    n560,
    n576,
    n475,
    n306
  );


  nand
  g740
  (
    n800,
    n375,
    n194,
    n265,
    n550
  );


  or
  g741
  (
    n848,
    n529,
    n544,
    n186,
    n522
  );


  xnor
  g742
  (
    n990,
    n505,
    n352,
    n515,
    n260
  );


  xnor
  g743
  (
    n1101,
    n467,
    n663,
    n419,
    n536
  );


  nor
  g744
  (
    n1033,
    n297,
    n654,
    n493,
    n507
  );


  and
  g745
  (
    n986,
    n590,
    n539,
    n201,
    n350
  );


  xor
  g746
  (
    n1051,
    n259,
    n164,
    n360,
    n518
  );


  xor
  g747
  (
    n776,
    n165,
    n601,
    n442,
    n592
  );


  xnor
  g748
  (
    n1031,
    n633,
    n516,
    n289,
    n237
  );


  nand
  g749
  (
    n810,
    n354,
    n455,
    n587,
    n536
  );


  nand
  g750
  (
    n902,
    n508,
    n400,
    n434,
    n203
  );


  nand
  g751
  (
    n891,
    n396,
    n516,
    n649,
    n332
  );


  xor
  g752
  (
    n998,
    n220,
    n347,
    n307,
    n462
  );


  and
  g753
  (
    n1126,
    n206,
    n311,
    n545,
    n524
  );


  xnor
  g754
  (
    n770,
    n523,
    n197,
    n340,
    n525
  );


  nor
  g755
  (
    n924,
    n631,
    n500,
    n267,
    n600
  );


  xnor
  g756
  (
    n823,
    n364,
    n312,
    n493,
    n512
  );


  and
  g757
  (
    n1021,
    n227,
    n225,
    n484,
    n430
  );


  xor
  g758
  (
    n1115,
    n513,
    n304,
    n253,
    n174
  );


  nand
  g759
  (
    n811,
    n284,
    n650,
    n563,
    n225
  );


  and
  g760
  (
    n967,
    n352,
    n666,
    n372,
    n242
  );


  nand
  g761
  (
    n932,
    n366,
    n596,
    n363,
    n665
  );


  xnor
  g762
  (
    n1181,
    n492,
    n512,
    n639,
    n599
  );


  xnor
  g763
  (
    n1047,
    n283,
    n301,
    n282,
    n452
  );


  nor
  g764
  (
    n771,
    n539,
    n544,
    n319,
    n615
  );


  nand
  g765
  (
    n905,
    n253,
    n301,
    n230,
    n597
  );


  nor
  g766
  (
    n1062,
    n495,
    n429,
    n482,
    n490
  );


  nor
  g767
  (
    n785,
    n205,
    n418,
    n619,
    n416
  );


  and
  g768
  (
    n1084,
    n414,
    n342,
    n434,
    n395
  );


  or
  g769
  (
    KeyWire_0_8,
    n376,
    n518,
    n401,
    n185
  );


  nor
  g770
  (
    n1170,
    n344,
    n202,
    n477,
    n600
  );


  xnor
  g771
  (
    n1154,
    n626,
    n439,
    n501,
    n381
  );


  and
  g772
  (
    n851,
    n614,
    n254,
    n603,
    n461
  );


  and
  g773
  (
    n936,
    n341,
    n309,
    n239,
    n255
  );


  nand
  g774
  (
    n728,
    n334,
    n501,
    n295,
    n239
  );


  or
  g775
  (
    n820,
    n647,
    n378,
    n622,
    n431
  );


  nor
  g776
  (
    n888,
    n490,
    n665,
    n644,
    n352
  );


  xnor
  g777
  (
    n1141,
    n446,
    n221,
    n502,
    n385
  );


  nor
  g778
  (
    n762,
    n663,
    n250,
    n612,
    n438
  );


  xor
  g779
  (
    n853,
    n668,
    n658,
    n610,
    n452
  );


  xnor
  g780
  (
    n931,
    n209,
    n223,
    n308,
    n302
  );


  and
  g781
  (
    n1136,
    n167,
    n161,
    n386,
    n336
  );


  xnor
  g782
  (
    n1148,
    n237,
    n319,
    n435,
    n229
  );


  nor
  g783
  (
    n675,
    n226,
    n321,
    n391,
    n401
  );


  nand
  g784
  (
    n974,
    n310,
    n388,
    n430,
    n369
  );


  xor
  g785
  (
    n999,
    n557,
    n273,
    n554,
    n167
  );


  xnor
  g786
  (
    n837,
    n462,
    n562,
    n344,
    n315
  );


  and
  g787
  (
    n1008,
    n609,
    n418,
    n666,
    n560
  );


  xnor
  g788
  (
    n754,
    n184,
    n166,
    n564,
    n636
  );


  or
  g789
  (
    n797,
    n185,
    n288,
    n394,
    n365
  );


  and
  g790
  (
    n1109,
    n583,
    n487,
    n217,
    n351
  );


  xor
  g791
  (
    n831,
    n242,
    n184,
    n487,
    n572
  );


  nor
  g792
  (
    n945,
    n215,
    n539,
    n579,
    n489
  );


  xnor
  g793
  (
    n686,
    n406,
    n441,
    n438,
    n629
  );


  xnor
  g794
  (
    n1160,
    n358,
    n666,
    n424,
    n485
  );


  and
  g795
  (
    n930,
    n384,
    n392,
    n527,
    n425
  );


  xor
  g796
  (
    n731,
    n367,
    n445,
    n392,
    n597
  );


  nand
  g797
  (
    n711,
    n263,
    n315,
    n168,
    n526
  );


  and
  g798
  (
    n947,
    n591,
    n411,
    n533,
    n637
  );


  xor
  g799
  (
    n1153,
    n483,
    n567,
    n508,
    n655
  );


  nor
  g800
  (
    n828,
    n608,
    n284,
    n439,
    n293
  );


  nor
  g801
  (
    n812,
    n235,
    n396,
    n278,
    n173
  );


  or
  g802
  (
    n916,
    n612,
    n399,
    n486,
    n198
  );


  xor
  g803
  (
    n912,
    n317,
    n541,
    n292,
    n403
  );


  nand
  g804
  (
    n732,
    n404,
    n163,
    n169,
    n632
  );


  and
  g805
  (
    n697,
    n183,
    n389,
    n552,
    n175
  );


  xnor
  g806
  (
    n1057,
    n542,
    n323,
    n226,
    n395
  );


  xnor
  g807
  (
    n755,
    n176,
    n390,
    n650,
    n550
  );


  and
  g808
  (
    n879,
    n627,
    n633,
    n244,
    n236
  );


  xor
  g809
  (
    n681,
    n210,
    n230,
    n411,
    n508
  );


  xnor
  g810
  (
    n1081,
    n610,
    n492,
    n635,
    n583
  );


  nand
  g811
  (
    n1094,
    n429,
    n239,
    n631,
    n257
  );


  nand
  g812
  (
    n744,
    n629,
    n495,
    n383,
    n447
  );


  or
  g813
  (
    n758,
    n467,
    n524,
    n497,
    n625
  );


  and
  g814
  (
    n1166,
    n205,
    n628,
    n284,
    n191
  );


  and
  g815
  (
    n918,
    n592,
    n565,
    n348,
    n630
  );


  nor
  g816
  (
    n1026,
    n567,
    n620,
    n479,
    n414
  );


  and
  g817
  (
    n688,
    n606,
    n227,
    n272,
    n266
  );


  nor
  g818
  (
    n739,
    n581,
    n192,
    n636,
    n276
  );


  xor
  g819
  (
    n1122,
    n320,
    n308,
    n507,
    n582
  );


  nor
  g820
  (
    n946,
    n606,
    n640,
    n404,
    n207
  );


  or
  g821
  (
    n907,
    n199,
    n236,
    n647,
    n626
  );


  xor
  g822
  (
    n987,
    n179,
    n163,
    n658,
    n259
  );


  xnor
  g823
  (
    n809,
    n575,
    n317,
    n201,
    n410
  );


  and
  g824
  (
    n1076,
    n553,
    n220,
    n515,
    n393
  );


  nand
  g825
  (
    n782,
    n633,
    n451,
    n660,
    n552
  );


  nand
  g826
  (
    n787,
    n327,
    n548,
    n608,
    n360
  );


  nor
  g827
  (
    n935,
    n193,
    n402,
    n374,
    n425
  );


  nor
  g828
  (
    n680,
    n508,
    n473,
    n448,
    n260
  );


  nand
  g829
  (
    n1074,
    n610,
    n268,
    n189,
    n206
  );


  xnor
  g830
  (
    n933,
    n219,
    n585,
    n565,
    n235
  );


  xor
  g831
  (
    n753,
    n607,
    n196,
    n362,
    n316
  );


  and
  g832
  (
    n982,
    n592,
    n330,
    n530,
    n474
  );


  xnor
  g833
  (
    n887,
    n545,
    n405,
    n383,
    n290
  );


  nor
  g834
  (
    n886,
    n222,
    n440,
    n176,
    n568
  );


  xnor
  g835
  (
    n1137,
    n314,
    n517,
    n359,
    n448
  );


  nor
  g836
  (
    n862,
    n185,
    n450,
    n472,
    n510
  );


  or
  g837
  (
    n704,
    n663,
    n536,
    n545,
    n585
  );


  or
  g838
  (
    n833,
    n302,
    n548,
    n386,
    n598
  );


  and
  g839
  (
    n759,
    n289,
    n497,
    n653,
    n199
  );


  nor
  g840
  (
    n1120,
    n382,
    n511,
    n657,
    n576
  );


  and
  g841
  (
    n876,
    n291,
    n302,
    n408,
    n631
  );


  or
  g842
  (
    n1065,
    n437,
    n371,
    n348,
    n239
  );


  nor
  g843
  (
    n801,
    n408,
    n424,
    n409,
    n453
  );


  xor
  g844
  (
    n1095,
    n235,
    n652,
    n231,
    n194
  );


  nor
  g845
  (
    n840,
    n412,
    n549,
    n460,
    n428
  );


  or
  g846
  (
    n1070,
    n327,
    n556,
    n495,
    n469
  );


  nor
  g847
  (
    n825,
    n528,
    n280,
    n377
  );


  nor
  g848
  (
    n1041,
    n247,
    n262,
    n449,
    n466
  );


  or
  g849
  (
    n708,
    n623,
    n400,
    n214,
    n547
  );


  xnor
  g850
  (
    n1088,
    n531,
    n568,
    n294,
    n275
  );


  nand
  g851
  (
    n1149,
    n354,
    n644,
    n546,
    n571
  );


  nand
  g852
  (
    n1171,
    n365,
    n339,
    n332,
    n367
  );


  or
  g853
  (
    n942,
    n471,
    n445,
    n657,
    n356
  );


  xnor
  g854
  (
    n789,
    n198,
    n357,
    n477,
    n334
  );


  nor
  g855
  (
    n1035,
    n398,
    n323,
    n209,
    n343
  );


  nand
  g856
  (
    n1037,
    n543,
    n361,
    n329,
    n358
  );


  xor
  g857
  (
    n964,
    n491,
    n511,
    n270,
    n282
  );


  nand
  g858
  (
    n1001,
    n277,
    n593,
    n616,
    n522
  );


  or
  g859
  (
    n1144,
    n193,
    n254,
    n192,
    n168
  );


  or
  g860
  (
    n1133,
    n226,
    n628,
    n447,
    n563
  );


  xor
  g861
  (
    n808,
    n276,
    n609,
    n208,
    n273
  );


  and
  g862
  (
    n751,
    n366,
    n443,
    n417,
    n441
  );


  nor
  g863
  (
    n804,
    n308,
    n384,
    n518,
    n172
  );


  and
  g864
  (
    n1032,
    n384,
    n439,
    n520,
    n423
  );


  and
  g865
  (
    n795,
    n645,
    n335,
    n225,
    n329
  );


  nor
  g866
  (
    n1106,
    n459,
    n266,
    n324,
    n444
  );


  xor
  g867
  (
    n906,
    n270,
    n361,
    n470,
    n396
  );


  nand
  g868
  (
    n861,
    n431,
    n668,
    n163,
    n594
  );


  nand
  g869
  (
    n1107,
    n400,
    n461,
    n258,
    n512
  );


  or
  g870
  (
    n683,
    n594,
    n169,
    n605,
    n655
  );


  nor
  g871
  (
    n1017,
    n561,
    n223,
    n190,
    n382
  );


  nand
  g872
  (
    n1118,
    n180,
    n643,
    n557,
    n490
  );


  nand
  g873
  (
    n730,
    n344,
    n648,
    n230,
    n405
  );


  and
  g874
  (
    n1058,
    n433,
    n163,
    n429,
    n581
  );


  and
  g875
  (
    n790,
    n609,
    n232,
    n388,
    n182
  );


  or
  g876
  (
    n940,
    n617,
    n547,
    n291,
    n187
  );


  or
  g877
  (
    n709,
    n295,
    n470,
    n166,
    n233
  );


  and
  g878
  (
    n1159,
    n449,
    n322,
    n463,
    n293
  );


  xor
  g879
  (
    n766,
    n606,
    n242,
    n181,
    n204
  );


  or
  g880
  (
    n698,
    n245,
    n393,
    n654,
    n517
  );


  xor
  g881
  (
    n894,
    n549,
    n566,
    n562,
    n169
  );


  or
  g882
  (
    n746,
    n534,
    n387,
    n544,
    n561
  );


  nor
  g883
  (
    n1108,
    n656,
    n499,
    n572,
    n556
  );


  nand
  g884
  (
    n951,
    n540,
    n268,
    n483,
    n203
  );


  or
  g885
  (
    n715,
    n207,
    n442,
    n288,
    n569
  );


  nand
  g886
  (
    n1175,
    n357,
    n202,
    n271,
    n219
  );


  xnor
  g887
  (
    n1105,
    n503,
    n421,
    n533,
    n188
  );


  xor
  g888
  (
    n871,
    n563,
    n248,
    n558,
    n530
  );


  xor
  g889
  (
    n1064,
    n471,
    n161,
    n553,
    n453
  );


  xor
  g890
  (
    n687,
    n638,
    n178,
    n403,
    n663
  );


  nand
  g891
  (
    n760,
    n555,
    n213,
    n371,
    n190
  );


  xor
  g892
  (
    n1090,
    n203,
    n384,
    n353,
    n602
  );


  and
  g893
  (
    n691,
    n591,
    n398,
    n468,
    n623
  );


  xnor
  g894
  (
    n956,
    n496,
    n198,
    n491,
    n526
  );


  xor
  g895
  (
    n1077,
    n283,
    n259,
    n425,
    n404
  );


  xnor
  g896
  (
    n719,
    n211,
    n505,
    n192,
    n473
  );


  xnor
  g897
  (
    n1158,
    n399,
    n527,
    n664,
    n340
  );


  nand
  g898
  (
    n928,
    n222,
    n397,
    n638,
    n461
  );


  nand
  g899
  (
    KeyWire_0_1,
    n209,
    n428,
    n652,
    n561
  );


  and
  g900
  (
    n872,
    n420,
    n528,
    n535,
    n174
  );


  nand
  g901
  (
    n1173,
    n476,
    n427,
    n306,
    n347
  );


  xor
  g902
  (
    n696,
    n595,
    n376,
    n598
  );


  xnor
  g903
  (
    n1092,
    n515,
    n300,
    n604,
    n628
  );


  xor
  g904
  (
    n1027,
    n377,
    n366,
    n238,
    n167
  );


  nand
  g905
  (
    n1103,
    n597,
    n309,
    n624,
    n591
  );


  nor
  g906
  (
    n814,
    n644,
    n521,
    n642,
    n220
  );


  nand
  g907
  (
    n1139,
    n619,
    n355,
    n443,
    n408
  );


  and
  g908
  (
    n1003,
    n206,
    n235,
    n161,
    n282
  );


  and
  g909
  (
    n856,
    n360,
    n242,
    n318,
    n173
  );


  or
  g910
  (
    n950,
    n238,
    n210,
    n428,
    n423
  );


  xor
  g911
  (
    n976,
    n456,
    n275,
    n169,
    n279
  );


  nand
  g912
  (
    n748,
    n359,
    n181,
    n253,
    n667
  );


  or
  g913
  (
    n743,
    n193,
    n371,
    n649,
    n572
  );


  xor
  g914
  (
    n1056,
    n181,
    n329,
    n458,
    n326
  );


  nand
  g915
  (
    n962,
    n500,
    n261,
    n476,
    n607
  );


  and
  g916
  (
    n1022,
    n320,
    n200,
    n392,
    n285
  );


  and
  g917
  (
    n684,
    n266,
    n298,
    n237,
    n243
  );


  nor
  g918
  (
    n961,
    n181,
    n253,
    n372,
    n602
  );


  nand
  g919
  (
    n726,
    n377,
    n409,
    n311,
    n433
  );


  or
  g920
  (
    n937,
    n417,
    n535,
    n532,
    n335
  );


  or
  g921
  (
    n1177,
    n166,
    n261,
    n205,
    n448
  );


  or
  g922
  (
    n818,
    n180,
    n357,
    n192,
    n595
  );


  xor
  g923
  (
    n957,
    n162,
    n458,
    n649,
    n574
  );


  xor
  g924
  (
    n773,
    n569,
    n639,
    n333,
    n337
  );


  xnor
  g925
  (
    n984,
    n614,
    n607,
    n489,
    n657
  );


  nand
  g926
  (
    n1082,
    n499,
    n512,
    n295,
    n623
  );


  xnor
  g927
  (
    n830,
    n208,
    n554,
    n243,
    n170
  );


  nand
  g928
  (
    n958,
    n442,
    n287,
    n592,
    n204
  );


  xnor
  g929
  (
    n737,
    n619,
    n252,
    n357,
    n173
  );


  xnor
  g930
  (
    n819,
    n621,
    n397,
    n210,
    n223
  );


  nand
  g931
  (
    n815,
    n271,
    n449,
    n273,
    n573
  );


  xor
  g932
  (
    n860,
    n195,
    n582,
    n380,
    n645
  );


  xnor
  g933
  (
    n798,
    n637,
    n640,
    n407,
    n331
  );


  or
  g934
  (
    n972,
    n351,
    n221,
    n454,
    n627
  );


  xor
  g935
  (
    n1172,
    n231,
    n333,
    n262,
    n464
  );


  xor
  g936
  (
    n725,
    n529,
    n187,
    n293,
    n486
  );


  xnor
  g937
  (
    n794,
    n272,
    n251,
    n586,
    n424
  );


  nor
  g938
  (
    n980,
    n303,
    n646,
    n260,
    n459
  );


  nor
  g939
  (
    n874,
    n191,
    n625,
    n642,
    n313
  );


  and
  g940
  (
    n775,
    n426,
    n190,
    n324,
    n172
  );


  or
  g941
  (
    n909,
    n342,
    n316,
    n286,
    n321
  );


  or
  g942
  (
    n724,
    n370,
    n597,
    n550,
    n462
  );


  nor
  g943
  (
    n884,
    n513,
    n581,
    n311,
    n614
  );


  and
  g944
  (
    n835,
    n217,
    n476,
    n391,
    n406
  );


  or
  g945
  (
    n788,
    n460,
    n424,
    n177,
    n620
  );


  and
  g946
  (
    n1055,
    n343,
    n336,
    n408,
    n307
  );


  or
  g947
  (
    n713,
    n370,
    n555,
    n288,
    n579
  );


  or
  g948
  (
    n921,
    n596,
    n504,
    n326,
    n421
  );


  nor
  g949
  (
    n1048,
    n531,
    n463,
    n504,
    n459
  );


  xor
  g950
  (
    n1086,
    n646,
    n286,
    n528
  );


  xnor
  g951
  (
    n842,
    n632,
    n299,
    n382,
    n279
  );


  or
  g952
  (
    n847,
    n651,
    n334,
    n243,
    n345
  );


  xor
  g953
  (
    n1096,
    n485,
    n267,
    n385,
    n625
  );


  nand
  g954
  (
    n824,
    n486,
    n202,
    n281,
    n661
  );


  nor
  g955
  (
    n707,
    n244,
    n209,
    n497,
    n240
  );


  nand
  g956
  (
    n839,
    n513,
    n376,
    n662,
    n529
  );


  and
  g957
  (
    n1176,
    n464,
    n437,
    n653,
    n489
  );


  xnor
  g958
  (
    n1049,
    n487,
    n660,
    n329,
    n237
  );


  nand
  g959
  (
    n1015,
    n306,
    n251,
    n374,
    n266
  );


  and
  g960
  (
    n803,
    n208,
    n643,
    n426,
    n487
  );


  xnor
  g961
  (
    n735,
    n522,
    n425,
    n615,
    n244
  );


  xor
  g962
  (
    n1000,
    n307,
    n273,
    n304,
    n285
  );


  xnor
  g963
  (
    n1142,
    n234,
    n527,
    n540,
    n639
  );


  xor
  g964
  (
    n703,
    n615,
    n652,
    n578,
    n488
  );


  and
  g965
  (
    n736,
    n650,
    n478,
    n584,
    n534
  );


  nor
  g966
  (
    n875,
    n665,
    n385,
    n542,
    n228
  );


  and
  g967
  (
    n1063,
    n316,
    n482,
    n587,
    n274
  );


  and
  g968
  (
    n720,
    n264,
    n661,
    n267,
    n368
  );


  and
  g969
  (
    n1002,
    n315,
    n358,
    n215,
    n394
  );


  nand
  g970
  (
    n1078,
    n174,
    n580,
    n211,
    n411
  );


  nand
  g971
  (
    n859,
    n230,
    n180,
    n456,
    n573
  );


  nand
  g972
  (
    n1127,
    n325,
    n349,
    n662,
    n542
  );


  xor
  g973
  (
    n821,
    n178,
    n372,
    n531,
    n461
  );


  nand
  g974
  (
    n692,
    n418,
    n278,
    n293,
    n201
  );


  or
  g975
  (
    n702,
    n634,
    n494,
    n496,
    n515
  );


  xor
  g976
  (
    n843,
    n175,
    n634,
    n465,
    n324
  );


  or
  g977
  (
    n712,
    n175,
    n229,
    n457,
    n582
  );


  nand
  g978
  (
    n846,
    n481,
    n342,
    n296,
    n403
  );


  xnor
  g979
  (
    n805,
    n331,
    n187,
    n246,
    n223
  );


  and
  g980
  (
    n749,
    n398,
    n350,
    n530,
    n373
  );


  or
  g981
  (
    n993,
    n453,
    n284,
    n249,
    n337
  );


  nor
  g982
  (
    n898,
    n299,
    n474,
    n560,
    n309
  );


  xor
  g983
  (
    n885,
    n247,
    n653,
    n228,
    n426
  );


  xnor
  g984
  (
    n834,
    n627,
    n587,
    n667,
    n543
  );


  xnor
  g985
  (
    n892,
    n415,
    n187,
    n216,
    n474
  );


  xor
  g986
  (
    n1029,
    n303,
    n333,
    n643,
    n604
  );


  xnor
  g987
  (
    n806,
    n534,
    n287,
    n256,
    n584
  );


  and
  g988
  (
    n852,
    n287,
    n332,
    n600,
    n617
  );


  nand
  g989
  (
    n791,
    n195,
    n488,
    n648,
    n373
  );


  nor
  g990
  (
    n981,
    n241,
    n660,
    n289,
    n602
  );


  nand
  g991
  (
    n926,
    n619,
    n328,
    n510,
    n589
  );


  nor
  g992
  (
    n878,
    n535,
    n231,
    n584,
    n277
  );


  xnor
  g993
  (
    n915,
    n381,
    n528,
    n319,
    n212
  );


  xor
  g994
  (
    n817,
    n336,
    n215,
    n170,
    n594
  );


  nand
  g995
  (
    n939,
    n474,
    n636,
    n348,
    n353
  );


  or
  g996
  (
    n1013,
    n218,
    n340,
    n499,
    n507
  );


  xor
  g997
  (
    n802,
    n570,
    n322,
    n176,
    n390
  );


  xor
  g998
  (
    n904,
    n338,
    n391,
    n179,
    n378
  );


  xnor
  g999
  (
    n1134,
    n649,
    n435,
    n213,
    n368
  );


  nand
  g1000
  (
    n816,
    n519,
    n394,
    n354,
    n382
  );


  nand
  g1001
  (
    n780,
    n483,
    n580,
    n214,
    n186
  );


  xnor
  g1002
  (
    n971,
    n166,
    n496,
    n420,
    n226
  );


  and
  g1003
  (
    n1110,
    n593,
    n593,
    n653,
    n603
  );


  nor
  g1004
  (
    n745,
    n503,
    n613,
    n471,
    n311
  );


  nand
  g1005
  (
    n870,
    n326,
    n343,
    n481,
    n498
  );


  nand
  g1006
  (
    n963,
    n604,
    n442,
    n466,
    n558
  );


  nor
  g1007
  (
    n1030,
    n255,
    n485,
    n505,
    n519
  );


  and
  g1008
  (
    n917,
    n162,
    n634,
    n389,
    n553
  );


  xor
  g1009
  (
    n973,
    n546,
    n314,
    n577,
    n410
  );


  xnor
  g1010
  (
    n838,
    n301,
    n246,
    n541,
    n379
  );


  or
  g1011
  (
    n996,
    n327,
    n255,
    n504,
    n547
  );


  nor
  g1012
  (
    n1099,
    n368,
    n614,
    n386,
    n599
  );


  or
  g1013
  (
    n1004,
    n599,
    n314,
    n188,
    n484
  );


  xnor
  g1014
  (
    n952,
    n413,
    n199,
    n568,
    n274
  );


  and
  g1015
  (
    n1050,
    n423,
    n238,
    n363,
    n523
  );


  and
  g1016
  (
    n1073,
    n184,
    n264,
    n330,
    n589
  );


  nand
  g1017
  (
    n910,
    n271,
    n558,
    n657,
    n281
  );


  or
  g1018
  (
    n994,
    n355,
    n491,
    n503,
    n328
  );


  and
  g1019
  (
    n822,
    n283,
    n196,
    n587,
    n616
  );


  and
  g1020
  (
    n1143,
    n341,
    n436,
    n440,
    n581
  );


  nand
  g1021
  (
    n941,
    n240,
    n655,
    n541,
    n245
  );


  and
  g1022
  (
    n883,
    n317,
    n356,
    n205,
    n203
  );


  xnor
  g1023
  (
    n750,
    n566,
    n246,
    n630,
    n262
  );


  nand
  g1024
  (
    n1104,
    n200,
    n340,
    n272,
    n217
  );


  and
  g1025
  (
    n1132,
    n501,
    n310,
    n407,
    n481
  );


  nand
  g1026
  (
    n900,
    n338,
    n537,
    n430,
    n388
  );


  xnor
  g1027
  (
    n718,
    n535,
    n326,
    n189,
    n164
  );


  xor
  g1028
  (
    n1071,
    n298,
    n521,
    n658,
    n261
  );


  xor
  g1029
  (
    n1087,
    n609,
    n577,
    n228,
    n529
  );


  and
  g1030
  (
    n1169,
    n661,
    n509,
    n473,
    n591
  );


  xor
  g1031
  (
    n1069,
    n598,
    n454,
    n272,
    n606
  );


  and
  g1032
  (
    n792,
    n483,
    n167,
    n380,
    n289
  );


  xnor
  g1033
  (
    n873,
    n320,
    n480,
    n636,
    n656
  );


  xnor
  g1034
  (
    n914,
    n440,
    n298,
    n588,
    n162
  );


  xnor
  g1035
  (
    n1028,
    n654,
    n475,
    n347,
    n320
  );


  nor
  g1036
  (
    n1179,
    n437,
    n419,
    n168,
    n218
  );


  and
  g1037
  (
    n850,
    n285,
    n514,
    n625,
    n224
  );


  nand
  g1038
  (
    n970,
    n612,
    n290,
    n263,
    n627
  );


  nand
  g1039
  (
    n920,
    n264,
    n214,
    n479,
    n336
  );


  nand
  g1040
  (
    n913,
    n637,
    n171,
    n227,
    n177
  );


  or
  g1041
  (
    n991,
    n540,
    n497,
    n556,
    n245
  );


  xnor
  g1042
  (
    n975,
    n400,
    n631,
    n182,
    n350
  );


  and
  g1043
  (
    n763,
    n264,
    n434,
    n406,
    n455
  );


  or
  g1044
  (
    n1114,
    n638,
    n514,
    n182,
    n411
  );


  xnor
  g1045
  (
    n1168,
    n161,
    n618,
    n526,
    n224
  );


  and
  g1046
  (
    n844,
    n392,
    n383,
    n559,
    n390
  );


  xor
  g1047
  (
    n740,
    n229,
    n516,
    n183,
    n556
  );


  xor
  g1048
  (
    n700,
    n580,
    n640,
    n559,
    n506
  );


  xnor
  g1049
  (
    n676,
    n365,
    n468,
    n165,
    n560
  );


  and
  g1050
  (
    n1038,
    n500,
    n637,
    n464,
    n629
  );


  nand
  g1051
  (
    n1147,
    n193,
    n546,
    n669,
    n579
  );


  and
  g1052
  (
    n1116,
    n519,
    n588,
    n247,
    n433
  );


  nand
  g1053
  (
    n689,
    n268,
    n168,
    n318,
    n666
  );


  xnor
  g1054
  (
    n882,
    n536,
    n280,
    n183,
    n312
  );


  xnor
  g1055
  (
    n779,
    n313,
    n467,
    n197
  );


  nor
  g1056
  (
    n1112,
    n296,
    n224,
    n406,
    n177
  );


  nor
  g1057
  (
    n1080,
    n359,
    n299,
    n586,
    n454
  );


  xnor
  g1058
  (
    n752,
    n493,
    n526,
    n574,
    n275
  );


  or
  g1059
  (
    n729,
    n559,
    n292,
    n438,
    n335
  );


  nor
  g1060
  (
    n1018,
    n312,
    n633,
    n387,
    n290
  );


  nor
  g1061
  (
    n948,
    n353,
    n616,
    n171,
    n322
  );


  and
  g1062
  (
    n1034,
    n566,
    n195,
    n475,
    n310
  );


  xnor
  g1063
  (
    n1123,
    n439,
    n647,
    n669,
    n456
  );


  xor
  g1064
  (
    n965,
    n385,
    n305,
    n469,
    n403
  );


  xor
  g1065
  (
    n783,
    n504,
    n171,
    n590,
    n520
  );


  xor
  g1066
  (
    n678,
    n521,
    n341,
    n291,
    n270
  );


  nand
  g1067
  (
    n1083,
    n446,
    n646,
    n583,
    n365
  );


  nor
  g1068
  (
    n765,
    n507,
    n328,
    n244,
    n422
  );


  nor
  g1069
  (
    n877,
    n213,
    n353,
    n314,
    n647
  );


  nand
  g1070
  (
    n1145,
    n305,
    n521,
    n537,
    n460
  );


  nand
  g1071
  (
    n922,
    n393,
    n335,
    n626,
    n635
  );


  nand
  g1072
  (
    n927,
    n297,
    n346,
    n481,
    n369
  );


  and
  g1073
  (
    n1165,
    n646,
    n197,
    n279,
    n555
  );


  or
  g1074
  (
    n1085,
    n668,
    n252,
    n202,
    n511
  );


  xnor
  g1075
  (
    n699,
    n626,
    n233,
    n574,
    n472
  );


  nor
  g1076
  (
    n1098,
    n541,
    n290,
    n584,
    n377
  );


  xnor
  g1077
  (
    n1014,
    n441,
    n283,
    n485,
    n257
  );


  nor
  g1078
  (
    n1135,
    n452,
    n303,
    n217,
    n500
  );


  nand
  g1079
  (
    n934,
    n294,
    n234,
    n189,
    n641
  );


  and
  g1080
  (
    n1075,
    n211,
    n520,
    n517,
    n449
  );


  or
  g1081
  (
    n723,
    n279,
    n378,
    n246,
    n540
  );


  nand
  g1082
  (
    n827,
    n373,
    n669,
    n398,
    n376
  );


  or
  g1083
  (
    n857,
    n664,
    n618,
    n249,
    n479
  );


  xor
  g1084
  (
    n1036,
    n438,
    n434,
    n623,
    n451
  );


  or
  g1085
  (
    n929,
    n605,
    n523,
    n174,
    n312
  );


  or
  g1086
  (
    n674,
    n341,
    n346,
    n488,
    n206
  );


  xor
  g1087
  (
    n968,
    n455,
    n362,
    n551,
    n617
  );


  xor
  g1088
  (
    n1155,
    n330,
    n656,
    n509,
    n562
  );


  xnor
  g1089
  (
    n694,
    n511,
    n370,
    n287,
    n185
  );


  and
  g1090
  (
    n925,
    n588,
    n221,
    n379,
    n220
  );


  nor
  g1091
  (
    n769,
    n232,
    n188,
    n509,
    n362
  );


  xnor
  g1092
  (
    n690,
    n412,
    n630,
    n374,
    n372
  );


  xnor
  g1093
  (
    n897,
    n624,
    n401,
    n610,
    n532
  );


  xor
  g1094
  (
    n983,
    n254,
    n644,
    n523,
    n482
  );


  or
  g1095
  (
    n799,
    n399,
    n380,
    n387,
    n583
  );


  and
  g1096
  (
    n1178,
    n402,
    n641,
    n634,
    n292
  );


  nand
  g1097
  (
    n733,
    n364,
    n648,
    n440,
    n321
  );


  or
  g1098
  (
    n943,
    n551,
    n658,
    n514,
    n563
  );


  xor
  g1099
  (
    n767,
    n478,
    n216,
    n245,
    n446
  );


  xor
  g1100
  (
    n1113,
    n241,
    n415,
    n664,
    n620
  );


  and
  g1101
  (
    n1131,
    n577,
    n395,
    n652,
    n207
  );


  nand
  g1102
  (
    n705,
    n502,
    n651,
    n254,
    n363
  );


  and
  g1103
  (
    n1067,
    n550,
    n232,
    n210,
    n325
  );


  nor
  g1104
  (
    n1150,
    n352,
    n460,
    n249,
    n645
  );


  and
  g1105
  (
    n768,
    n577,
    n532,
    n179,
    n349
  );


  nand
  g1106
  (
    n1046,
    n393,
    n346,
    n297,
    n437
  );


  nand
  g1107
  (
    n693,
    n208,
    n224,
    n505,
    n315
  );


  nor
  g1108
  (
    n1162,
    n197,
    n343,
    n221,
    n498
  );


  and
  g1109
  (
    n855,
    n324,
    n196,
    n635,
    n427
  );


  or
  g1110
  (
    n960,
    n379,
    n362,
    n292,
    n642
  );


  nor
  g1111
  (
    n889,
    n389,
    n659,
    n265,
    n222
  );


  xnor
  g1112
  (
    n1043,
    n453,
    n229,
    n502,
    n390
  );


  and
  g1113
  (
    n1019,
    n635,
    n274,
    n574,
    n459
  );


  xnor
  g1114
  (
    n796,
    n369,
    n615,
    n456,
    n256
  );


  and
  g1115
  (
    n953,
    n241,
    n370,
    n212,
    n519
  );


  or
  g1116
  (
    n832,
    n215,
    n304,
    n607,
    n422
  );


  xor
  g1117
  (
    n738,
    n624,
    n269,
    n228,
    n268
  );


  and
  g1118
  (
    n829,
    n532,
    n337,
    n354,
    n375
  );


  nand
  g1119
  (
    n865,
    n445,
    n659,
    n559,
    n419
  );


  or
  g1120
  (
    n1138,
    n436,
    n638,
    n513,
    n216
  );


  nor
  g1121
  (
    n1072,
    n468,
    n664,
    n407,
    n520
  );


  nor
  g1122
  (
    n706,
    n596,
    n317,
    n367,
    n445
  );


  xor
  g1123
  (
    n899,
    n240,
    n300,
    n323,
    n258
  );


  xnor
  g1124
  (
    n959,
    n570,
    n452,
    n243,
    n488
  );


  or
  g1125
  (
    n869,
    n478,
    n263,
    n277,
    n537
  );


  xor
  g1126
  (
    n895,
    n278,
    n501,
    n463,
    n175
  );


  nor
  g1127
  (
    n1012,
    n344,
    n388,
    n259,
    n570
  );


  or
  g1128
  (
    n1079,
    n538,
    n276,
    n269,
    n651
  );


  xnor
  g1129
  (
    n772,
    n514,
    n431,
    n386,
    n241
  );


  nor
  g1130
  (
    n710,
    n465,
    n594,
    n310,
    n482
  );


  xor
  g1131
  (
    n1011,
    n466,
    n369,
    n307,
    n250
  );


  nor
  g1132
  (
    n919,
    n178,
    n413,
    n640,
    n173
  );


  nor
  g1133
  (
    n1111,
    n433,
    n374,
    n413,
    n571
  );


  xor
  g1134
  (
    n1156,
    n305,
    n538,
    n269,
    n286
  );


  nor
  g1135
  (
    n854,
    n586,
    n345,
    n608
  );


  xor
  g1136
  (
    n1040,
    n525,
    n423,
    n650,
    n170
  );


  nand
  g1137
  (
    KeyWire_0_12,
    n503,
    n421,
    n464,
    n573
  );


  xor
  g1138
  (
    n781,
    n564,
    n446,
    n552,
    n539
  );


  xor
  g1139
  (
    n813,
    n186,
    n654,
    n431,
    n613
  );


  xnor
  g1140
  (
    n1010,
    n282,
    n572,
    n419,
    n371
  );


  nand
  g1141
  (
    n954,
    n274,
    n568,
    n430,
    n401
  );


  xor
  g1142
  (
    n845,
    n295,
    n351,
    n375,
    n327
  );


  nand
  g1143
  (
    n1089,
    n632,
    n571,
    n308,
    n212
  );


  xor
  g1144
  (
    n1097,
    n420,
    n189,
    n611,
    n435
  );


  nor
  g1145
  (
    n757,
    n225,
    n632,
    n313,
    n458
  );


  nand
  g1146
  (
    n1140,
    n366,
    n641,
    n538,
    n196
  );


  nor
  g1147
  (
    n1125,
    n669,
    n562,
    n180,
    n200
  );


  nor
  g1148
  (
    n881,
    n448,
    n318,
    n463,
    n234
  );


  not
  g1149
  (
    n1184,
    n698
  );


  not
  g1150
  (
    n1191,
    n700
  );


  not
  g1151
  (
    n1188,
    n692
  );


  buf
  g1152
  (
    n1193,
    n693
  );


  buf
  g1153
  (
    n1185,
    n677
  );


  buf
  g1154
  (
    n1195,
    n689
  );


  buf
  g1155
  (
    n1187,
    n679
  );


  buf
  g1156
  (
    n1199,
    n690
  );


  not
  g1157
  (
    n1186,
    n678
  );


  not
  g1158
  (
    n1194,
    n675
  );


  not
  g1159
  (
    n1198,
    n684
  );


  buf
  g1160
  (
    n1202,
    n694
  );


  not
  g1161
  (
    n1192,
    n688
  );


  buf
  g1162
  (
    n1190,
    n695
  );


  not
  g1163
  (
    n1182,
    n699
  );


  not
  g1164
  (
    n1189,
    n682
  );


  not
  g1165
  (
    n1197,
    n687
  );


  not
  g1166
  (
    n1200,
    n683
  );


  nand
  g1167
  (
    n1183,
    n680,
    n691
  );


  and
  g1168
  (
    n1196,
    n674,
    n681,
    n685,
    n697
  );


  nand
  g1169
  (
    n1201,
    n696,
    n686,
    n673,
    n676
  );


  buf
  g1170
  (
    n1203,
    n1182
  );


  buf
  g1171
  (
    n1204,
    n1182
  );


  not
  g1172
  (
    n1212,
    n1203
  );


  buf
  g1173
  (
    n1206,
    n1204
  );


  buf
  g1174
  (
    n1210,
    n1203
  );


  not
  g1175
  (
    n1205,
    n1204
  );


  buf
  g1176
  (
    n1209,
    n1204
  );


  not
  g1177
  (
    n1211,
    n701
  );


  not
  g1178
  (
    n1207,
    n1203
  );


  or
  g1179
  (
    n1208,
    n1204,
    n1203,
    n702
  );


  buf
  g1180
  (
    n1244,
    n1206
  );


  buf
  g1181
  (
    n1215,
    n1208
  );


  buf
  g1182
  (
    n1241,
    n1206
  );


  buf
  g1183
  (
    n1227,
    n1207
  );


  buf
  g1184
  (
    n1225,
    n1208
  );


  not
  g1185
  (
    n1218,
    n1207
  );


  buf
  g1186
  (
    n1242,
    n1211
  );


  not
  g1187
  (
    n1216,
    n1209
  );


  buf
  g1188
  (
    n1230,
    n1208
  );


  buf
  g1189
  (
    n1234,
    n1212
  );


  buf
  g1190
  (
    n1213,
    n1205
  );


  not
  g1191
  (
    n1222,
    n1209
  );


  not
  g1192
  (
    n1232,
    n1212
  );


  not
  g1193
  (
    n1214,
    n1205
  );


  buf
  g1194
  (
    n1224,
    n1210
  );


  buf
  g1195
  (
    n1243,
    n1205
  );


  buf
  g1196
  (
    n1235,
    n1211
  );


  not
  g1197
  (
    n1217,
    n1212
  );


  buf
  g1198
  (
    n1220,
    n1207
  );


  buf
  g1199
  (
    n1238,
    n1210
  );


  not
  g1200
  (
    n1240,
    n1209
  );


  buf
  g1201
  (
    n1226,
    n1207
  );


  not
  g1202
  (
    n1233,
    n1209
  );


  buf
  g1203
  (
    n1219,
    n1210
  );


  buf
  g1204
  (
    KeyWire_0_11,
    n1206
  );


  not
  g1205
  (
    n1229,
    n1211
  );


  not
  g1206
  (
    n1228,
    n1210
  );


  not
  g1207
  (
    n1239,
    n1206
  );


  not
  g1208
  (
    n1236,
    n1211
  );


  not
  g1209
  (
    n1231,
    n1208
  );


  not
  g1210
  (
    n1221,
    n1205
  );


  buf
  g1211
  (
    n1223,
    n1212
  );


  not
  g1212
  (
    n1245,
    n1216
  );


  buf
  g1213
  (
    n1253,
    n1216
  );


  not
  g1214
  (
    n1252,
    n1216
  );


  not
  g1215
  (
    n1248,
    n1214
  );


  buf
  g1216
  (
    n1251,
    n1215
  );


  buf
  g1217
  (
    n1254,
    n1214
  );


  not
  g1218
  (
    n1247,
    n1213
  );


  buf
  g1219
  (
    n1246,
    n1216
  );


  buf
  g1220
  (
    n1249,
    n1213
  );


  not
  g1221
  (
    n1250,
    n1215
  );


  not
  g1222
  (
    n1262,
    n1249
  );


  buf
  g1223
  (
    n1264,
    n1249
  );


  buf
  g1224
  (
    n1266,
    n1247
  );


  not
  g1225
  (
    n1268,
    n1250
  );


  not
  g1226
  (
    n1277,
    n1250
  );


  not
  g1227
  (
    n1260,
    n1246
  );


  not
  g1228
  (
    KeyWire_0_10,
    n1248
  );


  buf
  g1229
  (
    n1263,
    n1246
  );


  not
  g1230
  (
    n1273,
    n1249
  );


  buf
  g1231
  (
    n1278,
    n1247
  );


  not
  g1232
  (
    n1275,
    n1250
  );


  not
  g1233
  (
    n1276,
    n1248
  );


  not
  g1234
  (
    n1256,
    n1248
  );


  buf
  g1235
  (
    n1269,
    n1245
  );


  not
  g1236
  (
    n1272,
    n1246
  );


  not
  g1237
  (
    n1257,
    n1248
  );


  buf
  g1238
  (
    n1270,
    n1245
  );


  not
  g1239
  (
    n1255,
    n1247
  );


  buf
  g1240
  (
    n1271,
    n1245
  );


  buf
  g1241
  (
    n1259,
    n1249
  );


  buf
  g1242
  (
    n1258,
    n1246
  );


  buf
  g1243
  (
    n1274,
    n1245
  );


  not
  g1244
  (
    n1267,
    n1247
  );


  not
  g1245
  (
    n1265,
    n1250
  );


  not
  g1246
  (
    n1290,
    n1255
  );


  not
  g1247
  (
    n1293,
    n1255
  );


  buf
  g1248
  (
    n1283,
    n1255
  );


  buf
  g1249
  (
    n1296,
    n1261
  );


  not
  g1250
  (
    n1302,
    n1261
  );


  not
  g1251
  (
    n1295,
    n1258
  );


  buf
  g1252
  (
    n1304,
    n1258
  );


  not
  g1253
  (
    n1306,
    n1257
  );


  not
  g1254
  (
    n1279,
    n1262
  );


  buf
  g1255
  (
    n1280,
    n1256
  );


  not
  g1256
  (
    n1282,
    n1257
  );


  buf
  g1257
  (
    n1297,
    n1261
  );


  not
  g1258
  (
    n1281,
    n1262
  );


  not
  g1259
  (
    n1289,
    n1255
  );


  buf
  g1260
  (
    n1294,
    n1256
  );


  buf
  g1261
  (
    n1284,
    n1260
  );


  not
  g1262
  (
    n1303,
    n1259
  );


  not
  g1263
  (
    n1307,
    n1256
  );


  buf
  g1264
  (
    n1286,
    n1259
  );


  buf
  g1265
  (
    n1305,
    n1256
  );


  not
  g1266
  (
    n1287,
    n1260
  );


  buf
  g1267
  (
    n1298,
    n1260
  );


  buf
  g1268
  (
    n1299,
    n1258
  );


  not
  g1269
  (
    n1301,
    n1260
  );


  buf
  g1270
  (
    n1300,
    n1259
  );


  buf
  g1271
  (
    n1308,
    n1258
  );


  not
  g1272
  (
    n1291,
    n1257
  );


  not
  g1273
  (
    n1292,
    n1259
  );


  buf
  g1274
  (
    n1288,
    n1257
  );


  not
  g1275
  (
    n1285,
    n1261
  );


  xor
  g1276
  (
    n1309,
    n703,
    n704,
    n705,
    n1279
  );


  buf
  g1277
  (
    n1310,
    n1309
  );


  not
  g1278
  (
    n1311,
    n1309
  );


  or
  g1279
  (
    n1313,
    n1311,
    n706,
    n712,
    n1251
  );


  xnor
  g1280
  (
    n1312,
    n708,
    n1251
  );


  xnor
  g1281
  (
    n1315,
    n711,
    n714,
    n1253,
    n1310
  );


  or
  g1282
  (
    n1314,
    n1252,
    n1252,
    n1311,
    n1310
  );


  and
  g1283
  (
    n1317,
    n707,
    n710,
    n1252,
    n1253
  );


  and
  g1284
  (
    n1318,
    n713,
    n1253,
    n715,
    n709
  );


  xnor
  g1285
  (
    n1316,
    n1311,
    n1311,
    n1252,
    n1310
  );


  not
  g1286
  (
    n1327,
    n1312
  );


  buf
  g1287
  (
    n1328,
    n1313
  );


  buf
  g1288
  (
    n1325,
    n1313
  );


  not
  g1289
  (
    n1324,
    n1312
  );


  not
  g1290
  (
    n1322,
    n1314
  );


  buf
  g1291
  (
    n1320,
    n1315
  );


  not
  g1292
  (
    n1319,
    n1315
  );


  buf
  g1293
  (
    n1323,
    n1315
  );


  buf
  g1294
  (
    n1321,
    n1315
  );


  buf
  g1295
  (
    n1326,
    n1314
  );


  nor
  g1296
  (
    n1360,
    n734,
    n766,
    n1324
  );


  xnor
  g1297
  (
    n1357,
    n805,
    n756,
    n822,
    n754
  );


  nor
  g1298
  (
    n1365,
    n1326,
    n1325,
    n828,
    n719
  );


  xnor
  g1299
  (
    n1364,
    n1321,
    n731,
    n777,
    n797
  );


  nand
  g1300
  (
    n1330,
    n832,
    n1322,
    n816,
    n1326
  );


  and
  g1301
  (
    n1359,
    n736,
    n831,
    n818,
    n774
  );


  and
  g1302
  (
    n1340,
    n727,
    n765,
    n1321,
    n1328
  );


  or
  g1303
  (
    n1346,
    n770,
    n746,
    n758,
    n739
  );


  nor
  g1304
  (
    n1354,
    n1319,
    n763,
    n771,
    n761
  );


  xor
  g1305
  (
    n1347,
    n809,
    n718,
    n823,
    n716
  );


  or
  g1306
  (
    n1336,
    n721,
    n751,
    n795,
    n800
  );


  and
  g1307
  (
    n1352,
    n740,
    n729,
    n1328,
    n819
  );


  nor
  g1308
  (
    n1334,
    n742,
    n1323,
    n1324,
    n1320
  );


  or
  g1309
  (
    n1358,
    n829,
    n775,
    n807,
    n748
  );


  xnor
  g1310
  (
    n1333,
    n738,
    n735,
    n798,
    n1320
  );


  xnor
  g1311
  (
    n1338,
    n1325,
    n757,
    n722,
    n782
  );


  and
  g1312
  (
    n1335,
    n813,
    n737,
    n835,
    n827
  );


  nand
  g1313
  (
    n1368,
    n790,
    n785,
    n755,
    n783
  );


  or
  g1314
  (
    n1345,
    n744,
    n724,
    n747,
    n1327
  );


  xnor
  g1315
  (
    n1341,
    n825,
    n787,
    n812,
    n804
  );


  xnor
  g1316
  (
    KeyWire_0_3,
    n802,
    n814,
    n834,
    n1325
  );


  and
  g1317
  (
    n1356,
    n799,
    n817,
    n792,
    n801
  );


  and
  g1318
  (
    n1351,
    n796,
    n810,
    n1321,
    n1323
  );


  or
  g1319
  (
    n1332,
    n793,
    n772,
    n1327,
    n788
  );


  and
  g1320
  (
    n1329,
    n1322,
    n778,
    n1319,
    n1323
  );


  xnor
  g1321
  (
    n1344,
    n820,
    n1320,
    n773,
    n745
  );


  nor
  g1322
  (
    n1355,
    n764,
    n759,
    n743,
    n1319
  );


  or
  g1323
  (
    n1366,
    n768,
    n794,
    n833,
    n760
  );


  and
  g1324
  (
    n1363,
    n1321,
    n826,
    n1320,
    n1322
  );


  nor
  g1325
  (
    n1348,
    n769,
    n1327,
    n723,
    n803
  );


  xnor
  g1326
  (
    n1331,
    n815,
    n791,
    n780,
    n776
  );


  nand
  g1327
  (
    n1337,
    n1325,
    n730,
    n786,
    n779
  );


  xnor
  g1328
  (
    n1350,
    n789,
    n1327,
    n784,
    n1319
  );


  xor
  g1329
  (
    n1343,
    n1326,
    n749,
    n808,
    n753
  );


  xor
  g1330
  (
    n1342,
    n1324,
    n1322,
    n1326,
    n750
  );


  nor
  g1331
  (
    n1362,
    n1328,
    n811,
    n732,
    n830
  );


  nor
  g1332
  (
    n1361,
    n741,
    n733,
    n821,
    n781
  );


  xor
  g1333
  (
    n1349,
    n767,
    n806,
    n762,
    n717
  );


  and
  g1334
  (
    n1367,
    n752,
    n1328,
    n725,
    n728
  );


  xor
  g1335
  (
    n1339,
    n720,
    n726,
    n1323,
    n824
  );


  not
  g1336
  (
    n1370,
    n1330
  );


  not
  g1337
  (
    n1369,
    n1329
  );


  or
  g1338
  (
    n1371,
    n837,
    n836
  );


  and
  g1339
  (
    n1372,
    n849,
    n1369,
    n842,
    n845
  );


  xor
  g1340
  (
    n1373,
    n848,
    n847,
    n838,
    n843
  );


  and
  g1341
  (
    n1375,
    n1370,
    n844,
    n846,
    n841
  );


  xnor
  g1342
  (
    n1374,
    n839,
    n1371,
    n840
  );


  nor
  g1343
  (
    n1377,
    n670,
    n672,
    n860,
    n854
  );


  or
  g1344
  (
    n1385,
    n1375,
    n1373,
    n852
  );


  xor
  g1345
  (
    n1381,
    n670,
    n1372,
    n850,
    n1279
  );


  xnor
  g1346
  (
    n1384,
    n670,
    n1316,
    n857,
    n1375
  );


  xor
  g1347
  (
    n1379,
    n864,
    n1374,
    n670
  );


  xnor
  g1348
  (
    n1382,
    n671,
    n855,
    n1375,
    n1373
  );


  and
  g1349
  (
    n1386,
    n862,
    n1317,
    n1316,
    n1318
  );


  or
  g1350
  (
    n1376,
    n853,
    n671,
    n863,
    n1374
  );


  nand
  g1351
  (
    KeyWire_0_14,
    n1372,
    n1317,
    n858
  );


  and
  g1352
  (
    n1380,
    n1375,
    n672,
    n861,
    n1317
  );


  and
  g1353
  (
    n1378,
    n671,
    n859,
    n1374,
    n1316
  );


  xnor
  g1354
  (
    n1387,
    n1316,
    n851,
    n671,
    n856
  );


  not
  g1355
  (
    n1388,
    n1377
  );


  buf
  g1356
  (
    n1390,
    n1378
  );


  not
  g1357
  (
    n1392,
    n1380
  );


  not
  g1358
  (
    n1391,
    n1376
  );


  buf
  g1359
  (
    n1393,
    n1379
  );


  not
  g1360
  (
    n1389,
    n1381
  );


  not
  g1361
  (
    n1400,
    n1392
  );


  not
  g1362
  (
    n1413,
    n872
  );


  buf
  g1363
  (
    n1407,
    n1389
  );


  not
  g1364
  (
    n1409,
    n874
  );


  not
  g1365
  (
    n1401,
    n1390
  );


  not
  g1366
  (
    n1404,
    n1391
  );


  not
  g1367
  (
    n1396,
    n1392
  );


  buf
  g1368
  (
    n1405,
    n875
  );


  buf
  g1369
  (
    n1403,
    n871
  );


  buf
  g1370
  (
    n1416,
    n865
  );


  buf
  g1371
  (
    n1411,
    n1390
  );


  xor
  g1372
  (
    n1395,
    n901,
    n1391,
    n900
  );


  nand
  g1373
  (
    n1417,
    n866,
    n897,
    n1391,
    n882
  );


  and
  g1374
  (
    n1406,
    n1389,
    n881,
    n885,
    n889
  );


  and
  g1375
  (
    n1415,
    n888,
    n1388,
    n891,
    n1391
  );


  or
  g1376
  (
    n1399,
    n869,
    n1389,
    n1392,
    n1393
  );


  xor
  g1377
  (
    n1402,
    n902,
    n1390,
    n892,
    n880
  );


  xor
  g1378
  (
    n1412,
    n884,
    n873,
    n1393,
    n877
  );


  nor
  g1379
  (
    n1397,
    n870,
    n1388,
    n1390,
    n883
  );


  and
  g1380
  (
    n1398,
    n896,
    n1393,
    n887,
    n898
  );


  or
  g1381
  (
    n1410,
    n890,
    n878,
    n879,
    n867
  );


  xor
  g1382
  (
    n1408,
    n868,
    n886,
    n899,
    n876
  );


  nor
  g1383
  (
    n1394,
    n1393,
    n893,
    n1389,
    n895
  );


  nor
  g1384
  (
    n1414,
    n894,
    n1392,
    n1388
  );


  buf
  g1385
  (
    n1438,
    n1402
  );


  not
  g1386
  (
    n1506,
    n1400
  );


  buf
  g1387
  (
    n1468,
    n1404
  );


  buf
  g1388
  (
    n1502,
    n1201
  );


  not
  g1389
  (
    n1510,
    n1190
  );


  not
  g1390
  (
    n1507,
    n1197
  );


  not
  g1391
  (
    n1501,
    n1414
  );


  buf
  g1392
  (
    n1462,
    n1275
  );


  buf
  g1393
  (
    n1491,
    n1269
  );


  buf
  g1394
  (
    n1423,
    n1193
  );


  buf
  g1395
  (
    n1434,
    n1192
  );


  buf
  g1396
  (
    n1421,
    n1417
  );


  buf
  g1397
  (
    n1467,
    n1331
  );


  not
  g1398
  (
    n1483,
    n1273
  );


  not
  g1399
  (
    n1444,
    n1267
  );


  buf
  g1400
  (
    n1459,
    n1332
  );


  not
  g1401
  (
    n1500,
    n1196
  );


  not
  g1402
  (
    n1429,
    n1263
  );


  not
  g1403
  (
    n1439,
    n1195
  );


  buf
  g1404
  (
    n1498,
    n1412
  );


  buf
  g1405
  (
    n1503,
    n1399
  );


  not
  g1406
  (
    n1418,
    n1274
  );


  not
  g1407
  (
    n1494,
    n1333
  );


  not
  g1408
  (
    n1422,
    n1416
  );


  not
  g1409
  (
    n1505,
    n1411
  );


  buf
  g1410
  (
    n1458,
    n1415
  );


  not
  g1411
  (
    n1447,
    n1386
  );


  buf
  g1412
  (
    n1442,
    n1277
  );


  not
  g1413
  (
    n1497,
    n1271
  );


  buf
  g1414
  (
    n1449,
    n1200
  );


  not
  g1415
  (
    n1490,
    n1187
  );


  not
  g1416
  (
    n1476,
    n1200
  );


  buf
  g1417
  (
    n1493,
    n1409
  );


  not
  g1418
  (
    n1424,
    n1275
  );


  buf
  g1419
  (
    n1441,
    n1412
  );


  buf
  g1420
  (
    n1477,
    n1264
  );


  buf
  g1421
  (
    n1445,
    n1383
  );


  not
  g1422
  (
    n1482,
    n1398
  );


  buf
  g1423
  (
    n1457,
    n1218
  );


  not
  g1424
  (
    n1486,
    n1413
  );


  not
  g1425
  (
    n1426,
    n1272
  );


  not
  g1426
  (
    n1463,
    n1200
  );


  not
  g1427
  (
    n1443,
    n1335
  );


  xnor
  g1428
  (
    n1487,
    n1272,
    n1264
  );


  and
  g1429
  (
    n1455,
    n1403,
    n1191,
    n1264
  );


  and
  g1430
  (
    n1479,
    n1269,
    n1384,
    n1218
  );


  and
  g1431
  (
    n1472,
    n1267,
    n1275,
    n1218,
    n1406
  );


  and
  g1432
  (
    n1450,
    n1413,
    n1274,
    n1415,
    n1411
  );


  xor
  g1433
  (
    n1428,
    n1269,
    n1268,
    n1270,
    n1334
  );


  nand
  g1434
  (
    n1469,
    n1187,
    n1273,
    n1399,
    n1411
  );


  xnor
  g1435
  (
    n1478,
    n1395,
    n1401,
    n1417,
    n1382
  );


  xor
  g1436
  (
    n1466,
    n1184,
    n1334,
    n1412,
    n1395
  );


  xor
  g1437
  (
    n1465,
    n1394,
    n1401,
    n1272,
    n1269
  );


  and
  g1438
  (
    n1508,
    n1404,
    n1394,
    n1278,
    n1414
  );


  and
  g1439
  (
    n1437,
    n1404,
    n1263,
    n1202,
    n1417
  );


  or
  g1440
  (
    n1475,
    n1333,
    n1278,
    n1411,
    n1194
  );


  xor
  g1441
  (
    n1499,
    n1266,
    n1268,
    n1414,
    n1399
  );


  xor
  g1442
  (
    n1456,
    n1277,
    n1405,
    n1414,
    n1416
  );


  nand
  g1443
  (
    n1511,
    n1273,
    n1408,
    n1270,
    n1195
  );


  nor
  g1444
  (
    n1430,
    n1398,
    n1405,
    n1409,
    n1272
  );


  xor
  g1445
  (
    n1473,
    n1189,
    n1274,
    n1402,
    n1266
  );


  nand
  g1446
  (
    n1509,
    n1406,
    n1271,
    n1397,
    n1410
  );


  or
  g1447
  (
    n1420,
    n1413,
    n1413,
    n1202,
    n1416
  );


  or
  g1448
  (
    n1464,
    n1405,
    n1407,
    n1186,
    n1382
  );


  or
  g1449
  (
    n1454,
    n1188,
    n1267,
    n1217,
    n1394
  );


  xor
  g1450
  (
    n1432,
    n1186,
    n1276,
    n1397,
    n1396
  );


  or
  g1451
  (
    n1496,
    n1397,
    n1201,
    n1415,
    n1412
  );


  xnor
  g1452
  (
    n1433,
    n1194,
    n1266,
    n1398,
    n1415
  );


  xnor
  g1453
  (
    n1485,
    n1385,
    n1198,
    n1408,
    n1407
  );


  nand
  g1454
  (
    n1440,
    n1271,
    n1264,
    n1410,
    n1394
  );


  xnor
  g1455
  (
    KeyWire_0_13,
    n1263,
    n1265,
    n1318,
    n1266
  );


  nor
  g1456
  (
    n1446,
    n1200,
    n1403,
    n1278,
    n1400
  );


  and
  g1457
  (
    n1448,
    n1386,
    n1185,
    n1268,
    n1183
  );


  xnor
  g1458
  (
    n1480,
    n1401,
    n1196,
    n1277,
    n1397
  );


  and
  g1459
  (
    n1419,
    n1400,
    n1184,
    n1403,
    n1395
  );


  xor
  g1460
  (
    n1461,
    n1335,
    n1263,
    n1330,
    n1318
  );


  nor
  g1461
  (
    n1427,
    n1402,
    n1383,
    n1267,
    n1202
  );


  nand
  g1462
  (
    n1425,
    n1417,
    n1185,
    n1406,
    n1201
  );


  xor
  g1463
  (
    n1488,
    n1265,
    n1193,
    n1396,
    n1407
  );


  nor
  g1464
  (
    n1435,
    n1268,
    n1199,
    n1262
  );


  xor
  g1465
  (
    n1453,
    n1183,
    n1402,
    n1410,
    n1273
  );


  nor
  g1466
  (
    n1451,
    n1270,
    n1331,
    n1387,
    n1318
  );


  nor
  g1467
  (
    n1460,
    n1399,
    n1197,
    n1409,
    n1188
  );


  and
  g1468
  (
    n1484,
    n1262,
    n1407,
    n1332,
    n1192
  );


  nand
  g1469
  (
    n1431,
    n1409,
    n1265,
    n1189,
    n903
  );


  nand
  g1470
  (
    n1504,
    n1387,
    n1385,
    n1278,
    n1217
  );


  nand
  g1471
  (
    n1492,
    n1191,
    n1408,
    n1190,
    n1410
  );


  or
  g1472
  (
    n1436,
    n1217,
    n1416,
    n1276,
    n1274
  );


  xor
  g1473
  (
    n1489,
    n1395,
    n1270,
    n1217,
    n1276
  );


  xor
  g1474
  (
    n1495,
    n1398,
    n1275,
    n1271,
    n1406
  );


  xnor
  g1475
  (
    n1471,
    n1396,
    n1384,
    n1401,
    n1405
  );


  or
  g1476
  (
    n1452,
    n1218,
    n1404,
    n1408,
    n1265
  );


  nor
  g1477
  (
    n1474,
    n1396,
    n1403,
    n1198,
    n1276
  );


  nor
  g1478
  (
    n1470,
    n1202,
    n1400,
    n1277,
    n1201
  );


  xnor
  g1479
  (
    n1528,
    n907,
    n917,
    n1433,
    n921
  );


  xor
  g1480
  (
    n1525,
    n1430,
    n1421,
    n1426,
    n1447
  );


  xnor
  g1481
  (
    n1513,
    n923,
    n1418,
    n1423,
    n1443
  );


  nand
  g1482
  (
    n1526,
    n920,
    n925,
    n1442,
    n1428
  );


  nand
  g1483
  (
    n1523,
    n1432,
    n928,
    n1441,
    n1443
  );


  xnor
  g1484
  (
    n1518,
    n1429,
    n1431,
    n1446,
    n1436
  );


  or
  g1485
  (
    n1522,
    n1427,
    n1437,
    n1422
  );


  xnor
  g1486
  (
    n1527,
    n904,
    n1421,
    n1439,
    n1419
  );


  and
  g1487
  (
    n1514,
    n909,
    n1442,
    n911,
    n1438
  );


  xnor
  g1488
  (
    n1520,
    n1438,
    n1445,
    n1447,
    n931
  );


  or
  g1489
  (
    n1521,
    n1428,
    n1420,
    n1430,
    n1444
  );


  xor
  g1490
  (
    n1516,
    n924,
    n922,
    n1419,
    n1440
  );


  nor
  g1491
  (
    n1524,
    n1422,
    n1434,
    n905,
    n935
  );


  or
  g1492
  (
    n1515,
    n916,
    n1434,
    n1440,
    n919
  );


  xor
  g1493
  (
    n1533,
    n1446,
    n1431,
    n1436,
    n1445
  );


  and
  g1494
  (
    n1531,
    n1418,
    n906,
    n1420,
    n1435
  );


  xnor
  g1495
  (
    n1534,
    n1435,
    n913,
    n915,
    n1423
  );


  or
  g1496
  (
    n1512,
    n926,
    n1424,
    n908
  );


  xor
  g1497
  (
    n1517,
    n932,
    n912,
    n1427,
    n927
  );


  xnor
  g1498
  (
    n1529,
    n934,
    n1426,
    n1439,
    n933
  );


  or
  g1499
  (
    n1519,
    n910,
    n930,
    n1444,
    n918
  );


  xnor
  g1500
  (
    n1532,
    n1432,
    n1441,
    n914,
    n1425
  );


  nand
  g1501
  (
    n1530,
    n929,
    n1433,
    n1425,
    n1429
  );


  nand
  g1502
  (
    n1549,
    n972,
    n965,
    n959,
    n1523
  );


  nor
  g1503
  (
    n1547,
    n961,
    n950,
    n1534,
    n968
  );


  nand
  g1504
  (
    n1552,
    n1517,
    n1522,
    n980,
    n968
  );


  xnor
  g1505
  (
    n1536,
    n1532,
    n963,
    n967,
    n949
  );


  and
  g1506
  (
    n1542,
    n975,
    n1521,
    n943,
    n941
  );


  nor
  g1507
  (
    n1548,
    n1520,
    n971,
    n964,
    n979
  );


  nand
  g1508
  (
    n1545,
    n969,
    n955,
    n1525,
    n945
  );


  nor
  g1509
  (
    n1540,
    n948,
    n956,
    n962,
    n1529
  );


  xnor
  g1510
  (
    n1553,
    n944,
    n958,
    n1533,
    n1527
  );


  xnor
  g1511
  (
    n1539,
    n1526,
    n969,
    n1524,
    n967
  );


  nand
  g1512
  (
    n1535,
    n966,
    n978,
    n972,
    n975
  );


  and
  g1513
  (
    n1544,
    n946,
    n938,
    n942,
    n976
  );


  xnor
  g1514
  (
    n1537,
    n1530,
    n977,
    n954,
    n1518
  );


  xor
  g1515
  (
    n1554,
    n966,
    n952,
    n939,
    n937
  );


  nand
  g1516
  (
    n1551,
    n940,
    n957,
    n976,
    n1531
  );


  xnor
  g1517
  (
    n1538,
    n947,
    n974,
    n978,
    n960
  );


  nand
  g1518
  (
    n1550,
    n977,
    n953,
    n970,
    n1515
  );


  xor
  g1519
  (
    n1546,
    n979,
    n1528,
    n973,
    n1516
  );


  nand
  g1520
  (
    n1543,
    n971,
    n965,
    n936,
    n973
  );


  or
  g1521
  (
    n1541,
    n1519,
    n974,
    n970,
    n951
  );


  xnor
  g1522
  (
    n1583,
    n1488,
    n1504,
    n1535,
    n1546
  );


  nor
  g1523
  (
    n1602,
    n1458,
    n1238,
    n1490,
    n1497
  );


  nand
  g1524
  (
    n1564,
    n1493,
    n1464,
    n1219,
    n1536
  );


  or
  g1525
  (
    n1556,
    n1280,
    n1220,
    n1552,
    n1239
  );


  xor
  g1526
  (
    n1629,
    n1237,
    n1231,
    n1451,
    n1537
  );


  and
  g1527
  (
    n1620,
    n1470,
    n1230,
    n1550,
    n1448
  );


  or
  g1528
  (
    n1569,
    n1228,
    n1541,
    n1238,
    n981
  );


  or
  g1529
  (
    n1597,
    n1242,
    n1491,
    n1234,
    n1504
  );


  or
  g1530
  (
    n1580,
    n1225,
    n1465,
    n1461,
    n1227
  );


  xor
  g1531
  (
    n1560,
    n1473,
    n1501,
    n1228,
    n1225
  );


  nand
  g1532
  (
    n1598,
    n1455,
    n1243,
    n1454,
    n1551
  );


  nand
  g1533
  (
    n1603,
    n1487,
    n1550,
    n1229,
    n1462
  );


  or
  g1534
  (
    n1558,
    n1237,
    n1486,
    n1541,
    n1496
  );


  xnor
  g1535
  (
    n1586,
    n1552,
    n980,
    n1449,
    n1497
  );


  xnor
  g1536
  (
    n1605,
    n1236,
    n1551,
    n1550,
    n1337
  );


  or
  g1537
  (
    n1613,
    n1453,
    n1341,
    n1222,
    n1485
  );


  xnor
  g1538
  (
    n1610,
    n1234,
    n1474,
    n1336,
    n1468
  );


  xnor
  g1539
  (
    n1594,
    n1553,
    n1463,
    n1465,
    n1538
  );


  xnor
  g1540
  (
    n1608,
    n1220,
    n1547,
    n1242,
    n1552
  );


  and
  g1541
  (
    n1557,
    n1539,
    n1241,
    n1552,
    n1225
  );


  or
  g1542
  (
    n1596,
    n1503,
    n1229,
    n1494,
    n1538
  );


  xnor
  g1543
  (
    n1599,
    n1478,
    n1222,
    n1230,
    n1542
  );


  and
  g1544
  (
    n1614,
    n1535,
    n1478,
    n1543,
    n1233
  );


  or
  g1545
  (
    n1606,
    n1501,
    n1486,
    n1549,
    n1230
  );


  nor
  g1546
  (
    n1567,
    n1479,
    n1457,
    n1240,
    n1336
  );


  xor
  g1547
  (
    n1615,
    n1241,
    n1545,
    n1455,
    n1338
  );


  nor
  g1548
  (
    n1621,
    n1548,
    n1544,
    n1240
  );


  and
  g1549
  (
    n1625,
    n1541,
    n1448,
    n1227,
    n1468
  );


  and
  g1550
  (
    n1585,
    n1343,
    n1237,
    n1540,
    n1227
  );


  xnor
  g1551
  (
    n1633,
    n1224,
    n1461,
    n1537,
    n1547
  );


  and
  g1552
  (
    n1588,
    n1537,
    n1231,
    n1500,
    n1471
  );


  nand
  g1553
  (
    n1563,
    n1545,
    n1467,
    n1498,
    n1243
  );


  and
  g1554
  (
    n1581,
    n1543,
    n1475,
    n1459,
    n1240
  );


  nand
  g1555
  (
    n1611,
    n1484,
    n1229,
    n1554,
    n1502
  );


  nor
  g1556
  (
    KeyWire_0_5,
    n1449,
    n1537,
    n1238,
    n1477
  );


  nor
  g1557
  (
    n1573,
    n1499,
    n1340,
    n1226,
    n1221
  );


  nor
  g1558
  (
    n1570,
    n1502,
    n1219,
    n1551,
    n1340
  );


  xnor
  g1559
  (
    n1582,
    n1543,
    n1554,
    n1244,
    n1553
  );


  xor
  g1560
  (
    n1619,
    n1343,
    n1554,
    n1234,
    n1452
  );


  nand
  g1561
  (
    n1562,
    n1472,
    n1540,
    n1232,
    n1490
  );


  and
  g1562
  (
    n1577,
    n1550,
    n1223,
    n1231
  );


  xnor
  g1563
  (
    n1624,
    n1495,
    n1541,
    n1244,
    n1496
  );


  nor
  g1564
  (
    n1631,
    n1542,
    n1228,
    n1222,
    n1500
  );


  or
  g1565
  (
    n1604,
    n1548,
    n1482,
    n1227,
    n1236
  );


  xor
  g1566
  (
    n1571,
    n1339,
    n1456,
    n1481,
    n1548
  );


  nand
  g1567
  (
    n1575,
    n1458,
    n1553,
    n1491,
    n1239
  );


  or
  g1568
  (
    n1616,
    n1456,
    n1547,
    n1224,
    n1538
  );


  xnor
  g1569
  (
    n1600,
    n1549,
    n1228,
    n1476,
    n1232
  );


  xor
  g1570
  (
    n1630,
    n1244,
    n1553,
    n1235,
    n1453
  );


  xor
  g1571
  (
    n1555,
    n1536,
    n1235,
    n1244,
    n1494
  );


  or
  g1572
  (
    n1618,
    n1538,
    n1452,
    n1549,
    n1220
  );


  and
  g1573
  (
    n1609,
    n1482,
    n1457,
    n1239,
    n1226
  );


  and
  g1574
  (
    n1634,
    n1226,
    n1466,
    n1549,
    n1475
  );


  nand
  g1575
  (
    n1559,
    n1454,
    n1471,
    n1542
  );


  nand
  g1576
  (
    n1632,
    n1466,
    n1544,
    n1480,
    n1505
  );


  nand
  g1577
  (
    n1576,
    n1242,
    n1451,
    n1503,
    n1243
  );


  nor
  g1578
  (
    n1593,
    n1235,
    n1460,
    n1243,
    n1484
  );


  xor
  g1579
  (
    n1574,
    n1545,
    n1535,
    n1342,
    n1474
  );


  xnor
  g1580
  (
    n1622,
    n1221,
    n1477,
    n1223,
    n1495
  );


  nor
  g1581
  (
    n1565,
    n1535,
    n1498,
    n1479,
    n1222
  );


  nor
  g1582
  (
    n1578,
    n1470,
    n1551,
    n1480,
    n1539
  );


  and
  g1583
  (
    n1579,
    n1499,
    n1229,
    n672,
    n1337
  );


  nand
  g1584
  (
    n1584,
    n1536,
    n1242,
    n1492,
    n1221
  );


  xor
  g1585
  (
    n1572,
    n1493,
    n1546,
    n1232,
    n1224
  );


  nand
  g1586
  (
    n1623,
    n1489,
    n1241,
    n1481,
    n1544
  );


  and
  g1587
  (
    n1607,
    n1540,
    n1240,
    n1543,
    n1230
  );


  or
  g1588
  (
    n1591,
    n1232,
    n1459,
    n1338,
    n1223
  );


  or
  g1589
  (
    n1601,
    n1467,
    n1241,
    n1539,
    n1341
  );


  and
  g1590
  (
    n1592,
    n1473,
    n1239,
    n1476,
    n1463
  );


  or
  g1591
  (
    n1589,
    n1236,
    n1548,
    n1342,
    n1546
  );


  xnor
  g1592
  (
    n1568,
    n1536,
    n1483,
    n1238,
    n1450
  );


  and
  g1593
  (
    n1627,
    n1450,
    n1233,
    n1539,
    n1483
  );


  and
  g1594
  (
    n1628,
    n1487,
    n1488,
    n1221,
    n1231
  );


  and
  g1595
  (
    n1595,
    n1472,
    n1545,
    n1464,
    n1460
  );


  and
  g1596
  (
    n1590,
    n1219,
    n1492,
    n1462,
    n1220
  );


  and
  g1597
  (
    n1561,
    n1469,
    n1234,
    n1489,
    n1485
  );


  nand
  g1598
  (
    n1587,
    n1469,
    n1225,
    n1219,
    n1233
  );


  and
  g1599
  (
    n1612,
    n1546,
    n672,
    n1554,
    n1233
  );


  and
  g1600
  (
    n1566,
    n1224,
    n1236,
    n1540,
    n1226
  );


  nand
  g1601
  (
    n1617,
    n1547,
    n1339,
    n1235,
    n1237
  );


  not
  g1602
  (
    n1656,
    n1569
  );


  not
  g1603
  (
    n1660,
    n986
  );


  not
  g1604
  (
    n1671,
    n981
  );


  buf
  g1605
  (
    n1648,
    n1557
  );


  not
  g1606
  (
    n1642,
    n1562
  );


  not
  g1607
  (
    n1658,
    n1556
  );


  buf
  g1608
  (
    n1677,
    n1572
  );


  not
  g1609
  (
    n1649,
    n1570
  );


  buf
  g1610
  (
    n1657,
    n1555
  );


  not
  g1611
  (
    n1667,
    n1559
  );


  not
  g1612
  (
    n1652,
    n1573
  );


  buf
  g1613
  (
    n1636,
    n988
  );


  buf
  g1614
  (
    n1666,
    n1561
  );


  buf
  g1615
  (
    n1672,
    n1564
  );


  not
  g1616
  (
    n1640,
    n1571
  );


  not
  g1617
  (
    n1646,
    n989
  );


  not
  g1618
  (
    n1674,
    n1566
  );


  buf
  g1619
  (
    n1668,
    n1565
  );


  not
  g1620
  (
    n1654,
    n1558
  );


  buf
  g1621
  (
    n1673,
    n984
  );


  not
  g1622
  (
    n1639,
    n990
  );


  buf
  g1623
  (
    n1661,
    n987
  );


  not
  g1624
  (
    n1635,
    n986
  );


  not
  g1625
  (
    n1675,
    n1555
  );


  not
  g1626
  (
    n1647,
    n988
  );


  buf
  g1627
  (
    n1664,
    n1569
  );


  not
  g1628
  (
    n1645,
    n1558
  );


  not
  g1629
  (
    n1651,
    n1562
  );


  not
  g1630
  (
    n1659,
    n982
  );


  not
  g1631
  (
    n1637,
    n1574
  );


  buf
  g1632
  (
    n1663,
    n989
  );


  buf
  g1633
  (
    n1655,
    n983
  );


  buf
  g1634
  (
    n1641,
    n987
  );


  not
  g1635
  (
    n1669,
    n1576
  );


  not
  g1636
  (
    n1665,
    n1568
  );


  nand
  g1637
  (
    n1670,
    n1575,
    n1574,
    n1567
  );


  and
  g1638
  (
    n1676,
    n1567,
    n1572,
    n1571
  );


  xor
  g1639
  (
    n1650,
    n1573,
    n985,
    n1557
  );


  xor
  g1640
  (
    n1678,
    n984,
    n1575,
    n1576
  );


  nor
  g1641
  (
    n1638,
    n1563,
    n1565,
    n1564
  );


  nor
  g1642
  (
    n1644,
    n1568,
    n1570,
    n983
  );


  nand
  g1643
  (
    n1643,
    n982,
    n1563,
    n1560
  );


  nor
  g1644
  (
    n1653,
    n1556,
    n985,
    n1566
  );


  xor
  g1645
  (
    n1662,
    n1560,
    n1559,
    n1561
  );


  nand
  g1646
  (
    n1692,
    n1644,
    n1026,
    n1009,
    n993
  );


  nor
  g1647
  (
    n1694,
    n1036,
    n992,
    n1649,
    n994
  );


  and
  g1648
  (
    n1691,
    n1040,
    n1648,
    n994,
    n1022
  );


  xnor
  g1649
  (
    n1690,
    n1013,
    n1038,
    n1650,
    n1002
  );


  nor
  g1650
  (
    n1704,
    n1017,
    n1020,
    n1015,
    n1016
  );


  xnor
  g1651
  (
    n1703,
    n1639,
    n999,
    n1039,
    n997
  );


  xor
  g1652
  (
    n1710,
    n1003,
    n1642,
    n1008,
    n1640
  );


  xnor
  g1653
  (
    n1687,
    n1640,
    n1642,
    n1008,
    n1003
  );


  nand
  g1654
  (
    n1701,
    n1024,
    n1649,
    n1036,
    n1646
  );


  xor
  g1655
  (
    n1712,
    n993,
    n1002,
    n1010,
    n1037
  );


  xnor
  g1656
  (
    n1683,
    n1031,
    n999,
    n1636,
    n1011
  );


  nand
  g1657
  (
    n1679,
    n1012,
    n1647,
    n1022,
    n1637
  );


  xor
  g1658
  (
    n1707,
    n1035,
    n1032,
    n998
  );


  nand
  g1659
  (
    n1711,
    n1024,
    n1007,
    n1019,
    n1006
  );


  nand
  g1660
  (
    n1695,
    n1027,
    n990,
    n1011,
    n1641
  );


  nor
  g1661
  (
    n1686,
    n1001,
    n1643,
    n1021,
    n1030
  );


  nor
  g1662
  (
    n1682,
    n1016,
    n996,
    n1649,
    n1033
  );


  or
  g1663
  (
    n1684,
    n1031,
    n1018,
    n1004,
    n1015
  );


  xor
  g1664
  (
    n1689,
    n1006,
    n1635,
    n1010,
    n1644
  );


  nand
  g1665
  (
    n1681,
    n1638,
    n1001,
    n997,
    n1000
  );


  xnor
  g1666
  (
    n1702,
    n991,
    n1005,
    n1034,
    n1028
  );


  xnor
  g1667
  (
    n1700,
    n1636,
    n1637,
    n991,
    n1012
  );


  nand
  g1668
  (
    n1709,
    n1035,
    n1014,
    n1643,
    n995
  );


  nand
  g1669
  (
    n1708,
    n1041,
    n992,
    n1019,
    n1039
  );


  xnor
  g1670
  (
    n1685,
    n1026,
    n1000,
    n1025
  );


  and
  g1671
  (
    n1693,
    n1645,
    n1649,
    n1639,
    n1032
  );


  or
  g1672
  (
    n1688,
    n1021,
    n1638,
    n1005,
    n1028
  );


  xor
  g1673
  (
    n1680,
    n1650,
    n1017,
    n1029,
    n1645
  );


  or
  g1674
  (
    n1698,
    n1648,
    n1029,
    n1641,
    n995
  );


  xor
  g1675
  (
    n1706,
    n1004,
    n1635,
    n1009,
    n1646
  );


  xor
  g1676
  (
    n1705,
    n1027,
    n1007,
    n1023,
    n1034
  );


  nand
  g1677
  (
    n1699,
    n1038,
    n1023,
    n1040,
    n1033
  );


  nand
  g1678
  (
    n1696,
    n996,
    n1037,
    n1647,
    n1020
  );


  xor
  g1679
  (
    n1697,
    n1030,
    n1018,
    n1013,
    n1014
  );


  and
  g1680
  (
    n1719,
    n1685,
    n1358,
    n1290,
    n1712
  );


  and
  g1681
  (
    n1730,
    n1683,
    n1691,
    n1706,
    n1353
  );


  and
  g1682
  (
    n1723,
    n1352,
    n1298,
    n1346,
    n1702
  );


  nor
  g1683
  (
    n1714,
    n1297,
    n1303,
    n1357,
    n1286
  );


  xor
  g1684
  (
    n1721,
    n1682,
    n1346,
    n1301,
    n1306
  );


  xor
  g1685
  (
    n1727,
    n1351,
    n1284,
    n1359,
    n1293
  );


  or
  g1686
  (
    n1732,
    n1292,
    n1681,
    n1290,
    n1709
  );


  nand
  g1687
  (
    n1725,
    n1304,
    n1288,
    n1306,
    n1308
  );


  nor
  g1688
  (
    n1720,
    n1361,
    n1299,
    n1689,
    n1697
  );


  or
  g1689
  (
    n1737,
    n1042,
    n1345,
    n1308,
    n1693
  );


  nand
  g1690
  (
    n1746,
    n1304,
    n1284,
    n1291,
    n1345
  );


  xnor
  g1691
  (
    n1716,
    n1679,
    n1347,
    n1043,
    n1344
  );


  nand
  g1692
  (
    n1736,
    n1360,
    n1298,
    n1359,
    n1355
  );


  or
  g1693
  (
    n1739,
    n1291,
    n1686,
    n1353,
    n1280
  );


  xor
  g1694
  (
    n1741,
    n1043,
    n1283,
    n1699,
    n1297
  );


  nor
  g1695
  (
    n1743,
    n1688,
    n1700,
    n1349,
    n1306
  );


  nand
  g1696
  (
    n1731,
    n1687,
    n1293,
    n1710,
    n1360
  );


  xnor
  g1697
  (
    n1728,
    n1287,
    n1354,
    n1307
  );


  xor
  g1698
  (
    n1729,
    n1283,
    n1684,
    n1305,
    n1348
  );


  nor
  g1699
  (
    n1718,
    n1707,
    n1692,
    n1344,
    n1350
  );


  xor
  g1700
  (
    n1742,
    n1303,
    n1300,
    n1296,
    n1695
  );


  xnor
  g1701
  (
    n1747,
    n1705,
    n1650,
    n1711,
    n1042
  );


  nor
  g1702
  (
    n1745,
    n1351,
    n1289,
    n1282,
    n1307
  );


  nand
  g1703
  (
    n1744,
    n1281,
    n1302,
    n1294,
    n1295
  );


  nand
  g1704
  (
    n1740,
    n1289,
    n1305,
    n1698,
    n1299
  );


  or
  g1705
  (
    n1738,
    n1708,
    n1690,
    n1307,
    n1308
  );


  nand
  g1706
  (
    n1726,
    n1350,
    n1357,
    n1358,
    n1282
  );


  and
  g1707
  (
    n1713,
    n1712,
    n1704,
    n1696,
    n1286
  );


  nand
  g1708
  (
    n1715,
    n1292,
    n1356,
    n1285,
    n1348
  );


  xor
  g1709
  (
    n1717,
    n1349,
    n1044,
    n1356,
    n1703
  );


  and
  g1710
  (
    n1724,
    n1307,
    n1694,
    n1288,
    n1302
  );


  xor
  g1711
  (
    n1722,
    n1295,
    n1300,
    n1355,
    n1308
  );


  xnor
  g1712
  (
    n1734,
    n1352,
    n1281,
    n1294,
    n1347
  );


  nand
  g1713
  (
    n1733,
    n1287,
    n1701,
    n1044,
    n1285
  );


  and
  g1714
  (
    n1735,
    n1301,
    n1041,
    n1680,
    n1296
  );


  not
  g1715
  (
    n1872,
    n1659
  );


  buf
  g1716
  (
    n1815,
    n1731
  );


  buf
  g1717
  (
    n1881,
    n1672
  );


  buf
  g1718
  (
    n1852,
    n1621
  );


  buf
  g1719
  (
    n1846,
    n1584
  );


  not
  g1720
  (
    n1874,
    n1599
  );


  not
  g1721
  (
    n1779,
    n1725
  );


  not
  g1722
  (
    n1788,
    n1585
  );


  not
  g1723
  (
    n1842,
    n1362
  );


  not
  g1724
  (
    n1825,
    n1596
  );


  buf
  g1725
  (
    n1835,
    n1740
  );


  not
  g1726
  (
    n1878,
    n1737
  );


  not
  g1727
  (
    n1887,
    n1677
  );


  not
  g1728
  (
    n1804,
    n1660
  );


  buf
  g1729
  (
    n1829,
    n1594
  );


  not
  g1730
  (
    n1850,
    n1746
  );


  buf
  g1731
  (
    n1860,
    n1734
  );


  buf
  g1732
  (
    KeyWire_0_4,
    n1724
  );


  not
  g1733
  (
    n1751,
    n1593
  );


  buf
  g1734
  (
    n1856,
    n1579
  );


  buf
  g1735
  (
    n1799,
    n1580
  );


  not
  g1736
  (
    n1843,
    n1665
  );


  buf
  g1737
  (
    n1752,
    n1737
  );


  buf
  g1738
  (
    n1851,
    n1598
  );


  buf
  g1739
  (
    n1783,
    n1677
  );


  buf
  g1740
  (
    n1778,
    n1731
  );


  not
  g1741
  (
    n1816,
    n1659
  );


  not
  g1742
  (
    n1823,
    n1583
  );


  not
  g1743
  (
    n1848,
    n1667
  );


  buf
  g1744
  (
    n1865,
    n1590
  );


  and
  g1745
  (
    n1784,
    n1747,
    n1722,
    n1728,
    n1614
  );


  nand
  g1746
  (
    n1828,
    n1670,
    n1656,
    n1621,
    n1619
  );


  or
  g1747
  (
    n1885,
    n1598,
    n1585,
    n1673,
    n1593
  );


  nand
  g1748
  (
    n1786,
    n1584,
    n1651,
    n1599,
    n1594
  );


  or
  g1749
  (
    n1834,
    n1726,
    n1599,
    n1678,
    n1658
  );


  nand
  g1750
  (
    n1847,
    n1617,
    n1579,
    n1656,
    n1253
  );


  nand
  g1751
  (
    n1830,
    n1722,
    n1746,
    n1591,
    n1656
  );


  and
  g1752
  (
    n1812,
    n1622,
    n1612,
    n1587,
    n1590
  );


  xor
  g1753
  (
    n1871,
    n1740,
    n1673,
    n1666,
    n1587
  );


  xor
  g1754
  (
    n1781,
    n1723,
    n1605,
    n1604,
    n1603
  );


  xnor
  g1755
  (
    n1798,
    n1715,
    n1602,
    n1723,
    n1719
  );


  and
  g1756
  (
    n1800,
    n1739,
    n1601,
    n1604,
    n1738
  );


  nor
  g1757
  (
    n1775,
    n1595,
    n1652,
    n1593,
    n1713
  );


  xnor
  g1758
  (
    n1782,
    n1511,
    n1651,
    n1668,
    n1587
  );


  nor
  g1759
  (
    n1749,
    n1659,
    n1595,
    n1657,
    n1728
  );


  nor
  g1760
  (
    n1765,
    n1611,
    n1669,
    n1605,
    n1725
  );


  xnor
  g1761
  (
    n1794,
    n1653,
    n1615,
    n1743,
    n1597
  );


  or
  g1762
  (
    n1755,
    n1661,
    n1738,
    n1510,
    n1735
  );


  xor
  g1763
  (
    n1787,
    n1661,
    n1670,
    n1595,
    n1591
  );


  or
  g1764
  (
    n1813,
    n1721,
    n1651,
    n1731,
    n1677
  );


  and
  g1765
  (
    n1753,
    n1587,
    n1678,
    n1722,
    n1578
  );


  or
  g1766
  (
    n1831,
    n1719,
    n1589,
    n1361,
    n1577
  );


  and
  g1767
  (
    n1771,
    n1729,
    n1721,
    n1741,
    n1601
  );


  nor
  g1768
  (
    n1760,
    n1717,
    n1730,
    n1665,
    n1668
  );


  nand
  g1769
  (
    n1803,
    n1662,
    n1720,
    n1617,
    n1603
  );


  xnor
  g1770
  (
    n1886,
    n1579,
    n1667,
    n1670,
    n1606
  );


  xor
  g1771
  (
    n1821,
    n1592,
    n1658,
    n1650,
    n1713
  );


  xnor
  g1772
  (
    n1818,
    n1618,
    n1662,
    n1596,
    n1742
  );


  xor
  g1773
  (
    n1868,
    n1254,
    n1506,
    n1593,
    n1608
  );


  and
  g1774
  (
    n1777,
    n1724,
    n1677,
    n1582,
    n1590
  );


  xor
  g1775
  (
    n1884,
    n1715,
    n1599,
    n1655,
    n1718
  );


  xor
  g1776
  (
    n1845,
    n1617,
    n1747,
    n1676,
    n1507
  );


  nand
  g1777
  (
    n1750,
    n1662,
    n1715,
    n1586,
    n1727
  );


  xor
  g1778
  (
    n1841,
    n1747,
    n1601,
    n1734,
    n1727
  );


  xor
  g1779
  (
    n1795,
    n1616,
    n1663,
    n1747,
    n1364
  );


  and
  g1780
  (
    n1807,
    n1368,
    n1730,
    n1576,
    n1745
  );


  nand
  g1781
  (
    n1748,
    n1675,
    n1620,
    n1612,
    n1591
  );


  and
  g1782
  (
    n1801,
    n1718,
    n1743,
    n1717,
    n1746
  );


  xor
  g1783
  (
    n1849,
    n1676,
    n1611,
    n1608,
    n1509
  );


  or
  g1784
  (
    n1822,
    n1669,
    n1673,
    n1652,
    n1720
  );


  or
  g1785
  (
    n1776,
    n1713,
    n1744,
    n1607,
    n1254
  );


  and
  g1786
  (
    n1767,
    n1675,
    n1620,
    n1728,
    n1589
  );


  or
  g1787
  (
    n1817,
    n1614,
    n1589,
    n1676,
    n1714
  );


  xor
  g1788
  (
    n1757,
    n1672,
    n1727,
    n1740,
    n1678
  );


  xnor
  g1789
  (
    n1802,
    n1675,
    n1724,
    n1585,
    n1657
  );


  nor
  g1790
  (
    n1855,
    n1674,
    n1595,
    n1733,
    n1613
  );


  xnor
  g1791
  (
    n1797,
    n1662,
    n1658,
    n1580,
    n1741
  );


  and
  g1792
  (
    n1863,
    n1672,
    n1735,
    n1665,
    n1600
  );


  xor
  g1793
  (
    n1873,
    n1612,
    n1654,
    n1576,
    n1603
  );


  xor
  g1794
  (
    n1811,
    n1605,
    n1718,
    n1732,
    n1582
  );


  xor
  g1795
  (
    n1769,
    n1732,
    n1602,
    n1586,
    n1610
  );


  xor
  g1796
  (
    n1870,
    n1742,
    n1584,
    n1716,
    n1664
  );


  nor
  g1797
  (
    n1770,
    n1606,
    n1583,
    n1659
  );


  nor
  g1798
  (
    n1754,
    n1509,
    n1734,
    n1668,
    n1735
  );


  and
  g1799
  (
    n1790,
    n1602,
    n1658,
    n1678,
    n1508
  );


  xor
  g1800
  (
    n1862,
    n1724,
    n1614,
    n1620,
    n1507
  );


  or
  g1801
  (
    n1761,
    n1582,
    n1738,
    n1667,
    n1741
  );


  xor
  g1802
  (
    n1858,
    n1739,
    n1668,
    n1725,
    n1652
  );


  and
  g1803
  (
    n1806,
    n1588,
    n1745,
    n1616,
    n1729
  );


  nor
  g1804
  (
    n1796,
    n1666,
    n1592,
    n1598,
    n1743
  );


  or
  g1805
  (
    n1789,
    n1620,
    n1714,
    n1590,
    n1676
  );


  xor
  g1806
  (
    n1772,
    n1666,
    n1674,
    n1723,
    n1510
  );


  nor
  g1807
  (
    n1762,
    n1739,
    n1610,
    n1716
  );


  nor
  g1808
  (
    n1808,
    n1600,
    n1669,
    n1609,
    n1592
  );


  or
  g1809
  (
    n1832,
    n1664,
    n1743,
    n1615,
    n1657
  );


  and
  g1810
  (
    n1759,
    n1365,
    n1718,
    n1651,
    n1655
  );


  and
  g1811
  (
    n1861,
    n1733,
    n1732,
    n1614,
    n1586
  );


  nand
  g1812
  (
    n1864,
    n1671,
    n1654,
    n1665,
    n1669
  );


  xnor
  g1813
  (
    n1866,
    n1720,
    n1744,
    n1730,
    n1663
  );


  xor
  g1814
  (
    n1814,
    n1254,
    n1580,
    n1654,
    n1602
  );


  nand
  g1815
  (
    n1844,
    n1588,
    n1729,
    n1578,
    n1736
  );


  xnor
  g1816
  (
    n1826,
    n1745,
    n1615,
    n1732
  );


  xnor
  g1817
  (
    n1791,
    n1608,
    n1616,
    n1715,
    n1594
  );


  or
  g1818
  (
    n1840,
    n1672,
    n1613,
    n1674,
    n1621
  );


  and
  g1819
  (
    n1877,
    n1742,
    n1663,
    n1577,
    n1604
  );


  nand
  g1820
  (
    n1879,
    n1363,
    n1365,
    n1596,
    n1674
  );


  and
  g1821
  (
    n1763,
    n1607,
    n1612,
    n1606,
    n1740
  );


  nor
  g1822
  (
    n1827,
    n1581,
    n1607,
    n1654,
    n1652
  );


  nand
  g1823
  (
    n1854,
    n1733,
    n1661,
    n1577,
    n1585
  );


  nand
  g1824
  (
    n1766,
    n1577,
    n1367,
    n1363,
    n1741
  );


  and
  g1825
  (
    n1824,
    n1622,
    n1609,
    n1616,
    n1619
  );


  nor
  g1826
  (
    n1756,
    n1734,
    n1597,
    n1656,
    n1746
  );


  and
  g1827
  (
    n1838,
    n1738,
    n1719,
    n1739,
    n1609
  );


  and
  g1828
  (
    n1867,
    n1671,
    n1725,
    n1619,
    n1714
  );


  or
  g1829
  (
    n1792,
    n1506,
    n1610,
    n1663,
    n1660
  );


  nor
  g1830
  (
    n1880,
    n1596,
    n1254,
    n1736,
    n1597
  );


  xnor
  g1831
  (
    KeyWire_0_2,
    n1366,
    n1720,
    n1717,
    n1726
  );


  nor
  g1832
  (
    n1857,
    n1613,
    n1611,
    n1664,
    n1737
  );


  and
  g1833
  (
    n1819,
    n1600,
    n1723,
    n1735,
    n1714
  );


  xnor
  g1834
  (
    n1810,
    n1660,
    n1716,
    n1584,
    n1582
  );


  nand
  g1835
  (
    n1883,
    n1727,
    n1675,
    n1671,
    n1655
  );


  and
  g1836
  (
    n1809,
    n1673,
    n1578,
    n1744,
    n1742
  );


  xnor
  g1837
  (
    n1837,
    n1717,
    n1736,
    n1728,
    n1716
  );


  nor
  g1838
  (
    n1836,
    n1364,
    n1609,
    n1591,
    n1597
  );


  xnor
  g1839
  (
    n1820,
    n1580,
    n1617,
    n1729,
    n1598
  );


  xor
  g1840
  (
    n1882,
    n1594,
    n1621,
    n1653,
    n1613
  );


  or
  g1841
  (
    n1793,
    n1606,
    n1670,
    n1588,
    n1737
  );


  nand
  g1842
  (
    n1876,
    n1511,
    n1618,
    n1603,
    n1721
  );


  xor
  g1843
  (
    n1785,
    n1588,
    n1730,
    n1721,
    n1736
  );


  and
  g1844
  (
    n1869,
    n1666,
    n1618,
    n1719,
    n1722
  );


  xor
  g1845
  (
    n1780,
    n1367,
    n1592,
    n1726,
    n1366
  );


  nand
  g1846
  (
    n1853,
    n1661,
    n1508,
    n1586,
    n1505
  );


  or
  g1847
  (
    n1833,
    n1733,
    n1660,
    n1657,
    n1604
  );


  and
  g1848
  (
    n1764,
    n1745,
    n1671,
    n1619,
    n1368
  );


  and
  g1849
  (
    n1875,
    n1608,
    n1653,
    n1601,
    n1605
  );


  nor
  g1850
  (
    n1758,
    n1726,
    n1744,
    n1581,
    n1362
  );


  nor
  g1851
  (
    n1774,
    n1618,
    n1600,
    n1667,
    n1611
  );


  nor
  g1852
  (
    n1859,
    n1713,
    n1589,
    n1731,
    n1653
  );


  xor
  g1853
  (
    n1839,
    n1664,
    n1578,
    n1581
  );


  nor
  g1854
  (
    n1805,
    n1607,
    n1655,
    n1583,
    n1579
  );


  xor
  g1855
  (
    n1952,
    n1080,
    n1153,
    n1143,
    n1772
  );


  nand
  g1856
  (
    n1998,
    n1627,
    n1816,
    n1855,
    n1045
  );


  xor
  g1857
  (
    n1979,
    n1828,
    n1082,
    n1124,
    n1080
  );


  xor
  g1858
  (
    n1934,
    n1622,
    n1172,
    n1860,
    n1760
  );


  nand
  g1859
  (
    n1955,
    n1156,
    n1624,
    n1754,
    n1084
  );


  nor
  g1860
  (
    n1961,
    n1761,
    n1096,
    n1178,
    n1633
  );


  nand
  g1861
  (
    n1903,
    n1046,
    n1858,
    n1105,
    n1058
  );


  nand
  g1862
  (
    n1974,
    n1112,
    n1623,
    n1804,
    n1628
  );


  and
  g1863
  (
    n1990,
    n1166,
    n1775,
    n1631,
    n1849
  );


  or
  g1864
  (
    n1969,
    n1148,
    n1123,
    n1070,
    n1054
  );


  nand
  g1865
  (
    n1892,
    n1848,
    n1865,
    n1845,
    n1843
  );


  and
  g1866
  (
    n2001,
    n1134,
    n1164,
    n1630,
    n1048
  );


  and
  g1867
  (
    n1931,
    n1078,
    n1148,
    n1140,
    n1066
  );


  or
  g1868
  (
    n1929,
    n1814,
    n1624,
    n1864,
    n1626
  );


  and
  g1869
  (
    n2002,
    n1752,
    n1048,
    n1130,
    n1116
  );


  and
  g1870
  (
    n1935,
    n1085,
    n1881,
    n1629,
    n1105
  );


  or
  g1871
  (
    n1973,
    n1057,
    n1052,
    n1759,
    n1132
  );


  nor
  g1872
  (
    n1893,
    n1630,
    n1162,
    n1099,
    n1807
  );


  xnor
  g1873
  (
    n1991,
    n1825,
    n1079,
    n1126,
    n1869
  );


  xor
  g1874
  (
    n1959,
    n1076,
    n1175,
    n1832,
    n1120
  );


  nor
  g1875
  (
    n1986,
    n1853,
    n1096,
    n1846,
    n1109
  );


  or
  g1876
  (
    n1971,
    n1111,
    n1115,
    n1072,
    n1103
  );


  xor
  g1877
  (
    n1904,
    n1632,
    n1753,
    n1107,
    n1145
  );


  xnor
  g1878
  (
    n1932,
    n1762,
    n1049,
    n1167,
    n1854
  );


  xor
  g1879
  (
    n1949,
    n1113,
    n1622,
    n1070,
    n1075
  );


  nor
  g1880
  (
    n1890,
    n1887,
    n1780,
    n1133,
    n1122
  );


  xnor
  g1881
  (
    n1977,
    n1632,
    n1836,
    n1179,
    n1131
  );


  and
  g1882
  (
    n1916,
    n1063,
    n1093,
    n1626,
    n1176
  );


  or
  g1883
  (
    n1924,
    n1794,
    n1824,
    n1068,
    n1155
  );


  and
  g1884
  (
    n1936,
    n1058,
    n1169,
    n1086,
    n1758
  );


  xor
  g1885
  (
    n1976,
    n1790,
    n1177,
    n1136,
    n1059
  );


  nor
  g1886
  (
    n1941,
    n1776,
    n1162,
    n1090,
    n1151
  );


  xor
  g1887
  (
    n1913,
    n1088,
    n1050,
    n1630,
    n1808
  );


  xnor
  g1888
  (
    KeyWire_0_0,
    n1119,
    n1629,
    n1118,
    n1114
  );


  xor
  g1889
  (
    n1888,
    n1095,
    n1047,
    n1128,
    n1066
  );


  and
  g1890
  (
    n1915,
    n1628,
    n1781,
    n1081,
    n1885
  );


  nand
  g1891
  (
    n1899,
    n1166,
    n1108,
    n1065,
    n1149
  );


  nand
  g1892
  (
    n1950,
    n1053,
    n1139,
    n1101,
    n1176
  );


  nor
  g1893
  (
    n1997,
    n1763,
    n1160,
    n1073,
    n1154
  );


  and
  g1894
  (
    n1953,
    n1822,
    n1144,
    n1173,
    n1632
  );


  xnor
  g1895
  (
    n1962,
    n1631,
    n1099,
    n1883,
    n1076
  );


  nand
  g1896
  (
    n1920,
    n1631,
    n1150,
    n1815,
    n1056
  );


  nand
  g1897
  (
    n1907,
    n1121,
    n1056,
    n1112,
    n1633
  );


  and
  g1898
  (
    n1943,
    n1051,
    n1094,
    n1135,
    n1626
  );


  xnor
  g1899
  (
    n1895,
    n1168,
    n1059,
    n1634,
    n1764
  );


  or
  g1900
  (
    n1933,
    n1625,
    n1805,
    n1046,
    n1870
  );


  and
  g1901
  (
    n1967,
    n1767,
    n1175,
    n1130,
    n1095
  );


  or
  g1902
  (
    n1926,
    n1097,
    n1793,
    n1084,
    n1788
  );


  nand
  g1903
  (
    n1984,
    n1092,
    n1068,
    n1127,
    n1077
  );


  and
  g1904
  (
    n1921,
    n1871,
    n1147,
    n1629,
    n1069
  );


  xor
  g1905
  (
    n1958,
    n1072,
    n1167,
    n1135,
    n1139
  );


  nand
  g1906
  (
    n1889,
    n1839,
    n1784,
    n1811,
    n1057
  );


  xnor
  g1907
  (
    n1891,
    n1078,
    n1168,
    n1796,
    n1134
  );


  xor
  g1908
  (
    n1988,
    n1124,
    n1777,
    n1109,
    n1180
  );


  xor
  g1909
  (
    n1945,
    n1089,
    n1623,
    n1110,
    n1091
  );


  xnor
  g1910
  (
    n1951,
    n1097,
    n1876,
    n1129,
    n1170
  );


  xor
  g1911
  (
    n1939,
    n1165,
    n1868,
    n1633,
    n1768
  );


  nand
  g1912
  (
    n1938,
    n1053,
    n1098,
    n1144,
    n1074
  );


  xor
  g1913
  (
    n1906,
    n1634,
    n1071,
    n1102,
    n1833
  );


  nor
  g1914
  (
    n1937,
    n1067,
    n1156,
    n1789,
    n1061
  );


  and
  g1915
  (
    n1994,
    n1077,
    n1857,
    n1838,
    n1089
  );


  nor
  g1916
  (
    n2000,
    n1114,
    n1091,
    n1157,
    n1104
  );


  xnor
  g1917
  (
    n1970,
    n1803,
    n1823,
    n1634,
    n1103
  );


  or
  g1918
  (
    n2003,
    n1136,
    n1062,
    n1785,
    n1120
  );


  or
  g1919
  (
    n1894,
    n1625,
    n1161,
    n1791,
    n1840
  );


  nor
  g1920
  (
    KeyWire_0_9,
    n1797,
    n1131,
    n1141,
    n1847
  );


  or
  g1921
  (
    n1930,
    n1631,
    n1145,
    n1875,
    n1111
  );


  and
  g1922
  (
    n1978,
    n1169,
    n1122,
    n1164,
    n1809
  );


  or
  g1923
  (
    n1897,
    n1094,
    n1118,
    n1163,
    n1137
  );


  xor
  g1924
  (
    n1987,
    n1799,
    n1877,
    n1143,
    n1866
  );


  and
  g1925
  (
    n1908,
    n1829,
    n1123,
    n1770,
    n1159
  );


  and
  g1926
  (
    n1964,
    n1060,
    n1101,
    n1882,
    n1831
  );


  xnor
  g1927
  (
    n1914,
    n1082,
    n1125,
    n1117,
    n1088
  );


  xor
  g1928
  (
    n1972,
    n1750,
    n1792,
    n1063,
    n1627
  );


  and
  g1929
  (
    n1923,
    n1756,
    n1093,
    n1632,
    n1774
  );


  and
  g1930
  (
    n1960,
    n1142,
    n1087,
    n1100,
    n1121
  );


  and
  g1931
  (
    n1965,
    n1065,
    n1817,
    n1126,
    n1782
  );


  xnor
  g1932
  (
    n1925,
    n1152,
    n1067,
    n1051,
    n1138
  );


  and
  g1933
  (
    n1901,
    n1117,
    n1771,
    n1623,
    n1787
  );


  nor
  g1934
  (
    n1948,
    n1623,
    n1630,
    n1830,
    n1073
  );


  xor
  g1935
  (
    n1956,
    n1769,
    n1173,
    n1062,
    n1075
  );


  or
  g1936
  (
    n1980,
    n1624,
    n1872,
    n1826,
    n1625
  );


  nand
  g1937
  (
    n1902,
    n1874,
    n1154,
    n1060,
    n1172
  );


  nand
  g1938
  (
    n1968,
    n1102,
    n1125,
    n1628,
    n1174
  );


  and
  g1939
  (
    n1975,
    n1813,
    n1786,
    n1779,
    n1844
  );


  xnor
  g1940
  (
    n1989,
    n1879,
    n1778,
    n1810,
    n1146
  );


  and
  g1941
  (
    n1905,
    n1171,
    n1626,
    n1884,
    n1054
  );


  and
  g1942
  (
    n1940,
    n1069,
    n1064,
    n1147,
    n1106
  );


  nand
  g1943
  (
    n1900,
    n1087,
    n1064,
    n1181,
    n1174
  );


  and
  g1944
  (
    n1957,
    n1127,
    n1079,
    n1106,
    n1055
  );


  or
  g1945
  (
    n1954,
    n1100,
    n1842,
    n1783,
    n1165
  );


  nor
  g1946
  (
    n1942,
    n1812,
    n1146,
    n1878,
    n1170
  );


  nor
  g1947
  (
    n1985,
    n1798,
    n1801,
    n1757,
    n1116
  );


  or
  g1948
  (
    n1996,
    n1795,
    n1171,
    n1629,
    n1104
  );


  xor
  g1949
  (
    n1917,
    n1049,
    n1083,
    n1625,
    n1863
  );


  or
  g1950
  (
    n1898,
    n1153,
    n1110,
    n1755,
    n1841
  );


  xor
  g1951
  (
    n1928,
    n1634,
    n1806,
    n1050,
    n1862
  );


  or
  g1952
  (
    n1966,
    n1155,
    n1074,
    n1835,
    n1128
  );


  nand
  g1953
  (
    n1999,
    n1098,
    n1047,
    n1867,
    n1802
  );


  nor
  g1954
  (
    n1918,
    n1129,
    n1142,
    n1873,
    n1071
  );


  or
  g1955
  (
    n1912,
    n1751,
    n1137,
    n1819,
    n1851
  );


  xor
  g1956
  (
    n1963,
    n1800,
    n1765,
    n1119,
    n1180
  );


  nand
  g1957
  (
    n1927,
    n1179,
    n1856,
    n1820,
    n1052
  );


  and
  g1958
  (
    n1983,
    n1766,
    n1108,
    n1859,
    n1045
  );


  xnor
  g1959
  (
    n1919,
    n1083,
    n1627,
    n1161,
    n1749
  );


  xnor
  g1960
  (
    n1922,
    n1834,
    n1821,
    n1149,
    n1627
  );


  or
  g1961
  (
    n1982,
    n1886,
    n1133,
    n1132,
    n1138
  );


  xor
  g1962
  (
    n1944,
    n1055,
    n1141,
    n1061,
    n1178
  );


  nor
  g1963
  (
    n1947,
    n1090,
    n1181,
    n1151,
    n1818
  );


  xor
  g1964
  (
    n1981,
    n1850,
    n1107,
    n1159,
    n1773
  );


  nand
  g1965
  (
    n1909,
    n1086,
    n1633,
    n1092,
    n1628
  );


  and
  g1966
  (
    n1910,
    n1163,
    n1113,
    n1081,
    n1880
  );


  and
  g1967
  (
    n1993,
    n1150,
    n1152,
    n1748,
    n1158
  );


  nand
  g1968
  (
    n1992,
    n1160,
    n1827,
    n1115,
    n1861
  );


  and
  g1969
  (
    n1896,
    n1158,
    n1852,
    n1177,
    n1085
  );


  xnor
  g1970
  (
    n1995,
    n1837,
    n1624,
    n1140,
    n1157
  );


  xor
  g1971
  (
    n2030,
    n1991,
    n1897,
    n1893,
    n1894
  );


  or
  g1972
  (
    n2008,
    n1984,
    n1961,
    n1949,
    n1934
  );


  xnor
  g1973
  (
    n2032,
    n1924,
    n1977,
    n1923,
    n2002
  );


  xnor
  g1974
  (
    n2027,
    n1992,
    n1953,
    n1936,
    n1922
  );


  and
  g1975
  (
    n2025,
    n1948,
    n1963,
    n1909,
    n1969
  );


  nor
  g1976
  (
    n2020,
    n1906,
    n1929,
    n1890,
    n1899
  );


  or
  g1977
  (
    n2004,
    n1937,
    n1965,
    n1892,
    n1968
  );


  nor
  g1978
  (
    n2024,
    n1966,
    n1938,
    n1927,
    n1939
  );


  xnor
  g1979
  (
    n2022,
    n1935,
    n1970,
    n1898,
    n1981
  );


  xnor
  g1980
  (
    n2013,
    n1987,
    n1913,
    n1996,
    n1914
  );


  and
  g1981
  (
    n2023,
    n1978,
    n1976,
    n1955,
    n1960
  );


  nor
  g1982
  (
    n2016,
    n1990,
    n1988,
    n1904,
    n1905
  );


  nor
  g1983
  (
    n2012,
    n1980,
    n1989,
    n1896,
    n1926
  );


  nand
  g1984
  (
    n2006,
    n1907,
    n1947,
    n1908,
    n1903
  );


  and
  g1985
  (
    n2005,
    n1888,
    n1986,
    n1917,
    n1925
  );


  xor
  g1986
  (
    n2021,
    n1999,
    n1982,
    n1958,
    n1933
  );


  and
  g1987
  (
    n2010,
    n1891,
    n1983,
    n1997,
    n1956
  );


  nor
  g1988
  (
    n2026,
    n1943,
    n1951,
    n1971,
    n1920
  );


  xor
  g1989
  (
    n2017,
    n1889,
    n1918,
    n1952,
    n1957
  );


  and
  g1990
  (
    n2031,
    n1919,
    n1942,
    n1912,
    n1915
  );


  nand
  g1991
  (
    n2029,
    n1972,
    n1901,
    n2000,
    n1973
  );


  and
  g1992
  (
    n2009,
    n1946,
    n1979,
    n1944,
    n1985
  );


  xor
  g1993
  (
    n2015,
    n1967,
    n1998,
    n1930,
    n1964
  );


  xnor
  g1994
  (
    n2019,
    n1959,
    n1975,
    n1902,
    n1921
  );


  or
  g1995
  (
    n2018,
    n2003,
    n1932,
    n1974,
    n1940
  );


  nand
  g1996
  (
    n2014,
    n1931,
    n1995,
    n2001,
    n1916
  );


  nor
  g1997
  (
    n2007,
    n1910,
    n1950,
    n1962,
    n1994
  );


  nand
  g1998
  (
    n2011,
    n1928,
    n1945,
    n1954,
    n1941
  );


  xnor
  g1999
  (
    n2028,
    n1993,
    n1911,
    n1895,
    n1900
  );


  xor
  KeyGate_0_0
  (
    n1911,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n978,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1768,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1353,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1773,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1626,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n188,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n329,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1102,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1946,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1261,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1237,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1061,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1481,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1383,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n784,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule

