

module Stat_100_65
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n90,
  n122,
  n125,
  n128,
  n131,
  n108,
  n102,
  n120,
  n105,
  n130,
  n115,
  n112,
  n121,
  n107,
  n117,
  n114,
  n113,
  n126,
  n119,
  n124,
  n111,
  n106,
  n123,
  n127,
  n104,
  n118,
  n129,
  n132,
  n109,
  n110,
  n116,
  n103,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n90;
  output n122;
  output n125;
  output n128;
  output n131;
  output n108;
  output n102;
  output n120;
  output n105;
  output n130;
  output n115;
  output n112;
  output n121;
  output n107;
  output n117;
  output n114;
  output n113;
  output n126;
  output n119;
  output n124;
  output n111;
  output n106;
  output n123;
  output n127;
  output n104;
  output n118;
  output n129;
  output n132;
  output n109;
  output n110;
  output n116;
  output n103;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    n40,
    n25
  );


  not
  g1
  (
    KeyWire_0_17,
    n23
  );


  buf
  g2
  (
    KeyWire_0_3,
    n1
  );


  buf
  g3
  (
    n36,
    n6
  );


  buf
  g4
  (
    n38,
    n19
  );


  buf
  g5
  (
    KeyWire_0_8,
    n13
  );


  buf
  g6
  (
    n50,
    n31
  );


  buf
  g7
  (
    KeyWire_0_30,
    n30
  );


  not
  g8
  (
    n51,
    n21
  );


  buf
  g9
  (
    n33,
    n8
  );


  not
  g10
  (
    n42,
    n9
  );


  not
  g11
  (
    n45,
    n4
  );


  not
  g12
  (
    n35,
    n20
  );


  buf
  g13
  (
    n44,
    n7
  );


  and
  g14
  (
    n39,
    n26,
    n22
  );


  nor
  g15
  (
    KeyWire_0_23,
    n18,
    n32,
    n3,
    n24
  );


  and
  g16
  (
    n49,
    n11,
    n16,
    n29,
    n10
  );


  nand
  g17
  (
    KeyWire_0_18,
    n28,
    n27,
    n15,
    n17
  );


  xnor
  g18
  (
    n47,
    n14,
    n2,
    n12,
    n5
  );


  not
  g19
  (
    n58,
    n34
  );


  not
  g20
  (
    n81,
    n44
  );


  buf
  g21
  (
    KeyWire_0_26,
    n42
  );


  buf
  g22
  (
    n52,
    n41
  );


  not
  g23
  (
    n87,
    n39
  );


  not
  g24
  (
    n76,
    n42
  );


  not
  g25
  (
    n62,
    n46
  );


  buf
  g26
  (
    KeyWire_0_2,
    n48
  );


  not
  g27
  (
    n56,
    n44
  );


  buf
  g28
  (
    n66,
    n44
  );


  not
  g29
  (
    KeyWire_0_29,
    n45
  );


  buf
  g30
  (
    n83,
    n36
  );


  not
  g31
  (
    n57,
    n33
  );


  not
  g32
  (
    n86,
    n36
  );


  buf
  g33
  (
    n71,
    n39
  );


  not
  g34
  (
    n84,
    n40
  );


  buf
  g35
  (
    KeyWire_0_4,
    n46
  );


  buf
  g36
  (
    KeyWire_0_11,
    n47
  );


  not
  g37
  (
    n63,
    n40
  );


  buf
  g38
  (
    KeyWire_0_25,
    n36
  );


  buf
  g39
  (
    n88,
    n34
  );


  buf
  g40
  (
    KeyWire_0_13,
    n37
  );


  not
  g41
  (
    n73,
    n37
  );


  not
  g42
  (
    n53,
    n47
  );


  not
  g43
  (
    n77,
    n35
  );


  buf
  g44
  (
    n69,
    n38
  );


  not
  g45
  (
    n75,
    n43
  );


  not
  g46
  (
    n70,
    n38
  );


  buf
  g47
  (
    n54,
    n42
  );


  buf
  g48
  (
    KeyWire_0_22,
    n45
  );


  buf
  g49
  (
    n80,
    n33
  );


  not
  g50
  (
    n61,
    n34
  );


  not
  g51
  (
    n59,
    n38
  );


  not
  g52
  (
    KeyWire_0_28,
    n33
  );


  nand
  g53
  (
    n72,
    n45,
    n47,
    n41
  );


  xor
  g54
  (
    n79,
    n40,
    n35,
    n37,
    n39
  );


  and
  g55
  (
    n65,
    n35,
    n46,
    n43
  );


  not
  g56
  (
    KeyWire_0_0,
    n54
  );


  buf
  g57
  (
    n90,
    n53
  );


  nand
  g58
  (
    KeyWire_0_21,
    n52,
    n53
  );


  buf
  g59
  (
    n92,
    n91
  );


  not
  g60
  (
    KeyWire_0_10,
    n90
  );


  or
  g61
  (
    KeyWire_0_14,
    n57,
    n54
  );


  and
  g62
  (
    KeyWire_0_5,
    n51,
    n93,
    n55,
    n48
  );


  xnor
  g63
  (
    n100,
    n92,
    n57,
    n55,
    n54
  );


  and
  g64
  (
    n97,
    n49,
    n56,
    n50,
    n57
  );


  nor
  g65
  (
    KeyWire_0_15,
    n92,
    n51,
    n50,
    n55
  );


  xor
  g66
  (
    n95,
    n49,
    n49,
    n51,
    n50
  );


  xor
  g67
  (
    n101,
    n93,
    n92,
    n56
  );


  xor
  g68
  (
    n96,
    n56,
    n93,
    n48
  );


  nand
  g69
  (
    n109,
    n87,
    n71,
    n97,
    n72
  );


  or
  g70
  (
    n132,
    n100,
    n83,
    n68,
    n96
  );


  xnor
  g71
  (
    KeyWire_0_9,
    n58,
    n100,
    n67,
    n86
  );


  nor
  g72
  (
    n115,
    n95,
    n100,
    n66
  );


  nand
  g73
  (
    n121,
    n88,
    n84,
    n85,
    n74
  );


  and
  g74
  (
    n128,
    n98,
    n63,
    n101,
    n69
  );


  or
  g75
  (
    n107,
    n77,
    n71,
    n64,
    n62
  );


  and
  g76
  (
    KeyWire_0_24,
    n83,
    n65,
    n99,
    n95
  );


  xor
  g77
  (
    KeyWire_0_16,
    n72,
    n96,
    n95,
    n73
  );


  nor
  g78
  (
    n131,
    n80,
    n97,
    n70,
    n87
  );


  xor
  g79
  (
    n125,
    n101,
    n82,
    n86,
    n68
  );


  nor
  g80
  (
    n116,
    n77,
    n67,
    n78,
    n85
  );


  nor
  g81
  (
    KeyWire_0_7,
    n98,
    n97,
    n74,
    n76
  );


  xnor
  g82
  (
    n113,
    n86,
    n99,
    n59,
    n79
  );


  or
  g83
  (
    n111,
    n58,
    n58,
    n59,
    n88
  );


  or
  g84
  (
    KeyWire_0_12,
    n59,
    n74,
    n72,
    n65
  );


  nand
  g85
  (
    KeyWire_0_27,
    n61,
    n94,
    n80,
    n75
  );


  and
  g86
  (
    KeyWire_0_1,
    n71,
    n69,
    n65,
    n79
  );


  nor
  g87
  (
    n105,
    n94,
    n95,
    n82,
    n84
  );


  and
  g88
  (
    n106,
    n96,
    n94,
    n63,
    n87
  );


  xor
  g89
  (
    n119,
    n99,
    n61,
    n62,
    n81
  );


  xor
  g90
  (
    n102,
    n83,
    n78,
    n98,
    n77
  );


  xnor
  g91
  (
    KeyWire_0_19,
    n73,
    n78,
    n64,
    n70
  );


  xor
  g92
  (
    n114,
    n99,
    n76,
    n96,
    n88
  );


  nor
  g93
  (
    KeyWire_0_31,
    n84,
    n70,
    n101,
    n80
  );


  or
  g94
  (
    n118,
    n60,
    n68,
    n81
  );


  xnor
  g95
  (
    n122,
    n62,
    n75,
    n97,
    n82
  );


  xor
  g96
  (
    n110,
    n75,
    n67,
    n63,
    n79
  );


  or
  g97
  (
    KeyWire_0_20,
    n73,
    n66,
    n76,
    n64
  );


  xnor
  g98
  (
    n124,
    n85,
    n61,
    n101,
    n69
  );


  xor
  g99
  (
    KeyWire_0_6,
    n100,
    n60,
    n98
  );


  xnor
  KeyGate_0_0
  (
    n89,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n103,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n64,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n41,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n74,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n94,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n120,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n104,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n46,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n123,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n93,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n67,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n126,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n55,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n98,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n99,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n117,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n34,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n43,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n127,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n129,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n91,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n82,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n48,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n130,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n78,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n85,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n112,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n60,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n68,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n37,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n108,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

