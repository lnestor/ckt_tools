// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_201 written by SynthGen on 2021/04/05 11:08:35
module Stat_1000_201( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n871, n847, n863, n850, n858, n841, n854, n852,
 n955, n966, n943, n965, n957, n956, n952, n958,
 n954, n961, n968, n946, n950, n970, n976, n973,
 n1021, n1025, n1023, n1028, n1031, n1030, n1032, n1029);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n871, n847, n863, n850, n858, n841, n854, n852,
 n955, n966, n943, n965, n957, n956, n952, n958,
 n954, n961, n968, n946, n950, n970, n976, n973,
 n1021, n1025, n1023, n1028, n1031, n1030, n1032, n1029;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n842, n843, n844, n845, n846, n848, n849, n851,
 n853, n855, n856, n857, n859, n860, n861, n862,
 n864, n865, n866, n867, n868, n869, n870, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n944, n945,
 n947, n948, n949, n951, n953, n959, n960, n962,
 n963, n964, n967, n969, n971, n972, n974, n975,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1022, n1024, n1026, n1027;

buf  g0 (n51, n6);
not  g1 (n70, n31);
buf  g2 (n131, n12);
not  g3 (n154, n1);
buf  g4 (n110, n7);
not  g5 (n113, n3);
not  g6 (n77, n31);
not  g7 (n105, n17);
not  g8 (n145, n7);
not  g9 (n78, n15);
not  g10 (n148, n18);
buf  g11 (n129, n26);
buf  g12 (n33, n11);
not  g13 (n128, n21);
not  g14 (n104, n3);
buf  g15 (n119, n31);
not  g16 (n97, n2);
buf  g17 (n120, n17);
buf  g18 (n138, n29);
buf  g19 (n48, n6);
buf  g20 (n90, n26);
not  g21 (n92, n24);
not  g22 (n144, n8);
buf  g23 (n80, n22);
not  g24 (n137, n25);
buf  g25 (n108, n8);
not  g26 (n151, n18);
buf  g27 (n107, n8);
buf  g28 (n50, n22);
not  g29 (n63, n9);
not  g30 (n62, n27);
not  g31 (n140, n13);
not  g32 (n123, n19);
buf  g33 (n85, n19);
buf  g34 (n156, n25);
not  g35 (n44, n18);
not  g36 (n114, n12);
buf  g37 (n112, n22);
not  g38 (n117, n5);
not  g39 (n57, n28);
buf  g40 (n139, n23);
buf  g41 (n155, n11);
buf  g42 (n126, n23);
not  g43 (n40, n13);
buf  g44 (n74, n5);
buf  g45 (n106, n16);
buf  g46 (n135, n1);
buf  g47 (n149, n25);
not  g48 (n49, n7);
buf  g49 (n86, n11);
buf  g50 (n45, n10);
buf  g51 (n143, n3);
buf  g52 (n41, n18);
not  g53 (n71, n29);
buf  g54 (n73, n10);
buf  g55 (n141, n4);
buf  g56 (n121, n5);
not  g57 (n58, n23);
not  g58 (n94, n24);
not  g59 (n47, n9);
buf  g60 (n118, n19);
not  g61 (n66, n28);
buf  g62 (n95, n27);
not  g63 (n87, n20);
buf  g64 (n133, n28);
not  g65 (n52, n29);
buf  g66 (n124, n21);
not  g67 (n98, n19);
not  g68 (n43, n17);
buf  g69 (n103, n22);
buf  g70 (n56, n26);
buf  g71 (n82, n12);
buf  g72 (n38, n14);
not  g73 (n81, n2);
buf  g74 (n134, n17);
buf  g75 (n147, n30);
buf  g76 (n67, n15);
buf  g77 (n35, n29);
not  g78 (n152, n27);
not  g79 (n64, n25);
not  g80 (n96, n4);
not  g81 (n91, n7);
buf  g82 (n142, n24);
not  g83 (n36, n21);
buf  g84 (n61, n23);
buf  g85 (n54, n10);
buf  g86 (n39, n16);
not  g87 (n65, n10);
not  g88 (n59, n32);
not  g89 (n122, n28);
not  g90 (n132, n14);
buf  g91 (n88, n4);
not  g92 (n102, n20);
buf  g93 (n109, n15);
not  g94 (n76, n30);
not  g95 (n72, n5);
buf  g96 (n84, n15);
not  g97 (n69, n30);
buf  g98 (n127, n9);
not  g99 (n55, n31);
buf  g100 (n116, n12);
not  g101 (n111, n6);
not  g102 (n146, n13);
not  g103 (n34, n21);
buf  g104 (n89, n20);
buf  g105 (n93, n9);
not  g106 (n100, n11);
buf  g107 (n53, n4);
not  g108 (n60, n20);
not  g109 (n153, n1);
buf  g110 (n79, n13);
buf  g111 (n42, n2);
not  g112 (n125, n24);
buf  g113 (n46, n16);
not  g114 (n83, n6);
not  g115 (n101, n30);
buf  g116 (n136, n14);
buf  g117 (n37, n3);
not  g118 (n75, n16);
not  g119 (n115, n14);
not  g120 (n99, n26);
not  g121 (n130, n27);
not  g122 (n150, n8);
buf  g123 (n68, n2);
buf  g124 (n236, n89);
not  g125 (n399, n81);
buf  g126 (n410, n117);
buf  g127 (n374, n52);
buf  g128 (n322, n154);
buf  g129 (n407, n39);
not  g130 (n212, n121);
not  g131 (n288, n85);
not  g132 (n245, n49);
not  g133 (n224, n126);
not  g134 (n257, n58);
not  g135 (n246, n66);
not  g136 (n300, n110);
not  g137 (n433, n41);
buf  g138 (n427, n135);
not  g139 (n392, n36);
not  g140 (n178, n35);
buf  g141 (n317, n40);
buf  g142 (n183, n106);
buf  g143 (n185, n151);
not  g144 (n434, n102);
not  g145 (n237, n126);
not  g146 (n174, n108);
buf  g147 (n309, n143);
buf  g148 (n318, n61);
buf  g149 (n342, n44);
buf  g150 (n331, n50);
not  g151 (n351, n150);
buf  g152 (n321, n128);
not  g153 (n217, n34);
buf  g154 (n296, n80);
buf  g155 (n388, n97);
not  g156 (n378, n152);
not  g157 (n219, n141);
not  g158 (n370, n145);
buf  g159 (n250, n39);
not  g160 (n394, n128);
buf  g161 (n170, n109);
not  g162 (n166, n114);
not  g163 (n382, n142);
buf  g164 (n179, n83);
not  g165 (n232, n50);
not  g166 (n403, n81);
buf  g167 (n228, n51);
not  g168 (n314, n115);
not  g169 (n262, n116);
not  g170 (n160, n149);
buf  g171 (n171, n74);
not  g172 (n371, n55);
buf  g173 (n240, n94);
not  g174 (n199, n84);
not  g175 (n249, n111);
buf  g176 (n325, n114);
buf  g177 (n337, n39);
buf  g178 (n426, n98);
not  g179 (n428, n33);
not  g180 (n406, n38);
not  g181 (n276, n104);
buf  g182 (n226, n121);
not  g183 (n292, n47);
buf  g184 (n443, n56);
not  g185 (n369, n57);
buf  g186 (n400, n36);
not  g187 (n347, n38);
buf  g188 (n281, n67);
buf  g189 (n381, n76);
not  g190 (n188, n99);
buf  g191 (n377, n147);
not  g192 (n293, n141);
buf  g193 (n405, n113);
buf  g194 (n176, n103);
not  g195 (n303, n75);
buf  g196 (n338, n55);
not  g197 (n316, n34);
buf  g198 (n420, n136);
not  g199 (n366, n134);
buf  g200 (n215, n95);
buf  g201 (n299, n115);
not  g202 (n329, n33);
not  g203 (n326, n127);
not  g204 (n286, n144);
buf  g205 (n421, n154);
buf  g206 (n398, n122);
buf  g207 (n157, n73);
buf  g208 (n423, n49);
buf  g209 (n206, n60);
not  g210 (n162, n130);
buf  g211 (n290, n75);
not  g212 (n247, n130);
buf  g213 (n213, n82);
not  g214 (n356, n50);
buf  g215 (n235, n51);
not  g216 (n279, n153);
buf  g217 (n256, n139);
not  g218 (n163, n82);
not  g219 (n354, n71);
not  g220 (n208, n83);
buf  g221 (n308, n153);
not  g222 (n263, n104);
not  g223 (n319, n69);
buf  g224 (n415, n138);
buf  g225 (n436, n37);
not  g226 (n203, n102);
not  g227 (n209, n95);
not  g228 (n181, n47);
buf  g229 (n343, n53);
not  g230 (n190, n118);
buf  g231 (n417, n100);
buf  g232 (n275, n70);
not  g233 (n442, n111);
buf  g234 (n412, n41);
buf  g235 (n386, n83);
not  g236 (n207, n135);
buf  g237 (n327, n72);
buf  g238 (n201, n127);
not  g239 (n419, n142);
buf  g240 (n324, n153);
buf  g241 (n254, n57);
buf  g242 (n367, n148);
buf  g243 (n175, n62);
buf  g244 (n159, n68);
buf  g245 (n169, n54);
not  g246 (n221, n145);
buf  g247 (n204, n95);
not  g248 (n306, n72);
not  g249 (n233, n97);
buf  g250 (n211, n147);
not  g251 (n383, n35);
not  g252 (n258, n152);
not  g253 (n198, n66);
buf  g254 (n333, n46);
buf  g255 (n271, n71);
not  g256 (n267, n131);
not  g257 (n202, n94);
buf  g258 (n395, n151);
not  g259 (n380, n140);
not  g260 (n350, n48);
not  g261 (n283, n137);
not  g262 (n313, n143);
buf  g263 (n205, n93);
not  g264 (n251, n133);
buf  g265 (n365, n92);
not  g266 (n411, n147);
buf  g267 (n304, n52);
not  g268 (n172, n48);
buf  g269 (n298, n72);
buf  g270 (n429, n101);
buf  g271 (n297, n67);
buf  g272 (n241, n149);
not  g273 (n424, n129);
buf  g274 (n362, n146);
not  g275 (n242, n63);
not  g276 (n387, n122);
not  g277 (n282, n148);
not  g278 (n401, n68);
buf  g279 (n334, n129);
not  g280 (n260, n94);
buf  g281 (n345, n44);
not  g282 (n189, n140);
buf  g283 (n220, n86);
buf  g284 (n408, n52);
buf  g285 (n359, n105);
buf  g286 (n344, n132);
not  g287 (n280, n51);
not  g288 (n285, n55);
not  g289 (n200, n69);
not  g290 (n210, n42);
not  g291 (n158, n91);
buf  g292 (n268, n116);
not  g293 (n384, n133);
not  g294 (n244, n109);
buf  g295 (n368, n135);
not  g296 (n379, n128);
buf  g297 (n441, n107);
not  g298 (n252, n107);
buf  g299 (n349, n132);
not  g300 (n414, n113);
buf  g301 (n375, n96);
buf  g302 (n230, n146);
buf  g303 (n389, n108);
not  g304 (n278, n100);
not  g305 (n165, n42);
not  g306 (n358, n85);
not  g307 (n413, n149);
buf  g308 (n302, n34);
buf  g309 (n255, n119);
not  g310 (n301, n151);
buf  g311 (n216, n37);
buf  g312 (n161, n125);
not  g313 (n231, n87);
buf  g314 (n191, n86);
buf  g315 (n335, n59);
buf  g316 (n167, n58);
not  g317 (n346, n124);
buf  g318 (n432, n140);
not  g319 (n248, n40);
buf  g320 (n376, n88);
not  g321 (n409, n108);
buf  g322 (n364, n59);
buf  g323 (n438, n131);
not  g324 (n194, n117);
not  g325 (n284, n65);
not  g326 (n265, n56);
buf  g327 (n440, n61);
buf  g328 (n312, n38);
not  g329 (n402, n110);
buf  g330 (n239, n106);
buf  g331 (n273, n111);
not  g332 (n332, n154);
buf  g333 (n192, n133);
buf  g334 (n348, n124);
buf  g335 (n393, n91);
buf  g336 (n289, n112);
not  g337 (n307, n115);
not  g338 (n397, n35);
buf  g339 (n272, n91);
not  g340 (n270, n130);
not  g341 (n391, n137);
not  g342 (n363, n139);
buf  g343 (n404, n123);
buf  g344 (n339, n87);
buf  g345 (n336, n54);
buf  g346 (n385, n90);
buf  g347 (n253, n112);
not  g348 (n195, n126);
buf  g349 (n187, n141);
buf  g350 (n355, n88);
not  g351 (n291, n42);
buf  g352 (n164, n79);
not  g353 (n182, n86);
buf  g354 (n340, n106);
not  g355 (n277, n93);
buf  g356 (n180, n144);
not  g357 (n227, n74);
buf  g358 (n274, n110);
buf  g359 (n416, n58);
not  g360 (n444, n76);
not  g361 (n222, n81);
buf  g362 (n294, n129);
not  g363 (n218, n134);
not  g364 (n430, n87);
not  g365 (n320, n75);
not  g366 (n177, n98);
not  g367 (n431, n99);
buf  g368 (n184, n125);
not  g369 (n261, n103);
not  g370 (n341, n114);
not  g371 (n225, n132);
not  g372 (n305, n37);
not  g373 (n295, n48);
buf  g374 (n197, n136);
buf  g375 (n223, n155);
buf  g376 (n310, n80);
buf  g377 (n196, n46);
buf  g378 (n425, n57);
buf  g379 (n357, n134);
not  g380 (n259, n118);
buf  g381 (n396, n93);
buf  g382 (n373, n90);
buf  g383 (n243, n60);
buf  g384 (n186, n78);
xor  g385 (n353, n41, n60);
xnor g386 (n437, n117, n33, n77, n113);
nand g387 (n229, n98, n45, n138, n85);
xor  g388 (n193, n150, n36, n146, n88);
xnor g389 (n323, n70, n67, n62, n79);
xnor g390 (n435, n53, n64, n145, n70);
or   g391 (n264, n121, n90, n79, n120);
nor  g392 (n330, n77, n53, n54, n62);
nand g393 (n372, n74, n49, n66, n143);
nand g394 (n168, n112, n82, n123, n89);
xnor g395 (n238, n102, n43, n122, n107);
xnor g396 (n287, n116, n65, n105, n43);
or   g397 (n361, n68, n119, n127, n64);
nand g398 (n352, n101, n44, n45);
or   g399 (n234, n46, n59, n73, n84);
xor  g400 (n422, n92, n96, n100);
xor  g401 (n311, n152, n63, n43, n65);
nand g402 (n390, n71, n137, n47, n123);
nand g403 (n173, n89, n78, n109);
and  g404 (n214, n99, n73, n142, n77);
nand g405 (n266, n101, n148, n63, n80);
or   g406 (n439, n131, n76, n92, n105);
or   g407 (n315, n64, n104, n120, n97);
xor  g408 (n269, n118, n150, n136, n69);
xnor g409 (n360, n120, n84, n103, n144);
xnor g410 (n418, n56, n124, n139, n61);
nand g411 (n328, n40, n125, n119, n138);
xor  g412 (n553, n274, n365, n330, n288);
nor  g413 (n509, n390, n184, n320, n346);
xor  g414 (n554, n272, n191, n179, n366);
nor  g415 (n450, n322, n361, n365, n168);
and  g416 (n447, n283, n197, n316, n311);
or   g417 (n490, n278, n292, n386, n260);
xnor g418 (n488, n165, n232, n213, n247);
or   g419 (n558, n262, n299, n234, n386);
or   g420 (n599, n229, n354, n230, n351);
nand g421 (n526, n263, n362, n270, n230);
xor  g422 (n583, n335, n394, n244, n393);
xnor g423 (n592, n374, n178, n275, n285);
or   g424 (n533, n254, n232, n332, n290);
or   g425 (n454, n385, n212, n215, n331);
and  g426 (n517, n382, n308, n276, n252);
xnor g427 (n467, n392, n372, n274, n316);
xor  g428 (n458, n202, n291, n282, n381);
nand g429 (n564, n334, n306, n293, n195);
xor  g430 (n565, n312, n289, n320, n261);
nand g431 (n576, n201, n393, n333, n377);
nand g432 (n487, n182, n357, n342, n372);
nor  g433 (n544, n199, n301, n277, n276);
nand g434 (n597, n249, n236, n318, n182);
nand g435 (n469, n396, n396, n283, n180);
xor  g436 (n477, n171, n248, n395, n169);
or   g437 (n507, n368, n255, n277, n328);
nand g438 (n545, n217, n372, n315, n392);
nor  g439 (n522, n161, n288, n257, n211);
nand g440 (n459, n284, n395, n292, n307);
nor  g441 (n465, n300, n302, n364, n309);
and  g442 (n537, n259, n241, n173, n308);
nand g443 (n571, n352, n199, n190, n254);
nand g444 (n481, n363, n183, n394, n373);
and  g445 (n499, n345, n366, n390, n175);
xnor g446 (n505, n298, n253, n387, n187);
nor  g447 (n491, n297, n332, n388, n357);
xor  g448 (n542, n386, n267, n172, n266);
xnor g449 (n562, n231, n387, n296, n345);
nand g450 (n575, n279, n158, n185, n253);
and  g451 (n478, n242, n302, n387, n158);
or   g452 (n574, n157, n212, n368, n381);
xnor g453 (n483, n318, n286, n364, n383);
xor  g454 (n588, n258, n172, n162, n242);
nand g455 (n559, n338, n169, n240, n207);
and  g456 (n600, n220, n319, n163, n346);
xor  g457 (n446, n265, n175, n285, n223);
and  g458 (n540, n316, n350, n297, n166);
and  g459 (n535, n181, n185, n180, n384);
or   g460 (n510, n243, n270, n351, n353);
xnor g461 (n550, n167, n215, n268, n304);
nand g462 (n474, n289, n375, n234, n296);
or   g463 (n548, n360, n341, n373, n259);
xnor g464 (n513, n282, n334, n317, n319);
or   g465 (n561, n221, n251, n218, n241);
and  g466 (n568, n326, n318, n299, n164);
xnor g467 (n578, n320, n183, n225, n160);
and  g468 (n515, n378, n356, n210, n396);
and  g469 (n518, n330, n257, n173, n290);
nor  g470 (n536, n233, n379, n323);
xnor g471 (n464, n262, n359, n354, n310);
nor  g472 (n572, n267, n312, n245, n382);
nand g473 (n496, n343, n348, n222, n336);
and  g474 (n506, n192, n305, n166, n304);
and  g475 (n475, n355, n361, n250, n176);
xor  g476 (n557, n192, n293, n252, n321);
or   g477 (n460, n284, n294, n340, n303);
or   g478 (n586, n314, n236, n174, n258);
xor  g479 (n479, n295, n374, n174, n287);
nand g480 (n591, n378, n189, n295, n280);
xnor g481 (n589, n214, n296, n325, n339);
and  g482 (n525, n306, n397, n377, n328);
and  g483 (n551, n159, n321, n195, n293);
nand g484 (n449, n272, n206, n382, n246);
and  g485 (n529, n177, n339, n371, n163);
xnor g486 (n451, n209, n340, n251, n356);
xnor g487 (n471, n333, n268, n353, n346);
nand g488 (n470, n395, n184, n349, n295);
nor  g489 (n511, n325, n196, n377, n216);
nand g490 (n452, n304, n365, n221, n193);
nand g491 (n569, n392, n256, n362, n194);
xnor g492 (n566, n383, n275, n385, n343);
nand g493 (n555, n191, n312, n309, n314);
xnor g494 (n567, n351, n347, n266, n373);
nor  g495 (n519, n343, n287, n326, n194);
nor  g496 (n539, n264, n219, n335, n348);
or   g497 (n585, n269, n285, n203, n176);
or   g498 (n560, n235, n208, n266, n267);
xor  g499 (n579, n201, n376, n352, n247);
xnor g500 (n455, n281, n324, n352, n338);
and  g501 (n531, n347, n301, n336, n292);
xnor g502 (n527, n282, n389, n278, n193);
nor  g503 (n573, n273, n257, n186, n376);
or   g504 (n472, n181, n294, n337, n210);
nand g505 (n570, n367, n385, n324, n391);
and  g506 (n486, n313, n283, n381, n272);
and  g507 (n530, n256, n379, n190, n289);
xor  g508 (n594, n311, n356, n202, n238);
xnor g509 (n508, n237, n305, n342, n229);
nand g510 (n497, n369, n198, n349, n239);
nor  g511 (n514, n261, n369, n329, n393);
nor  g512 (n590, n275, n235, n279, n348);
nand g513 (n524, n265, n220, n269, n188);
nand g514 (n453, n265, n273, n164, n177);
and  g515 (n448, n228, n213, n286, n340);
or   g516 (n456, n345, n358, n363, n357);
xor  g517 (n543, n354, n313, n189, n226);
and  g518 (n484, n157, n271, n314, n281);
or   g519 (n556, n211, n350, n233, n256);
xor  g520 (n523, n170, n205, n206, n200);
nand g521 (n457, n380, n264, n227, n310);
xnor g522 (n463, n279, n325, n198, n291);
xnor g523 (n462, n287, n260, n331, n171);
nor  g524 (n596, n162, n226, n246, n294);
xor  g525 (n532, n336, n208, n355, n260);
xnor g526 (n587, n219, n204, n390, n239);
or   g527 (n503, n341, n300, n360, n259);
or   g528 (n445, n324, n248, n380, n326);
nand g529 (n521, n355, n167, n353, n306);
xor  g530 (n563, n187, n327, n376, n159);
xnor g531 (n528, n317, n337, n397, n244);
xnor g532 (n476, n261, n371, n209, n301);
xor  g533 (n495, n371, n364, n280, n310);
nand g534 (n500, n263, n268, n350, n224);
and  g535 (n582, n305, n297, n178, n307);
xnor g536 (n595, n245, n271, n224, n363);
nor  g537 (n498, n338, n335, n264, n391);
or   g538 (n473, n302, n327, n331, n328);
xnor g539 (n547, n160, n308, n231, n367);
xnor g540 (n502, n311, n374, n227, n378);
nor  g541 (n492, n339, n280, n360, n271);
xnor g542 (n512, n222, n298, n367);
and  g543 (n461, n375, n262, n223, n361);
and  g544 (n493, n362, n228, n379, n315);
or   g545 (n546, n237, n388, n359, n384);
xnor g546 (n549, n288, n214, n369, n286);
nand g547 (n552, n217, n258, n330, n225);
nor  g548 (n468, n370, n276, n329, n344);
xor  g549 (n501, n307, n165, n216, n290);
and  g550 (n494, n309, n315, n359, n334);
xnor g551 (n485, n196, n341, n300, n332);
nand g552 (n593, n263, n329, n388, n273);
xor  g553 (n489, n218, n370, n270, n333);
and  g554 (n482, n322, n358, n284, n375);
xnor g555 (n534, n368, n319, n383, n322);
and  g556 (n516, n207, n278, n274, n337);
xnor g557 (n577, n303, n281, n179, n391);
and  g558 (n466, n323, n317, n349, n389);
nand g559 (n480, n291, n250, n170, n168);
xor  g560 (n580, n321, n204, n370, n389);
or   g561 (n520, n344, n186, n238, n161);
nand g562 (n504, n240, n313, n344, n205);
and  g563 (n581, n200, n255, n384, n188);
nor  g564 (n538, n397, n394, n380, n327);
and  g565 (n598, n347, n358, n249, n269);
or   g566 (n584, n277, n203, n303, n342);
or   g567 (n541, n243, n366, n299, n197);
buf  g568 (n614, n480);
buf  g569 (n676, n471);
not  g570 (n632, n483);
not  g571 (n699, n577);
buf  g572 (n675, n531);
buf  g573 (n666, n530);
not  g574 (n636, n569);
not  g575 (n628, n551);
buf  g576 (n645, n524);
buf  g577 (n672, n523);
buf  g578 (n634, n596);
not  g579 (n613, n595);
not  g580 (n706, n487);
buf  g581 (n629, n538);
not  g582 (n667, n546);
not  g583 (n647, n591);
not  g584 (n607, n567);
not  g585 (n609, n518);
buf  g586 (n704, n495);
buf  g587 (n601, n593);
buf  g588 (n688, n453);
buf  g589 (n610, n552);
buf  g590 (n650, n579);
not  g591 (n651, n562);
not  g592 (n661, n535);
buf  g593 (n640, n541);
buf  g594 (n653, n593);
buf  g595 (n631, n595);
not  g596 (n633, n560);
not  g597 (n641, n555);
buf  g598 (n689, n527);
not  g599 (n649, n554);
not  g600 (n627, n546);
not  g601 (n707, n505);
buf  g602 (n696, n504);
buf  g603 (n700, n600);
buf  g604 (n665, n581);
not  g605 (n616, n597);
buf  g606 (n659, n538);
buf  g607 (n652, n577);
buf  g608 (n695, n525);
buf  g609 (n677, n581);
buf  g610 (n639, n510);
buf  g611 (n658, n584);
not  g612 (n657, n594);
buf  g613 (n617, n463);
buf  g614 (n680, n587);
not  g615 (n693, n502);
not  g616 (n626, n481);
buf  g617 (n606, n456);
not  g618 (n608, n490);
buf  g619 (n669, n455);
buf  g620 (n654, n573);
not  g621 (n690, n469);
buf  g622 (n674, n528);
not  g623 (n604, n568);
not  g624 (n670, n559);
buf  g625 (n687, n493);
not  g626 (n681, n494);
not  g627 (n698, n470);
not  g628 (n630, n547);
buf  g629 (n637, n497);
buf  g630 (n644, n592);
buf  g631 (n621, n457);
buf  g632 (n703, n565);
not  g633 (n622, n539);
buf  g634 (n663, n503);
not  g635 (n664, n561);
not  g636 (n710, n534);
buf  g637 (n643, n492);
not  g638 (n602, n553);
nor  g639 (n697, n563, n576, n543, n552);
xor  g640 (n611, n536, n600, n526, n554);
xnor g641 (n625, n501, n446, n474, n589);
or   g642 (n702, n567, n450, n566, n475);
nand g643 (n655, n516, n467, n485, n568);
nor  g644 (n671, n536, n520, n556, n569);
and  g645 (n684, n539, n541, n461, n599);
and  g646 (n692, n570, n556, n550, n540);
or   g647 (n642, n584, n543, n557, n445);
nor  g648 (n708, n589, n573, n590, n558);
nor  g649 (n660, n496, n508, n553, n537);
nor  g650 (n662, n563, n564, n557, n521);
or   g651 (n678, n533, n571, n580, n489);
xor  g652 (n615, n533, n507, n544, n560);
nor  g653 (n605, n500, n572, n545, n486);
or   g654 (n682, n462, n562, n561, n513);
or   g655 (n668, n534, n515, n590, n537);
nor  g656 (n691, n473, n449, n558, n571);
xnor g657 (n648, n594, n522, n548, n596);
and  g658 (n686, n532, n578, n452, n545);
nor  g659 (n701, n597, n551, n570, n565);
or   g660 (n673, n509, n465, n459, n550);
nor  g661 (n618, n466, n519, n476, n511);
nor  g662 (n635, n512, n542, n598, n549);
and  g663 (n603, n529, n588, n506, n464);
or   g664 (n612, n586, n532, n591, n542);
or   g665 (n679, n599, n549, n488, n448);
xnor g666 (n624, n559, n451, n530, n454);
xor  g667 (n620, n572, n583, n544, n535);
or   g668 (n694, n479, n585, n499, n468);
nand g669 (n646, n578, n472, n547, n484);
xnor g670 (n619, n566, n548, n517, n498);
or   g671 (n709, n586, n585, n582, n477);
or   g672 (n623, n576, n575, n540, n580);
and  g673 (n638, n514, n579, n598, n575);
and  g674 (n656, n460, n583, n491, n478);
or   g675 (n683, n587, n588, n458, n555);
or   g676 (n705, n582, n592, n574);
and  g677 (n685, n564, n482, n447, n531);
xnor g678 (n714, n613, n603, n610);
xnor g679 (n717, n616, n604, n607, n615);
xnor g680 (n715, n606, n613, n614, n608);
xnor g681 (n712, n617, n605, n613, n611);
nor  g682 (n716, n607, n612, n615, n602);
xnor g683 (n719, n603, n609, n605, n615);
or   g684 (n711, n602, n616, n612, n608);
nand g685 (n718, n602, n610, n604, n616);
xnor g686 (n720, n608, n611, n605, n609);
nand g687 (n713, n614, n606, n601, n611);
or   g688 (n722, n610, n614, n609, n601);
xor  g689 (n721, n612, n606, n607, n604);
not  g690 (n743, n716);
buf  g691 (n734, n716);
not  g692 (n730, n711);
not  g693 (n744, n714);
not  g694 (n729, n713);
not  g695 (n732, n719);
not  g696 (n727, n712);
not  g697 (n731, n717);
buf  g698 (n723, n713);
not  g699 (n726, n715);
not  g700 (n725, n717);
not  g701 (n735, n711);
not  g702 (n738, n718);
not  g703 (n737, n715);
buf  g704 (n733, n714);
buf  g705 (n742, n718);
not  g706 (n728, n714);
buf  g707 (n736, n716);
not  g708 (n741, n712);
not  g709 (n724, n718);
buf  g710 (n739, n715);
buf  g711 (n740, n717);
xnor g712 (n794, n742, n645, n681, n740);
or   g713 (n797, n631, n653, n744, n618);
or   g714 (n771, n650, n741, n623, n672);
nor  g715 (n747, n738, n734, n742, n732);
xnor g716 (n792, n634, n739, n665, n740);
xor  g717 (n767, n743, n636, n682, n639);
xor  g718 (n803, n737, n740, n617, n666);
and  g719 (n785, n644, n648, n637, n732);
nor  g720 (n796, n743, n653, n644, n737);
nand g721 (n802, n670, n739, n654, n678);
xor  g722 (n759, n677, n618, n647, n739);
nor  g723 (n775, n678, n641, n728, n741);
xnor g724 (n750, n736, n744, n652, n673);
nand g725 (n812, n729, n736, n656, n676);
xor  g726 (n799, n678, n617, n649, n645);
nand g727 (n774, n653, n732, n677, n734);
nand g728 (n795, n621, n650, n676, n636);
or   g729 (n763, n643, n657, n728, n641);
nor  g730 (n784, n655, n669, n640, n635);
or   g731 (n778, n736, n671, n723, n662);
or   g732 (n772, n668, n724, n674, n682);
nand g733 (n814, n657, n680, n740, n682);
nor  g734 (n748, n628, n621, n663, n726);
nor  g735 (n761, n735, n732, n658, n662);
xnor g736 (n758, n619, n731, n663, n659);
nor  g737 (n813, n643, n738, n648, n673);
nor  g738 (n782, n658, n628, n624, n672);
xor  g739 (n764, n661, n629, n664, n739);
nor  g740 (n769, n625, n629, n642, n622);
nor  g741 (n777, n731, n631, n671, n665);
or   g742 (n805, n727, n624, n652, n656);
or   g743 (n765, n730, n730, n669, n633);
nor  g744 (n745, n724, n656, n735, n727);
nand g745 (n756, n622, n681, n620, n632);
and  g746 (n789, n625, n658, n679, n743);
and  g747 (n800, n636, n730, n742, n735);
and  g748 (n760, n726, n651, n649, n741);
xor  g749 (n753, n670, n633, n651, n664);
or   g750 (n807, n637, n675, n627, n726);
and  g751 (n773, n667, n647, n729, n666);
xor  g752 (n801, n628, n632, n619, n625);
or   g753 (n798, n627, n660, n725, n646);
and  g754 (n762, n676, n669, n622, n634);
nor  g755 (n776, n677, n741, n734, n727);
or   g756 (n811, n723, n674, n635, n727);
and  g757 (n806, n674, n627, n743, n638);
and  g758 (n746, n733, n633, n623, n632);
xor  g759 (n752, n733, n725, n728, n626);
xnor g760 (n770, n737, n726, n629, n725);
nand g761 (n783, n670, n665, n639, n646);
or   g762 (n755, n634, n659, n650, n639);
xnor g763 (n766, n649, n654, n624, n734);
or   g764 (n768, n662, n642, n637, n652);
or   g765 (n780, n663, n666, n744, n630);
nor  g766 (n791, n661, n724, n644, n681);
nand g767 (n815, n630, n744, n672, n671);
and  g768 (n790, n731, n655, n646, n647);
nor  g769 (n779, n679, n648, n730, n620);
xor  g770 (n804, n651, n724, n728, n638);
nor  g771 (n793, n619, n738, n668, n729);
nor  g772 (n781, n630, n725, n723, n742);
xnor g773 (n749, n731, n660, n621, n733);
and  g774 (n754, n675, n664, n680, n642);
and  g775 (n810, n655, n626, n640, n673);
xor  g776 (n788, n631, n679, n729, n657);
nor  g777 (n809, n661, n626, n640, n735);
and  g778 (n751, n638, n618, n680, n635);
xor  g779 (n787, n623, n620, n737, n641);
nor  g780 (n757, n645, n667, n675);
xor  g781 (n808, n659, n733, n654, n660);
xnor g782 (n786, n738, n668, n736, n643);
nor  g783 (n823, n756, n748, n754, n745);
nor  g784 (n827, n757, n769, n760, n755);
xor  g785 (n820, n752, n775, n782, n767);
xor  g786 (n832, n766, n768, n767, n751);
or   g787 (n825, n776, n780, n781, n750);
nand g788 (n828, n779, n753, n764, n777);
nand g789 (n836, n758, n759, n753, n765);
and  g790 (n824, n773, n785, n745, n757);
or   g791 (n826, n754, n784, n749, n772);
xor  g792 (n822, n786, n747, n780, n768);
and  g793 (n821, n765, n762, n752, n774);
and  g794 (n817, n770, n784, n773, n772);
nand g795 (n829, n774, n776, n746, n781);
nand g796 (n816, n778, n783, n777, n747);
or   g797 (n834, n785, n760, n763, n746);
nand g798 (n819, n761, n759, n770, n766);
or   g799 (n830, n786, n762, n756, n771);
or   g800 (n831, n778, n750, n764, n763);
nor  g801 (n835, n783, n761, n771, n751);
xnor g802 (n818, n782, n748, n769, n755);
or   g803 (n833, n758, n779, n749, n775);
xnor g804 (n873, n816, n400);
xnor g805 (n862, n404, n835, n428, n414);
nor  g806 (n851, n685, n685, n823, n427);
and  g807 (n855, n424, n833, n421);
xor  g808 (n848, n401, n422, n410, n423);
nand g809 (n857, n410, n683, n828, n418);
nor  g810 (n838, n684, n402, n686, n407);
xnor g811 (n868, n427, n421, n823, n831);
and  g812 (n866, n400, n406, n420, n403);
nand g813 (n842, n818, n415, n422, n408);
and  g814 (n846, n420, n820, n422, n426);
nand g815 (n852, n820, n401, n417, n834);
nor  g816 (n840, n399, n412, n418, n684);
nor  g817 (n860, n414, n416, n817);
nand g818 (n853, n836, n822, n404, n423);
xnor g819 (n856, n419, n399, n428, n827);
nand g820 (n861, n411, n819, n818, n821);
or   g821 (n871, n825, n398, n417, n420);
or   g822 (n847, n414, n426, n835, n824);
xnor g823 (n843, n409, n819, n685, n418);
xor  g824 (n849, n413, n412, n683, n408);
xor  g825 (n869, n406, n424, n425);
or   g826 (n839, n417, n826, n425, n825);
nand g827 (n864, n832, n408, n683, n403);
and  g828 (n867, n426, n398, n830, n419);
and  g829 (n845, n415, n416, n413, n411);
and  g830 (n870, n427, n419, n826, n816);
nor  g831 (n837, n827, n684, n829, n410);
xor  g832 (n863, n404, n409, n424, n834);
nor  g833 (n850, n411, n405, n829, n407);
xor  g834 (n872, n406, n409, n423, n407);
nor  g835 (n844, n831, n399, n415, n402);
xor  g836 (n854, n821, n817, n830, n824);
and  g837 (n858, n828, n428, n833, n405);
xor  g838 (n859, n405, n403, n402, n398);
or   g839 (n865, n412, n413, n400, n401);
nand g840 (n841, n822, n836, n832, n429);
and  g841 (n894, n790, n433, n795, n793);
xnor g842 (n899, n802, n869, n859, n812);
or   g843 (n884, n800, n430, n796, n810);
nand g844 (n901, n795, n849, n845, n815);
nand g845 (n881, n806, n815, n804);
nor  g846 (n882, n811, n686, n793, n864);
and  g847 (n885, n852, n815, n814, n431);
or   g848 (n900, n796, n687, n871, n798);
nor  g849 (n878, n432, n690, n809, n807);
nand g850 (n886, n789, n431, n794, n867);
xnor g851 (n896, n813, n863, n799, n868);
or   g852 (n876, n792, n801, n787, n788);
or   g853 (n892, n431, n789, n794, n791);
xor  g854 (n897, n429, n851, n799, n858);
xor  g855 (n877, n432, n813, n429, n688);
nor  g856 (n888, n686, n687, n800, n432);
or   g857 (n880, n870, n802, n866, n808);
nor  g858 (n874, n814, n862, n801, n689);
or   g859 (n889, n814, n854, n810, n806);
nand g860 (n879, n812, n687, n847, n853);
xor  g861 (n891, n803, n811, n797, n430);
nor  g862 (n898, n788, n813, n787, n846);
xnor g863 (n875, n808, n803, n872, n850);
and  g864 (n895, n873, n855, n809, n688);
nor  g865 (n890, n812, n805, n861, n865);
xor  g866 (n887, n792, n805, n791, n798);
and  g867 (n883, n430, n857, n811, n860);
nor  g868 (n893, n807, n856, n689, n848);
or   g869 (n902, n689, n790, n797, n688);
nor  g870 (n907, n434, n702, n691, n899);
nand g871 (n904, n696, n882, n895, n700);
and  g872 (n916, n888, n876, n896, n900);
and  g873 (n915, n894, n875, n892, n886);
or   g874 (n937, n898, n891, n896, n893);
xor  g875 (n938, n698, n893, n693, n894);
xor  g876 (n914, n896, n695, n887, n155);
or   g877 (n936, n898, n891, n878, n889);
xor  g878 (n934, n884, n696, n435);
xor  g879 (n920, n892, n891, n32, n875);
and  g880 (n906, n691, n895, n719, n704);
nand g881 (n909, n693, n902, n880, n697);
xor  g882 (n940, n900, n880, n897, n888);
xor  g883 (n917, n895, n876, n890, n692);
xnor g884 (n913, n881, n879, n898, n874);
or   g885 (n935, n877, n701, n899, n875);
and  g886 (n933, n901, n882, n879, n435);
xnor g887 (n921, n902, n876, n698, n898);
xnor g888 (n942, n433, n435, n880, n702);
or   g889 (n912, n890, n720, n703, n694);
xor  g890 (n918, n878, n889, n697, n720);
and  g891 (n910, n721, n32, n894, n701);
xor  g892 (n930, n698, n889, n899, n878);
xor  g893 (n926, n883, n693, n884, n720);
xor  g894 (n919, n888, n702, n886, n883);
or   g895 (n908, n881, n704, n874, n691);
nor  g896 (n923, n692, n877, n884, n885);
xor  g897 (n925, n900, n694, n433, n877);
xor  g898 (n932, n897, n695, n700, n887);
or   g899 (n941, n902, n719, n882, n155);
nand g900 (n905, n879, n899, n156, n874);
and  g901 (n911, n900, n703, n901, n885);
xor  g902 (n928, n699, n902, n893, n897);
or   g903 (n924, n700, n434, n890, n692);
and  g904 (n929, n699, n32, n896, n721);
xor  g905 (n931, n434, n901, n697);
xor  g906 (n922, n721, n703, n881, n886);
nor  g907 (n903, n690, n885, n699, n887);
xnor g908 (n939, n897, n892, n694, n883);
nor  g909 (n927, n690, n701, n722, n695);
xor  g910 (n962, n921, n936, n928, n934);
nand g911 (n959, n923, n938, n937, n942);
nor  g912 (n952, n933, n919, n914, n930);
nand g913 (n943, n905, n922, n929, n927);
and  g914 (n960, n941, n926, n905, n939);
nor  g915 (n945, n924, n910, n937);
xor  g916 (n951, n926, n934, n925, n922);
nor  g917 (n967, n941, n908, n932);
nand g918 (n946, n939, n920, n942, n940);
xor  g919 (n958, n923, n935, n924, n939);
or   g920 (n957, n920, n935, n917, n922);
nand g921 (n956, n906, n912, n928, n909);
xor  g922 (n949, n929, n940, n436);
or   g923 (n964, n907, n936, n921, n931);
or   g924 (n969, n916, n935, n934, n156);
nand g925 (n953, n912, n929, n924, n903);
and  g926 (n961, n436, n936, n437, n909);
or   g927 (n944, n941, n916, n906, n921);
nor  g928 (n963, n914, n903, n931, n938);
xor  g929 (n947, n942, n931, n913, n938);
xor  g930 (n968, n911, n940, n933);
xor  g931 (n966, n918, n927, n913, n926);
or   g932 (n948, n919, n932, n911, n915);
or   g933 (n954, n937, n923, n930, n918);
nand g934 (n965, n928, n917, n908, n925);
and  g935 (n955, n904, n927, n907, n437);
or   g936 (n950, n930, n904, n915, n925);
not  g937 (n973, n959);
not  g938 (n972, n960);
buf  g939 (n976, n967);
not  g940 (n975, n966);
buf  g941 (n977, n965);
buf  g942 (n970, n962);
nand g943 (n974, n964, n956);
nand g944 (n971, n961, n963, n958, n957);
not  g945 (n978, n973);
buf  g946 (n981, n976);
not  g947 (n980, n974);
not  g948 (n979, n975);
not  g949 (n988, n980);
buf  g950 (n985, n980);
buf  g951 (n986, n978);
not  g952 (n983, n978);
buf  g953 (n984, n979);
not  g954 (n987, n981);
and  g955 (n982, n981, n979);
buf  g956 (n993, n441);
not  g957 (n990, n987);
not  g958 (n991, n986);
buf  g959 (n989, n438);
not  g960 (n992, n986);
buf  g961 (n1007, n983);
buf  g962 (n996, n437);
buf  g963 (n999, n982);
not  g964 (n1002, n441);
buf  g965 (n1000, n988);
buf  g966 (n1008, n983);
buf  g967 (n997, n984);
not  g968 (n1005, n977);
or   g969 (n1003, n438, n984, n440);
nor  g970 (n998, n442, n439, n984, n982);
nor  g971 (n995, n988, n441, n439, n985);
xnor g972 (n994, n440, n987, n985, n443);
nand g973 (n1004, n987, n442, n985, n988);
xnor g974 (n1001, n440, n986, n443, n438);
xnor g975 (n1006, n442, n983, n439, n443);
xnor g976 (n1015, n1007, n1000, n991, n1008);
nor  g977 (n1016, n1006, n1006, n995, n969);
or   g978 (n1014, n1001, n1003, n1004, n1002);
and  g979 (n1013, n998, n999, n1005, n989);
nor  g980 (n1009, n1008, n981, n994, n990);
or   g981 (n1012, n1004, n968, n1002, n1005);
nand g982 (n1017, n1007, n997, n993, n1003);
and  g983 (n1010, n1001, n998, n999, n1000);
or   g984 (n1011, n997, n156, n992, n996);
buf  g985 (n1019, n1009);
not  g986 (n1018, n1010);
xor  g987 (n1024, n1012, n1018, n1015);
xor  g988 (n1025, n1011, n1014, n1019);
nor  g989 (n1026, n1018, n707, n1010);
xnor g990 (n1021, n706, n722, n1018, n705);
and  g991 (n1020, n706, n722, n1015, n1013);
nor  g992 (n1023, n706, n1011, n1016, n707);
and  g993 (n1022, n704, n1012, n705, n1019);
nor  g994 (n1027, n1013, n1014, n705, n1019);
xor  g995 (n1028, n709, n708, n1017);
nand g996 (n1032, n1024, n444, n1025, n1016);
or   g997 (n1030, n710, n1027, n709, n1017);
xnor g998 (n1031, n1023, n444, n1026);
or   g999 (n1029, n708, n709, n710);
endmodule
