

module Stat_264_47
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n284,
  n273,
  n276,
  n283,
  n279,
  n278,
  n280,
  n274,
  n269,
  n277,
  n282,
  n267,
  n272,
  n285,
  n268,
  n270,
  n271,
  n275,
  n281
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n284;output n273;output n276;output n283;output n279;output n278;output n280;output n274;output n269;output n277;output n282;output n267;output n272;output n285;output n268;output n270;output n271;output n275;output n281;
  wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;

  not
  g0
  (
    n82,
    n9
  );


  not
  g1
  (
    n67,
    n14
  );


  buf
  g2
  (
    n77,
    n8
  );


  buf
  g3
  (
    n39,
    n1
  );


  buf
  g4
  (
    n84,
    n1
  );


  buf
  g5
  (
    n22,
    n13
  );


  not
  g6
  (
    n49,
    n15
  );


  buf
  g7
  (
    n63,
    n15
  );


  buf
  g8
  (
    n25,
    n6
  );


  buf
  g9
  (
    n28,
    n8
  );


  not
  g10
  (
    n57,
    n2
  );


  not
  g11
  (
    n30,
    n2
  );


  not
  g12
  (
    n83,
    n13
  );


  not
  g13
  (
    n42,
    n14
  );


  not
  g14
  (
    n35,
    n2
  );


  buf
  g15
  (
    n80,
    n6
  );


  buf
  g16
  (
    n79,
    n20
  );


  not
  g17
  (
    n47,
    n19
  );


  buf
  g18
  (
    n62,
    n21
  );


  not
  g19
  (
    n46,
    n5
  );


  buf
  g20
  (
    n74,
    n11
  );


  buf
  g21
  (
    n53,
    n9
  );


  not
  g22
  (
    n68,
    n15
  );


  not
  g23
  (
    n52,
    n3
  );


  buf
  g24
  (
    n50,
    n16
  );


  buf
  g25
  (
    n76,
    n10
  );


  buf
  g26
  (
    n44,
    n21
  );


  buf
  g27
  (
    n71,
    n19
  );


  buf
  g28
  (
    n66,
    n20
  );


  buf
  g29
  (
    n60,
    n16
  );


  buf
  g30
  (
    n45,
    n3
  );


  buf
  g31
  (
    n23,
    n21
  );


  buf
  g32
  (
    KeyWire_0_7,
    n1
  );


  buf
  g33
  (
    n38,
    n8
  );


  buf
  g34
  (
    n26,
    n14
  );


  not
  g35
  (
    n70,
    n4
  );


  buf
  g36
  (
    n32,
    n12
  );


  buf
  g37
  (
    n40,
    n17
  );


  not
  g38
  (
    n78,
    n17
  );


  not
  g39
  (
    n48,
    n18
  );


  not
  g40
  (
    n58,
    n12
  );


  buf
  g41
  (
    n37,
    n10
  );


  not
  g42
  (
    KeyWire_0_3,
    n12
  );


  buf
  g43
  (
    n73,
    n7
  );


  buf
  g44
  (
    n56,
    n7
  );


  buf
  g45
  (
    KeyWire_0_10,
    n5
  );


  not
  g46
  (
    n43,
    n16
  );


  buf
  g47
  (
    n69,
    n9
  );


  buf
  g48
  (
    n75,
    n20
  );


  buf
  g49
  (
    n41,
    n4
  );


  buf
  g50
  (
    n36,
    n18
  );


  buf
  g51
  (
    KeyWire_0_9,
    n19
  );


  buf
  g52
  (
    n72,
    n4
  );


  buf
  g53
  (
    n31,
    n18
  );


  buf
  g54
  (
    n59,
    n5
  );


  buf
  g55
  (
    n29,
    n3
  );


  not
  g56
  (
    n81,
    n11
  );


  buf
  g57
  (
    n54,
    n13
  );


  buf
  g58
  (
    n64,
    n17
  );


  buf
  g59
  (
    n65,
    n6
  );


  not
  g60
  (
    n33,
    n10
  );


  buf
  g61
  (
    n34,
    n11
  );


  buf
  g62
  (
    n61,
    n7
  );


  not
  g63
  (
    n162,
    n52
  );


  not
  g64
  (
    KeyWire_0_2,
    n47
  );


  not
  g65
  (
    n186,
    n80
  );


  buf
  g66
  (
    n120,
    n45
  );


  not
  g67
  (
    n135,
    n57
  );


  buf
  g68
  (
    n180,
    n70
  );


  buf
  g69
  (
    n104,
    n75
  );


  buf
  g70
  (
    KeyWire_0_5,
    n45
  );


  not
  g71
  (
    n102,
    n84
  );


  buf
  g72
  (
    n95,
    n67
  );


  buf
  g73
  (
    n114,
    n59
  );


  not
  g74
  (
    n127,
    n75
  );


  not
  g75
  (
    n154,
    n56
  );


  not
  g76
  (
    n134,
    n55
  );


  buf
  g77
  (
    n116,
    n66
  );


  not
  g78
  (
    n160,
    n59
  );


  not
  g79
  (
    n129,
    n70
  );


  not
  g80
  (
    n163,
    n60
  );


  not
  g81
  (
    n103,
    n69
  );


  buf
  g82
  (
    n158,
    n26
  );


  buf
  g83
  (
    n117,
    n67
  );


  not
  g84
  (
    n108,
    n69
  );


  buf
  g85
  (
    n132,
    n61
  );


  buf
  g86
  (
    n145,
    n39
  );


  not
  g87
  (
    n98,
    n28
  );


  not
  g88
  (
    n170,
    n42
  );


  not
  g89
  (
    n110,
    n51
  );


  buf
  g90
  (
    n131,
    n58
  );


  buf
  g91
  (
    n126,
    n66
  );


  not
  g92
  (
    n92,
    n40
  );


  not
  g93
  (
    n152,
    n65
  );


  not
  g94
  (
    n143,
    n43
  );


  buf
  g95
  (
    n93,
    n34
  );


  buf
  g96
  (
    n155,
    n29
  );


  not
  g97
  (
    n109,
    n43
  );


  not
  g98
  (
    n164,
    n28
  );


  buf
  g99
  (
    n87,
    n38
  );


  buf
  g100
  (
    n138,
    n53
  );


  buf
  g101
  (
    n130,
    n62
  );


  buf
  g102
  (
    n88,
    n67
  );


  buf
  g103
  (
    n153,
    n52
  );


  buf
  g104
  (
    n146,
    n68
  );


  not
  g105
  (
    n176,
    n31
  );


  buf
  g106
  (
    n141,
    n22
  );


  buf
  g107
  (
    KeyWire_0_14,
    n42
  );


  not
  g108
  (
    n125,
    n42
  );


  buf
  g109
  (
    n140,
    n43
  );


  buf
  g110
  (
    n128,
    n35
  );


  not
  g111
  (
    n169,
    n82
  );


  buf
  g112
  (
    n156,
    n36
  );


  not
  g113
  (
    n151,
    n25
  );


  buf
  g114
  (
    n171,
    n32
  );


  not
  g115
  (
    n119,
    n37
  );


  not
  g116
  (
    n178,
    n46
  );


  not
  g117
  (
    n86,
    n44
  );


  not
  g118
  (
    n121,
    n49
  );


  buf
  g119
  (
    n113,
    n29
  );


  buf
  g120
  (
    n188,
    n58
  );


  buf
  g121
  (
    n94,
    n50
  );


  buf
  g122
  (
    KeyWire_0_0,
    n74
  );


  buf
  g123
  (
    n115,
    n84
  );


  not
  g124
  (
    n147,
    n26
  );


  buf
  g125
  (
    n184,
    n53
  );


  buf
  g126
  (
    n107,
    n50
  );


  buf
  g127
  (
    n183,
    n61
  );


  buf
  g128
  (
    n142,
    n30
  );


  buf
  g129
  (
    KeyWire_0_12,
    n31
  );


  buf
  g130
  (
    n90,
    n23
  );


  not
  g131
  (
    n179,
    n46
  );


  not
  g132
  (
    n136,
    n70
  );


  not
  g133
  (
    n100,
    n29
  );


  buf
  g134
  (
    n175,
    n28
  );


  buf
  g135
  (
    n157,
    n45
  );


  not
  g136
  (
    n111,
    n23
  );


  buf
  g137
  (
    KeyWire_0_15,
    n37
  );


  buf
  g138
  (
    n91,
    n64
  );


  buf
  g139
  (
    n123,
    n77
  );


  not
  g140
  (
    KeyWire_0_11,
    n78
  );


  xnor
  g141
  (
    n124,
    n49,
    n33,
    n48
  );


  nand
  g142
  (
    n137,
    n50,
    n30,
    n71,
    n64
  );


  xnor
  g143
  (
    n101,
    n57,
    n53,
    n79,
    n56
  );


  xor
  g144
  (
    n177,
    n25,
    n54,
    n77,
    n73
  );


  xor
  g145
  (
    n167,
    n55,
    n73,
    n48,
    n54
  );


  or
  g146
  (
    n187,
    n30,
    n55,
    n46,
    n41
  );


  xor
  g147
  (
    n181,
    n25,
    n72,
    n51,
    n54
  );


  nand
  g148
  (
    n174,
    n63,
    n57,
    n79,
    n65
  );


  or
  g149
  (
    n96,
    n59,
    n80,
    n47,
    n68
  );


  nand
  g150
  (
    n122,
    n72,
    n68,
    n35,
    n33
  );


  nor
  g151
  (
    n148,
    n63,
    n41,
    n82,
    n80
  );


  xnor
  g152
  (
    n97,
    n47,
    n23,
    n76,
    n36
  );


  and
  g153
  (
    n172,
    n32,
    n84,
    n82,
    n44
  );


  xnor
  g154
  (
    n105,
    n71,
    n81,
    n69,
    n76
  );


  or
  g155
  (
    n85,
    n65,
    n34,
    n60,
    n37
  );


  nor
  g156
  (
    n149,
    n77,
    n39,
    n72,
    n83
  );


  nand
  g157
  (
    n159,
    n61,
    n48,
    n24
  );


  and
  g158
  (
    n99,
    n27,
    n40,
    n36,
    n35
  );


  xor
  g159
  (
    n182,
    n75,
    n26,
    n64,
    n63
  );


  xor
  g160
  (
    n189,
    n58,
    n78,
    n79,
    n24
  );


  nor
  g161
  (
    n173,
    n27,
    n52,
    n38,
    n76
  );


  xor
  g162
  (
    n106,
    n73,
    n32,
    n22,
    n51
  );


  nand
  g163
  (
    n144,
    n71,
    n83,
    n81,
    n49
  );


  nand
  g164
  (
    n150,
    n40,
    n38,
    n81,
    n62
  );


  nand
  g165
  (
    n190,
    n44,
    n56,
    n83,
    n31
  );


  nand
  g166
  (
    n118,
    n41,
    n74,
    n34
  );


  xor
  g167
  (
    n165,
    n33,
    n27,
    n39,
    n62
  );


  nor
  g168
  (
    n166,
    n60,
    n78,
    n22,
    n66
  );


  xor
  g169
  (
    n240,
    n106,
    n153,
    n177,
    n98
  );


  nand
  g170
  (
    n264,
    n150,
    n171,
    n185,
    n89
  );


  and
  g171
  (
    n202,
    n174,
    n159,
    n97,
    n152
  );


  and
  g172
  (
    n199,
    n139,
    n102,
    n161,
    n113
  );


  nor
  g173
  (
    n213,
    n94,
    n123,
    n95,
    n183
  );


  xor
  g174
  (
    n206,
    n158,
    n175,
    n102,
    n131
  );


  xor
  g175
  (
    n248,
    n136,
    n179,
    n127,
    n155
  );


  nand
  g176
  (
    n218,
    n128,
    n130,
    n96,
    n145
  );


  xnor
  g177
  (
    KeyWire_0_13,
    n145,
    n175,
    n172,
    n115
  );


  nand
  g178
  (
    n216,
    n104,
    n138,
    n175,
    n153
  );


  or
  g179
  (
    n196,
    n165,
    n132,
    n156,
    n102
  );


  nor
  g180
  (
    n200,
    n137,
    n97,
    n126,
    n143
  );


  nor
  g181
  (
    n219,
    n100,
    n148,
    n184,
    n132
  );


  or
  g182
  (
    n256,
    n172,
    n128,
    n150,
    n158
  );


  or
  g183
  (
    n229,
    n176,
    n180,
    n172,
    n160
  );


  or
  g184
  (
    n228,
    n133,
    n155,
    n106,
    n91
  );


  xnor
  g185
  (
    n192,
    n131,
    n177,
    n140,
    n134
  );


  or
  g186
  (
    n251,
    n125,
    n105,
    n142,
    n99
  );


  xor
  g187
  (
    n223,
    n165,
    n132,
    n113,
    n111
  );


  xnor
  g188
  (
    n211,
    n182,
    n93,
    n147,
    n164
  );


  nor
  g189
  (
    n266,
    n112,
    n159,
    n183,
    n95
  );


  xor
  g190
  (
    n241,
    n185,
    n188,
    n140,
    n162
  );


  or
  g191
  (
    n225,
    n125,
    n152,
    n178,
    n163
  );


  xnor
  g192
  (
    n226,
    n166,
    n155,
    n99,
    n128
  );


  xnor
  g193
  (
    n221,
    n96,
    n109,
    n147,
    n164
  );


  xor
  g194
  (
    n209,
    n157,
    n186,
    n159,
    n165
  );


  or
  g195
  (
    n210,
    n118,
    n123,
    n110,
    n127
  );


  xor
  g196
  (
    n194,
    n148,
    n119,
    n97,
    n95
  );


  nand
  g197
  (
    n197,
    n157,
    n103,
    n143,
    n116
  );


  xor
  g198
  (
    n232,
    n129,
    n138,
    n161,
    n122
  );


  nor
  g199
  (
    n246,
    n168,
    n108,
    n107,
    n135
  );


  xor
  g200
  (
    n201,
    n170,
    n92,
    n178,
    n119
  );


  xor
  g201
  (
    n208,
    n184,
    n142,
    n105,
    n176
  );


  nor
  g202
  (
    n205,
    n163,
    n189,
    n139,
    n88
  );


  nor
  g203
  (
    n257,
    n148,
    n109,
    n184,
    n181
  );


  and
  g204
  (
    n261,
    n118,
    n100,
    n166,
    n160
  );


  nor
  g205
  (
    n231,
    n124,
    n173,
    n158,
    n114
  );


  nor
  g206
  (
    n224,
    n125,
    n112,
    n136,
    n151
  );


  xor
  g207
  (
    n245,
    n94,
    n188,
    n186,
    n129
  );


  xnor
  g208
  (
    n265,
    n168,
    n161,
    n163,
    n120
  );


  and
  g209
  (
    n191,
    n117,
    n188,
    n171,
    n115
  );


  and
  g210
  (
    n203,
    n90,
    n112,
    n149,
    n182
  );


  and
  g211
  (
    n249,
    n104,
    n180,
    n116
  );


  or
  g212
  (
    n243,
    n135,
    n119,
    n129,
    n107
  );


  nand
  g213
  (
    n207,
    n169,
    n187,
    n133,
    n92
  );


  xnor
  g214
  (
    n242,
    n176,
    n173,
    n134,
    n167
  );


  and
  g215
  (
    n259,
    n141,
    n99,
    n121,
    n144
  );


  xor
  g216
  (
    n212,
    n145,
    n177,
    n136,
    n117
  );


  xor
  g217
  (
    n238,
    n115,
    n183,
    n166,
    n146
  );


  nor
  g218
  (
    n233,
    n189,
    n168,
    n152,
    n96
  );


  xnor
  g219
  (
    n262,
    n154,
    n179,
    n100,
    n126
  );


  and
  g220
  (
    n230,
    n123,
    n120,
    n85,
    n151
  );


  or
  g221
  (
    n254,
    n178,
    n156,
    n174,
    n140
  );


  nor
  g222
  (
    n222,
    n117,
    n146,
    n101,
    n133
  );


  or
  g223
  (
    n234,
    n106,
    n171,
    n131,
    n130
  );


  and
  g224
  (
    n227,
    n149,
    n137,
    n101,
    n174
  );


  nand
  g225
  (
    n198,
    n164,
    n181,
    n154,
    n130
  );


  xor
  g226
  (
    n247,
    n105,
    n141,
    n101
  );


  nand
  g227
  (
    n255,
    n104,
    n114,
    n162,
    n173
  );


  nor
  g228
  (
    n215,
    n118,
    n147,
    n162,
    n146
  );


  and
  g229
  (
    KeyWire_0_8,
    n93,
    n137,
    n189,
    n124
  );


  and
  g230
  (
    n195,
    n124,
    n187,
    n122
  );


  xor
  g231
  (
    n220,
    n135,
    n126,
    n157,
    n108
  );


  and
  g232
  (
    n250,
    n190,
    n169,
    n103,
    n151
  );


  and
  g233
  (
    n204,
    n139,
    n87,
    n98,
    n153
  );


  xor
  g234
  (
    n237,
    n170,
    n109,
    n142,
    n120
  );


  and
  g235
  (
    n193,
    n182,
    n149,
    n156,
    n113
  );


  and
  g236
  (
    n244,
    n181,
    n179,
    n121,
    n122
  );


  nand
  g237
  (
    n235,
    n110,
    n190,
    n154,
    n103
  );


  xor
  g238
  (
    n260,
    n167,
    n116,
    n150,
    n107
  );


  xor
  g239
  (
    n236,
    n111,
    n143,
    n94,
    n93
  );


  nor
  g240
  (
    n252,
    n167,
    n92,
    n190,
    n108
  );


  and
  g241
  (
    n263,
    n138,
    n160,
    n169,
    n110
  );


  xnor
  g242
  (
    n258,
    n144,
    n114,
    n98,
    n185
  );


  xnor
  g243
  (
    n214,
    n170,
    n186,
    n134,
    n111
  );


  nand
  g244
  (
    n253,
    n127,
    n144,
    n86,
    n121
  );


  or
  g245
  (
    n283,
    n211,
    n203,
    n231,
    n239
  );


  xnor
  g246
  (
    n267,
    n229,
    n226,
    n254,
    n222
  );


  nor
  g247
  (
    KeyWire_0_4,
    n206,
    n202,
    n197,
    n241
  );


  or
  g248
  (
    n281,
    n260,
    n198,
    n262,
    n194
  );


  xnor
  g249
  (
    n279,
    n244,
    n227,
    n196,
    n234
  );


  xor
  g250
  (
    n269,
    n216,
    n192,
    n232,
    n263
  );


  nor
  g251
  (
    n284,
    n240,
    n251,
    n228,
    n224
  );


  or
  g252
  (
    n282,
    n265,
    n246,
    n252,
    n249
  );


  and
  g253
  (
    n276,
    n210,
    n212,
    n214,
    n218
  );


  nor
  g254
  (
    n278,
    n253,
    n243,
    n248,
    n238
  );


  or
  g255
  (
    n272,
    n201,
    n264,
    n208,
    n209
  );


  and
  g256
  (
    KeyWire_0_1,
    n225,
    n199,
    n191,
    n205
  );


  xor
  g257
  (
    n280,
    n217,
    n250,
    n235,
    n242
  );


  or
  g258
  (
    n268,
    n261,
    n213,
    n219,
    n256
  );


  nor
  g259
  (
    n273,
    n233,
    n247,
    n257,
    n266
  );


  nor
  g260
  (
    n274,
    n236,
    n215,
    n259,
    n207
  );


  xor
  g261
  (
    n271,
    n223,
    n245,
    n200,
    n195
  );


  xnor
  g262
  (
    KeyWire_0_6,
    n220,
    n255,
    n258,
    n221
  );


  nor
  g263
  (
    n275,
    n204,
    n230,
    n193,
    n237
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n89,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n277,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n133,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n55,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n270,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n161,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n285,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n27,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n239,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n24,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n51,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n112,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n139,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n217,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n185,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n168,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


