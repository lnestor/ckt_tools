// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_175_832 written by SynthGen on 2021/05/24 19:46:51
module Stat_175_832( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21,
 n99, n113, n104, n108, n121, n116, n115, n109,
 n111, n107, n103, n120, n118, n185, n178, n188,
 n189, n192, n196, n186, n194, n193, n195, n187,
 n182, n179, n183, n181, n180, n190, n191, n184);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21;

output n99, n113, n104, n108, n121, n116, n115, n109,
 n111, n107, n103, n120, n118, n185, n178, n188,
 n189, n192, n196, n186, n194, n193, n195, n187,
 n182, n179, n183, n181, n180, n190, n191, n184;

wire n22, n23, n24, n25, n26, n27, n28, n29,
 n30, n31, n32, n33, n34, n35, n36, n37,
 n38, n39, n40, n41, n42, n43, n44, n45,
 n46, n47, n48, n49, n50, n51, n52, n53,
 n54, n55, n56, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n67, n68, n69,
 n70, n71, n72, n73, n74, n75, n76, n77,
 n78, n79, n80, n81, n82, n83, n84, n85,
 n86, n87, n88, n89, n90, n91, n92, n93,
 n94, n95, n96, n97, n98, n100, n101, n102,
 n105, n106, n110, n112, n114, n117, n119, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177;

buf  g0 (n47, n1);
buf  g1 (n34, n2);
not  g2 (n40, n2);
buf  g3 (n26, n3);
buf  g4 (n43, n3);
buf  g5 (n46, n1);
not  g6 (n32, n7);
buf  g7 (n35, n7);
not  g8 (n28, n5);
not  g9 (n42, n7);
buf  g10 (n50, n1);
buf  g11 (n45, n8);
buf  g12 (n25, n1);
buf  g13 (n23, n4);
buf  g14 (n30, n4);
buf  g15 (n38, n6);
buf  g16 (n44, n3);
buf  g17 (n27, n6);
buf  g18 (n36, n3);
buf  g19 (n41, n2);
not  g20 (n48, n4);
not  g21 (n37, n2);
not  g22 (n33, n5);
buf  g23 (n49, n5);
not  g24 (n51, n5);
buf  g25 (n31, n6);
not  g26 (n22, n4);
buf  g27 (n39, n7);
not  g28 (n29, n8);
not  g29 (n24, n6);
buf  g30 (n71, n24);
not  g31 (n57, n22);
nor  g32 (n55, n44, n42, n24, n45);
xnor g33 (n74, n34, n38, n37, n43);
and  g34 (n65, n46, n23, n39, n45);
and  g35 (n53, n24, n26, n22, n25);
nand g36 (n63, n30, n36, n46, n35);
nor  g37 (n76, n23, n41, n43, n25);
nand g38 (n75, n31, n23, n38, n29);
nand g39 (n68, n47, n25, n22, n27);
xnor g40 (n56, n32, n33, n44, n36);
or   g41 (n77, n26, n43, n35);
and  g42 (n72, n48, n28, n24, n39);
nor  g43 (n58, n39, n40, n47, n42);
nand g44 (n79, n30, n37, n42, n41);
and  g45 (n78, n45, n33, n38, n29);
xor  g46 (n52, n30, n26, n40, n36);
xnor g47 (n64, n48, n31, n36, n30);
or   g48 (n59, n38, n43, n41, n46);
xor  g49 (n54, n39, n31, n28, n22);
nand g50 (n61, n34, n27, n47, n23);
xnor g51 (n67, n47, n32, n33, n41);
nand g52 (n73, n44, n46, n28, n45);
xor  g53 (n70, n34, n44, n29, n37);
xor  g54 (n69, n31, n33, n27);
and  g55 (n60, n29, n34, n40, n32);
and  g56 (n66, n32, n28, n25, n37);
or   g57 (n62, n40, n26, n42, n35);
not  g58 (n84, n69);
buf  g59 (n99, n65);
not  g60 (n80, n52);
buf  g61 (n101, n67);
not  g62 (n90, n66);
not  g63 (n91, n64);
buf  g64 (n92, n59);
buf  g65 (n83, n68);
buf  g66 (n93, n60);
not  g67 (n85, n63);
not  g68 (n81, n69);
not  g69 (n86, n55);
not  g70 (n87, n67);
buf  g71 (n89, n56);
buf  g72 (n96, n62);
not  g73 (n95, n61);
buf  g74 (n97, n57);
buf  g75 (n98, n70);
buf  g76 (n100, n54);
not  g77 (n82, n53);
not  g78 (n88, n68);
buf  g79 (n94, n58);
not  g80 (n109, n49);
buf  g81 (n104, n49);
not  g82 (n121, n90);
not  g83 (n102, n96);
buf  g84 (n105, n89);
buf  g85 (n111, n101);
buf  g86 (n112, n100);
buf  g87 (n116, n48);
buf  g88 (n113, n92);
buf  g89 (n114, n99);
not  g90 (n115, n95);
not  g91 (n106, n50);
not  g92 (n110, n48);
buf  g93 (n119, n82);
not  g94 (n118, n85);
not  g95 (n120, n81);
not  g96 (n108, n98);
not  g97 (n122, n97);
xor  g98 (n103, n84, n49);
xor  g99 (n107, n83, n91, n93, n87);
and  g100 (n117, n94, n49, n86, n88);
not  g101 (n138, n70);
buf  g102 (n140, n8);
buf  g103 (n139, n102);
not  g104 (n135, n79);
buf  g105 (n123, n78);
not  g106 (n132, n106);
buf  g107 (n128, n118);
buf  g108 (n131, n76);
nor  g109 (n126, n78, n109, n77, n72);
or   g110 (n125, n10, n71, n107);
or   g111 (n127, n104, n112, n8, n10);
nor  g112 (n142, n120, n9);
nand g113 (n134, n73, n117, n75, n10);
xor  g114 (n130, n113, n78, n116, n77);
and  g115 (n133, n9, n76, n103, n115);
and  g116 (n141, n76, n76, n79, n111);
or   g117 (n129, n114, n79, n74, n121);
nor  g118 (n136, n77, n108, n78, n79);
and  g119 (n137, n73, n74, n72, n105);
and  g120 (n124, n75, n119, n77, n110);
buf  g121 (n144, n51);
nand g122 (n151, n50, n51, n140);
nor  g123 (n149, n136, n132, n135, n131);
and  g124 (n157, n140, n137, n130, n136);
xnor g125 (n148, n133, n51, n134, n138);
or   g126 (n153, n131, n132, n137, n130);
xnor g127 (n154, n131, n129, n51);
xnor g128 (n156, n50, n134, n139, n135);
xor  g129 (n145, n141, n137, n139, n127);
xor  g130 (n159, n134, n130, n138, n125);
or   g131 (n143, n137, n129, n139, n132);
xor  g132 (n152, n134, n133, n131);
nor  g133 (n146, n130, n123, n136, n141);
or   g134 (n155, n132, n124, n138, n141);
nand g135 (n147, n128, n135, n126);
or   g136 (n150, n136, n50, n141, n129);
xnor g137 (n158, n133, n140, n139, n138);
buf  g138 (n161, n157);
nor  g139 (n164, n151, n159, n21);
xnor g140 (n176, n18, n15, n17);
nand g141 (n173, n11, n150, n20);
xor  g142 (n177, n149, n143, n158, n148);
nor  g143 (n166, n155, n156, n157, n19);
nor  g144 (n165, n13, n11, n19, n155);
xor  g145 (n167, n14, n13, n21, n147);
xor  g146 (n170, n11, n12, n145);
or   g147 (n171, n14, n13, n20, n15);
xnor g148 (n174, n153, n19, n15, n16);
xnor g149 (n160, n159, n14, n18, n156);
nor  g150 (n169, n12, n16, n152, n21);
or   g151 (n172, n15, n158, n16, n12);
nand g152 (n175, n11, n19, n17, n13);
nand g153 (n163, n146, n16, n17, n21);
xor  g154 (n162, n10, n18, n122);
xnor g155 (n168, n144, n14, n20, n154);
nor  g156 (n180, n162, n167, n165, n170);
xor  g157 (n187, n177, n166, n163, n169);
or   g158 (n193, n169, n173, n174, n176);
and  g159 (n183, n162, n172, n164, n142);
xnor g160 (n186, n164, n167, n171, n174);
nor  g161 (n191, n162, n166, n175);
xor  g162 (n181, n176, n165, n177, n171);
nand g163 (n192, n163, n160, n167);
xor  g164 (n189, n175, n176, n171, n160);
nor  g165 (n195, n170, n165, n172, n142);
nor  g166 (n178, n174, n142, n170, n172);
nand g167 (n188, n171, n165, n168, n161);
xnor g168 (n196, n173, n160, n172, n175);
xnor g169 (n185, n168, n170, n169, n174);
or   g170 (n179, n173, n164, n168);
nand g171 (n182, n175, n177, n161, n167);
nand g172 (n194, n168, n162, n163, n173);
xor  g173 (n184, n161, n161, n166, n169);
nand g174 (n190, n177, n163, n176, n142);
endmodule
