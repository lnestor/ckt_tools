

module Stat_550_820
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n554,
  n557,
  n569,
  n572,
  n560,
  n555,
  n556,
  n553,
  n567,
  n574,
  n566,
  n559,
  n563,
  n568,
  n561,
  n573,
  n571,
  n565,
  n552,
  n558,
  n575,
  n570,
  n564,
  n562
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n554;output n557;output n569;output n572;output n560;output n555;output n556;output n553;output n567;output n574;output n566;output n559;output n563;output n568;output n561;output n573;output n571;output n565;output n552;output n558;output n575;output n570;output n564;output n562;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n31,
    n22
  );


  not
  g1
  (
    n33,
    n20
  );


  buf
  g2
  (
    n115,
    n3
  );


  not
  g3
  (
    KeyWire_0_17,
    n11
  );


  not
  g4
  (
    n118,
    n12
  );


  buf
  g5
  (
    n29,
    n11
  );


  buf
  g6
  (
    KeyWire_0_10,
    n13
  );


  not
  g7
  (
    n50,
    n24
  );


  buf
  g8
  (
    n123,
    n7
  );


  not
  g9
  (
    n97,
    n19
  );


  buf
  g10
  (
    n70,
    n4
  );


  buf
  g11
  (
    n42,
    n5
  );


  buf
  g12
  (
    n47,
    n5
  );


  not
  g13
  (
    n39,
    n1
  );


  buf
  g14
  (
    KeyWire_0_19,
    n14
  );


  buf
  g15
  (
    n99,
    n24
  );


  not
  g16
  (
    n85,
    n25
  );


  not
  g17
  (
    n56,
    n25
  );


  not
  g18
  (
    n65,
    n25
  );


  buf
  g19
  (
    n111,
    n16
  );


  buf
  g20
  (
    n83,
    n14
  );


  buf
  g21
  (
    n32,
    n2
  );


  not
  g22
  (
    n66,
    n4
  );


  not
  g23
  (
    n48,
    n23
  );


  buf
  g24
  (
    n101,
    n5
  );


  not
  g25
  (
    n38,
    n6
  );


  buf
  g26
  (
    n51,
    n1
  );


  buf
  g27
  (
    n116,
    n24
  );


  buf
  g28
  (
    n79,
    n6
  );


  buf
  g29
  (
    n58,
    n10
  );


  buf
  g30
  (
    n63,
    n18
  );


  buf
  g31
  (
    n84,
    n9
  );


  buf
  g32
  (
    n52,
    n11
  );


  buf
  g33
  (
    n34,
    n23
  );


  buf
  g34
  (
    KeyWire_0_6,
    n14
  );


  not
  g35
  (
    n80,
    n2
  );


  buf
  g36
  (
    n60,
    n21
  );


  not
  g37
  (
    n114,
    n8
  );


  buf
  g38
  (
    n110,
    n13
  );


  not
  g39
  (
    n37,
    n12
  );


  not
  g40
  (
    n92,
    n13
  );


  not
  g41
  (
    n105,
    n11
  );


  not
  g42
  (
    KeyWire_0_2,
    n7
  );


  buf
  g43
  (
    n76,
    n12
  );


  not
  g44
  (
    n108,
    n23
  );


  buf
  g45
  (
    n124,
    n14
  );


  not
  g46
  (
    n43,
    n22
  );


  buf
  g47
  (
    KeyWire_0_24,
    n20
  );


  not
  g48
  (
    n96,
    n15
  );


  not
  g49
  (
    n71,
    n16
  );


  buf
  g50
  (
    n73,
    n15
  );


  not
  g51
  (
    n59,
    n25
  );


  not
  g52
  (
    n55,
    n18
  );


  buf
  g53
  (
    n119,
    n18
  );


  not
  g54
  (
    n95,
    n21
  );


  not
  g55
  (
    n104,
    n24
  );


  buf
  g56
  (
    n69,
    n9
  );


  not
  g57
  (
    n68,
    n15
  );


  buf
  g58
  (
    n26,
    n17
  );


  not
  g59
  (
    n117,
    n20
  );


  not
  g60
  (
    n44,
    n3
  );


  buf
  g61
  (
    n40,
    n8
  );


  not
  g62
  (
    n94,
    n10
  );


  buf
  g63
  (
    n75,
    n19
  );


  not
  g64
  (
    n45,
    n10
  );


  not
  g65
  (
    n67,
    n2
  );


  buf
  g66
  (
    n113,
    n23
  );


  buf
  g67
  (
    n109,
    n16
  );


  not
  g68
  (
    n74,
    n6
  );


  not
  g69
  (
    n122,
    n3
  );


  not
  g70
  (
    n100,
    n12
  );


  not
  g71
  (
    n120,
    n18
  );


  not
  g72
  (
    n64,
    n16
  );


  buf
  g73
  (
    n91,
    n2
  );


  buf
  g74
  (
    n78,
    n13
  );


  not
  g75
  (
    n35,
    n19
  );


  buf
  g76
  (
    n88,
    n4
  );


  buf
  g77
  (
    n106,
    n20
  );


  buf
  g78
  (
    n53,
    n17
  );


  buf
  g79
  (
    n125,
    n1
  );


  buf
  g80
  (
    n86,
    n3
  );


  buf
  g81
  (
    n28,
    n8
  );


  buf
  g82
  (
    n82,
    n17
  );


  buf
  g83
  (
    n62,
    n8
  );


  not
  g84
  (
    n72,
    n22
  );


  not
  g85
  (
    n77,
    n5
  );


  not
  g86
  (
    n98,
    n9
  );


  buf
  g87
  (
    n49,
    n9
  );


  buf
  g88
  (
    n107,
    n10
  );


  not
  g89
  (
    n90,
    n21
  );


  not
  g90
  (
    n46,
    n19
  );


  not
  g91
  (
    n87,
    n17
  );


  not
  g92
  (
    n81,
    n6
  );


  not
  g93
  (
    n89,
    n7
  );


  buf
  g94
  (
    n112,
    n22
  );


  not
  g95
  (
    n61,
    n1
  );


  buf
  g96
  (
    n54,
    n15
  );


  not
  g97
  (
    n93,
    n7
  );


  not
  g98
  (
    n121,
    n21
  );


  buf
  g99
  (
    n57,
    n4
  );


  buf
  g100
  (
    n174,
    n27
  );


  not
  g101
  (
    n141,
    n28
  );


  buf
  g102
  (
    n137,
    n27
  );


  not
  g103
  (
    n151,
    n32
  );


  not
  g104
  (
    n145,
    n34
  );


  buf
  g105
  (
    n157,
    n31
  );


  buf
  g106
  (
    n165,
    n36
  );


  buf
  g107
  (
    n133,
    n27
  );


  buf
  g108
  (
    n131,
    n37
  );


  buf
  g109
  (
    n146,
    n28
  );


  not
  g110
  (
    n152,
    n35
  );


  not
  g111
  (
    n155,
    n33
  );


  not
  g112
  (
    n135,
    n26
  );


  not
  g113
  (
    n144,
    n34
  );


  buf
  g114
  (
    n168,
    n31
  );


  not
  g115
  (
    n147,
    n29
  );


  buf
  g116
  (
    KeyWire_0_5,
    n33
  );


  not
  g117
  (
    n156,
    n35
  );


  not
  g118
  (
    n158,
    n34
  );


  buf
  g119
  (
    n153,
    n26
  );


  not
  g120
  (
    n126,
    n32
  );


  buf
  g121
  (
    n128,
    n26
  );


  not
  g122
  (
    n172,
    n36
  );


  not
  g123
  (
    n142,
    n28
  );


  buf
  g124
  (
    n150,
    n37
  );


  buf
  g125
  (
    n130,
    n26
  );


  buf
  g126
  (
    n163,
    n36
  );


  not
  g127
  (
    n161,
    n33
  );


  buf
  g128
  (
    n162,
    n31
  );


  not
  g129
  (
    n166,
    n32
  );


  not
  g130
  (
    n148,
    n29
  );


  buf
  g131
  (
    n149,
    n29
  );


  buf
  g132
  (
    n164,
    n32
  );


  buf
  g133
  (
    n136,
    n29
  );


  buf
  g134
  (
    n143,
    n34
  );


  not
  g135
  (
    n169,
    n38
  );


  not
  g136
  (
    n134,
    n35
  );


  buf
  g137
  (
    n159,
    n31
  );


  not
  g138
  (
    n132,
    n30
  );


  not
  g139
  (
    KeyWire_0_12,
    n30
  );


  not
  g140
  (
    n170,
    n30
  );


  buf
  g141
  (
    n171,
    n28
  );


  buf
  g142
  (
    n173,
    n37
  );


  buf
  g143
  (
    n140,
    n36
  );


  buf
  g144
  (
    n139,
    n30
  );


  buf
  g145
  (
    n138,
    n27
  );


  buf
  g146
  (
    KeyWire_0_28,
    n37
  );


  buf
  g147
  (
    KeyWire_0_0,
    n35
  );


  not
  g148
  (
    n129,
    n33
  );


  buf
  g149
  (
    KeyWire_0_29,
    n142
  );


  not
  g150
  (
    n195,
    n146
  );


  not
  g151
  (
    n192,
    n147
  );


  not
  g152
  (
    n183,
    n127
  );


  not
  g153
  (
    n200,
    n153
  );


  not
  g154
  (
    n185,
    n128
  );


  not
  g155
  (
    n198,
    n149
  );


  buf
  g156
  (
    n199,
    n126
  );


  not
  g157
  (
    n177,
    n140
  );


  buf
  g158
  (
    n193,
    n132
  );


  buf
  g159
  (
    n190,
    n135
  );


  buf
  g160
  (
    n196,
    n141
  );


  not
  g161
  (
    n184,
    n145
  );


  not
  g162
  (
    n189,
    n134
  );


  not
  g163
  (
    n202,
    n133
  );


  not
  g164
  (
    n176,
    n150
  );


  buf
  g165
  (
    n178,
    n131
  );


  not
  g166
  (
    n186,
    n148
  );


  buf
  g167
  (
    n175,
    n139
  );


  not
  g168
  (
    KeyWire_0_23,
    n151
  );


  buf
  g169
  (
    n201,
    n136
  );


  buf
  g170
  (
    n179,
    n143
  );


  not
  g171
  (
    n197,
    n138
  );


  buf
  g172
  (
    n194,
    n137
  );


  not
  g173
  (
    n182,
    n130
  );


  not
  g174
  (
    n181,
    n152
  );


  not
  g175
  (
    n187,
    n129
  );


  buf
  g176
  (
    n191,
    n144
  );


  nor
  g177
  (
    n277,
    n114,
    n103,
    n94,
    n72
  );


  or
  g178
  (
    n276,
    n56,
    n66,
    n46,
    n48
  );


  xor
  g179
  (
    n263,
    n82,
    n107,
    n38,
    n178
  );


  xnor
  g180
  (
    n280,
    n42,
    n91,
    n184,
    n77
  );


  nor
  g181
  (
    n292,
    n57,
    n71,
    n64,
    n186
  );


  xnor
  g182
  (
    n211,
    n187,
    n53,
    n93,
    n196
  );


  or
  g183
  (
    n271,
    n90,
    n115,
    n102,
    n103
  );


  nor
  g184
  (
    n297,
    n69,
    n192,
    n97,
    n195
  );


  nor
  g185
  (
    n286,
    n187,
    n52,
    n41,
    n43
  );


  nor
  g186
  (
    n220,
    n95,
    n198,
    n103,
    n81
  );


  xnor
  g187
  (
    n256,
    n191,
    n72,
    n64,
    n86
  );


  nor
  g188
  (
    n212,
    n111,
    n44,
    n184,
    n114
  );


  xor
  g189
  (
    n281,
    n201,
    n60,
    n197,
    n75
  );


  and
  g190
  (
    n275,
    n77,
    n189,
    n64,
    n181
  );


  and
  g191
  (
    n229,
    n63,
    n80,
    n115,
    n65
  );


  and
  g192
  (
    n226,
    n76,
    n179,
    n199,
    n202
  );


  or
  g193
  (
    n261,
    n73,
    n81,
    n87,
    n93
  );


  xnor
  g194
  (
    n301,
    n178,
    n67,
    n90,
    n45
  );


  nand
  g195
  (
    n305,
    n62,
    n188,
    n113,
    n50
  );


  nand
  g196
  (
    n241,
    n187,
    n180,
    n109,
    n44
  );


  nor
  g197
  (
    n223,
    n58,
    n188,
    n83,
    n49
  );


  nor
  g198
  (
    n264,
    n182,
    n180,
    n54,
    n51
  );


  or
  g199
  (
    n296,
    n54,
    n87,
    n110,
    n114
  );


  nor
  g200
  (
    n295,
    n194,
    n115,
    n82
  );


  nor
  g201
  (
    n266,
    n194,
    n100,
    n117,
    n53
  );


  and
  g202
  (
    n274,
    n112,
    n189,
    n71,
    n183
  );


  or
  g203
  (
    n251,
    n42,
    n53,
    n185,
    n57
  );


  xor
  g204
  (
    n268,
    n77,
    n102,
    n52,
    n117
  );


  nand
  g205
  (
    n273,
    n96,
    n75,
    n175,
    n101
  );


  and
  g206
  (
    n240,
    n95,
    n199,
    n108,
    n75
  );


  or
  g207
  (
    n289,
    n45,
    n94,
    n78,
    n84
  );


  or
  g208
  (
    n283,
    n97,
    n39,
    n54,
    n116
  );


  and
  g209
  (
    n214,
    n89,
    n111,
    n48,
    n185
  );


  xor
  g210
  (
    n284,
    n62,
    n59,
    n55,
    n41
  );


  and
  g211
  (
    n205,
    n41,
    n64,
    n91,
    n101
  );


  xnor
  g212
  (
    n302,
    n192,
    n200,
    n191,
    n80
  );


  xnor
  g213
  (
    n259,
    n113,
    n182,
    n47,
    n193
  );


  nor
  g214
  (
    n225,
    n68,
    n44,
    n198,
    n55
  );


  xor
  g215
  (
    n213,
    n183,
    n79,
    n113,
    n112
  );


  or
  g216
  (
    n303,
    n176,
    n93,
    n196,
    n74
  );


  nand
  g217
  (
    n218,
    n178,
    n63,
    n74,
    n116
  );


  xnor
  g218
  (
    n232,
    n100,
    n42,
    n195,
    n102
  );


  nand
  g219
  (
    n279,
    n69,
    n201,
    n107,
    n175
  );


  xnor
  g220
  (
    n250,
    n90,
    n107,
    n85,
    n197
  );


  xnor
  g221
  (
    n227,
    n76,
    n65,
    n95,
    n67
  );


  nand
  g222
  (
    n239,
    n93,
    n108,
    n110
  );


  xnor
  g223
  (
    n293,
    n51,
    n58,
    n63,
    n117
  );


  or
  g224
  (
    n307,
    n67,
    n202,
    n80,
    n51
  );


  xor
  g225
  (
    n278,
    n102,
    n201,
    n43,
    n179
  );


  or
  g226
  (
    KeyWire_0_8,
    n50,
    n58,
    n105,
    n46
  );


  xor
  g227
  (
    n244,
    n108,
    n66,
    n109,
    n70
  );


  xor
  g228
  (
    n272,
    n111,
    n82,
    n51,
    n69
  );


  xor
  g229
  (
    n224,
    n104,
    n104,
    n192,
    n200
  );


  and
  g230
  (
    n267,
    n61,
    n92,
    n80,
    n188
  );


  or
  g231
  (
    n257,
    n39,
    n104,
    n66,
    n106
  );


  nand
  g232
  (
    n234,
    n61,
    n38,
    n189,
    n78
  );


  nor
  g233
  (
    n243,
    n191,
    n109,
    n62,
    n100
  );


  xnor
  g234
  (
    n287,
    n176,
    n85,
    n68,
    n81
  );


  and
  g235
  (
    n294,
    n190,
    n199,
    n70,
    n89
  );


  nor
  g236
  (
    n221,
    n190,
    n38,
    n92,
    n100
  );


  and
  g237
  (
    n265,
    n52,
    n113,
    n181,
    n116
  );


  or
  g238
  (
    n252,
    n177,
    n44,
    n184,
    n179
  );


  xor
  g239
  (
    n242,
    n191,
    n86,
    n61,
    n65
  );


  nand
  g240
  (
    n237,
    n52,
    n71,
    n55,
    n108
  );


  xor
  g241
  (
    n217,
    n95,
    n83,
    n81,
    n84
  );


  and
  g242
  (
    n210,
    n193,
    n60,
    n86,
    n91
  );


  xnor
  g243
  (
    n304,
    n99,
    n190,
    n50,
    n189
  );


  and
  g244
  (
    n254,
    n85,
    n48,
    n79,
    n88
  );


  nor
  g245
  (
    n230,
    n112,
    n40,
    n47,
    n92
  );


  nor
  g246
  (
    n216,
    n94,
    n56,
    n43
  );


  nand
  g247
  (
    n290,
    n89,
    n69,
    n188,
    n84
  );


  nor
  g248
  (
    n300,
    n88,
    n94,
    n92,
    n195
  );


  or
  g249
  (
    n246,
    n180,
    n183,
    n62,
    n71
  );


  nor
  g250
  (
    n285,
    n59,
    n107,
    n45,
    n73
  );


  xor
  g251
  (
    n238,
    n98,
    n65,
    n61,
    n106
  );


  nor
  g252
  (
    n207,
    n96,
    n60,
    n79,
    n58
  );


  xor
  g253
  (
    n222,
    n86,
    n97,
    n182
  );


  xnor
  g254
  (
    n255,
    n96,
    n74,
    n196,
    n41
  );


  or
  g255
  (
    n282,
    n101,
    n40,
    n105,
    n67
  );


  xor
  g256
  (
    n298,
    n185,
    n82,
    n68,
    n198
  );


  xnor
  g257
  (
    n288,
    n196,
    n76,
    n88,
    n70
  );


  xor
  g258
  (
    n233,
    n197,
    n187,
    n66,
    n87
  );


  or
  g259
  (
    n245,
    n111,
    n74,
    n181,
    n70
  );


  and
  g260
  (
    n308,
    n68,
    n114,
    n45,
    n49
  );


  nand
  g261
  (
    n249,
    n60,
    n56,
    n194,
    n180
  );


  xor
  g262
  (
    n209,
    n76,
    n87,
    n99,
    n49
  );


  nor
  g263
  (
    n215,
    n181,
    n105,
    n179,
    n39
  );


  nor
  g264
  (
    n269,
    n75,
    n90,
    n195,
    n112
  );


  xnor
  g265
  (
    n236,
    n193,
    n109,
    n54,
    n99
  );


  and
  g266
  (
    n228,
    n48,
    n202,
    n99,
    n192
  );


  xor
  g267
  (
    n248,
    n47,
    n49,
    n190,
    n43
  );


  xnor
  g268
  (
    n204,
    n63,
    n55,
    n42,
    n199
  );


  or
  g269
  (
    n253,
    n79,
    n105,
    n98,
    n186
  );


  xnor
  g270
  (
    n247,
    n200,
    n202,
    n57,
    n78
  );


  and
  g271
  (
    n208,
    n73,
    n85,
    n103,
    n193
  );


  xor
  g272
  (
    n235,
    n88,
    n200,
    n40,
    n91
  );


  nand
  g273
  (
    n262,
    n98,
    n201,
    n178,
    n59
  );


  or
  g274
  (
    n231,
    n57,
    n198,
    n197,
    n184
  );


  xor
  g275
  (
    n306,
    n50,
    n46,
    n186
  );


  xor
  g276
  (
    n291,
    n98,
    n101,
    n89,
    n78
  );


  xnor
  g277
  (
    n270,
    n116,
    n96,
    n40,
    n106
  );


  and
  g278
  (
    n258,
    n53,
    n84,
    n182,
    n110
  );


  xor
  g279
  (
    n260,
    n177,
    n47,
    n46,
    n73
  );


  nor
  g280
  (
    n206,
    n83,
    n106,
    n59,
    n183
  );


  nor
  g281
  (
    n219,
    n72,
    n77,
    n83,
    n39
  );


  nand
  g282
  (
    n299,
    n104,
    n194,
    n185,
    n72
  );


  buf
  g283
  (
    n378,
    n219
  );


  not
  g284
  (
    n361,
    n204
  );


  buf
  g285
  (
    n323,
    n214
  );


  buf
  g286
  (
    n327,
    n216
  );


  buf
  g287
  (
    n351,
    n207
  );


  buf
  g288
  (
    n359,
    n203
  );


  buf
  g289
  (
    n370,
    n220
  );


  buf
  g290
  (
    KeyWire_0_14,
    n203
  );


  buf
  g291
  (
    n357,
    n204
  );


  not
  g292
  (
    n311,
    n213
  );


  buf
  g293
  (
    n372,
    n210
  );


  not
  g294
  (
    n312,
    n205
  );


  not
  g295
  (
    n364,
    n205
  );


  not
  g296
  (
    n377,
    n216
  );


  buf
  g297
  (
    n355,
    n217
  );


  buf
  g298
  (
    n325,
    n219
  );


  buf
  g299
  (
    n352,
    n218
  );


  not
  g300
  (
    n337,
    n220
  );


  buf
  g301
  (
    n354,
    n215
  );


  not
  g302
  (
    n369,
    n208
  );


  not
  g303
  (
    n353,
    n205
  );


  not
  g304
  (
    n366,
    n154
  );


  buf
  g305
  (
    n321,
    n216
  );


  buf
  g306
  (
    n376,
    n203
  );


  not
  g307
  (
    n324,
    n209
  );


  buf
  g308
  (
    n356,
    n216
  );


  buf
  g309
  (
    KeyWire_0_27,
    n209
  );


  not
  g310
  (
    n348,
    n206
  );


  not
  g311
  (
    n342,
    n212
  );


  buf
  g312
  (
    n317,
    n207
  );


  buf
  g313
  (
    n335,
    n218
  );


  buf
  g314
  (
    n314,
    n212
  );


  buf
  g315
  (
    n374,
    n214
  );


  not
  g316
  (
    n346,
    n206
  );


  buf
  g317
  (
    n349,
    n208
  );


  buf
  g318
  (
    n334,
    n215
  );


  buf
  g319
  (
    n310,
    n213
  );


  not
  g320
  (
    n367,
    n211
  );


  buf
  g321
  (
    n328,
    n208
  );


  buf
  g322
  (
    n320,
    n204
  );


  buf
  g323
  (
    n345,
    n209
  );


  not
  g324
  (
    n329,
    n204
  );


  not
  g325
  (
    n331,
    n214
  );


  buf
  g326
  (
    n375,
    n205
  );


  not
  g327
  (
    n336,
    n217
  );


  buf
  g328
  (
    n365,
    n206
  );


  buf
  g329
  (
    n373,
    n208
  );


  buf
  g330
  (
    n313,
    n220
  );


  not
  g331
  (
    n315,
    n214
  );


  buf
  g332
  (
    n350,
    n209
  );


  buf
  g333
  (
    n322,
    n206
  );


  buf
  g334
  (
    n316,
    n213
  );


  not
  g335
  (
    n362,
    n211
  );


  buf
  g336
  (
    n363,
    n219
  );


  not
  g337
  (
    n319,
    n203
  );


  not
  g338
  (
    KeyWire_0_25,
    n217
  );


  not
  g339
  (
    n330,
    n219
  );


  buf
  g340
  (
    n371,
    n210
  );


  not
  g341
  (
    n318,
    n210
  );


  buf
  g342
  (
    n340,
    n212
  );


  buf
  g343
  (
    n309,
    n211
  );


  not
  g344
  (
    n339,
    n207
  );


  buf
  g345
  (
    n360,
    n215
  );


  buf
  g346
  (
    n347,
    n217
  );


  buf
  g347
  (
    n333,
    n207
  );


  buf
  g348
  (
    n358,
    n212
  );


  not
  g349
  (
    n344,
    n215
  );


  buf
  g350
  (
    n338,
    n210
  );


  buf
  g351
  (
    n341,
    n211
  );


  not
  g352
  (
    n379,
    n218
  );


  and
  g353
  (
    n343,
    n213,
    n218
  );


  and
  g354
  (
    n386,
    n368,
    n227,
    n224,
    n373
  );


  nor
  g355
  (
    n438,
    n319,
    n230,
    n372,
    n120
  );


  nor
  g356
  (
    n426,
    n242,
    n261,
    n245,
    n310
  );


  or
  g357
  (
    n396,
    n236,
    n263,
    n229,
    n269
  );


  xnor
  g358
  (
    n401,
    n221,
    n377,
    n230,
    n253
  );


  nand
  g359
  (
    n451,
    n253,
    n331,
    n361,
    n241
  );


  or
  g360
  (
    n403,
    n256,
    n246,
    n358,
    n250
  );


  nand
  g361
  (
    n434,
    n120,
    n120,
    n367,
    n247
  );


  and
  g362
  (
    n394,
    n264,
    n257,
    n231,
    n223
  );


  or
  g363
  (
    n397,
    n347,
    n235,
    n264,
    n226
  );


  nand
  g364
  (
    n417,
    n312,
    n363,
    n242,
    n125
  );


  and
  g365
  (
    n416,
    n235,
    n257,
    n121,
    n125
  );


  and
  g366
  (
    n445,
    n121,
    n238,
    n318,
    n125
  );


  or
  g367
  (
    n411,
    n330,
    n262,
    n265,
    n122
  );


  xor
  g368
  (
    KeyWire_0_22,
    n376,
    n222,
    n352,
    n264
  );


  nand
  g369
  (
    n380,
    n263,
    n233,
    n239,
    n320
  );


  or
  g370
  (
    n420,
    n260,
    n243,
    n378,
    n123
  );


  or
  g371
  (
    n408,
    n246,
    n227,
    n221,
    n124
  );


  xnor
  g372
  (
    n429,
    n236,
    n120,
    n376,
    n268
  );


  nor
  g373
  (
    n409,
    n228,
    n254,
    n236,
    n223
  );


  nand
  g374
  (
    n384,
    n235,
    n265,
    n252,
    n346
  );


  nand
  g375
  (
    n390,
    n263,
    n225,
    n266,
    n119
  );


  or
  g376
  (
    n407,
    n349,
    n258,
    n309,
    n243
  );


  and
  g377
  (
    n414,
    n232,
    n223,
    n328,
    n321
  );


  nand
  g378
  (
    n436,
    n240,
    n262,
    n344,
    n233
  );


  xor
  g379
  (
    KeyWire_0_3,
    n234,
    n222,
    n123,
    n258
  );


  xnor
  g380
  (
    n422,
    n234,
    n235,
    n266,
    n245
  );


  nand
  g381
  (
    n415,
    n221,
    n324,
    n247,
    n267
  );


  and
  g382
  (
    n425,
    n329,
    n228,
    n236,
    n248
  );


  or
  g383
  (
    n418,
    n234,
    n232,
    n342,
    n252
  );


  nand
  g384
  (
    n435,
    n314,
    n256,
    n249
  );


  or
  g385
  (
    n446,
    n228,
    n243,
    n375,
    n118
  );


  nor
  g386
  (
    n440,
    n247,
    n315,
    n226,
    n362
  );


  xor
  g387
  (
    n381,
    n123,
    n248,
    n243,
    n255
  );


  nand
  g388
  (
    n439,
    n241,
    n221,
    n341,
    n259
  );


  nor
  g389
  (
    KeyWire_0_9,
    n124,
    n224,
    n366,
    n229
  );


  or
  g390
  (
    n447,
    n254,
    n245,
    n226,
    n118
  );


  nand
  g391
  (
    n387,
    n123,
    n245,
    n327,
    n122
  );


  and
  g392
  (
    n441,
    n237,
    n230,
    n267,
    n255
  );


  xor
  g393
  (
    n437,
    n238,
    n226,
    n322,
    n268
  );


  or
  g394
  (
    n455,
    n244,
    n260,
    n124,
    n268
  );


  nor
  g395
  (
    n453,
    n227,
    n359,
    n125,
    n357
  );


  nor
  g396
  (
    n402,
    n355,
    n339,
    n374,
    n223
  );


  or
  g397
  (
    KeyWire_0_31,
    n316,
    n225,
    n119,
    n375
  );


  xor
  g398
  (
    n383,
    n354,
    n222,
    n119,
    n317
  );


  nand
  g399
  (
    n398,
    n253,
    n370,
    n256,
    n269
  );


  xnor
  g400
  (
    n432,
    n231,
    n232,
    n313,
    n345
  );


  and
  g401
  (
    n404,
    n254,
    n230,
    n260,
    n237
  );


  and
  g402
  (
    n454,
    n365,
    n220,
    n242,
    n258
  );


  or
  g403
  (
    n388,
    n122,
    n237,
    n360,
    n238
  );


  xnor
  g404
  (
    n448,
    n251,
    n251,
    n248,
    n257
  );


  and
  g405
  (
    n410,
    n231,
    n350,
    n249,
    n261
  );


  xor
  g406
  (
    n431,
    n124,
    n256,
    n121,
    n332
  );


  or
  g407
  (
    n442,
    n264,
    n356,
    n254,
    n351
  );


  and
  g408
  (
    n443,
    n250,
    n122,
    n244,
    n253
  );


  or
  g409
  (
    n413,
    n234,
    n117,
    n336,
    n340
  );


  nand
  g410
  (
    n444,
    n262,
    n252,
    n244,
    n250
  );


  xor
  g411
  (
    n423,
    n251,
    n259,
    n379,
    n239
  );


  xor
  g412
  (
    n412,
    n222,
    n323,
    n233,
    n251
  );


  xnor
  g413
  (
    n427,
    n246,
    n377,
    n119,
    n266
  );


  or
  g414
  (
    n385,
    n121,
    n241,
    n258,
    n240
  );


  xor
  g415
  (
    n389,
    n265,
    n343,
    n250,
    n337
  );


  and
  g416
  (
    n395,
    n338,
    n247,
    n232,
    n378
  );


  xnor
  g417
  (
    n399,
    n348,
    n261,
    n246,
    n248
  );


  nor
  g418
  (
    n430,
    n267,
    n239,
    n369,
    n231
  );


  nand
  g419
  (
    n400,
    n237,
    n364,
    n263,
    n225
  );


  xor
  g420
  (
    n452,
    n225,
    n335,
    n229,
    n240
  );


  nand
  g421
  (
    n433,
    n239,
    n333,
    n240,
    n224
  );


  nand
  g422
  (
    n421,
    n118,
    n353,
    n311,
    n260
  );


  or
  g423
  (
    n405,
    n371,
    n228,
    n227,
    n262
  );


  xor
  g424
  (
    n449,
    n241,
    n224,
    n242,
    n249
  );


  and
  g425
  (
    KeyWire_0_15,
    n379,
    n259,
    n334
  );


  nor
  g426
  (
    n428,
    n257,
    n261,
    n325,
    n326
  );


  xor
  g427
  (
    n392,
    n233,
    n238,
    n267,
    n265
  );


  nand
  g428
  (
    n450,
    n255,
    n266,
    n268,
    n252
  );


  nand
  g429
  (
    n382,
    n118,
    n229,
    n255,
    n244
  );


  xnor
  g430
  (
    n527,
    n455,
    n387,
    n450,
    n170
  );


  nor
  g431
  (
    n545,
    n303,
    n454,
    n306,
    n416
  );


  nand
  g432
  (
    n511,
    n277,
    n278,
    n432,
    n455
  );


  or
  g433
  (
    n490,
    n416,
    n428,
    n308,
    n295
  );


  nor
  g434
  (
    n458,
    n293,
    n419,
    n392,
    n300
  );


  or
  g435
  (
    n497,
    n423,
    n297,
    n279,
    n382
  );


  xor
  g436
  (
    n510,
    n426,
    n402,
    n452,
    n276
  );


  or
  g437
  (
    n475,
    n304,
    n441,
    n423,
    n163
  );


  or
  g438
  (
    n470,
    n278,
    n436,
    n302
  );


  nor
  g439
  (
    n509,
    n292,
    n269,
    n301,
    n441
  );


  nor
  g440
  (
    n495,
    n274,
    n284,
    n270,
    n296
  );


  nand
  g441
  (
    n476,
    n293,
    n453,
    n271,
    n283
  );


  xor
  g442
  (
    n494,
    n434,
    n438,
    n277,
    n279
  );


  xor
  g443
  (
    n547,
    n280,
    n271,
    n290,
    n453
  );


  xnor
  g444
  (
    n501,
    n441,
    n443,
    n174,
    n288
  );


  xor
  g445
  (
    n463,
    n164,
    n285,
    n298,
    n290
  );


  and
  g446
  (
    KeyWire_0_20,
    n297,
    n288,
    n301,
    n292
  );


  and
  g447
  (
    n479,
    n306,
    n161,
    n389,
    n393
  );


  or
  g448
  (
    n529,
    n439,
    n399,
    n275,
    n305
  );


  nand
  g449
  (
    n551,
    n291,
    n440,
    n276,
    n447
  );


  xnor
  g450
  (
    n461,
    n308,
    n282,
    n422,
    n412
  );


  nor
  g451
  (
    n505,
    n279,
    n278,
    n411,
    n440
  );


  xor
  g452
  (
    n456,
    n282,
    n412,
    n431,
    n408
  );


  or
  g453
  (
    n522,
    n272,
    n300,
    n420,
    n427
  );


  xor
  g454
  (
    n483,
    n454,
    n275,
    n444,
    n283
  );


  and
  g455
  (
    n467,
    n289,
    n307,
    n430
  );


  nand
  g456
  (
    n539,
    n287,
    n422,
    n433,
    n410
  );


  nor
  g457
  (
    n516,
    n413,
    n421,
    n451,
    n389
  );


  nor
  g458
  (
    n488,
    n273,
    n275,
    n293,
    n437
  );


  nor
  g459
  (
    KeyWire_0_30,
    n386,
    n396,
    n453,
    n280
  );


  xor
  g460
  (
    KeyWire_0_11,
    n304,
    n283,
    n398,
    n417
  );


  nand
  g461
  (
    n525,
    n419,
    n385,
    n454,
    n303
  );


  and
  g462
  (
    n496,
    n404,
    n162,
    n430,
    n290
  );


  xor
  g463
  (
    n519,
    n410,
    n442,
    n444,
    n446
  );


  xor
  g464
  (
    n524,
    n445,
    n442,
    n434,
    n302
  );


  nand
  g465
  (
    n486,
    n308,
    n302,
    n285,
    n440
  );


  xnor
  g466
  (
    n507,
    n438,
    n450,
    n439,
    n296
  );


  or
  g467
  (
    n538,
    n384,
    n429,
    n298,
    n382
  );


  or
  g468
  (
    n540,
    n421,
    n450,
    n282,
    n442
  );


  nor
  g469
  (
    n514,
    n286,
    n299,
    n391,
    n381
  );


  xor
  g470
  (
    n532,
    n296,
    n269,
    n435,
    n384
  );


  xor
  g471
  (
    n534,
    n301,
    n449,
    n414,
    n286
  );


  nand
  g472
  (
    n533,
    n438,
    n443,
    n431,
    n407
  );


  nor
  g473
  (
    n536,
    n290,
    n276,
    n284,
    n425
  );


  and
  g474
  (
    n512,
    n301,
    n405,
    n427,
    n407
  );


  nor
  g475
  (
    n518,
    n441,
    n281,
    n298,
    n284
  );


  xnor
  g476
  (
    n499,
    n438,
    n403,
    n437,
    n306
  );


  nand
  g477
  (
    n520,
    n272,
    n439,
    n432,
    n165
  );


  nor
  g478
  (
    n466,
    n284,
    n280,
    n390,
    n394
  );


  xor
  g479
  (
    n472,
    n432,
    n272,
    n455,
    n283
  );


  and
  g480
  (
    n484,
    n433,
    n388,
    n279,
    n383
  );


  nand
  g481
  (
    n537,
    n280,
    n277,
    n292,
    n380
  );


  xor
  g482
  (
    n459,
    n158,
    n426,
    n415,
    n424
  );


  xor
  g483
  (
    n550,
    n388,
    n285,
    n444,
    n434
  );


  xor
  g484
  (
    n542,
    n446,
    n386,
    n397,
    n444
  );


  and
  g485
  (
    n515,
    n400,
    n302,
    n418,
    n288
  );


  xnor
  g486
  (
    n477,
    n431,
    n455,
    n303,
    n452
  );


  xor
  g487
  (
    n474,
    n276,
    n281,
    n417,
    n437
  );


  xnor
  g488
  (
    n543,
    n387,
    n397,
    n409,
    n437
  );


  and
  g489
  (
    n481,
    n443,
    n299,
    n415
  );


  xor
  g490
  (
    n498,
    n270,
    n285,
    n448,
    n454
  );


  or
  g491
  (
    KeyWire_0_16,
    n396,
    n298,
    n304,
    n449
  );


  xnor
  g492
  (
    n480,
    n434,
    n270,
    n289,
    n160
  );


  and
  g493
  (
    n546,
    n445,
    n435,
    n381,
    n295
  );


  xor
  g494
  (
    n487,
    n278,
    n271,
    n411,
    n451
  );


  or
  g495
  (
    n521,
    n404,
    n287,
    n440,
    n294
  );


  and
  g496
  (
    n485,
    n296,
    n433,
    n307,
    n171
  );


  xnor
  g497
  (
    n506,
    n447,
    n156,
    n405,
    n297
  );


  nand
  g498
  (
    KeyWire_0_1,
    n425,
    n450,
    n398,
    n435
  );


  and
  g499
  (
    n502,
    n428,
    n447,
    n430,
    n432
  );


  nor
  g500
  (
    n541,
    n431,
    n451,
    n447,
    n270
  );


  xnor
  g501
  (
    n526,
    n406,
    n295,
    n430,
    n408
  );


  xor
  g502
  (
    n478,
    n297,
    n401,
    n288,
    n155
  );


  xnor
  g503
  (
    n535,
    n380,
    n289,
    n452
  );


  and
  g504
  (
    n492,
    n291,
    n452,
    n429,
    n273
  );


  xnor
  g505
  (
    n528,
    n169,
    n449,
    n273,
    n445
  );


  xnor
  g506
  (
    n482,
    n166,
    n392,
    n271,
    n304
  );


  and
  g507
  (
    n457,
    n453,
    n391,
    n443,
    n395
  );


  or
  g508
  (
    n523,
    n300,
    n394,
    n303,
    n448
  );


  or
  g509
  (
    n513,
    n305,
    n435,
    n395,
    n275
  );


  nor
  g510
  (
    n493,
    n293,
    n292,
    n295,
    n448
  );


  xnor
  g511
  (
    n544,
    n281,
    n157,
    n445,
    n433
  );


  nor
  g512
  (
    n491,
    n286,
    n449,
    n305,
    n291
  );


  xor
  g513
  (
    KeyWire_0_13,
    n414,
    n446,
    n306,
    n305
  );


  or
  g514
  (
    n500,
    n172,
    n274,
    n399,
    n442
  );


  xor
  g515
  (
    n465,
    n420,
    n168,
    n299,
    n272
  );


  or
  g516
  (
    n462,
    n294,
    n300,
    n403,
    n308
  );


  and
  g517
  (
    KeyWire_0_26,
    n286,
    n383,
    n436,
    n424
  );


  xor
  g518
  (
    n530,
    n385,
    n393,
    n274,
    n402
  );


  or
  g519
  (
    n464,
    n159,
    n436,
    n390,
    n281
  );


  nand
  g520
  (
    n503,
    n418,
    n451,
    n294,
    n406
  );


  nor
  g521
  (
    n468,
    n167,
    n273,
    n439,
    n429
  );


  or
  g522
  (
    n469,
    n173,
    n294,
    n413,
    n401
  );


  nand
  g523
  (
    KeyWire_0_4,
    n287,
    n282,
    n429,
    n400
  );


  or
  g524
  (
    n549,
    n274,
    n448,
    n287,
    n307
  );


  or
  g525
  (
    n517,
    n446,
    n409,
    n277,
    n291
  );


  and
  g526
  (
    KeyWire_0_18,
    n543,
    n538,
    n499,
    n472
  );


  xnor
  g527
  (
    n557,
    n507,
    n508,
    n509,
    n534
  );


  nand
  g528
  (
    n563,
    n487,
    n475,
    n473,
    n551
  );


  xor
  g529
  (
    n559,
    n527,
    n535,
    n512,
    n469
  );


  or
  g530
  (
    n556,
    n529,
    n496,
    n541,
    n511
  );


  xnor
  g531
  (
    KeyWire_0_7,
    n470,
    n471,
    n549,
    n460
  );


  nor
  g532
  (
    n552,
    n531,
    n518,
    n528,
    n484
  );


  or
  g533
  (
    n575,
    n486,
    n515,
    n546,
    n474
  );


  nor
  g534
  (
    n564,
    n466,
    n514,
    n524,
    n495
  );


  or
  g535
  (
    n565,
    n545,
    n467,
    n492,
    n482
  );


  xor
  g536
  (
    KeyWire_0_21,
    n533,
    n491,
    n498,
    n516
  );


  nor
  g537
  (
    n558,
    n456,
    n468,
    n540,
    n513
  );


  xor
  g538
  (
    n554,
    n458,
    n536,
    n525,
    n526
  );


  and
  g539
  (
    n562,
    n510,
    n521,
    n547,
    n542
  );


  and
  g540
  (
    n560,
    n483,
    n493,
    n502,
    n457
  );


  and
  g541
  (
    n569,
    n501,
    n490,
    n530,
    n464
  );


  or
  g542
  (
    n571,
    n480,
    n519,
    n503,
    n459
  );


  xor
  g543
  (
    n573,
    n465,
    n517,
    n505,
    n478
  );


  nand
  g544
  (
    n561,
    n488,
    n544,
    n548,
    n494
  );


  xor
  g545
  (
    n568,
    n532,
    n479,
    n506,
    n477
  );


  xor
  g546
  (
    n555,
    n489,
    n463,
    n504,
    n523
  );


  nor
  g547
  (
    n553,
    n537,
    n461,
    n500,
    n481
  );


  nand
  g548
  (
    n574,
    n520,
    n485,
    n462,
    n497
  );


  xor
  g549
  (
    n572,
    n476,
    n539,
    n550,
    n522
  );


  xor
  KeyGate_0_0
  (
    n167,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n508,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n103,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n391,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n489,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n160,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n27,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n566,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n203,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n424,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n30,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n504,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n127,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n548,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n368,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n419,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n531,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n41,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n570,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n36,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n471,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n567,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n406,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n188,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n102,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n332,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n460,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n326,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n154,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n180,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n473,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n393,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


