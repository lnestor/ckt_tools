// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_913_268 written by SynthGen on 2021/05/24 19:48:31
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_913_268 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n681, n686, n684, n682, n690, n693, n696, n692,
 n691, n699, n695, n698, n865, n943, n938, n945,
 n941, n940, n937, n942, n935, n936, n939, n944);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n681, n686, n684, n682, n690, n693, n696, n692,
 n691, n699, n695, n698, n865, n943, n938, n945,
 n941, n940, n937, n942, n935, n936, n939, n944;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n683, n685, n687, n688, n689, n694, n697, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n758, n759, n760, n761, n762, n763, n764,
 n765, n766, n767, n768, n769, n770, n771, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n866, n867, n868, n869,
 n870, n871, n872, n873, n874, n875, n876, n877,
 n878, n879, n880, n881, n882, n883, n884, n885,
 n886, n887, n888, n889, n890, n891, n892, n893,
 n894, n895, n896, n897, n898, n899, n900, n901,
 n902, n903, n904, n905, n906, n907, n908, n909,
 n910, n911, n912, n913, n914, n915, n916, n917,
 n918, n919, n920, n921, n922, n923, n924, n925,
 n926, n927, n928, n929, n930, n931, n932, n933,
 n934;

buf  g0 (n157, n10);
not  g1 (n94, n26);
buf  g2 (n121, n1);
not  g3 (n125, n21);
buf  g4 (n47, n27);
buf  g5 (n151, n15);
not  g6 (n37, n29);
buf  g7 (n111, n25);
buf  g8 (n80, n18);
not  g9 (n84, n31);
not  g10 (n128, n28);
not  g11 (n103, n30);
not  g12 (n150, n14);
not  g13 (n38, n5);
not  g14 (n105, n23);
not  g15 (n132, n15);
buf  g16 (n152, n6);
not  g17 (n137, n26);
not  g18 (n41, n24);
not  g19 (n81, n12);
not  g20 (n99, n4);
not  g21 (n88, n23);
not  g22 (n71, n32);
not  g23 (n139, n15);
not  g24 (n146, n6);
buf  g25 (n98, n28);
buf  g26 (n122, n3);
buf  g27 (n54, n29);
buf  g28 (n113, n21);
not  g29 (n66, n11);
buf  g30 (n119, n25);
not  g31 (n69, n16);
buf  g32 (n110, n7);
not  g33 (n72, n14);
buf  g34 (n44, n10);
buf  g35 (n90, n28);
buf  g36 (n148, n19);
not  g37 (n63, n22);
buf  g38 (n67, n28);
buf  g39 (n89, n12);
not  g40 (n97, n31);
not  g41 (n65, n31);
not  g42 (n142, n10);
not  g43 (n33, n18);
buf  g44 (n159, n9);
buf  g45 (n73, n1);
not  g46 (n87, n9);
not  g47 (n149, n5);
buf  g48 (n102, n14);
not  g49 (n61, n24);
not  g50 (n147, n13);
buf  g51 (n108, n7);
buf  g52 (n124, n13);
buf  g53 (n93, n5);
not  g54 (n43, n25);
not  g55 (n153, n29);
not  g56 (n145, n21);
not  g57 (n130, n11);
buf  g58 (n135, n32);
buf  g59 (n158, n14);
not  g60 (n64, n8);
not  g61 (n106, n27);
buf  g62 (n136, n8);
buf  g63 (n129, n3);
not  g64 (n50, n30);
not  g65 (n49, n15);
not  g66 (n144, n20);
buf  g67 (n74, n27);
not  g68 (n82, n18);
not  g69 (n95, n24);
buf  g70 (n115, n4);
not  g71 (n116, n32);
not  g72 (n83, n7);
not  g73 (n48, n18);
not  g74 (n91, n8);
not  g75 (n101, n26);
buf  g76 (n117, n27);
not  g77 (n59, n31);
not  g78 (n127, n17);
buf  g79 (n52, n23);
buf  g80 (n155, n16);
not  g81 (n160, n22);
not  g82 (n36, n26);
not  g83 (n78, n32);
not  g84 (n70, n2);
buf  g85 (n141, n9);
buf  g86 (n34, n1);
not  g87 (n143, n25);
buf  g88 (n56, n30);
buf  g89 (n68, n13);
not  g90 (n60, n16);
buf  g91 (n120, n2);
buf  g92 (n77, n12);
buf  g93 (n112, n19);
not  g94 (n86, n3);
buf  g95 (n51, n4);
not  g96 (n55, n20);
buf  g97 (n109, n1);
not  g98 (n75, n23);
not  g99 (n42, n17);
buf  g100 (n46, n11);
buf  g101 (n85, n4);
not  g102 (n126, n29);
buf  g103 (n39, n22);
not  g104 (n62, n20);
not  g105 (n76, n12);
buf  g106 (n57, n17);
not  g107 (n92, n10);
buf  g108 (n45, n3);
not  g109 (n134, n30);
buf  g110 (n138, n21);
not  g111 (n114, n22);
not  g112 (n58, n19);
not  g113 (n53, n2);
not  g114 (n100, n9);
buf  g115 (n154, n6);
buf  g116 (n140, n7);
not  g117 (n131, n16);
not  g118 (n107, n24);
not  g119 (n133, n13);
buf  g120 (n79, n17);
not  g121 (n123, n19);
buf  g122 (n40, n8);
not  g123 (n156, n11);
buf  g124 (n35, n20);
not  g125 (n96, n6);
not  g126 (n104, n5);
not  g127 (n118, n2);
not  g128 (n392, n33);
buf  g129 (n213, n142);
not  g130 (n306, n75);
not  g131 (n202, n51);
buf  g132 (n182, n67);
buf  g133 (n429, n45);
not  g134 (n442, n61);
buf  g135 (n178, n117);
buf  g136 (n322, n56);
buf  g137 (n342, n144);
not  g138 (n169, n148);
buf  g139 (n179, n136);
not  g140 (n247, n128);
buf  g141 (n210, n74);
not  g142 (n272, n137);
not  g143 (n197, n99);
buf  g144 (n358, n136);
not  g145 (n257, n35);
buf  g146 (n294, n46);
buf  g147 (n302, n50);
not  g148 (n451, n145);
not  g149 (n377, n47);
buf  g150 (n224, n147);
buf  g151 (n414, n122);
not  g152 (n276, n126);
not  g153 (n323, n107);
not  g154 (n352, n84);
buf  g155 (n223, n68);
buf  g156 (n399, n53);
not  g157 (n436, n37);
not  g158 (n419, n91);
buf  g159 (n263, n113);
not  g160 (n389, n56);
buf  g161 (n232, n76);
not  g162 (n295, n91);
not  g163 (n362, n42);
not  g164 (n338, n91);
not  g165 (n382, n108);
buf  g166 (n349, n90);
buf  g167 (n471, n72);
buf  g168 (n261, n146);
buf  g169 (n446, n140);
not  g170 (n353, n113);
not  g171 (n395, n94);
not  g172 (n415, n88);
buf  g173 (n273, n147);
not  g174 (n423, n82);
buf  g175 (n312, n91);
not  g176 (n246, n147);
not  g177 (n435, n81);
not  g178 (n360, n132);
not  g179 (n409, n142);
not  g180 (n385, n65);
not  g181 (n404, n145);
buf  g182 (n443, n129);
buf  g183 (n198, n86);
buf  g184 (n420, n120);
not  g185 (n229, n142);
buf  g186 (n316, n118);
buf  g187 (n344, n96);
buf  g188 (n403, n37);
not  g189 (n278, n34);
buf  g190 (n464, n126);
buf  g191 (n196, n38);
buf  g192 (n245, n48);
buf  g193 (n175, n97);
not  g194 (n287, n49);
not  g195 (n288, n39);
not  g196 (n274, n116);
not  g197 (n383, n72);
buf  g198 (n172, n150);
not  g199 (n215, n122);
not  g200 (n356, n124);
buf  g201 (n239, n88);
not  g202 (n265, n106);
not  g203 (n454, n115);
buf  g204 (n388, n138);
not  g205 (n386, n135);
not  g206 (n290, n84);
buf  g207 (n235, n69);
not  g208 (n381, n95);
not  g209 (n199, n124);
not  g210 (n244, n107);
buf  g211 (n359, n81);
not  g212 (n298, n47);
buf  g213 (n397, n43);
not  g214 (n343, n123);
not  g215 (n328, n128);
buf  g216 (n194, n126);
buf  g217 (n432, n109);
buf  g218 (n363, n34);
not  g219 (n333, n117);
not  g220 (n228, n71);
not  g221 (n309, n92);
buf  g222 (n268, n49);
not  g223 (n410, n88);
buf  g224 (n264, n154);
not  g225 (n424, n34);
not  g226 (n472, n89);
buf  g227 (n440, n66);
buf  g228 (n171, n102);
not  g229 (n254, n127);
not  g230 (n369, n40);
not  g231 (n260, n67);
buf  g232 (n332, n114);
buf  g233 (n334, n37);
buf  g234 (n370, n148);
buf  g235 (n315, n103);
buf  g236 (n378, n45);
buf  g237 (n475, n66);
not  g238 (n405, n151);
buf  g239 (n325, n60);
buf  g240 (n321, n79);
buf  g241 (n307, n46);
buf  g242 (n331, n77);
buf  g243 (n310, n96);
not  g244 (n296, n36);
buf  g245 (n350, n120);
buf  g246 (n188, n74);
not  g247 (n367, n92);
not  g248 (n402, n111);
not  g249 (n262, n83);
buf  g250 (n324, n69);
not  g251 (n366, n65);
not  g252 (n418, n79);
buf  g253 (n167, n69);
buf  g254 (n201, n124);
not  g255 (n177, n127);
not  g256 (n444, n55);
buf  g257 (n200, n125);
not  g258 (n463, n122);
buf  g259 (n212, n152);
buf  g260 (n161, n41);
not  g261 (n162, n106);
not  g262 (n303, n47);
not  g263 (n330, n76);
not  g264 (n434, n83);
not  g265 (n391, n38);
buf  g266 (n291, n131);
buf  g267 (n227, n41);
not  g268 (n318, n36);
buf  g269 (n368, n43);
not  g270 (n271, n115);
not  g271 (n340, n78);
buf  g272 (n433, n150);
not  g273 (n181, n84);
not  g274 (n209, n136);
buf  g275 (n412, n40);
not  g276 (n237, n94);
not  g277 (n173, n148);
buf  g278 (n455, n44);
buf  g279 (n190, n104);
buf  g280 (n374, n131);
not  g281 (n259, n53);
buf  g282 (n365, n105);
buf  g283 (n417, n67);
not  g284 (n279, n107);
not  g285 (n217, n85);
not  g286 (n241, n151);
buf  g287 (n195, n134);
buf  g288 (n207, n95);
not  g289 (n387, n102);
not  g290 (n300, n152);
not  g291 (n460, n103);
not  g292 (n336, n68);
buf  g293 (n269, n63);
not  g294 (n456, n59);
buf  g295 (n408, n59);
buf  g296 (n345, n141);
buf  g297 (n170, n114);
not  g298 (n165, n143);
buf  g299 (n219, n129);
buf  g300 (n281, n35);
not  g301 (n384, n100);
buf  g302 (n208, n100);
buf  g303 (n448, n98);
not  g304 (n411, n44);
not  g305 (n441, n38);
buf  g306 (n252, n52);
not  g307 (n299, n40);
not  g308 (n308, n121);
not  g309 (n248, n87);
not  g310 (n311, n109);
not  g311 (n327, n89);
buf  g312 (n275, n134);
buf  g313 (n166, n110);
buf  g314 (n314, n76);
buf  g315 (n192, n108);
not  g316 (n204, n75);
not  g317 (n430, n80);
buf  g318 (n355, n65);
not  g319 (n267, n127);
not  g320 (n280, n119);
not  g321 (n428, n90);
buf  g322 (n230, n98);
not  g323 (n465, n80);
buf  g324 (n238, n134);
buf  g325 (n211, n62);
buf  g326 (n317, n56);
buf  g327 (n461, n133);
not  g328 (n250, n101);
not  g329 (n220, n50);
buf  g330 (n176, n105);
not  g331 (n185, n109);
buf  g332 (n351, n139);
not  g333 (n187, n149);
not  g334 (n427, n102);
buf  g335 (n186, n122);
buf  g336 (n270, n56);
not  g337 (n469, n82);
not  g338 (n406, n124);
not  g339 (n214, n71);
buf  g340 (n329, n76);
buf  g341 (n297, n84);
not  g342 (n462, n140);
not  g343 (n304, n139);
buf  g344 (n163, n78);
not  g345 (n354, n55);
not  g346 (n305, n86);
buf  g347 (n242, n73);
buf  g348 (n277, n68);
not  g349 (n174, n52);
not  g350 (n326, n89);
not  g351 (n470, n152);
not  g352 (n438, n107);
buf  g353 (n337, n146);
not  g354 (n361, n120);
not  g355 (n218, n139);
buf  g356 (n205, n82);
not  g357 (n400, n60);
buf  g358 (n286, n64);
buf  g359 (n236, n80);
buf  g360 (n258, n94);
not  g361 (n206, n78);
not  g362 (n347, n146);
buf  g363 (n289, n114);
not  g364 (n180, n61);
not  g365 (n203, n121);
buf  g366 (n293, n132);
not  g367 (n393, n63);
not  g368 (n221, n136);
buf  g369 (n466, n120);
buf  g370 (n346, n70);
not  g371 (n447, n55);
not  g372 (n253, n106);
buf  g373 (n425, n135);
not  g374 (n422, n60);
buf  g375 (n401, n111);
buf  g376 (n183, n109);
buf  g377 (n283, n39);
buf  g378 (n474, n47);
buf  g379 (n292, n73);
not  g380 (n375, n113);
not  g381 (n320, n51);
not  g382 (n473, n73);
not  g383 (n467, n64);
buf  g384 (n371, n125);
not  g385 (n284, n42);
nor  g386 (n357, n62, n137, n59);
xor  g387 (n439, n51, n39, n42, n103);
or   g388 (n431, n110, n39, n137, n64);
and  g389 (n376, n118, n45, n44, n104);
xor  g390 (n233, n70, n133, n75, n130);
nand g391 (n421, n137, n74, n115, n57);
xnor g392 (n164, n58, n99, n121, n110);
xor  g393 (n226, n87, n61, n96, n101);
xnor g394 (n319, n135, n141, n112, n134);
nand g395 (n450, n112, n57, n104, n138);
xor  g396 (n168, n104, n121, n48, n41);
and  g397 (n243, n149, n85, n111, n130);
and  g398 (n416, n132, n85, n118, n130);
or   g399 (n453, n38, n49, n98, n130);
xor  g400 (n407, n149, n138, n147, n69);
xnor g401 (n234, n149, n75, n60, n140);
nand g402 (n458, n116, n145, n153, n72);
and  g403 (n437, n92, n95, n67, n62);
xnor g404 (n282, n81, n52, n79, n53);
and  g405 (n189, n112, n119, n64, n68);
or   g406 (n255, n62, n113, n105, n36);
nand g407 (n364, n123, n117, n111, n131);
xnor g408 (n348, n96, n94, n140, n63);
nor  g409 (n452, n135, n33, n119, n143);
or   g410 (n313, n141, n70, n34, n108);
xor  g411 (n426, n78, n44, n98, n77);
xor  g412 (n339, n101, n43, n99, n61);
nor  g413 (n240, n37, n86, n41, n152);
nand g414 (n222, n114, n93, n106, n82);
nor  g415 (n398, n89, n46, n97, n73);
nor  g416 (n468, n151, n87, n116, n153);
nor  g417 (n301, n123, n139, n50, n142);
or   g418 (n193, n129, n51, n133, n59);
xor  g419 (n372, n48, n48, n54, n63);
nand g420 (n459, n126, n112, n93, n153);
or   g421 (n445, n43, n97, n74, n110);
or   g422 (n390, n144, n58, n80, n33);
xor  g423 (n231, n58, n151, n93, n70);
and  g424 (n256, n35, n128, n85, n86);
and  g425 (n449, n58, n148, n146, n55);
xnor g426 (n373, n77, n100, n145, n57);
and  g427 (n285, n52, n35, n88, n99);
nor  g428 (n379, n54, n66, n138, n117);
xor  g429 (n380, n131, n118, n81, n144);
and  g430 (n266, n132, n79, n54, n108);
xor  g431 (n184, n93, n153, n115, n150);
xor  g432 (n216, n123, n66, n87, n105);
and  g433 (n341, n72, n71, n102, n83);
xor  g434 (n225, n133, n144, n129, n97);
nor  g435 (n335, n45, n150, n116, n71);
xor  g436 (n249, n57, n119, n125, n143);
xnor g437 (n191, n83, n128, n65, n92);
or   g438 (n413, n127, n77, n33, n90);
and  g439 (n457, n143, n49, n125, n50);
nand g440 (n251, n53, n103, n100, n101);
nand g441 (n394, n90, n36, n40, n141);
nand g442 (n396, n95, n42, n46, n54);
nand g443 (n491, n178, n181, n220, n222);
or   g444 (n490, n162, n170, n217, n200);
nand g445 (n484, n212, n186, n184, n227);
nor  g446 (n492, n183, n205, n175, n190);
xor  g447 (n478, n214, n196, n163, n216);
or   g448 (n476, n179, n191, n206, n164);
xnor g449 (n488, n177, n172, n182, n161);
nor  g450 (n493, n180, n202, n174, n219);
xor  g451 (n479, n204, n228, n171, n207);
xor  g452 (n483, n213, n209, n169, n166);
nor  g453 (n477, n185, n195, n199, n229);
xnor g454 (n481, n197, n173, n225, n232);
nand g455 (n489, n176, n230, n189, n211);
xnor g456 (n485, n165, n223, n188, n194);
xor  g457 (n486, n208, n167, n201, n224);
xor  g458 (n482, n226, n192, n210, n218);
xor  g459 (n487, n168, n193, n198, n203);
xnor g460 (n480, n231, n187, n215, n221);
not  g461 (n494, n155);
buf  g462 (n501, n156);
buf  g463 (n502, n154);
buf  g464 (n495, n481);
not  g465 (n505, n485);
buf  g466 (n497, n479);
or   g467 (n496, n487, n157);
or   g468 (n498, n484, n478, n155, n156);
xnor g469 (n500, n480, n158, n482, n157);
or   g470 (n499, n486, n155, n156);
or   g471 (n504, n157, n155, n154);
nand g472 (n503, n477, n476, n483, n157);
not  g473 (n507, n495);
buf  g474 (n515, n495);
buf  g475 (n509, n494);
not  g476 (n508, n496);
buf  g477 (n511, n494);
buf  g478 (n513, n496);
buf  g479 (n512, n496);
buf  g480 (n506, n495);
buf  g481 (n516, n495);
buf  g482 (n514, n494);
not  g483 (n510, n494);
buf  g484 (n531, n508);
not  g485 (n532, n489);
buf  g486 (n521, n507);
buf  g487 (n527, n508);
not  g488 (n523, n506);
not  g489 (n526, n506);
buf  g490 (n517, n509);
not  g491 (n518, n509);
buf  g492 (n530, n507);
not  g493 (n522, n509);
buf  g494 (n520, n509);
buf  g495 (n525, n507);
not  g496 (n519, n507);
not  g497 (n529, n506);
not  g498 (n524, n508);
or   g499 (n528, n506, n488, n508, n490);
not  g500 (n536, n497);
not  g501 (n537, n519);
not  g502 (n539, n518);
buf  g503 (n541, n500);
nor  g504 (n533, n499, n497);
nand g505 (n538, n491, n518, n500);
or   g506 (n534, n501, n498, n518);
or   g507 (n540, n499, n497, n498, n518);
xnor g508 (n535, n499, n497, n517);
nor  g509 (n543, n498, n519, n517);
and  g510 (n542, n500, n519, n499, n496);
not  g511 (n546, n503);
buf  g512 (n566, n543);
not  g513 (n564, n542);
buf  g514 (n548, n540);
not  g515 (n568, n543);
buf  g516 (n559, n504);
buf  g517 (n565, n537);
not  g518 (n553, n510);
not  g519 (n561, n503);
buf  g520 (n558, n503);
buf  g521 (n551, n505);
buf  g522 (n545, n535);
buf  g523 (n544, n541);
buf  g524 (n569, n510);
buf  g525 (n560, n539);
not  g526 (n555, n511);
nand g527 (n557, n542, n501, n543);
xor  g528 (n552, n504, n539, n501, n505);
xnor g529 (n567, n511, n234, n502, n235);
xnor g530 (n547, n533, n502, n501, n504);
or   g531 (n562, n541, n504, n502, n511);
nor  g532 (n549, n540, n503, n542, n233);
xnor g533 (n563, n502, n541, n539, n534);
and  g534 (n550, n505, n536, n538, n511);
nand g535 (n554, n540, n510);
and  g536 (n556, n541, n542, n539, n505);
not  g537 (n575, n547);
buf  g538 (n585, n545);
buf  g539 (n589, n520);
buf  g540 (n572, n548);
not  g541 (n588, n520);
buf  g542 (n571, n521);
buf  g543 (n578, n547);
buf  g544 (n590, n546);
not  g545 (n576, n545);
not  g546 (n574, n520);
buf  g547 (n570, n549);
buf  g548 (n573, n548);
buf  g549 (n587, n548);
not  g550 (n580, n544);
buf  g551 (n584, n546);
buf  g552 (n581, n544);
not  g553 (n577, n548);
not  g554 (n579, n521);
or   g555 (n582, n544, n519);
or   g556 (n586, n522, n544, n545);
xnor g557 (n591, n547, n521, n520);
or   g558 (n583, n547, n546, n549);
buf  g559 (n613, n572);
buf  g560 (n596, n572);
not  g561 (n611, n570);
buf  g562 (n603, n573);
buf  g563 (n593, n574);
not  g564 (n595, n528);
not  g565 (n601, n527);
not  g566 (n614, n528);
not  g567 (n592, n528);
not  g568 (n597, n570);
not  g569 (n604, n526);
not  g570 (n608, n574);
not  g571 (n609, n523);
and  g572 (n612, n573, n525);
and  g573 (n602, n529, n570, n522, n524);
nand g574 (n598, n523, n571, n574, n573);
nand g575 (n607, n528, n573, n574, n572);
nor  g576 (n606, n525, n570, n575, n571);
nand g577 (n605, n571, n572, n575, n524);
nor  g578 (n615, n524, n529, n571, n527);
nand g579 (n610, n523, n529, n522, n526);
and  g580 (n594, n530, n524, n526);
or   g581 (n599, n525, n527, n529, n575);
nor  g582 (n600, n523, n522, n527, n575);
or   g583 (n629, n594, n236, n558, n593);
nor  g584 (n628, n597, n595, n554, n549);
xor  g585 (n637, n558, n564, n563, n592);
xor  g586 (n643, n594, n515, n557);
and  g587 (n618, n514, n595, n554);
xor  g588 (n630, n599, n564, n596, n600);
xnor g589 (n639, n562, n565, n239, n563);
xor  g590 (n640, n515, n562, n595, n592);
nor  g591 (n634, n563, n513, n554);
xnor g592 (n616, n551, n598, n600, n564);
xor  g593 (n649, n561, n557, n562, n237);
nor  g594 (n624, n514, n569, n592, n566);
nor  g595 (n617, n559, n564, n599);
nor  g596 (n632, n550, n552, n599, n566);
xnor g597 (n642, n556, n555, n563, n242);
or   g598 (n625, n566, n562, n550, n560);
nor  g599 (n648, n559, n550, n567, n568);
and  g600 (n644, n596, n561, n559, n594);
xnor g601 (n635, n555, n569, n596, n592);
nor  g602 (n631, n553, n569, n551, n243);
xnor g603 (n623, n552, n559, n240, n514);
xnor g604 (n645, n558, n568, n551, n512);
nor  g605 (n650, n569, n513, n593, n556);
xnor g606 (n641, n597, n568, n560);
and  g607 (n646, n555, n565, n552, n566);
and  g608 (n619, n512, n551, n600, n560);
or   g609 (n626, n561, n241, n554, n512);
and  g610 (n633, n244, n553, n598, n512);
xnor g611 (n621, n594, n552, n567, n513);
nor  g612 (n647, n514, n598, n567, n565);
xor  g613 (n622, n567, n597, n556, n555);
nor  g614 (n620, n553, n593, n565, n556);
nor  g615 (n638, n561, n557, n550, n598);
nand g616 (n627, n596, n553, n558, n560);
xor  g617 (n636, n549, n593, n597, n238);
xnor g618 (n652, n581, n581, n578, n623);
xnor g619 (n656, n618, n582, n577, n621);
and  g620 (n655, n622, n579, n576);
xnor g621 (n657, n580, n577, n581);
xor  g622 (n659, n582, n578, n580);
nor  g623 (n658, n624, n582, n580, n577);
xor  g624 (n651, n581, n576, n578);
xor  g625 (n654, n619, n576, n620, n616);
xor  g626 (n653, n617, n580, n579);
not  g627 (n669, n654);
buf  g628 (n667, n653);
buf  g629 (n665, n652);
not  g630 (n668, n653);
not  g631 (n679, n651);
not  g632 (n660, n654);
not  g633 (n672, n652);
buf  g634 (n671, n600);
buf  g635 (n675, n651);
buf  g636 (n673, n652);
buf  g637 (n677, n653);
not  g638 (n674, n601);
buf  g639 (n666, n601);
not  g640 (n661, n601);
buf  g641 (n662, n651);
buf  g642 (n663, n653);
not  g643 (n664, n602);
buf  g644 (n676, n654);
nor  g645 (n678, n651, n655);
xor  g646 (n670, n652, n601, n655, n654);
nor  g647 (n686, n625, n603, n660);
xnor g648 (n685, n605, n604, n603, n661);
xnor g649 (n682, n660, n604, n602, n606);
and  g650 (n680, n602, n605, n604, n661);
nand g651 (n684, n604, n606, n603, n605);
xor  g652 (n681, n627, n605, n603, n660);
xor  g653 (n683, n661, n626, n606, n602);
nand g654 (n689, n631, n632, n684, n630);
and  g655 (n688, n629, n635, n628, n636);
xor  g656 (n687, n633, n634, n685, n686);
xnor g657 (n701, n669, n689, n665, n662);
or   g658 (n691, n663, n669, n687);
or   g659 (n697, n670, n668, n666, n664);
or   g660 (n693, n668, n688, n665, n662);
xor  g661 (n698, n662, n689, n670, n666);
nor  g662 (n692, n667, n666, n687);
nor  g663 (n694, n670, n664, n667, n665);
and  g664 (n699, n662, n666, n689, n663);
xor  g665 (n690, n661, n688, n664, n669);
and  g666 (n696, n669, n688, n664, n665);
or   g667 (n700, n663, n689, n668);
nor  g668 (n695, n663, n688, n667);
nand g669 (n705, n671, n672, n673);
nand g670 (n703, n701, n672, n670);
xnor g671 (n704, n671, n673, n699);
nand g672 (n702, n671, n671, n698, n700);
nor  g673 (n707, n704, n656, n609, n608);
nand g674 (n714, n609, n585, n640, n644);
or   g675 (n719, n608, n608, n515, n584);
xor  g676 (n718, n607, n702, n583, n639);
and  g677 (n715, n705, n638, n703, n704);
nor  g678 (n712, n656, n606, n637, n607);
nand g679 (n711, n610, n583, n656, n643);
nor  g680 (n716, n656, n642, n612, n702);
xnor g681 (n717, n583, n705, n607, n611);
nor  g682 (n706, n609, n582, n611, n607);
xnor g683 (n721, n611, n608, n703, n609);
xnor g684 (n710, n516, n515, n703, n610);
nor  g685 (n709, n704, n702, n584);
xnor g686 (n720, n611, n610, n705, n702);
xnor g687 (n708, n704, n641, n703, n705);
or   g688 (n713, n584, n610, n612, n583);
not  g689 (n742, n710);
buf  g690 (n734, n706);
not  g691 (n745, n706);
not  g692 (n726, n708);
not  g693 (n747, n708);
not  g694 (n744, n711);
buf  g695 (n746, n707);
not  g696 (n727, n709);
not  g697 (n739, n707);
buf  g698 (n724, n710);
not  g699 (n735, n712);
not  g700 (n725, n706);
not  g701 (n738, n706);
not  g702 (n731, n709);
not  g703 (n736, n707);
not  g704 (n737, n711);
not  g705 (n740, n710);
buf  g706 (n730, n711);
not  g707 (n723, n712);
not  g708 (n729, n708);
buf  g709 (n741, n708);
buf  g710 (n733, n710);
buf  g711 (n728, n707);
not  g712 (n743, n711);
buf  g713 (n722, n709);
not  g714 (n732, n709);
xor  g715 (n780, n726, n741, n673);
xnor g716 (n766, n727, n461, n159, n349);
nor  g717 (n797, n736, n727, n399, n739);
xnor g718 (n807, n730, n614, n740, n376);
xnor g719 (n816, n587, n467, n746, n423);
xnor g720 (n764, n739, n585, n471, n492);
or   g721 (n753, n379, n472, n160, n587);
or   g722 (n817, n733, n417, n732, n470);
xnor g723 (n790, n462, n329, n269, n734);
or   g724 (n782, n158, n442, n273, n675);
and  g725 (n837, n254, n263, n590, n431);
nand g726 (n819, n308, n374, n403, n460);
xor  g727 (n841, n428, n742, n588, n586);
xnor g728 (n788, n388, n474, n355, n331);
and  g729 (n781, n313, n725, n372, n456);
xnor g730 (n755, n474, n464, n415, n412);
and  g731 (n750, n418, n457, n675, n470);
or   g732 (n846, n741, n731, n251, n726);
xnor g733 (n825, n395, n435, n304, n358);
and  g734 (n751, n317, n336, n407, n436);
xnor g735 (n834, n587, n275, n531, n590);
nor  g736 (n770, n250, n339, n409, n327);
nor  g737 (n773, n742, n290, n466, n738);
nand g738 (n802, n745, n475, n253);
xnor g739 (n769, n341, n159, n274, n326);
nor  g740 (n848, n258, n448, n724, n314);
or   g741 (n811, n402, n398, n743, n255);
and  g742 (n795, n366, n383, n247, n282);
nand g743 (n784, n674, n345, n588, n731);
nor  g744 (n789, n324, n724, n293, n734);
or   g745 (n844, n265, n350, n472, n449);
xor  g746 (n815, n472, n722, n411, n249);
xor  g747 (n809, n260, n318, n424, n724);
xnor g748 (n783, n733, n419, n737, n248);
nor  g749 (n775, n335, n433, n322, n589);
nor  g750 (n771, n320, n421, n730, n347);
and  g751 (n785, n729, n158, n441, n740);
xor  g752 (n831, n729, n590, n589, n312);
xor  g753 (n828, n444, n286, n256, n453);
nor  g754 (n799, n408, n585, n613, n473);
and  g755 (n761, n612, n728, n735, n473);
and  g756 (n787, n300, n723, n385, n724);
nand g757 (n804, n741, n261, n160, n739);
and  g758 (n835, n471, n343, n532, n591);
xor  g759 (n774, n746, n381, n736, n323);
xor  g760 (n845, n726, n295, n737, n272);
xor  g761 (n779, n392, n373, n731, n727);
xor  g762 (n801, n420, n612, n732, n585);
xnor g763 (n850, n746, n405, n438, n397);
or   g764 (n810, n369, n287, n736, n303);
nor  g765 (n759, n382, n736, n340, n354);
or   g766 (n752, n674, n396, n586, n365);
nor  g767 (n760, n443, n613, n380, n262);
xnor g768 (n793, n288, n743, n451, n298);
xnor g769 (n765, n532, n257, n353, n375);
xor  g770 (n851, n384, n416, n732, n531);
nor  g771 (n824, n296, n377, n734, n268);
nor  g772 (n756, n747, n352, n738, n252);
xor  g773 (n826, n281, n731, n342, n474);
and  g774 (n822, n276, n446, n725, n469);
nor  g775 (n832, n746, n356, n306, n271);
or   g776 (n827, n390, n738, n472, n413);
nor  g777 (n758, n739, n733, n246, n292);
nand g778 (n805, n159, n589, n289, n735);
nand g779 (n767, n532, n730, n747, n325);
and  g780 (n838, n470, n674, n530, n744);
xnor g781 (n768, n725, n294, n676, n359);
nor  g782 (n763, n722, n455, n264, n747);
xnor g783 (n791, n410, n588, n330, n307);
or   g784 (n833, n590, n742, n722, n591);
and  g785 (n820, n302, n465, n471, n735);
xnor g786 (n748, n473, n531, n351, n160);
xor  g787 (n849, n645, n309, n328, n371);
or   g788 (n840, n743, n440, n474, n277);
or   g789 (n754, n463, n744, n266, n613);
xor  g790 (n772, n728, n725, n473, n425);
nor  g791 (n806, n723, n338, n445, n422);
nor  g792 (n762, n297, n737, n728, n259);
xnor g793 (n808, n439, n387, n319, n613);
and  g794 (n839, n738, n735, n159, n301);
xor  g795 (n792, n344, n400, n391, n311);
or   g796 (n794, n740, n727, n316, n279);
nor  g797 (n778, n468, n426, n434, n406);
or   g798 (n796, n429, n722, n675, n432);
nor  g799 (n818, n733, n437, n321, n742);
and  g800 (n803, n732, n357, n530, n283);
and  g801 (n800, n745, n346, n530, n452);
nand g802 (n798, n404, n299, n378, n160);
and  g803 (n776, n734, n587, n245, n723);
or   g804 (n823, n348, n740, n459, n393);
or   g805 (n786, n744, n267, n728, n729);
xnor g806 (n821, n367, n532, n729, n414);
xnor g807 (n749, n386, n447, n270, n744);
and  g808 (n842, n285, n360, n743, n745);
and  g809 (n829, n747, n370, n586, n458);
and  g810 (n812, n401, n280, n361, n589);
and  g811 (n814, n531, n368, n586, n475);
xnor g812 (n843, n394, n745, n315, n450);
nor  g813 (n777, n334, n332, n364, n284);
nor  g814 (n813, n427, n737, n291, n675);
xor  g815 (n847, n730, n278, n362, n310);
xor  g816 (n830, n389, n363, n726, n454);
nand g817 (n836, n333, n158, n337, n430);
and  g818 (n757, n674, n588, n305, n723);
and  g819 (n854, n713, n754);
xor  g820 (n852, n714, n716, n713, n750);
xnor g821 (n855, n753, n749, n715, n712);
and  g822 (n858, n717, n716, n714, n713);
xor  g823 (n857, n716, n715, n717);
xnor g824 (n853, n715, n748, n714, n716);
xor  g825 (n859, n755, n752, n717);
nor  g826 (n856, n714, n751, n713, n712);
xor  g827 (n863, n718, n719, n591, n721);
xor  g828 (n864, n591, n721, n855);
nor  g829 (n860, n855, n719);
nor  g830 (n861, n718, n720, n853, n855);
xnor g831 (n865, n854, n720, n721);
xnor g832 (n862, n852, n718, n720);
or   g833 (n866, n757, n759, n766, n762);
xnor g834 (n867, n863, n862, n768, n770);
xnor g835 (n870, n758, n769, n865, n861);
or   g836 (n869, n767, n760, n764, n763);
nor  g837 (n868, n765, n756, n761, n864);
and  g838 (n876, n789, n867, n779, n787);
and  g839 (n890, n797, n783, n784, n788);
and  g840 (n882, n870, n830, n866, n828);
nor  g841 (n883, n870, n804, n829, n816);
nand g842 (n874, n802, n867, n866);
xor  g843 (n871, n818, n793, n819, n782);
or   g844 (n887, n869, n866, n868, n780);
xor  g845 (n879, n800, n795, n796, n869);
nand g846 (n886, n791, n812, n823, n870);
and  g847 (n885, n867, n868, n821);
xnor g848 (n878, n799, n810, n808, n794);
or   g849 (n881, n775, n869, n820, n814);
xor  g850 (n880, n869, n807, n822, n785);
xnor g851 (n875, n773, n798, n781, n774);
nor  g852 (n884, n824, n790, n866, n803);
nand g853 (n877, n815, n827, n771, n811);
xnor g854 (n872, n813, n778, n801, n868);
nand g855 (n889, n817, n825, n809, n772);
xnor g856 (n888, n792, n805, n777, n776);
or   g857 (n873, n786, n826, n806, n870);
nand g858 (n907, n837, n850, n856, n843);
xnor g859 (n903, n678, n887, n832, n657);
xor  g860 (n928, n840, n834, n657, n516);
nand g861 (n902, n659, n848, n858, n658);
and  g862 (n892, n658, n887, n882, n614);
or   g863 (n926, n835, n851, n882, n847);
nand g864 (n904, n843, n849, n887, n879);
or   g865 (n906, n881, n844, n883, n677);
and  g866 (n909, n856, n659, n615, n475);
nand g867 (n893, n657, n886, n648, n888);
xor  g868 (n921, n840, n840, n659, n646);
nor  g869 (n923, n841, n885, n872, n850);
or   g870 (n918, n833, n881, n851, n859);
or   g871 (n898, n845, n878, n676, n842);
nand g872 (n894, n880, n859, n849, n841);
xnor g873 (n934, n846, n844, n881, n885);
and  g874 (n891, n846, n848, n856, n658);
xnor g875 (n905, n886, n846, n890, n883);
or   g876 (n930, n880, n881, n839, n858);
nand g877 (n915, n615, n838, n845, n884);
nand g878 (n927, n848, n851, n884);
xor  g879 (n908, n879, n845, n871, n840);
nand g880 (n901, n882, n858, n873);
nand g881 (n931, n888, n890, n847, n883);
nand g882 (n929, n676, n831, n847, n845);
and  g883 (n911, n676, n659, n857, n877);
nand g884 (n920, n883, n882, n890, n842);
nand g885 (n895, n844, n842, n857, n884);
or   g886 (n913, n677, n649, n859, n847);
xnor g887 (n912, n851, n677, n678, n679);
nand g888 (n925, n887, n876, n890, n889);
or   g889 (n924, n889, n647, n839, n855);
nor  g890 (n916, n842, n850, n886, n889);
xnor g891 (n914, n493, n885, n857, n657);
xnor g892 (n900, n857, n849, n516, n678);
xor  g893 (n897, n856, n874, n516, n614);
nor  g894 (n919, n886, n679, n880, n615);
or   g895 (n933, n879, n614, n885, n679);
xor  g896 (n896, n839, n888, n849, n880);
and  g897 (n910, n679, n888, n848, n650);
xnor g898 (n922, n843, n875, n841, n836);
nand g899 (n932, n859, n841, n844, n846);
nand g900 (n917, n678, n658, n889, n850);
nor  g901 (n899, n677, n615, n839, n843);
nand g902 (n939, n931, n891, n933, n929);
nand g903 (n937, n906, n927, n896, n893);
xnor g904 (n935, n923, n932, n897, n904);
xnor g905 (n940, n912, n902, n921, n908);
or   g906 (n942, n913, n895, n918, n920);
and  g907 (n943, n930, n911, n907, n901);
xor  g908 (n936, n892, n925, n915, n934);
nor  g909 (n941, n924, n894, n899, n898);
xor  g910 (n944, n903, n916, n905, n909);
nor  g911 (n945, n900, n914, n917, n928);
nor  g912 (n938, n910, n922, n919, n926);
endmodule
