

module Stat_2000_227
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1359,
  n1419,
  n1325,
  n1408,
  n1365,
  n1394,
  n1405,
  n1399,
  n1380,
  n1363,
  n1389,
  n1313,
  n1308,
  n1367,
  n1348,
  n1366,
  n1407,
  n1396,
  n2022,
  n2024,
  n2021,
  n2029,
  n2028,
  n2023,
  n2025,
  n2026,
  n2027,
  n2030,
  n2019,
  n2020,
  n2032,
  n2031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1359;
  output n1419;
  output n1325;
  output n1408;
  output n1365;
  output n1394;
  output n1405;
  output n1399;
  output n1380;
  output n1363;
  output n1389;
  output n1313;
  output n1308;
  output n1367;
  output n1348;
  output n1366;
  output n1407;
  output n1396;
  output n2022;
  output n2024;
  output n2021;
  output n2029;
  output n2028;
  output n2023;
  output n2025;
  output n2026;
  output n2027;
  output n2030;
  output n2019;
  output n2020;
  output n2032;
  output n2031;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1364;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1395;
  wire n1397;
  wire n1398;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1406;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n57,
    n8
  );


  buf
  g1
  (
    n64,
    n1
  );


  not
  g2
  (
    n42,
    n2
  );


  buf
  g3
  (
    n67,
    n4
  );


  buf
  g4
  (
    n60,
    n7
  );


  not
  g5
  (
    n48,
    n1
  );


  not
  g6
  (
    n46,
    n1
  );


  buf
  g7
  (
    n37,
    n2
  );


  buf
  g8
  (
    n63,
    n7
  );


  buf
  g9
  (
    n33,
    n5
  );


  not
  g10
  (
    n34,
    n6
  );


  not
  g11
  (
    n54,
    n6
  );


  not
  g12
  (
    n50,
    n8
  );


  not
  g13
  (
    n66,
    n9
  );


  not
  g14
  (
    n56,
    n9
  );


  buf
  g15
  (
    n36,
    n2
  );


  not
  g16
  (
    n68,
    n9
  );


  not
  g17
  (
    n58,
    n4
  );


  not
  g18
  (
    n53,
    n8
  );


  buf
  g19
  (
    n52,
    n7
  );


  not
  g20
  (
    n39,
    n5
  );


  not
  g21
  (
    n49,
    n4
  );


  buf
  g22
  (
    n51,
    n3
  );


  buf
  g23
  (
    n43,
    n3
  );


  buf
  g24
  (
    n38,
    n1
  );


  buf
  g25
  (
    n62,
    n6
  );


  buf
  g26
  (
    n65,
    n7
  );


  buf
  g27
  (
    n44,
    n2
  );


  buf
  g28
  (
    n35,
    n6
  );


  buf
  g29
  (
    n61,
    n5
  );


  not
  g30
  (
    n41,
    n5
  );


  buf
  g31
  (
    n47,
    n9
  );


  not
  g32
  (
    n40,
    n4
  );


  not
  g33
  (
    n55,
    n8
  );


  buf
  g34
  (
    n45,
    n3
  );


  not
  g35
  (
    n59,
    n3
  );


  buf
  g36
  (
    n148,
    n51
  );


  not
  g37
  (
    n132,
    n39
  );


  buf
  g38
  (
    n104,
    n41
  );


  buf
  g39
  (
    n163,
    n36
  );


  not
  g40
  (
    n183,
    n48
  );


  buf
  g41
  (
    n128,
    n61
  );


  not
  g42
  (
    n140,
    n58
  );


  buf
  g43
  (
    n113,
    n52
  );


  buf
  g44
  (
    n76,
    n42
  );


  not
  g45
  (
    n151,
    n48
  );


  not
  g46
  (
    n185,
    n59
  );


  not
  g47
  (
    n155,
    n34
  );


  buf
  g48
  (
    n139,
    n33
  );


  buf
  g49
  (
    n170,
    n63
  );


  not
  g50
  (
    n180,
    n60
  );


  buf
  g51
  (
    n95,
    n61
  );


  not
  g52
  (
    n172,
    n52
  );


  buf
  g53
  (
    n111,
    n51
  );


  buf
  g54
  (
    n77,
    n63
  );


  buf
  g55
  (
    n102,
    n57
  );


  buf
  g56
  (
    n190,
    n54
  );


  buf
  g57
  (
    n78,
    n46
  );


  not
  g58
  (
    n165,
    n51
  );


  not
  g59
  (
    n130,
    n45
  );


  not
  g60
  (
    n81,
    n41
  );


  buf
  g61
  (
    n84,
    n36
  );


  not
  g62
  (
    n97,
    n43
  );


  not
  g63
  (
    n193,
    n54
  );


  not
  g64
  (
    n120,
    n46
  );


  not
  g65
  (
    n150,
    n45
  );


  buf
  g66
  (
    n94,
    n55
  );


  buf
  g67
  (
    n116,
    n49
  );


  buf
  g68
  (
    n149,
    n61
  );


  not
  g69
  (
    n74,
    n55
  );


  not
  g70
  (
    n160,
    n50
  );


  buf
  g71
  (
    n112,
    n35
  );


  buf
  g72
  (
    n184,
    n43
  );


  not
  g73
  (
    n106,
    n40
  );


  buf
  g74
  (
    n101,
    n60
  );


  not
  g75
  (
    n147,
    n42
  );


  not
  g76
  (
    n88,
    n37
  );


  buf
  g77
  (
    n131,
    n49
  );


  buf
  g78
  (
    n173,
    n50
  );


  not
  g79
  (
    n91,
    n42
  );


  buf
  g80
  (
    n100,
    n35
  );


  buf
  g81
  (
    n152,
    n44
  );


  buf
  g82
  (
    n98,
    n59
  );


  not
  g83
  (
    n189,
    n39
  );


  not
  g84
  (
    n82,
    n51
  );


  not
  g85
  (
    n187,
    n62
  );


  not
  g86
  (
    n182,
    n44
  );


  not
  g87
  (
    n157,
    n62
  );


  not
  g88
  (
    n127,
    n59
  );


  not
  g89
  (
    n166,
    n62
  );


  not
  g90
  (
    n79,
    n53
  );


  not
  g91
  (
    n123,
    n53
  );


  not
  g92
  (
    n137,
    n47
  );


  not
  g93
  (
    n192,
    n40
  );


  buf
  g94
  (
    n118,
    n56
  );


  buf
  g95
  (
    n121,
    n46
  );


  buf
  g96
  (
    n134,
    n48
  );


  buf
  g97
  (
    n161,
    n47
  );


  not
  g98
  (
    n73,
    n60
  );


  buf
  g99
  (
    n129,
    n34
  );


  not
  g100
  (
    n186,
    n53
  );


  not
  g101
  (
    n144,
    n42
  );


  buf
  g102
  (
    n85,
    n34
  );


  not
  g103
  (
    n110,
    n58
  );


  not
  g104
  (
    n158,
    n36
  );


  not
  g105
  (
    n136,
    n52
  );


  buf
  g106
  (
    n105,
    n43
  );


  buf
  g107
  (
    n75,
    n38
  );


  not
  g108
  (
    n174,
    n52
  );


  buf
  g109
  (
    n176,
    n44
  );


  not
  g110
  (
    n175,
    n39
  );


  buf
  g111
  (
    n159,
    n45
  );


  buf
  g112
  (
    n162,
    n58
  );


  not
  g113
  (
    n154,
    n59
  );


  not
  g114
  (
    n145,
    n38
  );


  not
  g115
  (
    n171,
    n56
  );


  buf
  g116
  (
    n117,
    n60
  );


  not
  g117
  (
    n86,
    n40
  );


  buf
  g118
  (
    n133,
    n35
  );


  buf
  g119
  (
    n167,
    n57
  );


  buf
  g120
  (
    n90,
    n37
  );


  buf
  g121
  (
    n177,
    n62
  );


  buf
  g122
  (
    n181,
    n35
  );


  not
  g123
  (
    n80,
    n53
  );


  not
  g124
  (
    n103,
    n56
  );


  not
  g125
  (
    n146,
    n56
  );


  buf
  g126
  (
    n178,
    n50
  );


  not
  g127
  (
    n87,
    n37
  );


  not
  g128
  (
    n93,
    n33
  );


  not
  g129
  (
    n143,
    n45
  );


  buf
  g130
  (
    n142,
    n55
  );


  buf
  g131
  (
    n71,
    n54
  );


  buf
  g132
  (
    n191,
    n47
  );


  not
  g133
  (
    n107,
    n40
  );


  not
  g134
  (
    n89,
    n43
  );


  not
  g135
  (
    n126,
    n63
  );


  buf
  g136
  (
    n122,
    n38
  );


  buf
  g137
  (
    n72,
    n33
  );


  buf
  g138
  (
    n135,
    n54
  );


  not
  g139
  (
    n115,
    n58
  );


  buf
  g140
  (
    n153,
    n57
  );


  not
  g141
  (
    n108,
    n38
  );


  buf
  g142
  (
    n168,
    n47
  );


  buf
  g143
  (
    n138,
    n63
  );


  not
  g144
  (
    n141,
    n49
  );


  not
  g145
  (
    n114,
    n41
  );


  not
  g146
  (
    n109,
    n64
  );


  not
  g147
  (
    n83,
    n34
  );


  buf
  g148
  (
    n96,
    n39
  );


  not
  g149
  (
    n164,
    n57
  );


  not
  g150
  (
    n119,
    n46
  );


  not
  g151
  (
    n188,
    n49
  );


  not
  g152
  (
    n124,
    n33
  );


  buf
  g153
  (
    n92,
    n61
  );


  buf
  g154
  (
    n169,
    n44
  );


  buf
  g155
  (
    n179,
    n37
  );


  buf
  g156
  (
    n156,
    n55
  );


  not
  g157
  (
    n69,
    n50
  );


  not
  g158
  (
    n70,
    n41
  );


  buf
  g159
  (
    n125,
    n48
  );


  buf
  g160
  (
    n99,
    n36
  );


  buf
  g161
  (
    n200,
    n90
  );


  not
  g162
  (
    n360,
    n75
  );


  not
  g163
  (
    n667,
    n171
  );


  buf
  g164
  (
    n660,
    n117
  );


  not
  g165
  (
    n248,
    n167
  );


  buf
  g166
  (
    n295,
    n91
  );


  buf
  g167
  (
    n212,
    n180
  );


  buf
  g168
  (
    n607,
    n187
  );


  not
  g169
  (
    n328,
    n167
  );


  not
  g170
  (
    n516,
    n143
  );


  not
  g171
  (
    n428,
    n129
  );


  not
  g172
  (
    n491,
    n171
  );


  buf
  g173
  (
    n327,
    n161
  );


  not
  g174
  (
    n333,
    n125
  );


  not
  g175
  (
    n261,
    n172
  );


  not
  g176
  (
    n269,
    n173
  );


  buf
  g177
  (
    n355,
    n134
  );


  not
  g178
  (
    n549,
    n123
  );


  not
  g179
  (
    n488,
    n160
  );


  not
  g180
  (
    n563,
    n181
  );


  not
  g181
  (
    n278,
    n78
  );


  buf
  g182
  (
    n474,
    n76
  );


  not
  g183
  (
    n394,
    n137
  );


  not
  g184
  (
    n230,
    n169
  );


  not
  g185
  (
    n338,
    n157
  );


  not
  g186
  (
    n303,
    n144
  );


  not
  g187
  (
    n460,
    n149
  );


  buf
  g188
  (
    n531,
    n92
  );


  not
  g189
  (
    n341,
    n92
  );


  not
  g190
  (
    n229,
    n159
  );


  buf
  g191
  (
    n283,
    n116
  );


  buf
  g192
  (
    n376,
    n88
  );


  buf
  g193
  (
    n464,
    n179
  );


  not
  g194
  (
    n207,
    n122
  );


  buf
  g195
  (
    n445,
    n137
  );


  not
  g196
  (
    n571,
    n79
  );


  buf
  g197
  (
    n424,
    n180
  );


  buf
  g198
  (
    n511,
    n112
  );


  not
  g199
  (
    n223,
    n130
  );


  buf
  g200
  (
    n203,
    n103
  );


  buf
  g201
  (
    n490,
    n117
  );


  not
  g202
  (
    n357,
    n91
  );


  not
  g203
  (
    n354,
    n158
  );


  buf
  g204
  (
    n621,
    n69
  );


  buf
  g205
  (
    n425,
    n154
  );


  buf
  g206
  (
    n290,
    n104
  );


  buf
  g207
  (
    n204,
    n169
  );


  not
  g208
  (
    n572,
    n124
  );


  buf
  g209
  (
    n492,
    n185
  );


  buf
  g210
  (
    n400,
    n121
  );


  not
  g211
  (
    n663,
    n147
  );


  buf
  g212
  (
    n397,
    n166
  );


  buf
  g213
  (
    n321,
    n74
  );


  not
  g214
  (
    n444,
    n134
  );


  buf
  g215
  (
    n244,
    n163
  );


  not
  g216
  (
    n661,
    n114
  );


  buf
  g217
  (
    n461,
    n146
  );


  not
  g218
  (
    n466,
    n87
  );


  not
  g219
  (
    n544,
    n118
  );


  not
  g220
  (
    n391,
    n100
  );


  buf
  g221
  (
    n503,
    n91
  );


  buf
  g222
  (
    n301,
    n89
  );


  not
  g223
  (
    n656,
    n156
  );


  buf
  g224
  (
    n545,
    n132
  );


  not
  g225
  (
    n489,
    n167
  );


  buf
  g226
  (
    n282,
    n114
  );


  buf
  g227
  (
    n206,
    n118
  );


  buf
  g228
  (
    n243,
    n79
  );


  buf
  g229
  (
    n615,
    n105
  );


  not
  g230
  (
    n408,
    n140
  );


  not
  g231
  (
    n378,
    n185
  );


  buf
  g232
  (
    n548,
    n172
  );


  not
  g233
  (
    n584,
    n174
  );


  not
  g234
  (
    n335,
    n93
  );


  not
  g235
  (
    n476,
    n166
  );


  buf
  g236
  (
    n276,
    n116
  );


  not
  g237
  (
    n440,
    n80
  );


  buf
  g238
  (
    n326,
    n158
  );


  buf
  g239
  (
    n628,
    n77
  );


  buf
  g240
  (
    n277,
    n166
  );


  buf
  g241
  (
    n366,
    n126
  );


  not
  g242
  (
    n219,
    n106
  );


  not
  g243
  (
    n310,
    n171
  );


  not
  g244
  (
    n271,
    n160
  );


  buf
  g245
  (
    n604,
    n113
  );


  not
  g246
  (
    n518,
    n123
  );


  not
  g247
  (
    n555,
    n113
  );


  buf
  g248
  (
    n483,
    n103
  );


  not
  g249
  (
    n287,
    n174
  );


  not
  g250
  (
    n241,
    n94
  );


  not
  g251
  (
    n343,
    n168
  );


  not
  g252
  (
    n612,
    n95
  );


  not
  g253
  (
    n336,
    n70
  );


  not
  g254
  (
    n600,
    n120
  );


  buf
  g255
  (
    n666,
    n172
  );


  not
  g256
  (
    n650,
    n147
  );


  not
  g257
  (
    n358,
    n86
  );


  not
  g258
  (
    n627,
    n165
  );


  not
  g259
  (
    n245,
    n104
  );


  buf
  g260
  (
    n586,
    n71
  );


  not
  g261
  (
    n448,
    n73
  );


  not
  g262
  (
    n349,
    n133
  );


  not
  g263
  (
    n232,
    n107
  );


  buf
  g264
  (
    n469,
    n180
  );


  not
  g265
  (
    n579,
    n99
  );


  not
  g266
  (
    n569,
    n181
  );


  not
  g267
  (
    n194,
    n106
  );


  buf
  g268
  (
    n673,
    n76
  );


  not
  g269
  (
    n345,
    n141
  );


  buf
  g270
  (
    n657,
    n156
  );


  not
  g271
  (
    n455,
    n184
  );


  not
  g272
  (
    n538,
    n181
  );


  not
  g273
  (
    n613,
    n164
  );


  buf
  g274
  (
    n573,
    n111
  );


  not
  g275
  (
    n529,
    n126
  );


  not
  g276
  (
    n433,
    n186
  );


  not
  g277
  (
    n286,
    n87
  );


  not
  g278
  (
    n554,
    n114
  );


  buf
  g279
  (
    n553,
    n102
  );


  buf
  g280
  (
    n668,
    n184
  );


  buf
  g281
  (
    n582,
    n153
  );


  buf
  g282
  (
    n356,
    n125
  );


  not
  g283
  (
    n551,
    n139
  );


  not
  g284
  (
    n405,
    n128
  );


  buf
  g285
  (
    n399,
    n137
  );


  not
  g286
  (
    n209,
    n149
  );


  buf
  g287
  (
    n198,
    n86
  );


  buf
  g288
  (
    n373,
    n119
  );


  buf
  g289
  (
    n382,
    n72
  );


  not
  g290
  (
    n350,
    n175
  );


  not
  g291
  (
    n616,
    n103
  );


  not
  g292
  (
    n514,
    n182
  );


  not
  g293
  (
    n467,
    n149
  );


  buf
  g294
  (
    n452,
    n145
  );


  buf
  g295
  (
    n258,
    n99
  );


  not
  g296
  (
    n380,
    n147
  );


  not
  g297
  (
    n435,
    n108
  );


  not
  g298
  (
    n498,
    n116
  );


  not
  g299
  (
    n669,
    n109
  );


  buf
  g300
  (
    n386,
    n78
  );


  buf
  g301
  (
    n524,
    n156
  );


  buf
  g302
  (
    n462,
    n182
  );


  not
  g303
  (
    n449,
    n186
  );


  not
  g304
  (
    n426,
    n69
  );


  buf
  g305
  (
    n251,
    n78
  );


  buf
  g306
  (
    n504,
    n135
  );


  not
  g307
  (
    n395,
    n183
  );


  buf
  g308
  (
    n371,
    n176
  );


  buf
  g309
  (
    n337,
    n101
  );


  buf
  g310
  (
    n527,
    n136
  );


  buf
  g311
  (
    n329,
    n158
  );


  buf
  g312
  (
    n369,
    n96
  );


  not
  g313
  (
    n353,
    n97
  );


  buf
  g314
  (
    n617,
    n126
  );


  not
  g315
  (
    n671,
    n110
  );


  buf
  g316
  (
    n635,
    n111
  );


  buf
  g317
  (
    n332,
    n104
  );


  buf
  g318
  (
    n305,
    n127
  );


  not
  g319
  (
    KeyWire_0_1,
    n148
  );


  buf
  g320
  (
    n252,
    n100
  );


  buf
  g321
  (
    n540,
    n89
  );


  not
  g322
  (
    n228,
    n94
  );


  not
  g323
  (
    n453,
    n85
  );


  buf
  g324
  (
    n606,
    n136
  );


  buf
  g325
  (
    n331,
    n176
  );


  buf
  g326
  (
    n249,
    n178
  );


  buf
  g327
  (
    n471,
    n79
  );


  buf
  g328
  (
    n609,
    n94
  );


  not
  g329
  (
    n562,
    n132
  );


  buf
  g330
  (
    n221,
    n122
  );


  not
  g331
  (
    n642,
    n170
  );


  not
  g332
  (
    n383,
    n76
  );


  not
  g333
  (
    n222,
    n164
  );


  not
  g334
  (
    n557,
    n82
  );


  buf
  g335
  (
    n523,
    n73
  );


  not
  g336
  (
    n525,
    n83
  );


  not
  g337
  (
    n259,
    n99
  );


  not
  g338
  (
    n289,
    n154
  );


  not
  g339
  (
    n316,
    n108
  );


  not
  g340
  (
    n575,
    n135
  );


  buf
  g341
  (
    n659,
    n157
  );


  buf
  g342
  (
    n239,
    n161
  );


  not
  g343
  (
    n567,
    n168
  );


  buf
  g344
  (
    n414,
    n70
  );


  not
  g345
  (
    n296,
    n82
  );


  not
  g346
  (
    n497,
    n177
  );


  buf
  g347
  (
    n533,
    n181
  );


  buf
  g348
  (
    n412,
    n110
  );


  not
  g349
  (
    n318,
    n185
  );


  buf
  g350
  (
    n547,
    n101
  );


  buf
  g351
  (
    n284,
    n150
  );


  buf
  g352
  (
    n515,
    n134
  );


  buf
  g353
  (
    n417,
    n74
  );


  not
  g354
  (
    n441,
    n77
  );


  not
  g355
  (
    n274,
    n159
  );


  not
  g356
  (
    n570,
    n119
  );


  buf
  g357
  (
    n348,
    n74
  );


  buf
  g358
  (
    n447,
    n87
  );


  buf
  g359
  (
    n247,
    n141
  );


  buf
  g360
  (
    n298,
    n186
  );


  buf
  g361
  (
    n513,
    n76
  );


  not
  g362
  (
    n205,
    n131
  );


  not
  g363
  (
    n493,
    n84
  );


  not
  g364
  (
    n478,
    n138
  );


  buf
  g365
  (
    n392,
    n75
  );


  not
  g366
  (
    n377,
    n98
  );


  not
  g367
  (
    n655,
    n141
  );


  not
  g368
  (
    n208,
    n141
  );


  buf
  g369
  (
    n402,
    n112
  );


  buf
  g370
  (
    n591,
    n113
  );


  buf
  g371
  (
    n398,
    n153
  );


  not
  g372
  (
    n450,
    n124
  );


  not
  g373
  (
    n262,
    n178
  );


  not
  g374
  (
    n431,
    n169
  );


  not
  g375
  (
    n599,
    n164
  );


  not
  g376
  (
    n368,
    n168
  );


  not
  g377
  (
    n451,
    n119
  );


  buf
  g378
  (
    n534,
    n144
  );


  not
  g379
  (
    n496,
    n140
  );


  buf
  g380
  (
    n566,
    n94
  );


  buf
  g381
  (
    n434,
    n99
  );


  not
  g382
  (
    n253,
    n95
  );


  not
  g383
  (
    n519,
    n179
  );


  not
  g384
  (
    n201,
    n120
  );


  buf
  g385
  (
    n564,
    n130
  );


  buf
  g386
  (
    n611,
    n128
  );


  not
  g387
  (
    n304,
    n73
  );


  not
  g388
  (
    n587,
    n160
  );


  buf
  g389
  (
    n257,
    n148
  );


  buf
  g390
  (
    n280,
    n165
  );


  buf
  g391
  (
    n231,
    n154
  );


  not
  g392
  (
    n535,
    n172
  );


  not
  g393
  (
    n281,
    n152
  );


  not
  g394
  (
    n324,
    n145
  );


  buf
  g395
  (
    n499,
    n109
  );


  not
  g396
  (
    n211,
    n95
  );


  not
  g397
  (
    n308,
    n79
  );


  not
  g398
  (
    n639,
    n152
  );


  not
  g399
  (
    n517,
    n128
  );


  not
  g400
  (
    n279,
    n89
  );


  not
  g401
  (
    n552,
    n72
  );


  not
  g402
  (
    n605,
    n175
  );


  not
  g403
  (
    n658,
    n188
  );


  not
  g404
  (
    n456,
    n97
  );


  not
  g405
  (
    n590,
    n102
  );


  buf
  g406
  (
    n352,
    n187
  );


  not
  g407
  (
    n665,
    n165
  );


  buf
  g408
  (
    n215,
    n110
  );


  not
  g409
  (
    n195,
    n157
  );


  not
  g410
  (
    n236,
    n90
  );


  buf
  g411
  (
    n644,
    n127
  );


  buf
  g412
  (
    n422,
    n121
  );


  not
  g413
  (
    n472,
    n170
  );


  buf
  g414
  (
    n311,
    n96
  );


  not
  g415
  (
    n463,
    n186
  );


  buf
  g416
  (
    n265,
    n187
  );


  buf
  g417
  (
    n521,
    n122
  );


  buf
  g418
  (
    n436,
    n140
  );


  not
  g419
  (
    n646,
    n188
  );


  buf
  g420
  (
    n539,
    n182
  );


  not
  g421
  (
    n411,
    n75
  );


  buf
  g422
  (
    n583,
    n142
  );


  buf
  g423
  (
    n415,
    n163
  );


  buf
  g424
  (
    n292,
    n105
  );


  buf
  g425
  (
    n420,
    n83
  );


  buf
  g426
  (
    n662,
    n110
  );


  buf
  g427
  (
    n477,
    n149
  );


  not
  g428
  (
    n625,
    n182
  );


  not
  g429
  (
    n294,
    n82
  );


  buf
  g430
  (
    n409,
    n143
  );


  not
  g431
  (
    n473,
    n139
  );


  buf
  g432
  (
    n626,
    n144
  );


  buf
  g433
  (
    n390,
    n130
  );


  buf
  g434
  (
    n220,
    n70
  );


  not
  g435
  (
    n217,
    n146
  );


  not
  g436
  (
    n254,
    n155
  );


  buf
  g437
  (
    n647,
    n85
  );


  buf
  g438
  (
    n481,
    n97
  );


  buf
  g439
  (
    n593,
    n174
  );


  not
  g440
  (
    n653,
    n140
  );


  buf
  g441
  (
    n559,
    n118
  );


  not
  g442
  (
    n260,
    n169
  );


  buf
  g443
  (
    n214,
    n74
  );


  buf
  g444
  (
    n196,
    n171
  );


  buf
  g445
  (
    n300,
    n73
  );


  not
  g446
  (
    n293,
    n81
  );


  not
  g447
  (
    n313,
    n142
  );


  buf
  g448
  (
    n375,
    n107
  );


  not
  g449
  (
    n597,
    n88
  );


  buf
  g450
  (
    n307,
    n183
  );


  not
  g451
  (
    n317,
    n115
  );


  buf
  g452
  (
    n225,
    n125
  );


  buf
  g453
  (
    n309,
    n134
  );


  not
  g454
  (
    n407,
    n162
  );


  buf
  g455
  (
    n631,
    n111
  );


  buf
  g456
  (
    n643,
    n162
  );


  buf
  g457
  (
    n624,
    n150
  );


  buf
  g458
  (
    n528,
    n109
  );


  buf
  g459
  (
    n351,
    n86
  );


  not
  g460
  (
    n306,
    n84
  );


  not
  g461
  (
    n379,
    n78
  );


  buf
  g462
  (
    n648,
    n167
  );


  buf
  g463
  (
    n581,
    n152
  );


  not
  g464
  (
    n346,
    n83
  );


  buf
  g465
  (
    n413,
    n152
  );


  not
  g466
  (
    n427,
    n80
  );


  not
  g467
  (
    n442,
    n123
  );


  not
  g468
  (
    n510,
    n173
  );


  not
  g469
  (
    n410,
    n183
  );


  not
  g470
  (
    n325,
    n111
  );


  buf
  g471
  (
    n598,
    n162
  );


  not
  g472
  (
    n601,
    n153
  );


  not
  g473
  (
    n637,
    n176
  );


  buf
  g474
  (
    n363,
    n139
  );


  buf
  g475
  (
    n302,
    n75
  );


  buf
  g476
  (
    n330,
    n116
  );


  buf
  g477
  (
    n319,
    n177
  );


  not
  g478
  (
    n418,
    n165
  );


  not
  g479
  (
    n640,
    n154
  );


  not
  g480
  (
    n250,
    n183
  );


  buf
  g481
  (
    n482,
    n170
  );


  not
  g482
  (
    n256,
    n101
  );


  not
  g483
  (
    n585,
    n129
  );


  buf
  g484
  (
    n384,
    n102
  );


  buf
  g485
  (
    n588,
    n95
  );


  not
  g486
  (
    n416,
    n127
  );


  not
  g487
  (
    n213,
    n115
  );


  buf
  g488
  (
    n266,
    n129
  );


  buf
  g489
  (
    n475,
    n131
  );


  buf
  g490
  (
    n288,
    n71
  );


  not
  g491
  (
    n505,
    n187
  );


  not
  g492
  (
    n234,
    n131
  );


  not
  g493
  (
    n634,
    n142
  );


  not
  g494
  (
    n226,
    n151
  );


  not
  g495
  (
    n273,
    n184
  );


  not
  g496
  (
    n340,
    n112
  );


  not
  g497
  (
    n596,
    n174
  );


  not
  g498
  (
    n501,
    n91
  );


  not
  g499
  (
    n536,
    n119
  );


  not
  g500
  (
    n361,
    n161
  );


  not
  g501
  (
    n320,
    n123
  );


  buf
  g502
  (
    n419,
    n166
  );


  not
  g503
  (
    n314,
    n93
  );


  not
  g504
  (
    n439,
    n144
  );


  not
  g505
  (
    n502,
    n179
  );


  not
  g506
  (
    n430,
    n109
  );


  not
  g507
  (
    n454,
    n178
  );


  buf
  g508
  (
    n537,
    n104
  );


  buf
  g509
  (
    n576,
    n98
  );


  buf
  g510
  (
    n216,
    n86
  );


  buf
  g511
  (
    n423,
    n118
  );


  not
  g512
  (
    n610,
    n136
  );


  buf
  g513
  (
    n465,
    n147
  );


  buf
  g514
  (
    n556,
    n122
  );


  buf
  g515
  (
    n396,
    n163
  );


  buf
  g516
  (
    n494,
    n132
  );


  buf
  g517
  (
    n237,
    n173
  );


  not
  g518
  (
    n568,
    n170
  );


  not
  g519
  (
    n602,
    n115
  );


  not
  g520
  (
    n458,
    n146
  );


  not
  g521
  (
    n334,
    n163
  );


  buf
  g522
  (
    n509,
    n162
  );


  not
  g523
  (
    n651,
    n80
  );


  not
  g524
  (
    n297,
    n71
  );


  buf
  g525
  (
    n485,
    n132
  );


  not
  g526
  (
    n654,
    n83
  );


  buf
  g527
  (
    n470,
    n179
  );


  not
  g528
  (
    n622,
    n69
  );


  buf
  g529
  (
    n227,
    n131
  );


  buf
  g530
  (
    n370,
    n84
  );


  not
  g531
  (
    n636,
    n106
  );


  not
  g532
  (
    n242,
    n176
  );


  not
  g533
  (
    n233,
    n145
  );


  not
  g534
  (
    n393,
    n126
  );


  buf
  g535
  (
    n255,
    n112
  );


  buf
  g536
  (
    n620,
    n92
  );


  buf
  g537
  (
    n339,
    n173
  );


  not
  g538
  (
    n558,
    n97
  );


  not
  g539
  (
    n438,
    n150
  );


  not
  g540
  (
    n486,
    n69
  );


  buf
  g541
  (
    n578,
    n160
  );


  buf
  g542
  (
    n546,
    n155
  );


  buf
  g543
  (
    n672,
    n184
  );


  not
  g544
  (
    n526,
    n77
  );


  not
  g545
  (
    n291,
    n77
  );


  not
  g546
  (
    n421,
    n159
  );


  not
  g547
  (
    n389,
    n138
  );


  buf
  g548
  (
    n520,
    n138
  );


  not
  g549
  (
    n388,
    n130
  );


  not
  g550
  (
    n268,
    n177
  );


  buf
  g551
  (
    n315,
    n88
  );


  not
  g552
  (
    n618,
    n71
  );


  buf
  g553
  (
    n652,
    n81
  );


  not
  g554
  (
    n638,
    n178
  );


  not
  g555
  (
    n580,
    n106
  );


  not
  g556
  (
    n312,
    n98
  );


  not
  g557
  (
    n614,
    n72
  );


  buf
  g558
  (
    n322,
    n127
  );


  buf
  g559
  (
    n574,
    n142
  );


  not
  g560
  (
    n630,
    n143
  );


  not
  g561
  (
    n344,
    n96
  );


  not
  g562
  (
    n238,
    n129
  );


  buf
  g563
  (
    n565,
    n151
  );


  not
  g564
  (
    n364,
    n72
  );


  not
  g565
  (
    n495,
    n100
  );


  not
  g566
  (
    n619,
    n107
  );


  not
  g567
  (
    n365,
    n177
  );


  buf
  g568
  (
    n542,
    n180
  );


  not
  g569
  (
    n210,
    n136
  );


  buf
  g570
  (
    n272,
    n84
  );


  buf
  g571
  (
    n595,
    n137
  );


  buf
  g572
  (
    n506,
    n135
  );


  buf
  g573
  (
    n632,
    n175
  );


  buf
  g574
  (
    n374,
    n81
  );


  buf
  g575
  (
    n432,
    n105
  );


  not
  g576
  (
    n664,
    n156
  );


  not
  g577
  (
    n670,
    n90
  );


  buf
  g578
  (
    n246,
    n159
  );


  buf
  g579
  (
    n459,
    n133
  );


  not
  g580
  (
    n649,
    n80
  );


  not
  g581
  (
    n385,
    n185
  );


  not
  g582
  (
    n508,
    n85
  );


  not
  g583
  (
    n347,
    n155
  );


  buf
  g584
  (
    n468,
    n89
  );


  buf
  g585
  (
    n641,
    n146
  );


  not
  g586
  (
    n264,
    n108
  );


  not
  g587
  (
    n629,
    n108
  );


  not
  g588
  (
    n530,
    n103
  );


  buf
  g589
  (
    n543,
    n120
  );


  buf
  g590
  (
    n267,
    n93
  );


  not
  g591
  (
    n603,
    n133
  );


  buf
  g592
  (
    n199,
    n150
  );


  buf
  g593
  (
    n359,
    n124
  );


  not
  g594
  (
    n406,
    n138
  );


  buf
  g595
  (
    n577,
    n135
  );


  buf
  g596
  (
    n479,
    n121
  );


  buf
  g597
  (
    n263,
    n100
  );


  not
  g598
  (
    n197,
    n164
  );


  buf
  g599
  (
    n429,
    n120
  );


  buf
  g600
  (
    n323,
    n139
  );


  not
  g601
  (
    n457,
    n113
  );


  buf
  g602
  (
    n608,
    n82
  );


  not
  g603
  (
    n561,
    n98
  );


  not
  g604
  (
    n594,
    n125
  );


  buf
  g605
  (
    n372,
    n124
  );


  buf
  g606
  (
    n522,
    n90
  );


  not
  g607
  (
    n270,
    n107
  );


  not
  g608
  (
    n403,
    n175
  );


  not
  g609
  (
    n592,
    n128
  );


  buf
  g610
  (
    n387,
    n188
  );


  not
  g611
  (
    n240,
    n81
  );


  not
  g612
  (
    n550,
    n105
  );


  not
  g613
  (
    n401,
    n85
  );


  buf
  g614
  (
    n512,
    n145
  );


  not
  g615
  (
    n560,
    n70
  );


  buf
  g616
  (
    n487,
    n87
  );


  not
  g617
  (
    n224,
    n117
  );


  buf
  g618
  (
    n532,
    n158
  );


  buf
  g619
  (
    n541,
    n121
  );


  not
  g620
  (
    n235,
    n115
  );


  not
  g621
  (
    n645,
    n102
  );


  not
  g622
  (
    n342,
    n148
  );


  buf
  g623
  (
    n285,
    n117
  );


  not
  g624
  (
    n437,
    n157
  );


  buf
  g625
  (
    n443,
    n143
  );


  buf
  g626
  (
    n633,
    n161
  );


  buf
  g627
  (
    n507,
    n101
  );


  not
  g628
  (
    n589,
    n88
  );


  buf
  g629
  (
    n202,
    n92
  );


  buf
  g630
  (
    n480,
    n148
  );


  not
  g631
  (
    n218,
    n151
  );


  buf
  g632
  (
    n484,
    n93
  );


  buf
  g633
  (
    n299,
    n114
  );


  buf
  g634
  (
    n623,
    n188
  );


  not
  g635
  (
    n362,
    n151
  );


  buf
  g636
  (
    n500,
    n155
  );


  buf
  g637
  (
    n381,
    n168
  );


  not
  g638
  (
    n275,
    n96
  );


  not
  g639
  (
    n367,
    n153
  );


  not
  g640
  (
    n404,
    n133
  );


  buf
  g641
  (
    n1204,
    n662
  );


  buf
  g642
  (
    n1147,
    n616
  );


  not
  g643
  (
    n1073,
    n488
  );


  not
  g644
  (
    KeyWire_0_0,
    n662
  );


  not
  g645
  (
    n1067,
    n631
  );


  buf
  g646
  (
    n1274,
    n326
  );


  buf
  g647
  (
    n880,
    n379
  );


  buf
  g648
  (
    n1223,
    n441
  );


  not
  g649
  (
    n1183,
    n510
  );


  not
  g650
  (
    n775,
    n431
  );


  not
  g651
  (
    n822,
    n255
  );


  not
  g652
  (
    n1170,
    n302
  );


  buf
  g653
  (
    n1031,
    n285
  );


  buf
  g654
  (
    n942,
    n269
  );


  buf
  g655
  (
    n732,
    n491
  );


  buf
  g656
  (
    n953,
    n259
  );


  buf
  g657
  (
    n800,
    n489
  );


  not
  g658
  (
    n1015,
    n292
  );


  not
  g659
  (
    n864,
    n248
  );


  buf
  g660
  (
    n1236,
    n583
  );


  buf
  g661
  (
    n1174,
    n370
  );


  buf
  g662
  (
    n714,
    n643
  );


  buf
  g663
  (
    n674,
    n593
  );


  buf
  g664
  (
    n1024,
    n545
  );


  not
  g665
  (
    n939,
    n327
  );


  buf
  g666
  (
    n769,
    n562
  );


  not
  g667
  (
    n934,
    n488
  );


  buf
  g668
  (
    n1007,
    n537
  );


  buf
  g669
  (
    n1190,
    n360
  );


  not
  g670
  (
    n1257,
    n547
  );


  not
  g671
  (
    n761,
    n251
  );


  buf
  g672
  (
    n831,
    n272
  );


  not
  g673
  (
    n998,
    n602
  );


  buf
  g674
  (
    n947,
    n530
  );


  not
  g675
  (
    n1180,
    n385
  );


  not
  g676
  (
    n794,
    n481
  );


  not
  g677
  (
    n1193,
    n353
  );


  buf
  g678
  (
    n772,
    n252
  );


  buf
  g679
  (
    n1254,
    n548
  );


  not
  g680
  (
    n1019,
    n432
  );


  buf
  g681
  (
    n784,
    n432
  );


  not
  g682
  (
    n1033,
    n544
  );


  not
  g683
  (
    n1296,
    n490
  );


  buf
  g684
  (
    n1112,
    n313
  );


  buf
  g685
  (
    n811,
    n526
  );


  not
  g686
  (
    n711,
    n485
  );


  buf
  g687
  (
    n762,
    n449
  );


  buf
  g688
  (
    n684,
    n448
  );


  buf
  g689
  (
    n720,
    n483
  );


  not
  g690
  (
    n1069,
    n591
  );


  not
  g691
  (
    n861,
    n340
  );


  buf
  g692
  (
    n1277,
    n327
  );


  not
  g693
  (
    n1253,
    n585
  );


  not
  g694
  (
    n1087,
    n278
  );


  not
  g695
  (
    n1111,
    n572
  );


  not
  g696
  (
    n1049,
    n568
  );


  not
  g697
  (
    n773,
    n474
  );


  buf
  g698
  (
    n923,
    n461
  );


  not
  g699
  (
    n853,
    n212
  );


  buf
  g700
  (
    n1068,
    n619
  );


  not
  g701
  (
    n882,
    n380
  );


  not
  g702
  (
    n1238,
    n300
  );


  buf
  g703
  (
    n1187,
    n386
  );


  buf
  g704
  (
    n1098,
    n418
  );


  not
  g705
  (
    n850,
    n664
  );


  not
  g706
  (
    n1205,
    n436
  );


  buf
  g707
  (
    n852,
    n422
  );


  not
  g708
  (
    n1215,
    n533
  );


  not
  g709
  (
    n890,
    n457
  );


  buf
  g710
  (
    n685,
    n526
  );


  not
  g711
  (
    n1272,
    n531
  );


  buf
  g712
  (
    n952,
    n261
  );


  buf
  g713
  (
    n1291,
    n527
  );


  buf
  g714
  (
    n870,
    n349
  );


  not
  g715
  (
    n983,
    n366
  );


  buf
  g716
  (
    n1262,
    n550
  );


  buf
  g717
  (
    n807,
    n380
  );


  buf
  g718
  (
    n962,
    n524
  );


  not
  g719
  (
    n1000,
    n344
  );


  buf
  g720
  (
    n1138,
    n503
  );


  not
  g721
  (
    n678,
    n413
  );


  not
  g722
  (
    n957,
    n468
  );


  not
  g723
  (
    n989,
    n483
  );


  buf
  g724
  (
    n1171,
    n594
  );


  buf
  g725
  (
    n965,
    n507
  );


  not
  g726
  (
    n716,
    n308
  );


  not
  g727
  (
    n888,
    n237
  );


  not
  g728
  (
    n1284,
    n373
  );


  not
  g729
  (
    n1305,
    n307
  );


  buf
  g730
  (
    n1212,
    n576
  );


  not
  g731
  (
    n1189,
    n460
  );


  buf
  g732
  (
    n781,
    n357
  );


  not
  g733
  (
    n1036,
    n509
  );


  buf
  g734
  (
    n1157,
    n534
  );


  buf
  g735
  (
    n845,
    n618
  );


  not
  g736
  (
    n854,
    n260
  );


  buf
  g737
  (
    n1026,
    n547
  );


  not
  g738
  (
    n1139,
    n575
  );


  not
  g739
  (
    n1005,
    n548
  );


  buf
  g740
  (
    n742,
    n664
  );


  buf
  g741
  (
    n1158,
    n549
  );


  buf
  g742
  (
    n1041,
    n371
  );


  not
  g743
  (
    n760,
    n583
  );


  buf
  g744
  (
    n1125,
    n260
  );


  buf
  g745
  (
    n747,
    n552
  );


  not
  g746
  (
    n1283,
    n581
  );


  not
  g747
  (
    n1259,
    n456
  );


  not
  g748
  (
    n844,
    n396
  );


  buf
  g749
  (
    n799,
    n385
  );


  buf
  g750
  (
    n791,
    n534
  );


  not
  g751
  (
    n1050,
    n601
  );


  not
  g752
  (
    n897,
    n461
  );


  not
  g753
  (
    n839,
    n633
  );


  not
  g754
  (
    n1129,
    n226
  );


  not
  g755
  (
    n721,
    n241
  );


  not
  g756
  (
    n901,
    n419
  );


  buf
  g757
  (
    n1163,
    n546
  );


  buf
  g758
  (
    n833,
    n651
  );


  buf
  g759
  (
    n886,
    n516
  );


  not
  g760
  (
    n1270,
    n258
  );


  not
  g761
  (
    n1121,
    n498
  );


  not
  g762
  (
    n1248,
    n340
  );


  buf
  g763
  (
    n1235,
    n590
  );


  not
  g764
  (
    n697,
    n194
  );


  not
  g765
  (
    n1148,
    n561
  );


  buf
  g766
  (
    n1232,
    n359
  );


  buf
  g767
  (
    n765,
    n194
  );


  buf
  g768
  (
    n759,
    n417
  );


  buf
  g769
  (
    n1243,
    n567
  );


  not
  g770
  (
    n806,
    n433
  );


  buf
  g771
  (
    n948,
    n379
  );


  buf
  g772
  (
    n1058,
    n630
  );


  not
  g773
  (
    n702,
    n245
  );


  not
  g774
  (
    n1197,
    n350
  );


  buf
  g775
  (
    n1079,
    n355
  );


  not
  g776
  (
    n986,
    n347
  );


  buf
  g777
  (
    n1292,
    n356
  );


  not
  g778
  (
    n745,
    n497
  );


  not
  g779
  (
    n1159,
    n480
  );


  not
  g780
  (
    n744,
    n457
  );


  not
  g781
  (
    n804,
    n603
  );


  buf
  g782
  (
    n1186,
    n569
  );


  not
  g783
  (
    n676,
    n394
  );


  not
  g784
  (
    n730,
    n300
  );


  not
  g785
  (
    n900,
    n576
  );


  not
  g786
  (
    n715,
    n403
  );


  not
  g787
  (
    n1255,
    n211
  );


  buf
  g788
  (
    n988,
    n455
  );


  buf
  g789
  (
    n1208,
    n661
  );


  buf
  g790
  (
    n1293,
    n500
  );


  buf
  g791
  (
    n696,
    n555
  );


  not
  g792
  (
    n1221,
    n342
  );


  not
  g793
  (
    n1302,
    n506
  );


  buf
  g794
  (
    n894,
    n639
  );


  not
  g795
  (
    n1074,
    n580
  );


  buf
  g796
  (
    n798,
    n561
  );


  buf
  g797
  (
    n1128,
    n428
  );


  buf
  g798
  (
    n812,
    n433
  );


  not
  g799
  (
    n788,
    n202
  );


  buf
  g800
  (
    n736,
    n405
  );


  buf
  g801
  (
    n1055,
    n558
  );


  not
  g802
  (
    n891,
    n662
  );


  not
  g803
  (
    n789,
    n209
  );


  not
  g804
  (
    n1018,
    n527
  );


  buf
  g805
  (
    n825,
    n548
  );


  not
  g806
  (
    n985,
    n587
  );


  not
  g807
  (
    n677,
    n303
  );


  not
  g808
  (
    n1169,
    n382
  );


  buf
  g809
  (
    n937,
    n475
  );


  not
  g810
  (
    n940,
    n538
  );


  buf
  g811
  (
    n921,
    n326
  );


  not
  g812
  (
    n1116,
    n558
  );


  not
  g813
  (
    n733,
    n327
  );


  buf
  g814
  (
    n911,
    n605
  );


  buf
  g815
  (
    n691,
    n210
  );


  buf
  g816
  (
    n1165,
    n508
  );


  buf
  g817
  (
    n1027,
    n204
  );


  buf
  g818
  (
    n731,
    n472
  );


  buf
  g819
  (
    n1273,
    n227
  );


  buf
  g820
  (
    n680,
    n287
  );


  buf
  g821
  (
    n1130,
    n638
  );


  buf
  g822
  (
    n1135,
    n201
  );


  buf
  g823
  (
    n686,
    n278
  );


  buf
  g824
  (
    n1146,
    n436
  );


  not
  g825
  (
    n1084,
    n557
  );


  not
  g826
  (
    n776,
    n637
  );


  buf
  g827
  (
    n1249,
    n646
  );


  not
  g828
  (
    n902,
    n606
  );


  not
  g829
  (
    n840,
    n220
  );


  buf
  g830
  (
    n1075,
    n331
  );


  not
  g831
  (
    n1188,
    n393
  );


  buf
  g832
  (
    n1127,
    n320
  );


  not
  g833
  (
    n1141,
    n649
  );


  buf
  g834
  (
    n1006,
    n665
  );


  not
  g835
  (
    n827,
    n500
  );


  buf
  g836
  (
    n1251,
    n264
  );


  not
  g837
  (
    n1017,
    n612
  );


  not
  g838
  (
    n1252,
    n641
  );


  not
  g839
  (
    n1172,
    n450
  );


  not
  g840
  (
    n828,
    n446
  );


  not
  g841
  (
    n824,
    n509
  );


  not
  g842
  (
    n1306,
    n487
  );


  not
  g843
  (
    n1271,
    n614
  );


  not
  g844
  (
    n1056,
    n610
  );


  not
  g845
  (
    n838,
    n357
  );


  not
  g846
  (
    n797,
    n234
  );


  not
  g847
  (
    n914,
    n521
  );


  not
  g848
  (
    n846,
    n412
  );


  not
  g849
  (
    n1207,
    n459
  );


  buf
  g850
  (
    n991,
    n536
  );


  not
  g851
  (
    n1156,
    n218
  );


  buf
  g852
  (
    n754,
    n359
  );


  not
  g853
  (
    n1016,
    n625
  );


  not
  g854
  (
    n767,
    n393
  );


  buf
  g855
  (
    n785,
    n301
  );


  buf
  g856
  (
    n1229,
    n287
  );


  not
  g857
  (
    n735,
    n258
  );


  not
  g858
  (
    n1288,
    n508
  );


  not
  g859
  (
    n1009,
    n383
  );


  not
  g860
  (
    n1126,
    n663
  );


  buf
  g861
  (
    n866,
    n453
  );


  not
  g862
  (
    n1286,
    n508
  );


  not
  g863
  (
    n813,
    n362
  );


  not
  g864
  (
    n972,
    n646
  );


  buf
  g865
  (
    n927,
    n617
  );


  not
  g866
  (
    n1168,
    n659
  );


  not
  g867
  (
    n1118,
    n473
  );


  buf
  g868
  (
    n995,
    n570
  );


  not
  g869
  (
    n943,
    n537
  );


  not
  g870
  (
    n1195,
    n590
  );


  not
  g871
  (
    n787,
    n354
  );


  buf
  g872
  (
    n1011,
    n510
  );


  not
  g873
  (
    KeyWire_0_3,
    n532
  );


  not
  g874
  (
    n830,
    n318
  );


  not
  g875
  (
    n795,
    n554
  );


  buf
  g876
  (
    n909,
    n373
  );


  not
  g877
  (
    n1029,
    n573
  );


  buf
  g878
  (
    n722,
    n549
  );


  not
  g879
  (
    n1176,
    n467
  );


  not
  g880
  (
    n1136,
    n513
  );


  not
  g881
  (
    n1153,
    n434
  );


  buf
  g882
  (
    n1088,
    n631
  );


  buf
  g883
  (
    n1239,
    n429
  );


  buf
  g884
  (
    n1061,
    n606
  );


  not
  g885
  (
    n1131,
    n504
  );


  buf
  g886
  (
    n1103,
    n585
  );


  not
  g887
  (
    n763,
    n376
  );


  not
  g888
  (
    n757,
    n590
  );


  not
  g889
  (
    n878,
    n652
  );


  buf
  g890
  (
    n1117,
    n620
  );


  not
  g891
  (
    n933,
    n655
  );


  buf
  g892
  (
    n1295,
    n350
  );


  not
  g893
  (
    n1150,
    n641
  );


  buf
  g894
  (
    n1234,
    n529
  );


  not
  g895
  (
    n837,
    n198
  );


  not
  g896
  (
    n1053,
    n494
  );


  buf
  g897
  (
    n961,
    n435
  );


  not
  g898
  (
    n1022,
    n299
  );


  not
  g899
  (
    n1166,
    n408
  );


  buf
  g900
  (
    n1216,
    n316
  );


  not
  g901
  (
    KeyWire_0_5,
    n537
  );


  not
  g902
  (
    n1185,
    n608
  );


  not
  g903
  (
    n1267,
    n361
  );


  buf
  g904
  (
    n768,
    n536
  );


  not
  g905
  (
    n1045,
    n597
  );


  not
  g906
  (
    n774,
    n619
  );


  not
  g907
  (
    n826,
    n376
  );


  buf
  g908
  (
    n1093,
    n279
  );


  not
  g909
  (
    n930,
    n235
  );


  not
  g910
  (
    n740,
    n271
  );


  buf
  g911
  (
    n792,
    n268
  );


  buf
  g912
  (
    n1104,
    n659
  );


  not
  g913
  (
    n692,
    n552
  );


  not
  g914
  (
    n1242,
    n235
  );


  not
  g915
  (
    n750,
    n581
  );


  not
  g916
  (
    n741,
    n376
  );


  not
  g917
  (
    n949,
    n652
  );


  buf
  g918
  (
    n1012,
    n284
  );


  buf
  g919
  (
    n1108,
    n564
  );


  not
  g920
  (
    n1096,
    n451
  );


  buf
  g921
  (
    n938,
    n411
  );


  not
  g922
  (
    n867,
    n371
  );


  buf
  g923
  (
    n778,
    n493
  );


  not
  g924
  (
    n908,
    n495
  );


  buf
  g925
  (
    n1099,
    n466
  );


  buf
  g926
  (
    n1113,
    n223
  );


  buf
  g927
  (
    n782,
    n666
  );


  not
  g928
  (
    n1210,
    n584
  );


  not
  g929
  (
    n1301,
    n563
  );


  buf
  g930
  (
    n1294,
    n543
  );


  not
  g931
  (
    n910,
    n336
  );


  buf
  g932
  (
    n1278,
    n499
  );


  not
  g933
  (
    n1280,
    n575
  );


  buf
  g934
  (
    n941,
    n311
  );


  not
  g935
  (
    n1032,
    n422
  );


  not
  g936
  (
    n1155,
    n280
  );


  buf
  g937
  (
    n1137,
    n242
  );


  not
  g938
  (
    n887,
    n334
  );


  not
  g939
  (
    n699,
    n665
  );


  not
  g940
  (
    n956,
    n563
  );


  not
  g941
  (
    n1152,
    n505
  );


  not
  g942
  (
    n1192,
    n265
  );


  not
  g943
  (
    n1124,
    n497
  );


  buf
  g944
  (
    n932,
    n646
  );


  not
  g945
  (
    n1132,
    n229
  );


  not
  g946
  (
    n918,
    n221
  );


  buf
  g947
  (
    n1106,
    n567
  );


  or
  g948
  (
    n821,
    n487,
    n565
  );


  xor
  g949
  (
    n996,
    n427,
    n613,
    n642,
    n640
  );


  xnor
  g950
  (
    n1091,
    n529,
    n495,
    n580,
    n334
  );


  and
  g951
  (
    n803,
    n622,
    n375,
    n205,
    n525
  );


  nand
  g952
  (
    n1085,
    n615,
    n565,
    n457,
    n362
  );


  xor
  g953
  (
    n734,
    n625,
    n532,
    n339,
    n542
  );


  xnor
  g954
  (
    n1082,
    n227,
    n614,
    n242,
    n586
  );


  and
  g955
  (
    n1025,
    n245,
    n473,
    n656,
    n210
  );


  or
  g956
  (
    n1122,
    n421,
    n424,
    n535,
    n338
  );


  and
  g957
  (
    n977,
    n424,
    n574,
    n541,
    n324
  );


  and
  g958
  (
    n1162,
    n476,
    n597,
    n647,
    n617
  );


  or
  g959
  (
    n1244,
    n372,
    n451,
    n201,
    n540
  );


  or
  g960
  (
    n1179,
    n529,
    n463,
    n526,
    n258
  );


  and
  g961
  (
    n703,
    n312,
    n462,
    n530,
    n636
  );


  xor
  g962
  (
    n975,
    n208,
    n402,
    n454,
    n533
  );


  nand
  g963
  (
    n1037,
    n319,
    n635,
    n648,
    n580
  );


  nor
  g964
  (
    n951,
    n553,
    n348,
    n278,
    n496
  );


  or
  g965
  (
    n842,
    n356,
    n539,
    n357,
    n566
  );


  nand
  g966
  (
    n694,
    n507,
    n489,
    n562,
    n661
  );


  nand
  g967
  (
    n907,
    n621,
    n615,
    n539,
    n656
  );


  nand
  g968
  (
    n978,
    n232,
    n455,
    n238,
    n513
  );


  xor
  g969
  (
    n1047,
    n654,
    n294,
    n265,
    n414
  );


  xnor
  g970
  (
    n992,
    n216,
    n465,
    n643,
    n320
  );


  nor
  g971
  (
    n832,
    n296,
    n572,
    n281,
    n314
  );


  xor
  g972
  (
    n1028,
    n396,
    n471,
    n435,
    n264
  );


  xor
  g973
  (
    n1203,
    n663,
    n553,
    n384,
    n574
  );


  xnor
  g974
  (
    n1034,
    n607,
    n513,
    n341,
    n617
  );


  nor
  g975
  (
    n857,
    n288,
    n595,
    n637,
    n262
  );


  nand
  g976
  (
    n718,
    n522,
    n657,
    n399,
    n263
  );


  and
  g977
  (
    n805,
    n557,
    n661,
    n587,
    n406
  );


  or
  g978
  (
    n1241,
    n577,
    n427,
    n621,
    n472
  );


  xor
  g979
  (
    n979,
    n593,
    n219,
    n560,
    n259
  );


  and
  g980
  (
    n698,
    n305,
    n622,
    n498,
    n542
  );


  or
  g981
  (
    n823,
    n499,
    n337,
    n524,
    n571
  );


  xor
  g982
  (
    n871,
    n494,
    n415,
    n525,
    n523
  );


  nor
  g983
  (
    n1289,
    n374,
    n284,
    n481,
    n582
  );


  xor
  g984
  (
    n879,
    n667,
    n407,
    n316,
    n578
  );


  or
  g985
  (
    n1133,
    n213,
    n443,
    n520,
    n308
  );


  nand
  g986
  (
    n884,
    n405,
    n502,
    n601,
    n249
  );


  nor
  g987
  (
    n1281,
    n197,
    n212,
    n564,
    n341
  );


  or
  g988
  (
    n755,
    n344,
    n540,
    n616,
    n409
  );


  or
  g989
  (
    n1003,
    n416,
    n592,
    n391,
    n559
  );


  and
  g990
  (
    n1200,
    n570,
    n471,
    n220,
    n636
  );


  xor
  g991
  (
    KeyWire_0_13,
    n381,
    n618,
    n206,
    n636
  );


  xor
  g992
  (
    n1237,
    n512,
    n280,
    n629,
    n616
  );


  xnor
  g993
  (
    n1268,
    n426,
    n378,
    n507,
    n562
  );


  nor
  g994
  (
    n847,
    n377,
    n198,
    n369,
    n365
  );


  xnor
  g995
  (
    n924,
    n276,
    n640,
    n516,
    n253
  );


  or
  g996
  (
    n1102,
    n632,
    n361,
    n288,
    n245
  );


  or
  g997
  (
    n1094,
    n453,
    n386,
    n352,
    n635
  );


  xnor
  g998
  (
    n1202,
    n624,
    n414,
    n527,
    n574
  );


  or
  g999
  (
    n1046,
    n332,
    n597,
    n415,
    n544
  );


  xnor
  g1000
  (
    n958,
    n626,
    n239,
    n506,
    n627
  );


  nand
  g1001
  (
    n1266,
    n390,
    n476,
    n450,
    n647
  );


  or
  g1002
  (
    n1043,
    n390,
    n283,
    n249,
    n506
  );


  xor
  g1003
  (
    n920,
    n464,
    n528,
    n293,
    n484
  );


  nor
  g1004
  (
    n1004,
    n372,
    n465,
    n454,
    n664
  );


  nor
  g1005
  (
    n1107,
    n530,
    n639,
    n657,
    n465
  );


  xnor
  g1006
  (
    n916,
    n511,
    n223,
    n404,
    n668
  );


  or
  g1007
  (
    n877,
    n195,
    n477,
    n325,
    n575
  );


  xnor
  g1008
  (
    n849,
    n217,
    n501,
    n210,
    n459
  );


  xor
  g1009
  (
    n802,
    n346,
    n207,
    n596,
    n446
  );


  or
  g1010
  (
    n1057,
    n282,
    n292,
    n248,
    n440
  );


  xnor
  g1011
  (
    n751,
    n338,
    n516,
    n573,
    n217
  );


  xnor
  g1012
  (
    n896,
    n346,
    n631,
    n588,
    n603
  );


  and
  g1013
  (
    n1245,
    n293,
    n502,
    n215,
    n574
  );


  nand
  g1014
  (
    n1123,
    n491,
    n659,
    n242,
    n401
  );


  xor
  g1015
  (
    n1178,
    n195,
    n602,
    n598,
    n224
  );


  xor
  g1016
  (
    n841,
    n227,
    n214,
    n662,
    n234
  );


  and
  g1017
  (
    n818,
    n230,
    n218,
    n556,
    n231
  );


  and
  g1018
  (
    n967,
    n420,
    n269,
    n318,
    n215
  );


  nor
  g1019
  (
    n708,
    n428,
    n304,
    n467,
    n642
  );


  and
  g1020
  (
    n1071,
    n462,
    n272,
    n664,
    n283
  );


  xor
  g1021
  (
    n1065,
    n244,
    n600,
    n650,
    n496
  );


  and
  g1022
  (
    n860,
    n241,
    n543,
    n458,
    n304
  );


  xnor
  g1023
  (
    n1051,
    n640,
    n347,
    n433,
    n487
  );


  xor
  g1024
  (
    n1140,
    n214,
    n305,
    n228,
    n430
  );


  nand
  g1025
  (
    n1228,
    n564,
    n290,
    n307,
    n288
  );


  xnor
  g1026
  (
    n873,
    n613,
    n480,
    n651,
    n605
  );


  xor
  g1027
  (
    n1224,
    n617,
    n497,
    n246,
    n535
  );


  nor
  g1028
  (
    n1149,
    n388,
    n482,
    n598,
    n266
  );


  nor
  g1029
  (
    n1142,
    n352,
    n531,
    n292,
    n403
  );


  xor
  g1030
  (
    n1198,
    n250,
    n626,
    n651,
    n211
  );


  xnor
  g1031
  (
    n710,
    n524,
    n271,
    n360,
    n269
  );


  xor
  g1032
  (
    n1115,
    n200,
    n594,
    n367,
    n503
  );


  or
  g1033
  (
    n926,
    n594,
    n622,
    n641,
    n539
  );


  and
  g1034
  (
    n881,
    n382,
    n213,
    n592,
    n419
  );


  and
  g1035
  (
    n971,
    n667,
    n295,
    n324,
    n235
  );


  nor
  g1036
  (
    n816,
    n570,
    n351,
    n466,
    n301
  );


  and
  g1037
  (
    n1021,
    n343,
    n485,
    n569,
    n321
  );


  xnor
  g1038
  (
    n994,
    n222,
    n525,
    n440,
    n252
  );


  and
  g1039
  (
    n1039,
    n398,
    n427,
    n409,
    n544
  );


  or
  g1040
  (
    n981,
    n391,
    n632,
    n563,
    n634
  );


  or
  g1041
  (
    n898,
    n576,
    n528,
    n483,
    n253
  );


  nand
  g1042
  (
    n915,
    n445,
    n517,
    n225,
    n470
  );


  nor
  g1043
  (
    n738,
    n601,
    n642,
    n520,
    n266
  );


  and
  g1044
  (
    n1077,
    n630,
    n343,
    n541,
    n656
  );


  nor
  g1045
  (
    n817,
    n328,
    n612,
    n576,
    n444
  );


  xnor
  g1046
  (
    n683,
    n443,
    n234,
    n379,
    n349
  );


  and
  g1047
  (
    n700,
    n416,
    n440,
    n265,
    n231
  );


  nand
  g1048
  (
    n843,
    n554,
    n492,
    n238,
    n384
  );


  or
  g1049
  (
    n976,
    n665,
    n639,
    n501,
    n577
  );


  or
  g1050
  (
    n709,
    n322,
    n481,
    n639,
    n398
  );


  nor
  g1051
  (
    n1044,
    n255,
    n623,
    n587
  );


  nand
  g1052
  (
    n969,
    n332,
    n203,
    n489,
    n545
  );


  xor
  g1053
  (
    n728,
    n374,
    n513,
    n626,
    n416
  );


  xor
  g1054
  (
    n1062,
    n584,
    n231,
    n389,
    n289
  );


  nand
  g1055
  (
    n945,
    n502,
    n545,
    n546,
    n666
  );


  xnor
  g1056
  (
    n743,
    n279,
    n628,
    n203,
    n579
  );


  nand
  g1057
  (
    n1089,
    n287,
    n423,
    n552,
    n318
  );


  and
  g1058
  (
    n1191,
    n609,
    n549,
    n222,
    n610
  );


  xnor
  g1059
  (
    n1109,
    n455,
    n420,
    n607,
    n402
  );


  and
  g1060
  (
    n793,
    n658,
    n660,
    n566,
    n530
  );


  nor
  g1061
  (
    n689,
    n275,
    n511,
    n356,
    n239
  );


  xnor
  g1062
  (
    n913,
    n322,
    n631,
    n573,
    n329
  );


  xnor
  g1063
  (
    n869,
    n392,
    n325,
    n538,
    n536
  );


  nor
  g1064
  (
    n770,
    n329,
    n589,
    n644,
    n246
  );


  or
  g1065
  (
    n893,
    n567,
    n529,
    n363,
    n298
  );


  or
  g1066
  (
    n928,
    n474,
    n232,
    n374,
    n406
  );


  or
  g1067
  (
    n1164,
    n358,
    n390,
    n644,
    n490
  );


  or
  g1068
  (
    n987,
    n509,
    n510,
    n531,
    n309
  );


  xor
  g1069
  (
    n829,
    n330,
    n603,
    n550,
    n657
  );


  nor
  g1070
  (
    n1101,
    n615,
    n519,
    n448,
    n508
  );


  xor
  g1071
  (
    n705,
    n236,
    n444,
    n492,
    n611
  );


  nor
  g1072
  (
    n1260,
    n368,
    n568,
    n205,
    n605
  );


  or
  g1073
  (
    n1080,
    n666,
    n479,
    n599,
    n504
  );


  or
  g1074
  (
    n865,
    n303,
    n488,
    n425,
    n498
  );


  nand
  g1075
  (
    n1048,
    n279,
    n521,
    n533,
    n397
  );


  nor
  g1076
  (
    n858,
    n503,
    n504,
    n600,
    n247
  );


  nor
  g1077
  (
    n1086,
    n290,
    n438,
    n600,
    n451
  );


  nor
  g1078
  (
    n964,
    n226,
    n647,
    n404,
    n634
  );


  nor
  g1079
  (
    n695,
    n586,
    n604,
    n616,
    n353
  );


  xor
  g1080
  (
    n1052,
    n475,
    n493,
    n435,
    n309
  );


  xor
  g1081
  (
    n1010,
    n239,
    n645,
    n442,
    n262
  );


  xor
  g1082
  (
    n1290,
    n456,
    n445,
    n407,
    n270
  );


  xnor
  g1083
  (
    n1144,
    n406,
    n439,
    n313,
    n216
  );


  xnor
  g1084
  (
    n1298,
    n518,
    n593,
    n423,
    n408
  );


  or
  g1085
  (
    n723,
    n371,
    n609,
    n360,
    n370
  );


  and
  g1086
  (
    n999,
    n246,
    n241,
    n546,
    n355
  );


  nand
  g1087
  (
    n1184,
    n591,
    n472,
    n522,
    n314
  );


  xor
  g1088
  (
    n856,
    n335,
    n559,
    n629,
    n200
  );


  or
  g1089
  (
    n906,
    n620,
    n468,
    n375,
    n667
  );


  nor
  g1090
  (
    n1275,
    n467,
    n436,
    n524,
    n586
  );


  xnor
  g1091
  (
    n1240,
    n389,
    n577,
    n237,
    n589
  );


  and
  g1092
  (
    n727,
    n658,
    n302,
    n291,
    n648
  );


  nor
  g1093
  (
    n790,
    n654,
    n375,
    n306,
    n476
  );


  nand
  g1094
  (
    n968,
    n233,
    n640,
    n614,
    n295
  );


  or
  g1095
  (
    n1120,
    n250,
    n447,
    n251,
    n648
  );


  xnor
  g1096
  (
    n779,
    n553,
    n518,
    n495,
    n470
  );


  xor
  g1097
  (
    n859,
    n470,
    n458,
    n229,
    n273
  );


  and
  g1098
  (
    n820,
    n583,
    n607,
    n599,
    n262
  );


  nor
  g1099
  (
    n1160,
    n211,
    n257,
    n196,
    n395
  );


  xnor
  g1100
  (
    n931,
    n315,
    n633,
    n500,
    n654
  );


  xor
  g1101
  (
    n681,
    n502,
    n625,
    n547,
    n453
  );


  nor
  g1102
  (
    n1269,
    n571,
    n326,
    n342,
    n652
  );


  or
  g1103
  (
    n1219,
    n335,
    n447,
    n229,
    n532
  );


  nor
  g1104
  (
    n835,
    n209,
    n209,
    n256,
    n604
  );


  nor
  g1105
  (
    n726,
    n517,
    n348,
    n388,
    n395
  );


  and
  g1106
  (
    n980,
    n535,
    n303,
    n491,
    n512
  );


  or
  g1107
  (
    n868,
    n382,
    n422,
    n385,
    n541
  );


  xnor
  g1108
  (
    n693,
    n215,
    n638,
    n421,
    n297
  );


  nor
  g1109
  (
    n737,
    n222,
    n543,
    n459,
    n412
  );


  nand
  g1110
  (
    n758,
    n207,
    n660,
    n523,
    n315
  );


  xnor
  g1111
  (
    n1217,
    n514,
    n638,
    n458,
    n238
  );


  nor
  g1112
  (
    n1173,
    n598,
    n236,
    n311,
    n558
  );


  or
  g1113
  (
    n724,
    n243,
    n346,
    n333,
    n214
  );


  or
  g1114
  (
    n1285,
    n487,
    n264,
    n256,
    n551
  );


  nor
  g1115
  (
    n1070,
    n466,
    n635,
    n663,
    n282
  );


  xor
  g1116
  (
    n706,
    n352,
    n620,
    n545,
    n413
  );


  nor
  g1117
  (
    n1035,
    n339,
    n399,
    n198,
    n197
  );


  nand
  g1118
  (
    n766,
    n381,
    n469,
    n417,
    n637
  );


  and
  g1119
  (
    n1211,
    n368,
    n590,
    n283,
    n627
  );


  xnor
  g1120
  (
    n936,
    n329,
    n270,
    n551,
    n354
  );


  xnor
  g1121
  (
    n1276,
    n469,
    n650,
    n626,
    n212
  );


  and
  g1122
  (
    n1233,
    n366,
    n527,
    n522,
    n606
  );


  or
  g1123
  (
    n717,
    n392,
    n557,
    n645,
    n471
  );


  nand
  g1124
  (
    n1076,
    n525,
    n349,
    n655,
    n537
  );


  and
  g1125
  (
    n780,
    n341,
    n253,
    n217,
    n409
  );


  and
  g1126
  (
    n1090,
    n539,
    n478,
    n595,
    n582
  );


  xnor
  g1127
  (
    n912,
    n598,
    n339,
    n514,
    n237
  );


  nand
  g1128
  (
    n810,
    n332,
    n263,
    n257,
    n522
  );


  and
  g1129
  (
    n771,
    n503,
    n653,
    n331,
    n420
  );


  xnor
  g1130
  (
    n1078,
    n547,
    n397,
    n314,
    n496
  );


  and
  g1131
  (
    n1063,
    n500,
    n532,
    n490,
    n542
  );


  or
  g1132
  (
    n917,
    n649,
    n606,
    n568,
    n267
  );


  nand
  g1133
  (
    n929,
    n304,
    n634,
    n504,
    n610
  );


  xnor
  g1134
  (
    n752,
    n270,
    n347,
    n251,
    n591
  );


  nand
  g1135
  (
    n1002,
    n443,
    n306,
    n589,
    n659
  );


  xnor
  g1136
  (
    n1227,
    n200,
    n228,
    n225,
    n540
  );


  nor
  g1137
  (
    n713,
    n660,
    n280,
    n232,
    n515
  );


  nor
  g1138
  (
    n834,
    n653,
    n423,
    n493,
    n482
  );


  or
  g1139
  (
    n707,
    n611,
    n308,
    n244,
    n560
  );


  xor
  g1140
  (
    n1054,
    n515,
    n650,
    n431,
    n534
  );


  nor
  g1141
  (
    n960,
    n597,
    n483,
    n560,
    n413
  );


  or
  g1142
  (
    n1110,
    n315,
    n351,
    n604,
    n286
  );


  and
  g1143
  (
    n1299,
    n400,
    n337,
    n646,
    n355
  );


  nor
  g1144
  (
    n1161,
    n464,
    n494,
    n381,
    n387
  );


  xor
  g1145
  (
    n1175,
    n260,
    n498,
    n521,
    n195
  );


  xor
  g1146
  (
    n756,
    n310,
    n515,
    n311,
    n600
  );


  and
  g1147
  (
    n1100,
    n577,
    n221,
    n199,
    n444
  );


  or
  g1148
  (
    n970,
    n437,
    n328,
    n221,
    n225
  );


  and
  g1149
  (
    n872,
    n439,
    n594,
    n383,
    n549
  );


  nor
  g1150
  (
    n1226,
    n307,
    n401,
    n516,
    n561
  );


  nand
  g1151
  (
    n863,
    n384,
    n634,
    n243,
    n538
  );


  and
  g1152
  (
    n899,
    n573,
    n492,
    n336,
    n319
  );


  xor
  g1153
  (
    n712,
    n223,
    n592,
    n257,
    n452
  );


  xnor
  g1154
  (
    n749,
    n410,
    n219,
    n555,
    n660
  );


  or
  g1155
  (
    n984,
    n644,
    n507,
    n296,
    n541
  );


  or
  g1156
  (
    n959,
    n557,
    n570,
    n480,
    n236
  );


  or
  g1157
  (
    n1038,
    n430,
    n358,
    n528,
    n563
  );


  xnor
  g1158
  (
    KeyWire_0_9,
    n250,
    n395,
    n201,
    n578
  );


  and
  g1159
  (
    n1279,
    n625,
    n254,
    n521,
    n648
  );


  and
  g1160
  (
    n704,
    n627,
    n194,
    n448,
    n266
  );


  xnor
  g1161
  (
    n719,
    n407,
    n367,
    n589,
    n274
  );


  and
  g1162
  (
    n801,
    n559,
    n197,
    n437,
    n377
  );


  xor
  g1163
  (
    n876,
    n658,
    n593,
    n560,
    n431
  );


  xnor
  g1164
  (
    n1300,
    n285,
    n544,
    n401,
    n585
  );


  xor
  g1165
  (
    n883,
    n608,
    n555,
    n484,
    n567
  );


  and
  g1166
  (
    n1119,
    n556,
    n474,
    n566,
    n249
  );


  nor
  g1167
  (
    n950,
    n581,
    n542,
    n636,
    n267
  );


  or
  g1168
  (
    n1167,
    n477,
    n628,
    n603,
    n526
  );


  nor
  g1169
  (
    n1040,
    n400,
    n312,
    n515,
    n389
  );


  nand
  g1170
  (
    n1023,
    n338,
    n643,
    n322,
    n632
  );


  nor
  g1171
  (
    n796,
    n571,
    n365,
    n437,
    n647
  );


  and
  g1172
  (
    n1097,
    n538,
    n601,
    n226,
    n482
  );


  xor
  g1173
  (
    n725,
    n452,
    n429,
    n216,
    n599
  );


  xnor
  g1174
  (
    n1134,
    n334,
    n224,
    n272,
    n312
  );


  xnor
  g1175
  (
    n1247,
    n536,
    n452,
    n313,
    n403
  );


  xor
  g1176
  (
    n1209,
    n386,
    n321,
    n377,
    n621
  );


  nand
  g1177
  (
    n851,
    n387,
    n240,
    n464,
    n319
  );


  xnor
  g1178
  (
    n903,
    n276,
    n333,
    n495,
    n584
  );


  xor
  g1179
  (
    n1145,
    n438,
    n316,
    n587,
    n410
  );


  xnor
  g1180
  (
    n889,
    n275,
    n337,
    n551,
    n494
  );


  or
  g1181
  (
    n1114,
    n579,
    n578,
    n552,
    n460
  );


  nor
  g1182
  (
    n954,
    n364,
    n613,
    n259,
    n233
  );


  and
  g1183
  (
    n836,
    n298,
    n614,
    n441,
    n657
  );


  nor
  g1184
  (
    n922,
    n628,
    n432,
    n310,
    n429
  );


  and
  g1185
  (
    n748,
    n393,
    n363,
    n203,
    n523
  );


  or
  g1186
  (
    n777,
    n290,
    n608,
    n419,
    n641
  );


  or
  g1187
  (
    n815,
    n535,
    n665,
    n588,
    n348
  );


  and
  g1188
  (
    n1042,
    n445,
    n363,
    n405,
    n196
  );


  xor
  g1189
  (
    n679,
    n629,
    n533,
    n492,
    n294
  );


  or
  g1190
  (
    n855,
    n276,
    n298,
    n596,
    n421
  );


  nor
  g1191
  (
    n1066,
    n378,
    n565,
    n543
  );


  xor
  g1192
  (
    n1081,
    n621,
    n268,
    n309,
    n302
  );


  xor
  g1193
  (
    n1287,
    n633,
    n612,
    n463,
    n486
  );


  xor
  g1194
  (
    n966,
    n497,
    n398,
    n450,
    n619
  );


  nand
  g1195
  (
    n687,
    n428,
    n323,
    n592,
    n568
  );


  or
  g1196
  (
    n753,
    n218,
    n638,
    n449,
    n252
  );


  or
  g1197
  (
    n1264,
    n628,
    n208,
    n425,
    n330
  );


  or
  g1198
  (
    n1013,
    n528,
    n281,
    n369,
    n284
  );


  nand
  g1199
  (
    n809,
    n499,
    n637,
    n324,
    n299
  );


  nor
  g1200
  (
    n997,
    n642,
    n645,
    n305,
    n478
  );


  and
  g1201
  (
    n990,
    n282,
    n268,
    n359,
    n501
  );


  and
  g1202
  (
    n955,
    n248,
    n206,
    n604,
    n486
  );


  xor
  g1203
  (
    n1014,
    n566,
    n512,
    n317,
    n571
  );


  xor
  g1204
  (
    n1256,
    n442,
    n596,
    n572,
    n294
  );


  xnor
  g1205
  (
    n1220,
    n556,
    n418,
    n651,
    n479
  );


  and
  g1206
  (
    n1230,
    n297,
    n514,
    n486,
    n582
  );


  xor
  g1207
  (
    n1231,
    n523,
    n364,
    n372,
    n417
  );


  xnor
  g1208
  (
    n786,
    n618,
    n373,
    n654,
    n519
  );


  nor
  g1209
  (
    n1154,
    n475,
    n383,
    n402,
    n623
  );


  xnor
  g1210
  (
    n1143,
    n430,
    n345,
    n354,
    n666
  );


  xnor
  g1211
  (
    n1095,
    n286,
    n342,
    n425,
    n202
  );


  nand
  g1212
  (
    n1263,
    n622,
    n220,
    n564,
    n244
  );


  xor
  g1213
  (
    n885,
    n653,
    n396,
    n485,
    n608
  );


  xor
  g1214
  (
    n701,
    n439,
    n602,
    n496
  );


  nand
  g1215
  (
    n1265,
    n519,
    n387,
    n649,
    n572
  );


  or
  g1216
  (
    n1282,
    n579,
    n473,
    n620,
    n551
  );


  nor
  g1217
  (
    n1303,
    n478,
    n520,
    n291,
    n412
  );


  xor
  g1218
  (
    n904,
    n584,
    n619,
    n205,
    n643
  );


  xor
  g1219
  (
    n848,
    n331,
    n358,
    n414,
    n596
  );


  or
  g1220
  (
    n1258,
    n335,
    n548,
    n463,
    n493
  );


  xnor
  g1221
  (
    n1206,
    n350,
    n267,
    n394,
    n295
  );


  and
  g1222
  (
    n1199,
    n306,
    n505,
    n661,
    n461
  );


  xor
  g1223
  (
    n1225,
    n399,
    n449,
    n207,
    n580
  );


  nand
  g1224
  (
    n1072,
    n477,
    n658,
    n274,
    n514
  );


  xor
  g1225
  (
    n892,
    n196,
    n274,
    n208,
    n578
  );


  nor
  g1226
  (
    n1177,
    n456,
    n519,
    n273,
    n479
  );


  nor
  g1227
  (
    n935,
    n366,
    n599,
    n289,
    n362
  );


  nand
  g1228
  (
    n1196,
    n273,
    n635,
    n650,
    n663
  );


  or
  g1229
  (
    n982,
    n554,
    n394,
    n489,
    n441
  );


  nor
  g1230
  (
    n819,
    n369,
    n345,
    n275,
    n228
  );


  xor
  g1231
  (
    n1020,
    n240,
    n581,
    n410,
    n645
  );


  xor
  g1232
  (
    n963,
    n501,
    n325,
    n404,
    n277
  );


  xor
  g1233
  (
    n974,
    n591,
    n505,
    n585,
    n468
  );


  nor
  g1234
  (
    n690,
    n368,
    n286,
    n615,
    n323
  );


  and
  g1235
  (
    n814,
    n630,
    n534,
    n199,
    n484
  );


  xor
  g1236
  (
    n973,
    n277,
    n595,
    n353,
    n378
  );


  nand
  g1237
  (
    n1304,
    n301,
    n240,
    n609,
    n575
  );


  and
  g1238
  (
    n946,
    n562,
    n462,
    n219,
    n388
  );


  nor
  g1239
  (
    n783,
    n520,
    n469,
    n300,
    n655
  );


  xor
  g1240
  (
    n1214,
    n488,
    n293,
    n365,
    n484
  );


  or
  g1241
  (
    n925,
    n649,
    n559,
    n460,
    n490
  );


  nand
  g1242
  (
    n1008,
    n263,
    n632,
    n391,
    n446
  );


  xnor
  g1243
  (
    n874,
    n408,
    n442,
    n434,
    n328
  );


  xor
  g1244
  (
    n688,
    n340,
    n509,
    n624,
    n482
  );


  nor
  g1245
  (
    n1064,
    n296,
    n254,
    n285,
    n202
  );


  nor
  g1246
  (
    n1105,
    n411,
    n361,
    n629,
    n281
  );


  or
  g1247
  (
    n1297,
    n555,
    n644,
    n392,
    n518
  );


  and
  g1248
  (
    n1261,
    n511,
    n204,
    n553,
    n582
  );


  xor
  g1249
  (
    n895,
    n230,
    n561,
    n618,
    n554
  );


  xor
  g1250
  (
    n1030,
    n299,
    n485,
    n247,
    n310
  );


  and
  g1251
  (
    n808,
    n655,
    n486,
    n605,
    n344
  );


  xor
  g1252
  (
    n1092,
    n277,
    n297,
    n517,
    n511
  );


  nor
  g1253
  (
    n944,
    n424,
    n595,
    n336,
    n438
  );


  and
  g1254
  (
    n875,
    n512,
    n579,
    n330,
    n633
  );


  nor
  g1255
  (
    n1218,
    n204,
    n623,
    n627,
    n426
  );


  and
  g1256
  (
    n764,
    n556,
    n323,
    n317,
    n247
  );


  nand
  g1257
  (
    n1246,
    n367,
    n351,
    n611,
    n447
  );


  xnor
  g1258
  (
    n1060,
    n558,
    n426,
    n540,
    n454
  );


  nand
  g1259
  (
    n1001,
    n434,
    n652,
    n624,
    n233
  );


  and
  g1260
  (
    n729,
    n499,
    n255,
    n291,
    n317
  );


  and
  g1261
  (
    n1222,
    n611,
    n320,
    n415,
    n199
  );


  nand
  g1262
  (
    n682,
    n370,
    n491,
    n612,
    n380
  );


  nand
  g1263
  (
    n905,
    n256,
    n550,
    n243,
    n506
  );


  xor
  g1264
  (
    n675,
    n343,
    n230,
    n289,
    n411
  );


  xnor
  g1265
  (
    n1181,
    n588,
    n546,
    n364,
    n518
  );


  nor
  g1266
  (
    n1059,
    n656,
    n624,
    n224,
    n418
  );


  and
  g1267
  (
    n746,
    n345,
    n254,
    n531,
    n653
  );


  nand
  g1268
  (
    n1194,
    n588,
    n321,
    n510,
    n569
  );


  and
  g1269
  (
    n1213,
    n667,
    n397,
    n505,
    n213
  );


  nand
  g1270
  (
    n993,
    n569,
    n550,
    n517,
    n271
  );


  nand
  g1271
  (
    n919,
    n609,
    n610,
    n400,
    n630
  );


  xnor
  g1272
  (
    n1250,
    n261,
    n607,
    n613,
    n206
  );


  or
  g1273
  (
    n739,
    n333,
    n583,
    n261,
    n586
  );


  nand
  g1274
  (
    n1387,
    n1035,
    n1008,
    n889,
    n851
  );


  and
  g1275
  (
    n1321,
    n908,
    n676,
    n1144,
    n1190
  );


  or
  g1276
  (
    n1360,
    n795,
    n785,
    n801,
    n1033
  );


  nand
  g1277
  (
    n1423,
    n1101,
    n996,
    n997,
    n1169
  );


  and
  g1278
  (
    n1372,
    n727,
    n780,
    n1106,
    n781
  );


  xor
  g1279
  (
    n1431,
    n755,
    n1052,
    n933,
    n1181
  );


  xor
  g1280
  (
    n1370,
    n721,
    n811,
    n765,
    n715
  );


  nor
  g1281
  (
    n1369,
    n698,
    n834,
    n748,
    n965
  );


  nor
  g1282
  (
    n1402,
    n1125,
    n799,
    n1166,
    n1150
  );


  nor
  g1283
  (
    n1361,
    n978,
    n1107,
    n722,
    n754
  );


  or
  g1284
  (
    n1343,
    n1063,
    n905,
    n1177,
    n869
  );


  nand
  g1285
  (
    n1324,
    n890,
    n1149,
    n880,
    n803
  );


  nand
  g1286
  (
    n1359,
    n1090,
    n903,
    n1045,
    n995
  );


  xor
  g1287
  (
    n1331,
    n981,
    n777,
    n720,
    n1104
  );


  and
  g1288
  (
    n1334,
    n974,
    n1119,
    n952,
    n861
  );


  xor
  g1289
  (
    n1325,
    n929,
    n1178,
    n1188,
    n967
  );


  nand
  g1290
  (
    n1404,
    n953,
    n912,
    n973,
    n787
  );


  or
  g1291
  (
    n1437,
    n977,
    n1088,
    n691,
    n984
  );


  or
  g1292
  (
    n1337,
    n1124,
    n959,
    n1185,
    n1162
  );


  or
  g1293
  (
    n1385,
    n769,
    n1015,
    n1157,
    n809
  );


  xnor
  g1294
  (
    n1340,
    n700,
    n876,
    n778,
    n786
  );


  xor
  g1295
  (
    n1384,
    n1198,
    n773,
    n1002,
    n800
  );


  or
  g1296
  (
    n1418,
    n897,
    n838,
    n1103,
    n1203
  );


  xnor
  g1297
  (
    n1414,
    n979,
    n687,
    n1174,
    n716
  );


  or
  g1298
  (
    n1347,
    n1086,
    n839,
    n1018,
    n1006
  );


  nor
  g1299
  (
    n1427,
    n775,
    n848,
    n1175,
    n833
  );


  and
  g1300
  (
    n1394,
    n919,
    n1095,
    n988,
    n759
  );


  and
  g1301
  (
    n1438,
    n1154,
    n925,
    n793,
    n751
  );


  and
  g1302
  (
    n1326,
    n1102,
    n852,
    n1099,
    n990
  );


  or
  g1303
  (
    n1401,
    n961,
    n744,
    n1130,
    n1011
  );


  and
  g1304
  (
    n1426,
    n900,
    n766,
    n746,
    n872
  );


  or
  g1305
  (
    n1390,
    n709,
    n918,
    n1205,
    n937
  );


  nand
  g1306
  (
    n1311,
    n854,
    n936,
    n960,
    n914
  );


  nor
  g1307
  (
    n1417,
    n1009,
    n1065,
    n899,
    n845
  );


  xnor
  g1308
  (
    n1318,
    n949,
    n1056,
    n913,
    n926
  );


  xnor
  g1309
  (
    n1429,
    n1025,
    n1084,
    n734,
    n843
  );


  nor
  g1310
  (
    n1351,
    n1014,
    n794,
    n837,
    n817
  );


  or
  g1311
  (
    n1395,
    n946,
    n901,
    n878,
    n1127
  );


  xor
  g1312
  (
    n1408,
    n1078,
    n868,
    n860,
    n823
  );


  and
  g1313
  (
    n1368,
    n761,
    n699,
    n1165,
    n1044
  );


  nor
  g1314
  (
    n1333,
    n1028,
    n694,
    n808,
    n742
  );


  xnor
  g1315
  (
    n1435,
    n948,
    n877,
    n713,
    n920
  );


  and
  g1316
  (
    n1422,
    n1022,
    n941,
    n1168,
    n1030
  );


  xor
  g1317
  (
    n1355,
    n940,
    n688,
    n681,
    n1024
  );


  nand
  g1318
  (
    n1350,
    n1046,
    n782,
    n832,
    n856
  );


  and
  g1319
  (
    n1400,
    n1121,
    n1069,
    n682,
    n1191
  );


  nand
  g1320
  (
    n1354,
    n1094,
    n745,
    n1032,
    n791
  );


  xnor
  g1321
  (
    n1389,
    n1019,
    n911,
    n675,
    n693
  );


  and
  g1322
  (
    n1412,
    n760,
    n772,
    n1079,
    n1055
  );


  xnor
  g1323
  (
    n1439,
    n1036,
    n708,
    n707,
    n870
  );


  and
  g1324
  (
    n1348,
    n1195,
    n1058,
    n1005,
    n942
  );


  and
  g1325
  (
    n1339,
    n1096,
    n1135,
    n1012,
    n1139
  );


  xor
  g1326
  (
    n1344,
    n1070,
    n739,
    n1117,
    n726
  );


  nand
  g1327
  (
    n1425,
    n762,
    n714,
    n1161,
    n1097
  );


  nand
  g1328
  (
    n1378,
    n1176,
    n1129,
    n1179,
    n767
  );


  xor
  g1329
  (
    n1397,
    n1192,
    n758,
    n821,
    n686
  );


  nor
  g1330
  (
    n1317,
    n874,
    n1141,
    n1077,
    n902
  );


  xnor
  g1331
  (
    n1399,
    n898,
    n969,
    n1193,
    n805
  );


  nor
  g1332
  (
    n1428,
    n887,
    n1093,
    n1082,
    n704
  );


  xnor
  g1333
  (
    n1380,
    n1145,
    n958,
    n830,
    n1120
  );


  nand
  g1334
  (
    n1433,
    n740,
    n999,
    n696,
    n951
  );


  or
  g1335
  (
    n1379,
    n944,
    n964,
    n807,
    n1039
  );


  and
  g1336
  (
    n1349,
    n1142,
    n1118,
    n883,
    n757
  );


  xnor
  g1337
  (
    n1329,
    n1110,
    n895,
    n1187,
    n894
  );


  and
  g1338
  (
    n1430,
    n994,
    n1051,
    n678,
    n1076
  );


  nand
  g1339
  (
    n1403,
    n982,
    n975,
    n692,
    n892
  );


  nor
  g1340
  (
    n1320,
    n886,
    n683,
    n989,
    n1038
  );


  nor
  g1341
  (
    n1367,
    n1074,
    n737,
    n863,
    n966
  );


  nand
  g1342
  (
    n1406,
    n1001,
    n1000,
    n1137,
    n827
  );


  and
  g1343
  (
    n1352,
    n888,
    n1010,
    n702,
    n935
  );


  nor
  g1344
  (
    n1328,
    n1172,
    n1072,
    n1043,
    n1153
  );


  nand
  g1345
  (
    n1420,
    n938,
    n836,
    n1048,
    n743
  );


  nor
  g1346
  (
    n1377,
    n738,
    n904,
    n906,
    n1171
  );


  xnor
  g1347
  (
    n1407,
    n1136,
    n840,
    n701,
    n1059
  );


  and
  g1348
  (
    n1312,
    n985,
    n1004,
    n1021,
    n814
  );


  or
  g1349
  (
    n1313,
    n689,
    n828,
    n1003,
    n818
  );


  nand
  g1350
  (
    n1410,
    n865,
    n790,
    n789,
    n1123
  );


  nand
  g1351
  (
    n1436,
    n1204,
    n1112,
    n719,
    n1116
  );


  xnor
  g1352
  (
    n1373,
    n695,
    n1156,
    n764,
    n1049
  );


  or
  g1353
  (
    n1366,
    n857,
    n813,
    n1054,
    n932
  );


  nand
  g1354
  (
    n1323,
    n1023,
    n939,
    n806,
    n690
  );


  nand
  g1355
  (
    n1388,
    n1183,
    n879,
    n776,
    n1068
  );


  and
  g1356
  (
    n1382,
    n835,
    n788,
    n991,
    n1133
  );


  xnor
  g1357
  (
    n1332,
    n752,
    n712,
    n1199,
    n923
  );


  xnor
  g1358
  (
    n1358,
    n674,
    n1131,
    n916,
    n1189
  );


  and
  g1359
  (
    n1346,
    n822,
    n1031,
    n1053,
    n749
  );


  nor
  g1360
  (
    n1357,
    n987,
    n921,
    n1075,
    n680
  );


  xnor
  g1361
  (
    n1413,
    n1115,
    n797,
    n1186,
    n972
  );


  xnor
  g1362
  (
    n1322,
    n1138,
    n980,
    n1151,
    n1085
  );


  nor
  g1363
  (
    n1335,
    n779,
    n710,
    n774,
    n1066
  );


  or
  g1364
  (
    n1396,
    n1146,
    n1060,
    n677,
    n829
  );


  nand
  g1365
  (
    n1307,
    n1184,
    n1197,
    n810,
    n1122
  );


  or
  g1366
  (
    n1381,
    n1167,
    n1170,
    n842,
    n763
  );


  and
  g1367
  (
    n1386,
    n1100,
    n697,
    n873,
    n1108
  );


  nor
  g1368
  (
    n1336,
    n922,
    n907,
    n893,
    n846
  );


  nor
  g1369
  (
    n1375,
    n957,
    n1113,
    n867,
    n986
  );


  xor
  g1370
  (
    n1392,
    n1109,
    n825,
    n705,
    n849
  );


  xnor
  g1371
  (
    n1393,
    n1182,
    n1062,
    n956,
    n1041
  );


  or
  g1372
  (
    n1341,
    n1147,
    n1134,
    n924,
    n768
  );


  and
  g1373
  (
    n1308,
    n750,
    n819,
    n1201,
    n882
  );


  nor
  g1374
  (
    n1416,
    n753,
    n1020,
    n816,
    n862
  );


  nand
  g1375
  (
    n1314,
    n1126,
    n1037,
    n812,
    n934
  );


  or
  g1376
  (
    n1310,
    n1029,
    n1026,
    n1180,
    n864
  );


  or
  g1377
  (
    n1316,
    n844,
    n1089,
    n1061,
    n1111
  );


  or
  g1378
  (
    n1365,
    n747,
    n885,
    n976,
    n815
  );


  or
  g1379
  (
    n1345,
    n729,
    n1105,
    n733,
    n1158
  );


  nor
  g1380
  (
    n1371,
    n1091,
    n928,
    n1027,
    n1071
  );


  nand
  g1381
  (
    n1424,
    n1160,
    n855,
    n728,
    n1114
  );


  xnor
  g1382
  (
    n1309,
    n820,
    n871,
    n968,
    n1163
  );


  xor
  g1383
  (
    n1376,
    n884,
    n947,
    n826,
    n943
  );


  nor
  g1384
  (
    n1364,
    n998,
    n684,
    n1057,
    n756
  );


  or
  g1385
  (
    n1432,
    n804,
    n917,
    n910,
    n1098
  );


  and
  g1386
  (
    n1391,
    n770,
    n1047,
    n1007,
    n792
  );


  nor
  g1387
  (
    n1315,
    n927,
    n1132,
    n1155,
    n1140
  );


  nand
  g1388
  (
    n1419,
    n703,
    n711,
    n881,
    n824
  );


  and
  g1389
  (
    n1353,
    n741,
    n679,
    n1128,
    n718
  );


  nor
  g1390
  (
    n1330,
    n1196,
    n1092,
    n1200,
    n963
  );


  xnor
  g1391
  (
    n1374,
    n970,
    n850,
    n1159,
    n1202
  );


  nand
  g1392
  (
    n1434,
    n1016,
    n1017,
    n930,
    n1081
  );


  xor
  g1393
  (
    n1319,
    n841,
    n796,
    n993,
    n802
  );


  nor
  g1394
  (
    n1383,
    n866,
    n847,
    n706,
    n1067
  );


  xor
  g1395
  (
    n1421,
    n771,
    n945,
    n1173,
    n1073
  );


  and
  g1396
  (
    n1363,
    n1064,
    n950,
    n915,
    n831
  );


  or
  g1397
  (
    n1398,
    n955,
    n723,
    n731,
    n1083
  );


  or
  g1398
  (
    n1405,
    n962,
    n1042,
    n730,
    n732
  );


  xor
  g1399
  (
    n1362,
    n859,
    n1087,
    n725,
    n1148
  );


  xnor
  g1400
  (
    n1411,
    n853,
    n1040,
    n1164,
    n1080
  );


  nor
  g1401
  (
    n1415,
    n784,
    n798,
    n1013,
    n1034
  );


  and
  g1402
  (
    n1356,
    n992,
    n875,
    n1152,
    n896
  );


  or
  g1403
  (
    n1342,
    n736,
    n954,
    n983,
    n891
  );


  nor
  g1404
  (
    n1327,
    n783,
    n717,
    n858,
    n1050
  );


  nand
  g1405
  (
    n1409,
    n1194,
    n931,
    n685,
    n1143
  );


  xnor
  g1406
  (
    n1338,
    n735,
    n724,
    n909,
    n971
  );


  not
  g1407
  (
    n1445,
    n1316
  );


  not
  g1408
  (
    n1450,
    n1313
  );


  buf
  g1409
  (
    n1448,
    n1318
  );


  buf
  g1410
  (
    n1453,
    n1315
  );


  buf
  g1411
  (
    n1447,
    n1321
  );


  buf
  g1412
  (
    n1454,
    n1314
  );


  not
  g1413
  (
    n1441,
    n1319
  );


  buf
  g1414
  (
    n1452,
    n1312
  );


  buf
  g1415
  (
    n1451,
    n1320
  );


  buf
  g1416
  (
    n1449,
    n1317
  );


  buf
  g1417
  (
    n1440,
    n1309
  );


  buf
  g1418
  (
    n1442,
    n1323
  );


  not
  g1419
  (
    n1443,
    n1310
  );


  not
  g1420
  (
    n1455,
    n1311
  );


  buf
  g1421
  (
    n1446,
    n1322
  );


  buf
  g1422
  (
    n1444,
    n1324
  );


  nand
  g1423
  (
    n1457,
    n1446,
    n1252,
    n1275,
    n1229
  );


  nand
  g1424
  (
    n1472,
    n1227,
    n1254,
    n1286,
    n1277
  );


  or
  g1425
  (
    n1465,
    n1239,
    n1238,
    n1220,
    n1206
  );


  nor
  g1426
  (
    n1470,
    n1283,
    n1442,
    n1251,
    n1273
  );


  and
  g1427
  (
    n1474,
    n1233,
    n1221,
    n1266,
    n1215
  );


  or
  g1428
  (
    n1466,
    n1207,
    n1228,
    n1237,
    n1281
  );


  or
  g1429
  (
    n1456,
    n1257,
    n1282,
    n1443,
    n1211
  );


  xor
  g1430
  (
    n1461,
    n1270,
    n1224,
    n1263,
    n1267
  );


  xor
  g1431
  (
    n1478,
    n1440,
    n1249,
    n1250,
    n1242
  );


  xnor
  g1432
  (
    n1476,
    n1441,
    n1280,
    n1446,
    n1271
  );


  xnor
  g1433
  (
    n1460,
    n1272,
    n1231,
    n1285,
    n1265
  );


  or
  g1434
  (
    n1480,
    n1258,
    n1261,
    n1244,
    n1445
  );


  or
  g1435
  (
    n1481,
    n1274,
    n1218,
    n1222,
    n1278
  );


  nand
  g1436
  (
    n1458,
    n1216,
    n1245,
    n1225,
    n1284
  );


  nor
  g1437
  (
    n1469,
    n1443,
    n1441,
    n1241,
    n1243
  );


  nor
  g1438
  (
    n1464,
    n1445,
    n1441,
    n1255,
    n1259
  );


  nand
  g1439
  (
    n1479,
    n1269,
    n1445,
    n1276,
    n1444
  );


  nand
  g1440
  (
    n1473,
    n1219,
    n1440,
    n1208,
    n1246
  );


  nand
  g1441
  (
    n1462,
    n1446,
    n1232,
    n1440,
    n1230
  );


  and
  g1442
  (
    n1463,
    n1444,
    n1442,
    n1235,
    n1264
  );


  and
  g1443
  (
    n1477,
    n1226,
    n1268,
    n1240,
    n1223
  );


  or
  g1444
  (
    n1468,
    n1279,
    n1442,
    n1213,
    n1253
  );


  xor
  g1445
  (
    n1471,
    n1210,
    n1444,
    n1445,
    n1256
  );


  and
  g1446
  (
    n1475,
    n1443,
    n1442,
    n1236,
    n1247
  );


  xnor
  g1447
  (
    n1459,
    n1443,
    n1262,
    n1212,
    n1217
  );


  nand
  g1448
  (
    n1482,
    n1214,
    n1444,
    n1440,
    n1209
  );


  xor
  g1449
  (
    n1467,
    n1260,
    n1248,
    n1234,
    n1441
  );


  and
  g1450
  (
    n1485,
    n1381,
    n1458,
    n1379,
    n1386
  );


  xnor
  g1451
  (
    n1510,
    n1392,
    n1341,
    n1367,
    n1345
  );


  nand
  g1452
  (
    n1488,
    n1359,
    n1460,
    n1344,
    n1374
  );


  xor
  g1453
  (
    KeyWire_0_15,
    n1457,
    n1399,
    n1372,
    n1401
  );


  xor
  g1454
  (
    n1508,
    n1460,
    n1395,
    n1360,
    n1380
  );


  or
  g1455
  (
    n1489,
    n1403,
    n1327,
    n1349,
    n1456
  );


  xnor
  g1456
  (
    n1506,
    n1394,
    n1456,
    n1350,
    n1337
  );


  nor
  g1457
  (
    n1492,
    n1370,
    n1414,
    n1354,
    n1463
  );


  or
  g1458
  (
    n1486,
    n1365,
    n1389,
    n1364,
    n1405
  );


  xnor
  g1459
  (
    n1496,
    n1413,
    n1407,
    n1368,
    n1366
  );


  nand
  g1460
  (
    n1505,
    n1390,
    n1397,
    n1460,
    n1457
  );


  nor
  g1461
  (
    n1512,
    n1362,
    n1339,
    n1459,
    n1461
  );


  and
  g1462
  (
    n1497,
    n1373,
    n1347,
    n1356,
    n1334
  );


  nand
  g1463
  (
    n1495,
    n1343,
    n1363,
    n1329,
    n1353
  );


  nand
  g1464
  (
    n1483,
    n1402,
    n1382,
    n1383,
    n1378
  );


  or
  g1465
  (
    n1498,
    n1459,
    n1338,
    n1351,
    n1461
  );


  xnor
  g1466
  (
    n1511,
    n1461,
    n1336,
    n1400,
    n1462
  );


  nor
  g1467
  (
    n1491,
    n1328,
    n1342,
    n1325,
    n1398
  );


  xnor
  g1468
  (
    n1494,
    n1369,
    n1457,
    n1375,
    n1396
  );


  or
  g1469
  (
    n1504,
    n1459,
    n1332,
    n1411,
    n1333
  );


  and
  g1470
  (
    n1502,
    n1461,
    n1387,
    n1404,
    n1410
  );


  and
  g1471
  (
    KeyWire_0_14,
    n1409,
    n1412,
    n1456,
    n1331
  );


  and
  g1472
  (
    n1500,
    n1458,
    n1330,
    n1335,
    n1462
  );


  and
  g1473
  (
    n1503,
    n1459,
    n1376,
    n1361,
    n1348
  );


  xnor
  g1474
  (
    n1501,
    n1457,
    n1458,
    n1391,
    n1326
  );


  xor
  g1475
  (
    n1490,
    n1355,
    n1460,
    n1358,
    n1340
  );


  nor
  g1476
  (
    n1507,
    n1352,
    n1357,
    n1377,
    n1384
  );


  and
  g1477
  (
    n1487,
    n1462,
    n1458,
    n1463,
    n1456
  );


  xor
  g1478
  (
    n1484,
    n1385,
    n1393,
    n1346,
    n1371
  );


  xor
  g1479
  (
    n1499,
    n1408,
    n1388,
    n1462,
    n1406
  );


  not
  g1480
  (
    n1552,
    n192
  );


  not
  g1481
  (
    n1527,
    n11
  );


  not
  g1482
  (
    n1526,
    n190
  );


  buf
  g1483
  (
    n1531,
    n1464
  );


  nor
  g1484
  (
    n1548,
    n1486,
    n1455
  );


  and
  g1485
  (
    n1513,
    n1506,
    n1451,
    n1511,
    n193
  );


  xnor
  g1486
  (
    n1514,
    n1295,
    n1448,
    n1511,
    n1505
  );


  and
  g1487
  (
    n1539,
    n668,
    n1449,
    n193,
    n1464
  );


  and
  g1488
  (
    n1550,
    n1501,
    n1466,
    n1465,
    n1447
  );


  or
  g1489
  (
    n1537,
    n1484,
    n1508,
    n1453,
    n1507
  );


  nor
  g1490
  (
    n1542,
    n1450,
    n1503,
    n1485,
    n1449
  );


  or
  g1491
  (
    n1524,
    n1512,
    n1292,
    n1450,
    n1509
  );


  xnor
  g1492
  (
    n1547,
    n191,
    n1448,
    n1453,
    n1492
  );


  nor
  g1493
  (
    n1519,
    n1491,
    n1504,
    n1502,
    n1510
  );


  nor
  g1494
  (
    n1518,
    n64,
    n11,
    n1490,
    n1448
  );


  nor
  g1495
  (
    n1515,
    n1466,
    n668,
    n10,
    n1287
  );


  xor
  g1496
  (
    n1535,
    n1487,
    n668,
    n10,
    n1504
  );


  xor
  g1497
  (
    n1525,
    n1464,
    n669,
    n1512,
    n1415
  );


  nand
  g1498
  (
    KeyWire_0_7,
    n190,
    n1483,
    n1464,
    n1451
  );


  and
  g1499
  (
    n1520,
    n192,
    n190,
    n669,
    n189
  );


  xnor
  g1500
  (
    n1540,
    n11,
    n65,
    n1465,
    n189
  );


  xnor
  g1501
  (
    n1541,
    n64,
    n191,
    n1453,
    n1455
  );


  nand
  g1502
  (
    n1532,
    n191,
    n1454,
    n1499,
    n1505
  );


  xnor
  g1503
  (
    n1538,
    n1450,
    n1495,
    n1289,
    n1452
  );


  or
  g1504
  (
    n1529,
    n1455,
    n192,
    n11,
    n1497
  );


  nor
  g1505
  (
    n1536,
    n10,
    n1452,
    n1489,
    n1291
  );


  or
  g1506
  (
    n1528,
    n1510,
    n1509,
    n1508,
    n1452
  );


  and
  g1507
  (
    n1543,
    n1447,
    n1500,
    n1506,
    n1296
  );


  nand
  g1508
  (
    n1517,
    n1496,
    n1290,
    n12,
    n1455
  );


  and
  g1509
  (
    n1533,
    n65,
    n189,
    n1449,
    n1507
  );


  nand
  g1510
  (
    n1549,
    n1493,
    n1299,
    n1463,
    n1450
  );


  nor
  g1511
  (
    n1551,
    n1297,
    n1298,
    n1453,
    n1498
  );


  xor
  g1512
  (
    n1523,
    n669,
    n1463,
    n1451,
    n1300
  );


  or
  g1513
  (
    n1516,
    n1301,
    n1454,
    n1446,
    n1447
  );


  xnor
  g1514
  (
    n1546,
    n1452,
    n1503,
    n10,
    n1449
  );


  or
  g1515
  (
    n1545,
    n64,
    n1293,
    n1288,
    n1465
  );


  or
  g1516
  (
    n1522,
    n189,
    n1451,
    n1302,
    n191
  );


  or
  g1517
  (
    n1521,
    n1465,
    n1454,
    n1294,
    n65
  );


  xor
  g1518
  (
    n1544,
    n192,
    n1494,
    n190,
    n1488
  );


  nand
  g1519
  (
    n1530,
    n65,
    n1447,
    n1454,
    n1448
  );


  buf
  g1520
  (
    n1575,
    n1547
  );


  buf
  g1521
  (
    n1665,
    n1537
  );


  not
  g1522
  (
    n1708,
    n1548
  );


  buf
  g1523
  (
    n1693,
    n1527
  );


  buf
  g1524
  (
    n1650,
    n30
  );


  not
  g1525
  (
    n1689,
    n1540
  );


  buf
  g1526
  (
    n1660,
    n17
  );


  buf
  g1527
  (
    n1561,
    n1551
  );


  buf
  g1528
  (
    n1656,
    n1469
  );


  buf
  g1529
  (
    n1620,
    n1536
  );


  not
  g1530
  (
    n1574,
    n1470
  );


  not
  g1531
  (
    n1572,
    n29
  );


  buf
  g1532
  (
    n1566,
    n21
  );


  not
  g1533
  (
    n1648,
    n1524
  );


  buf
  g1534
  (
    n1638,
    n22
  );


  buf
  g1535
  (
    n1647,
    n1478
  );


  buf
  g1536
  (
    n1663,
    n1478
  );


  not
  g1537
  (
    n1707,
    n1532
  );


  not
  g1538
  (
    n1587,
    n1479
  );


  not
  g1539
  (
    n1674,
    n1516
  );


  buf
  g1540
  (
    n1629,
    n31
  );


  not
  g1541
  (
    n1664,
    n19
  );


  not
  g1542
  (
    n1591,
    n1541
  );


  buf
  g1543
  (
    n1560,
    n28
  );


  buf
  g1544
  (
    n1642,
    n32
  );


  buf
  g1545
  (
    n1576,
    n24
  );


  not
  g1546
  (
    n1617,
    n1514
  );


  buf
  g1547
  (
    n1643,
    n1524
  );


  not
  g1548
  (
    n1634,
    n1467
  );


  buf
  g1549
  (
    n1652,
    n1542
  );


  buf
  g1550
  (
    n1627,
    n1547
  );


  buf
  g1551
  (
    n1631,
    n1523
  );


  not
  g1552
  (
    n1635,
    n1470
  );


  buf
  g1553
  (
    n1659,
    n1531
  );


  buf
  g1554
  (
    n1622,
    n25
  );


  buf
  g1555
  (
    n1555,
    n1538
  );


  not
  g1556
  (
    KeyWire_0_4,
    n1475
  );


  buf
  g1557
  (
    KeyWire_0_11,
    n16
  );


  buf
  g1558
  (
    n1640,
    n21
  );


  buf
  g1559
  (
    n1625,
    n1517
  );


  buf
  g1560
  (
    KeyWire_0_10,
    n31
  );


  buf
  g1561
  (
    n1711,
    n14
  );


  not
  g1562
  (
    n1583,
    n1518
  );


  buf
  g1563
  (
    n1600,
    n1548
  );


  not
  g1564
  (
    n1585,
    n1544
  );


  buf
  g1565
  (
    n1614,
    n22
  );


  not
  g1566
  (
    n1559,
    n1518
  );


  buf
  g1567
  (
    n1691,
    n16
  );


  buf
  g1568
  (
    n1655,
    n19
  );


  buf
  g1569
  (
    n1662,
    n1543
  );


  buf
  g1570
  (
    n1606,
    n28
  );


  not
  g1571
  (
    n1694,
    n1477
  );


  buf
  g1572
  (
    n1666,
    n20
  );


  buf
  g1573
  (
    n1658,
    n1546
  );


  not
  g1574
  (
    n1599,
    n1530
  );


  buf
  g1575
  (
    n1564,
    n29
  );


  buf
  g1576
  (
    n1688,
    n1526
  );


  buf
  g1577
  (
    n1567,
    n17
  );


  buf
  g1578
  (
    n1613,
    n30
  );


  buf
  g1579
  (
    n1710,
    n1517
  );


  not
  g1580
  (
    n1675,
    n1477
  );


  buf
  g1581
  (
    n1582,
    n1530
  );


  buf
  g1582
  (
    n1651,
    n1473
  );


  buf
  g1583
  (
    n1624,
    n1480
  );


  buf
  g1584
  (
    n1702,
    n24
  );


  buf
  g1585
  (
    n1667,
    n1474
  );


  buf
  g1586
  (
    n1712,
    n1546
  );


  not
  g1587
  (
    n1696,
    n26
  );


  buf
  g1588
  (
    n1657,
    n1468
  );


  buf
  g1589
  (
    n1578,
    n1538
  );


  not
  g1590
  (
    n1581,
    n1548
  );


  buf
  g1591
  (
    n1679,
    n66
  );


  buf
  g1592
  (
    n1593,
    n1532
  );


  not
  g1593
  (
    n1568,
    n1471
  );


  buf
  g1594
  (
    n1597,
    n1533
  );


  buf
  g1595
  (
    n1706,
    n32
  );


  buf
  g1596
  (
    n1616,
    n22
  );


  buf
  g1597
  (
    n1698,
    n26
  );


  buf
  g1598
  (
    n1697,
    n1479
  );


  buf
  g1599
  (
    n1601,
    n15
  );


  not
  g1600
  (
    n1681,
    n1541
  );


  buf
  g1601
  (
    n1586,
    n18
  );


  not
  g1602
  (
    n1579,
    n1547
  );


  buf
  g1603
  (
    n1569,
    n1515
  );


  buf
  g1604
  (
    n1670,
    n1552
  );


  not
  g1605
  (
    n1612,
    n1521
  );


  buf
  g1606
  (
    n1703,
    n1519
  );


  not
  g1607
  (
    n1577,
    n15
  );


  not
  g1608
  (
    n1595,
    n12
  );


  buf
  g1609
  (
    n1628,
    n1536
  );


  not
  g1610
  (
    n1654,
    n1530
  );


  not
  g1611
  (
    KeyWire_0_8,
    n1531
  );


  not
  g1612
  (
    n1641,
    n29
  );


  buf
  g1613
  (
    n1686,
    n1516
  );


  not
  g1614
  (
    n1678,
    n19
  );


  not
  g1615
  (
    n1623,
    n1531
  );


  buf
  g1616
  (
    n1604,
    n1468
  );


  buf
  g1617
  (
    n1699,
    n27
  );


  not
  g1618
  (
    n1690,
    n1533
  );


  not
  g1619
  (
    n1671,
    n1544
  );


  buf
  g1620
  (
    n1571,
    n1537
  );


  buf
  g1621
  (
    n1639,
    n13
  );


  not
  g1622
  (
    n1632,
    n1551
  );


  not
  g1623
  (
    n1589,
    n14
  );


  not
  g1624
  (
    n1645,
    n1525
  );


  buf
  g1625
  (
    n1615,
    n66
  );


  not
  g1626
  (
    n1621,
    n1466
  );


  buf
  g1627
  (
    n1683,
    n1480
  );


  nand
  g1628
  (
    n1704,
    n1552,
    n1546,
    n1472,
    n1521
  );


  xnor
  g1629
  (
    n1562,
    n1552,
    n1544,
    n1533,
    n1479
  );


  or
  g1630
  (
    n1669,
    n1532,
    n1476,
    n1536,
    n67
  );


  and
  g1631
  (
    n1598,
    n1545,
    n1531,
    n1539,
    n1520
  );


  nand
  g1632
  (
    n1556,
    n26,
    n1532,
    n1467,
    n1471
  );


  xor
  g1633
  (
    n1580,
    n30,
    n20,
    n32,
    n67
  );


  xor
  g1634
  (
    n1676,
    n1528,
    n23,
    n1539,
    n1517
  );


  xor
  g1635
  (
    n1611,
    n1515,
    n1518,
    n1539,
    n1523
  );


  xnor
  g1636
  (
    n1653,
    n1551,
    n18,
    n1524,
    n1545
  );


  nand
  g1637
  (
    n1588,
    n1545,
    n31,
    n1549,
    n1473
  );


  xor
  g1638
  (
    n1677,
    n1470,
    n1480,
    n1529
  );


  nor
  g1639
  (
    n1705,
    n1520,
    n1475,
    n1473,
    n1469
  );


  xnor
  g1640
  (
    n1610,
    n1545,
    n21,
    n14,
    n25
  );


  nor
  g1641
  (
    n1633,
    n1481,
    n1514,
    n1542,
    n1534
  );


  and
  g1642
  (
    n1672,
    n17,
    n15,
    n1550,
    n1538
  );


  or
  g1643
  (
    n1685,
    n1477,
    n1526,
    n1533,
    n13
  );


  nand
  g1644
  (
    n1609,
    n24,
    n1514,
    n1544,
    n18
  );


  or
  g1645
  (
    n1668,
    n23,
    n1528,
    n1540,
    n1542
  );


  xnor
  g1646
  (
    n1626,
    n1551,
    n18,
    n1539,
    n29
  );


  and
  g1647
  (
    n1590,
    n1467,
    n1522,
    n1473,
    n24
  );


  xnor
  g1648
  (
    n1558,
    n1472,
    n15,
    n1524,
    n1482
  );


  or
  g1649
  (
    n1673,
    n1518,
    n19,
    n1482,
    n1535
  );


  or
  g1650
  (
    n1630,
    n1527,
    n1534,
    n23,
    n1535
  );


  and
  g1651
  (
    n1554,
    n1550,
    n1543,
    n1481,
    n16
  );


  xor
  g1652
  (
    n1602,
    n66,
    n1474,
    n1513,
    n1476
  );


  nor
  g1653
  (
    n1584,
    n1550,
    n1528,
    n1516,
    n25
  );


  xor
  g1654
  (
    n1637,
    n1535,
    n66,
    n1475,
    n1478
  );


  xor
  g1655
  (
    n1573,
    n1467,
    n1536,
    n1519,
    n1475
  );


  nand
  g1656
  (
    n1644,
    n1519,
    n1530,
    n25,
    n1549
  );


  xor
  g1657
  (
    n1687,
    n1468,
    n28,
    n1534,
    n1472
  );


  and
  g1658
  (
    n1594,
    n17,
    n1529,
    n1522,
    n1474
  );


  or
  g1659
  (
    n1684,
    n1525,
    n1478,
    n1481,
    n1482
  );


  xnor
  g1660
  (
    n1619,
    n1547,
    n1543,
    n1529,
    n1542
  );


  nor
  g1661
  (
    n1709,
    n1525,
    n1527,
    n1481,
    n1482
  );


  nand
  g1662
  (
    KeyWire_0_2,
    n1538,
    n1521,
    n1517,
    n1468
  );


  nor
  g1663
  (
    n1636,
    n1522,
    n1540,
    n1476,
    n1477
  );


  xor
  g1664
  (
    n1553,
    n1516,
    n1541,
    n1469,
    n1550
  );


  xnor
  g1665
  (
    n1557,
    n30,
    n1525,
    n1527,
    n1546
  );


  and
  g1666
  (
    n1592,
    n1523,
    n21,
    n20,
    n1549
  );


  xor
  g1667
  (
    n1695,
    n20,
    n1526,
    n1537,
    n1471
  );


  nand
  g1668
  (
    n1692,
    n22,
    n1552,
    n26,
    n1540
  );


  and
  g1669
  (
    n1570,
    n32,
    n27,
    n1522,
    n1479
  );


  nor
  g1670
  (
    n1596,
    n1466,
    n1470,
    n1515,
    n14
  );


  or
  g1671
  (
    n1565,
    n31,
    n1513,
    n12,
    n1514
  );


  nand
  g1672
  (
    n1607,
    n1521,
    n1474,
    n1513,
    n28
  );


  nor
  g1673
  (
    n1682,
    n1534,
    n1471,
    n1537,
    n27
  );


  and
  g1674
  (
    n1680,
    n16,
    n13,
    n1513,
    n1476
  );


  nor
  g1675
  (
    n1605,
    n1549,
    n13,
    n1520
  );


  nor
  g1676
  (
    n1608,
    n1469,
    n23,
    n1526,
    n1528
  );


  or
  g1677
  (
    n1661,
    n12,
    n1523,
    n1472,
    n1543
  );


  and
  g1678
  (
    n1649,
    n27,
    n1548,
    n67,
    n1519
  );


  xor
  g1679
  (
    n1618,
    n1529,
    n1541,
    n1535,
    n1515
  );


  xor
  g1680
  (
    n1771,
    n1622,
    n1575,
    n1557,
    n1612
  );


  and
  g1681
  (
    n1756,
    n1579,
    n1670,
    n1583,
    n1573
  );


  xor
  g1682
  (
    n1774,
    n1644,
    n1665,
    n1566,
    n1652
  );


  nor
  g1683
  (
    n1777,
    n1554,
    n1631,
    n1582,
    n1651
  );


  or
  g1684
  (
    n1744,
    n1627,
    n1576,
    n1560,
    n1618
  );


  xor
  g1685
  (
    n1793,
    n1602,
    n1632,
    n1585,
    n1665
  );


  xor
  g1686
  (
    n1788,
    n1599,
    n1646,
    n1615,
    n1604
  );


  nor
  g1687
  (
    n1729,
    n1573,
    n1632,
    n1584,
    n1628
  );


  nand
  g1688
  (
    n1751,
    n1559,
    n1658,
    n1617,
    n1645
  );


  nand
  g1689
  (
    n1769,
    n1603,
    n1625,
    n1650,
    n1651
  );


  nand
  g1690
  (
    n1736,
    n1568,
    n1568,
    n1604,
    n1605
  );


  and
  g1691
  (
    n1734,
    n1635,
    n1647,
    n1667,
    n1596
  );


  xnor
  g1692
  (
    n1783,
    n1662,
    n1584,
    n1620,
    n1646
  );


  and
  g1693
  (
    n1801,
    n1628,
    n1594,
    n1635,
    n1571
  );


  and
  g1694
  (
    n1779,
    n1588,
    n1648,
    n1611,
    n1612
  );


  xor
  g1695
  (
    n1721,
    n1610,
    n1661,
    n1567,
    n1657
  );


  nor
  g1696
  (
    n1764,
    n1609,
    n1577,
    n1660,
    n1644
  );


  xnor
  g1697
  (
    n1730,
    n1594,
    n1663,
    n1646,
    n1658
  );


  xor
  g1698
  (
    n1775,
    n1616,
    n1663,
    n1654,
    n1664
  );


  nand
  g1699
  (
    n1767,
    n1672,
    n1648,
    n1624,
    n1615
  );


  and
  g1700
  (
    n1718,
    n1594,
    n1607,
    n1591,
    n1569
  );


  xnor
  g1701
  (
    n1761,
    n1636,
    n1624,
    n1625,
    n1607
  );


  nor
  g1702
  (
    n1713,
    n1655,
    n1558,
    n1587,
    n1610
  );


  xor
  g1703
  (
    n1726,
    n1622,
    n1640,
    n1645,
    n1653
  );


  nor
  g1704
  (
    n1762,
    n1555,
    n1634,
    n1581,
    n1606
  );


  and
  g1705
  (
    n1765,
    n1622,
    n1603,
    n1633,
    n1627
  );


  xor
  g1706
  (
    n1768,
    n1644,
    n1611,
    n1629,
    n1660
  );


  xnor
  g1707
  (
    n1731,
    n1586,
    n1617,
    n1565,
    n1663
  );


  xor
  g1708
  (
    n1716,
    n1565,
    n1563,
    n1557,
    n1609
  );


  nand
  g1709
  (
    n1732,
    n1561,
    n1655,
    n1595,
    n1562
  );


  nand
  g1710
  (
    n1720,
    n1592,
    n1595,
    n1580
  );


  xor
  g1711
  (
    n1778,
    n1566,
    n1574,
    n1596,
    n1632
  );


  xnor
  g1712
  (
    n1727,
    n1563,
    n1619,
    n1581,
    n1659
  );


  nor
  g1713
  (
    n1766,
    n1613,
    n1553,
    n1592,
    n1669
  );


  and
  g1714
  (
    n1750,
    n1607,
    n1558,
    n1591,
    n1608
  );


  nand
  g1715
  (
    n1745,
    n1601,
    n1627,
    n1617,
    n1609
  );


  nand
  g1716
  (
    n1757,
    n1567,
    n1588,
    n1579,
    n1666
  );


  xor
  g1717
  (
    n1780,
    n1561,
    n1642,
    n1569,
    n1611
  );


  xor
  g1718
  (
    n1752,
    n1571,
    n1637,
    n1642,
    n1640
  );


  nor
  g1719
  (
    n1743,
    n1643,
    n1621,
    n1638,
    n1624
  );


  nor
  g1720
  (
    n1795,
    n1638,
    n1621,
    n1595,
    n1648
  );


  nor
  g1721
  (
    n1776,
    n1600,
    n1568,
    n1564,
    n1639
  );


  nor
  g1722
  (
    n1738,
    n1571,
    n1623,
    n1638,
    n1588
  );


  xor
  g1723
  (
    n1749,
    n1572,
    n1625,
    n1652,
    n1618
  );


  and
  g1724
  (
    n1737,
    n1605,
    n1585,
    n1637,
    n1657
  );


  xor
  g1725
  (
    n1794,
    n1560,
    n1664,
    n1599,
    n1575
  );


  xor
  g1726
  (
    n1799,
    n1559,
    n1596,
    n1634,
    n1572
  );


  or
  g1727
  (
    n1770,
    n1629,
    n1641,
    n1586,
    n1667
  );


  and
  g1728
  (
    n1787,
    n1654,
    n1650,
    n1626,
    n1583
  );


  and
  g1729
  (
    n1785,
    n1601,
    n1649,
    n1598,
    n1615
  );


  nand
  g1730
  (
    n1758,
    n1660,
    n1554,
    n1636,
    n1572
  );


  xor
  g1731
  (
    n1733,
    n1656,
    n1556,
    n1619,
    n1672
  );


  xnor
  g1732
  (
    n1724,
    n1619,
    n1658,
    n1579,
    n1636
  );


  nor
  g1733
  (
    n1763,
    n1661,
    n1593,
    n1567,
    n1604
  );


  and
  g1734
  (
    n1796,
    n1612,
    n1671,
    n1647,
    n1645
  );


  and
  g1735
  (
    n1791,
    n1601,
    n1643,
    n1562,
    n1578
  );


  nand
  g1736
  (
    n1797,
    n1587,
    n1582,
    n1635,
    n1637
  );


  xor
  g1737
  (
    n1754,
    n1664,
    n1651,
    n1653,
    n1643
  );


  nand
  g1738
  (
    n1717,
    n1600,
    n1672,
    n1606,
    n1613
  );


  nand
  g1739
  (
    n1782,
    n1583,
    n1661,
    n1671,
    n1564
  );


  nor
  g1740
  (
    n1781,
    n1620,
    n1593,
    n1614,
    n1566
  );


  xor
  g1741
  (
    n1798,
    n1621,
    n1563,
    n1591,
    n1598
  );


  xnor
  g1742
  (
    n1740,
    n1662,
    n1629,
    n1597,
    n1577
  );


  nand
  g1743
  (
    n1728,
    n1650,
    n1616,
    n1633,
    n1555
  );


  nand
  g1744
  (
    n1725,
    n1593,
    n1578,
    n1597,
    n1576
  );


  or
  g1745
  (
    n1715,
    n1630,
    n1641,
    n1589,
    n1631
  );


  or
  g1746
  (
    n1735,
    n1580,
    n1590,
    n1608,
    n1570
  );


  xnor
  g1747
  (
    n1748,
    n1589,
    n1565,
    n1630,
    n1639
  );


  nand
  g1748
  (
    n1747,
    n1559,
    n1561,
    n1556,
    n1655
  );


  xnor
  g1749
  (
    n1786,
    n1669,
    n1574,
    n1626,
    n1647
  );


  xnor
  g1750
  (
    n1784,
    n1603,
    n1659,
    n1640,
    n1558
  );


  xor
  g1751
  (
    n1742,
    n1641,
    n1631,
    n1628,
    n1575
  );


  or
  g1752
  (
    n1746,
    n1560,
    n1584,
    n1614,
    n1618
  );


  nor
  g1753
  (
    n1790,
    n1573,
    n1670,
    n1639,
    n1582
  );


  xnor
  g1754
  (
    n1739,
    n1620,
    n1668,
    n1666,
    n1587
  );


  nor
  g1755
  (
    n1741,
    n1614,
    n1562,
    n1574,
    n1606
  );


  and
  g1756
  (
    n1792,
    n1585,
    n1557,
    n1608,
    n1570
  );


  or
  g1757
  (
    n1772,
    n1553,
    n1667,
    n1605,
    n1626
  );


  xor
  g1758
  (
    n1800,
    n1576,
    n1581,
    n1592,
    n1671
  );


  and
  g1759
  (
    n1753,
    n1666,
    n1654,
    n1564,
    n1590
  );


  or
  g1760
  (
    n1789,
    n1669,
    n1623,
    n1613,
    n1662
  );


  nor
  g1761
  (
    n1723,
    n1586,
    n1656,
    n1602,
    n1642
  );


  nand
  g1762
  (
    n1714,
    n1649,
    n1599,
    n1590,
    n1623
  );


  nand
  g1763
  (
    n1719,
    n1656,
    n1630,
    n1602,
    n1600
  );


  nor
  g1764
  (
    n1755,
    n1668,
    n1653,
    n1649,
    n1652
  );


  xor
  g1765
  (
    n1722,
    n1589,
    n1665,
    n1657,
    n1578
  );


  xor
  g1766
  (
    n1759,
    n1616,
    n1633,
    n1577,
    n1570
  );


  nor
  g1767
  (
    n1773,
    n1668,
    n1569,
    n1670,
    n1634
  );


  nor
  g1768
  (
    n1760,
    n1597,
    n1610,
    n1598,
    n1659
  );


  buf
  g1769
  (
    n1803,
    n1722
  );


  buf
  g1770
  (
    n1804,
    n1720
  );


  not
  g1771
  (
    n1807,
    n1724
  );


  buf
  g1772
  (
    n1806,
    n1713
  );


  and
  g1773
  (
    n1802,
    n1717,
    n1723,
    n1714,
    n1721
  );


  and
  g1774
  (
    n1805,
    n1715,
    n1718,
    n1719,
    n1716
  );


  not
  g1775
  (
    n1819,
    n1804
  );


  buf
  g1776
  (
    n1810,
    n1804
  );


  buf
  g1777
  (
    n1812,
    n1805
  );


  not
  g1778
  (
    n1809,
    n1802
  );


  buf
  g1779
  (
    n1818,
    n1803
  );


  not
  g1780
  (
    n1808,
    n1804
  );


  not
  g1781
  (
    n1814,
    n1806
  );


  not
  g1782
  (
    n1811,
    n1805
  );


  buf
  g1783
  (
    n1813,
    n1803
  );


  not
  g1784
  (
    n1815,
    n1803
  );


  not
  g1785
  (
    n1817,
    n1805
  );


  not
  g1786
  (
    n1816,
    n1802
  );


  not
  g1787
  (
    n1821,
    n1808
  );


  not
  g1788
  (
    n1822,
    n1809
  );


  not
  g1789
  (
    n1823,
    n1303
  );


  not
  g1790
  (
    n1825,
    n1808
  );


  buf
  g1791
  (
    n1820,
    n1809
  );


  not
  g1792
  (
    n1826,
    n1808
  );


  xnor
  g1793
  (
    n1824,
    n1809,
    n1808
  );


  buf
  g1794
  (
    n1831,
    n1822
  );


  buf
  g1795
  (
    n1835,
    n1823
  );


  buf
  g1796
  (
    n1841,
    n1821
  );


  buf
  g1797
  (
    n1827,
    n1826
  );


  buf
  g1798
  (
    n1844,
    n1824
  );


  not
  g1799
  (
    n1850,
    n1825
  );


  buf
  g1800
  (
    n1853,
    n1821
  );


  buf
  g1801
  (
    n1854,
    n1821
  );


  buf
  g1802
  (
    n1834,
    n1823
  );


  buf
  g1803
  (
    KeyWire_0_6,
    n1825
  );


  not
  g1804
  (
    n1838,
    n1826
  );


  not
  g1805
  (
    n1832,
    n1820
  );


  not
  g1806
  (
    n1836,
    n1825
  );


  not
  g1807
  (
    n1846,
    n1820
  );


  buf
  g1808
  (
    n1848,
    n1824
  );


  not
  g1809
  (
    n1845,
    n1825
  );


  not
  g1810
  (
    n1852,
    n1824
  );


  buf
  g1811
  (
    n1830,
    n1822
  );


  not
  g1812
  (
    n1839,
    n1822
  );


  not
  g1813
  (
    n1833,
    n1820
  );


  buf
  g1814
  (
    n1829,
    n1826
  );


  buf
  g1815
  (
    n1837,
    n1823
  );


  buf
  g1816
  (
    n1842,
    n1822
  );


  buf
  g1817
  (
    n1849,
    n1823
  );


  buf
  g1818
  (
    n1847,
    n1821
  );


  buf
  g1819
  (
    n1828,
    n1826
  );


  buf
  g1820
  (
    n1851,
    n1820
  );


  buf
  g1821
  (
    n1843,
    n1824
  );


  not
  g1822
  (
    n1869,
    n1833
  );


  xnor
  g1823
  (
    n1855,
    n1846,
    n1828,
    n1833
  );


  and
  g1824
  (
    n1882,
    n1813,
    n1844,
    n1838,
    n1819
  );


  and
  g1825
  (
    n1871,
    n1819,
    n1846,
    n1831,
    n1827
  );


  or
  g1826
  (
    KeyWire_0_12,
    n1833,
    n1840,
    n1416
  );


  and
  g1827
  (
    n1868,
    n1829,
    n1814,
    n1815,
    n1843
  );


  and
  g1828
  (
    n1877,
    n1827,
    n1839,
    n1818,
    n1842
  );


  nor
  g1829
  (
    n1883,
    n1839,
    n1845,
    n1848,
    n1838
  );


  or
  g1830
  (
    n1890,
    n1832,
    n1819,
    n1818,
    n1834
  );


  and
  g1831
  (
    n1864,
    n1811,
    n1851,
    n1849,
    n1847
  );


  and
  g1832
  (
    n1875,
    n1815,
    n1838,
    n1850,
    n1837
  );


  xnor
  g1833
  (
    n1862,
    n1835,
    n1842,
    n1844,
    n1839
  );


  nor
  g1834
  (
    n1873,
    n1846,
    n1840,
    n1816,
    n1837
  );


  nand
  g1835
  (
    n1879,
    n1813,
    n1811,
    n1827,
    n1836
  );


  xnor
  g1836
  (
    n1874,
    n1847,
    n1849,
    n1836
  );


  nand
  g1837
  (
    n1866,
    n1811,
    n1850,
    n1831,
    n1817
  );


  xor
  g1838
  (
    n1861,
    n1835,
    n1841,
    n1814,
    n1817
  );


  xnor
  g1839
  (
    n1867,
    n1814,
    n1818,
    n1417,
    n1816
  );


  nand
  g1840
  (
    n1888,
    n1830,
    n1816,
    n1829
  );


  and
  g1841
  (
    n1857,
    n1848,
    n1813,
    n1837,
    n1845
  );


  xnor
  g1842
  (
    n1859,
    n1841,
    n1843,
    n1847,
    n1832
  );


  xnor
  g1843
  (
    n1884,
    n1831,
    n1810,
    n1818,
    n1834
  );


  and
  g1844
  (
    n1886,
    n1848,
    n1830,
    n1833,
    n1840
  );


  xnor
  g1845
  (
    n1872,
    n1842,
    n1814,
    n1810,
    n1831
  );


  xnor
  g1846
  (
    n1860,
    n1809,
    n1827,
    n1836,
    n1835
  );


  or
  g1847
  (
    n1870,
    n1845,
    n1830,
    n1841,
    n1811
  );


  nor
  g1848
  (
    n1881,
    n1850,
    n1842,
    n1832,
    n1836
  );


  nand
  g1849
  (
    n1887,
    n1830,
    n1816,
    n1817
  );


  xnor
  g1850
  (
    n1863,
    n1844,
    n1848,
    n1812,
    n1834
  );


  or
  g1851
  (
    n1889,
    n1829,
    n1847,
    n1843,
    n1810
  );


  or
  g1852
  (
    n1876,
    n1828,
    n1835,
    n1844,
    n1841
  );


  and
  g1853
  (
    n1858,
    n1834,
    n1812,
    n1837
  );


  or
  g1854
  (
    n1878,
    n1810,
    n1812,
    n1849,
    n1828
  );


  or
  g1855
  (
    n1856,
    n1828,
    n1815,
    n1819,
    n1845
  );


  xnor
  g1856
  (
    n1885,
    n1846,
    n1839,
    n1843,
    n1850
  );


  nand
  g1857
  (
    n1880,
    n1832,
    n1813,
    n1838,
    n1815
  );


  not
  g1858
  (
    n1894,
    n1856
  );


  buf
  g1859
  (
    n1892,
    n1858
  );


  buf
  g1860
  (
    n1893,
    n1855
  );


  not
  g1861
  (
    n1891,
    n1857
  );


  and
  g1862
  (
    n1902,
    n671,
    n1853,
    n1428,
    n670
  );


  xor
  g1863
  (
    n1898,
    n672,
    n1894,
    n1893,
    n1432
  );


  and
  g1864
  (
    n1905,
    n1851,
    n1854,
    n1427,
    n1433
  );


  xnor
  g1865
  (
    n1904,
    n1854,
    n1892,
    n1851,
    n1421
  );


  nand
  g1866
  (
    n1907,
    n1853,
    n1893,
    n1422
  );


  xnor
  g1867
  (
    n1895,
    n673,
    n1425,
    n1853,
    n670
  );


  and
  g1868
  (
    n1909,
    n672,
    n1424,
    n1891,
    n1852
  );


  xnor
  g1869
  (
    n1901,
    n1420,
    n670,
    n1431,
    n1852
  );


  or
  g1870
  (
    n1903,
    n1304,
    n1853,
    n1419,
    n1418
  );


  nor
  g1871
  (
    n1908,
    n1893,
    n1891,
    n1434
  );


  xor
  g1872
  (
    n1910,
    n669,
    n1852,
    n672,
    n1429
  );


  xnor
  g1873
  (
    n1896,
    n671,
    n1852,
    n1854,
    n672
  );


  xor
  g1874
  (
    n1897,
    n1894,
    n673,
    n1891,
    n1423
  );


  xor
  g1875
  (
    n1900,
    n1894,
    n1426,
    n671,
    n1854
  );


  or
  g1876
  (
    n1899,
    n670,
    n1892,
    n1894
  );


  nand
  g1877
  (
    n1906,
    n1851,
    n671,
    n1892,
    n1430
  );


  nor
  g1878
  (
    n1919,
    n68,
    n1910,
    n1906
  );


  xnor
  g1879
  (
    n1918,
    n1437,
    n1861,
    n1869
  );


  nor
  g1880
  (
    n1923,
    n1435,
    n1863,
    n1884
  );


  and
  g1881
  (
    n1922,
    n1905,
    n1910,
    n1867
  );


  and
  g1882
  (
    n1913,
    n1874,
    n1877,
    n1909
  );


  nor
  g1883
  (
    n1926,
    n1864,
    n1900,
    n1885
  );


  nor
  g1884
  (
    n1927,
    n1876,
    n1865,
    n1887
  );


  nor
  g1885
  (
    n1921,
    n1872,
    n1878,
    n1883
  );


  xnor
  g1886
  (
    n1912,
    n1860,
    n1908,
    n68
  );


  nand
  g1887
  (
    n1924,
    n1890,
    n193,
    n68
  );


  xor
  g1888
  (
    n1925,
    n1898,
    n1880,
    n1895
  );


  or
  g1889
  (
    n1929,
    n1907,
    n1899,
    n1889
  );


  and
  g1890
  (
    n1914,
    n1902,
    n1908,
    n1868
  );


  xnor
  g1891
  (
    n1915,
    n1866,
    n1879,
    n1862
  );


  and
  g1892
  (
    n1917,
    n1901,
    n1909,
    n1439
  );


  xnor
  g1893
  (
    n1911,
    n1896,
    n1897,
    n1859
  );


  nor
  g1894
  (
    n1928,
    n1873,
    n1903,
    n1875,
    n1882
  );


  xnor
  g1895
  (
    n1916,
    n1871,
    n1886,
    n1870,
    n67
  );


  xor
  g1896
  (
    n1920,
    n193,
    n68,
    n1888,
    n1438
  );


  nor
  g1897
  (
    n1930,
    n1881,
    n1907,
    n1904,
    n1436
  );


  or
  g1898
  (
    n1967,
    n1694,
    n1700,
    n1921,
    n1928
  );


  nor
  g1899
  (
    n1944,
    n1682,
    n1693,
    n1705,
    n1695
  );


  and
  g1900
  (
    n1960,
    n1683,
    n1912,
    n1694,
    n1681
  );


  xor
  g1901
  (
    n1933,
    n1711,
    n1673,
    n1929,
    n1690
  );


  xor
  g1902
  (
    n1958,
    n1688,
    n1701,
    n1920,
    n1673
  );


  or
  g1903
  (
    n1968,
    n1676,
    n1916,
    n1696,
    n1701
  );


  nor
  g1904
  (
    n1964,
    n1923,
    n1675,
    n1928,
    n1698
  );


  nand
  g1905
  (
    n1950,
    n1687,
    n1926,
    n1674,
    n1673
  );


  xnor
  g1906
  (
    n1954,
    n1923,
    n1680,
    n1699,
    n1708
  );


  nor
  g1907
  (
    n1965,
    n1679,
    n1710,
    n1915
  );


  nand
  g1908
  (
    n1936,
    n1916,
    n1924,
    n1680,
    n1697
  );


  xor
  g1909
  (
    n1959,
    n1688,
    n1930,
    n1681,
    n1693
  );


  or
  g1910
  (
    n1962,
    n1696,
    n1682,
    n1674,
    n1683
  );


  nor
  g1911
  (
    n1955,
    n1929,
    n1700,
    n1702,
    n1926
  );


  nand
  g1912
  (
    n1956,
    n1922,
    n1911,
    n1913
  );


  nand
  g1913
  (
    n1945,
    n1921,
    n1685,
    n1696,
    n1707
  );


  xnor
  g1914
  (
    n1951,
    n1925,
    n1703,
    n1677,
    n1919
  );


  xor
  g1915
  (
    n1952,
    n1686,
    n1708,
    n1914,
    n1694
  );


  and
  g1916
  (
    n1961,
    n1684,
    n1706,
    n1693,
    n1678
  );


  or
  g1917
  (
    n1963,
    n1709,
    n1699,
    n1686,
    n1691
  );


  xor
  g1918
  (
    n1946,
    n1917,
    n1689,
    n1703,
    n1709
  );


  or
  g1919
  (
    n1932,
    n1680,
    n1929,
    n1706,
    n1927
  );


  nor
  g1920
  (
    n1937,
    n1684,
    n1695,
    n1918,
    n1682
  );


  nor
  g1921
  (
    n1935,
    n1681,
    n1706,
    n1703,
    n1690
  );


  nand
  g1922
  (
    n1942,
    n1684,
    n1702,
    n1697,
    n1920
  );


  xnor
  g1923
  (
    n1966,
    n1704,
    n1924,
    n1918,
    n1697
  );


  nor
  g1924
  (
    n1949,
    n1686,
    n1927,
    n1683,
    n1679
  );


  xnor
  g1925
  (
    n1934,
    n1712,
    n1914,
    n1704,
    n1701
  );


  or
  g1926
  (
    n1943,
    n1687,
    n1687,
    n1700,
    n1702
  );


  and
  g1927
  (
    n1939,
    n1692,
    n1689,
    n1691,
    n1925
  );


  xnor
  g1928
  (
    n1948,
    n1699,
    n1691,
    n1705,
    n1710
  );


  nor
  g1929
  (
    n1947,
    n1709,
    n1930,
    n1698,
    n1688
  );


  or
  g1930
  (
    n1941,
    n1679,
    n1919,
    n1917,
    n1707
  );


  xnor
  g1931
  (
    n1957,
    n1922,
    n1711,
    n1698,
    n1677
  );


  and
  g1932
  (
    n1970,
    n1675,
    n1915,
    n1707,
    n1678
  );


  or
  g1933
  (
    n1969,
    n1695,
    n1676,
    n1930,
    n1708
  );


  or
  g1934
  (
    n1938,
    n1689,
    n1678,
    n1705,
    n1676
  );


  xor
  g1935
  (
    n1931,
    n1704,
    n1677,
    n1692,
    n1712
  );


  nand
  g1936
  (
    n1953,
    n1690,
    n1674,
    n1711,
    n1675
  );


  xor
  g1937
  (
    n1940,
    n1685,
    n1685,
    n1712,
    n1692
  );


  and
  g1938
  (
    n1985,
    n1730,
    n1959,
    n1946,
    n1962
  );


  or
  g1939
  (
    n2005,
    n1777,
    n1965,
    n1800
  );


  nor
  g1940
  (
    n1977,
    n1933,
    n1725,
    n1757,
    n1944
  );


  xor
  g1941
  (
    n2009,
    n1955,
    n1958,
    n1942,
    n1774
  );


  nor
  g1942
  (
    n1986,
    n673,
    n1745,
    n1969,
    n1779
  );


  nand
  g1943
  (
    n2000,
    n1732,
    n1769,
    n1948,
    n1947
  );


  or
  g1944
  (
    n1998,
    n1945,
    n1750,
    n1969
  );


  or
  g1945
  (
    n1993,
    n1932,
    n1739,
    n1953,
    n1934
  );


  xnor
  g1946
  (
    n1976,
    n1776,
    n1944,
    n1966,
    n1941
  );


  xor
  g1947
  (
    n1987,
    n1738,
    n1962,
    n1788,
    n1787
  );


  xor
  g1948
  (
    n1979,
    n1963,
    n1952,
    n1939,
    n1957
  );


  xor
  g1949
  (
    n2010,
    n1764,
    n1970,
    n1763,
    n1933
  );


  nor
  g1950
  (
    n2002,
    n1784,
    n1749,
    n1940,
    n1798
  );


  xor
  g1951
  (
    n2018,
    n1786,
    n1947,
    n1746,
    n1968
  );


  xnor
  g1952
  (
    n2007,
    n1939,
    n1729,
    n1942,
    n1781
  );


  nor
  g1953
  (
    n1997,
    n1940,
    n1968,
    n1736,
    n1943
  );


  xor
  g1954
  (
    n2004,
    n1943,
    n1743,
    n1951,
    n1963
  );


  nor
  g1955
  (
    n1984,
    n1956,
    n1950,
    n1958,
    n1935
  );


  nand
  g1956
  (
    n2006,
    n1759,
    n1946,
    n1937,
    n1748
  );


  or
  g1957
  (
    n1980,
    n1961,
    n1948,
    n1744
  );


  xnor
  g1958
  (
    n2003,
    n1791,
    n1964,
    n1959,
    n1954
  );


  and
  g1959
  (
    n1972,
    n1931,
    n1954,
    n1951,
    n1956
  );


  nor
  g1960
  (
    n1988,
    n1735,
    n1967,
    n1726,
    n1953
  );


  or
  g1961
  (
    n1992,
    n1967,
    n1932,
    n1961,
    n1797
  );


  xor
  g1962
  (
    n1982,
    n1773,
    n1944,
    n1772,
    n1767
  );


  xor
  g1963
  (
    n1990,
    n1782,
    n1742,
    n1949
  );


  xor
  g1964
  (
    n1991,
    n1790,
    n1943,
    n1799,
    n1728
  );


  xor
  g1965
  (
    n2013,
    n1970,
    n1747,
    n1952,
    n1958
  );


  xor
  g1966
  (
    n2017,
    n1938,
    n1795,
    n1771,
    n1964
  );


  xnor
  g1967
  (
    n2011,
    n1952,
    n1931,
    n1960,
    n1789
  );


  or
  g1968
  (
    n1978,
    n1794,
    n1966,
    n1945,
    n1960
  );


  and
  g1969
  (
    n1973,
    n1796,
    n1951,
    n1938,
    n1970
  );


  or
  g1970
  (
    n2016,
    n1942,
    n1783,
    n1954,
    n1792
  );


  nor
  g1971
  (
    n2001,
    n1936,
    n1727,
    n1955,
    n1934
  );


  nand
  g1972
  (
    n1975,
    n1737,
    n1955,
    n1785,
    n1741
  );


  nand
  g1973
  (
    n1995,
    n1961,
    n1939,
    n1766,
    n1966
  );


  nand
  g1974
  (
    n1996,
    n1964,
    n1960,
    n1770,
    n1936
  );


  nand
  g1975
  (
    n1974,
    n1778,
    n1793,
    n1967,
    n1947
  );


  xor
  g1976
  (
    n2008,
    n1753,
    n1957,
    n1761,
    n1963
  );


  or
  g1977
  (
    n2012,
    n1941,
    n1953,
    n1956,
    n1775
  );


  nand
  g1978
  (
    n1989,
    n1765,
    n1937,
    n1755,
    n1962
  );


  nand
  g1979
  (
    n2015,
    n1938,
    n1945,
    n1965,
    n1959
  );


  nor
  g1980
  (
    n1999,
    n1968,
    n1937,
    n1950,
    n1801
  );


  or
  g1981
  (
    n1983,
    n1751,
    n1768,
    n1758,
    n1957
  );


  and
  g1982
  (
    n1981,
    n1780,
    n1754,
    n1733,
    n1946
  );


  nand
  g1983
  (
    n1971,
    n1949,
    n1760,
    n1950,
    n1941
  );


  nand
  g1984
  (
    n2014,
    n1740,
    n1762,
    n1734,
    n1756
  );


  or
  g1985
  (
    n1994,
    n1940,
    n1935,
    n1731,
    n1752
  );


  and
  g1986
  (
    n2020,
    n1993,
    n1807,
    n2000,
    n1991
  );


  xor
  g1987
  (
    n2024,
    n2004,
    n673,
    n2006,
    n1806
  );


  xnor
  g1988
  (
    n2025,
    n1992,
    n1997,
    n1990,
    n2011
  );


  or
  g1989
  (
    n2023,
    n2010,
    n1994,
    n1999,
    n2007
  );


  xor
  g1990
  (
    n2027,
    n1806,
    n2003,
    n2008,
    n1979
  );


  xnor
  g1991
  (
    n2029,
    n2017,
    n1974,
    n2002,
    n1995
  );


  xor
  g1992
  (
    n2031,
    n1980,
    n1305,
    n2016,
    n2012
  );


  nor
  g1993
  (
    n2021,
    n1998,
    n1996,
    n1984,
    n1972
  );


  and
  g1994
  (
    n2032,
    n1807,
    n1985,
    n1982,
    n1987
  );


  or
  g1995
  (
    n2022,
    n1306,
    n1978,
    n2009,
    n1973
  );


  and
  g1996
  (
    n2026,
    n1989,
    n1976,
    n1986,
    n1977
  );


  and
  g1997
  (
    n2030,
    n2001,
    n1981,
    n1988,
    n2015
  );


  nor
  g1998
  (
    n2028,
    n1971,
    n1983,
    n2014,
    n2013
  );


  and
  g1999
  (
    n2019,
    n2005,
    n2018,
    n1807,
    n1975
  );


  xor
  KeyGate_0_0
  (
    n1201,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n446,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1701,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1083,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1646,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n862,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1840,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1534,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1603,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1182,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n1563,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1700,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n1865,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1151,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1493,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1509,
    KeyNOTWire_0_15
  );


endmodule

