

module Stat_1000_341
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n900,
  n901,
  n903,
  n905,
  n909,
  n904,
  n910,
  n922,
  n924,
  n926,
  n927,
  n933,
  n936,
  n1032,
  n1018,
  n1021,
  n1015,
  n1029,
  n1023,
  n1019,
  n1020,
  n1022,
  n1030,
  n1027,
  n1014,
  n1028,
  n1025,
  n1026,
  n1016,
  n1024,
  n1017,
  n1031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n900;
  output n901;
  output n903;
  output n905;
  output n909;
  output n904;
  output n910;
  output n922;
  output n924;
  output n926;
  output n927;
  output n933;
  output n936;
  output n1032;
  output n1018;
  output n1021;
  output n1015;
  output n1029;
  output n1023;
  output n1019;
  output n1020;
  output n1022;
  output n1030;
  output n1027;
  output n1014;
  output n1028;
  output n1025;
  output n1026;
  output n1016;
  output n1024;
  output n1017;
  output n1031;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n902;
  wire n906;
  wire n907;
  wire n908;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n923;
  wire n925;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n934;
  wire n935;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n37,
    n5
  );


  buf
  g1
  (
    n81,
    n4
  );


  buf
  g2
  (
    KeyWire_0_43,
    n11
  );


  buf
  g3
  (
    n48,
    n6
  );


  buf
  g4
  (
    n34,
    n11
  );


  buf
  g5
  (
    n42,
    n2
  );


  buf
  g6
  (
    n51,
    n8
  );


  buf
  g7
  (
    n66,
    n3
  );


  buf
  g8
  (
    n64,
    n3
  );


  buf
  g9
  (
    n68,
    n2
  );


  not
  g10
  (
    n63,
    n13
  );


  not
  g11
  (
    n82,
    n10
  );


  buf
  g12
  (
    n59,
    n3
  );


  not
  g13
  (
    KeyWire_0_57,
    n1
  );


  buf
  g14
  (
    KeyWire_0_9,
    n6
  );


  buf
  g15
  (
    n47,
    n14
  );


  not
  g16
  (
    n79,
    n6
  );


  not
  g17
  (
    n70,
    n4
  );


  buf
  g18
  (
    n65,
    n10
  );


  buf
  g19
  (
    n78,
    n8
  );


  not
  g20
  (
    n44,
    n12
  );


  not
  g21
  (
    n85,
    n12
  );


  buf
  g22
  (
    n54,
    n4
  );


  not
  g23
  (
    n88,
    n5
  );


  not
  g24
  (
    n49,
    n8
  );


  buf
  g25
  (
    n55,
    n4
  );


  not
  g26
  (
    n76,
    n14
  );


  not
  g27
  (
    n73,
    n1
  );


  not
  g28
  (
    n62,
    n13
  );


  not
  g29
  (
    n87,
    n7
  );


  not
  g30
  (
    n35,
    n3
  );


  buf
  g31
  (
    n41,
    n9
  );


  not
  g32
  (
    n33,
    n9
  );


  buf
  g33
  (
    KeyWire_0_18,
    n5
  );


  not
  g34
  (
    n77,
    n2
  );


  not
  g35
  (
    n39,
    n7
  );


  not
  g36
  (
    n45,
    n12
  );


  not
  g37
  (
    n75,
    n7
  );


  not
  g38
  (
    n86,
    n8
  );


  buf
  g39
  (
    n56,
    n10
  );


  buf
  g40
  (
    n53,
    n1
  );


  not
  g41
  (
    n52,
    n6
  );


  not
  g42
  (
    n80,
    n9
  );


  buf
  g43
  (
    n43,
    n14
  );


  not
  g44
  (
    n61,
    n13
  );


  not
  g45
  (
    n46,
    n10
  );


  buf
  g46
  (
    n71,
    n9
  );


  buf
  g47
  (
    n58,
    n2
  );


  buf
  g48
  (
    n38,
    n1
  );


  not
  g49
  (
    n67,
    n12
  );


  not
  g50
  (
    n40,
    n5
  );


  not
  g51
  (
    n60,
    n14
  );


  not
  g52
  (
    n72,
    n11
  );


  buf
  g53
  (
    n84,
    n11
  );


  buf
  g54
  (
    n74,
    n13
  );


  not
  g55
  (
    n50,
    n7
  );


  not
  g56
  (
    KeyWire_0_24,
    n36
  );


  buf
  g57
  (
    n149,
    n71
  );


  not
  g58
  (
    n97,
    n50
  );


  buf
  g59
  (
    n120,
    n67
  );


  not
  g60
  (
    n175,
    n60
  );


  not
  g61
  (
    n130,
    n44
  );


  buf
  g62
  (
    KeyWire_0_33,
    n38
  );


  not
  g63
  (
    n116,
    n77
  );


  buf
  g64
  (
    KeyWire_0_1,
    n68
  );


  not
  g65
  (
    n143,
    n69
  );


  not
  g66
  (
    n234,
    n47
  );


  buf
  g67
  (
    n259,
    n49
  );


  not
  g68
  (
    n166,
    n33
  );


  buf
  g69
  (
    n121,
    n35
  );


  not
  g70
  (
    n157,
    n46
  );


  not
  g71
  (
    n119,
    n70
  );


  buf
  g72
  (
    n192,
    n72
  );


  not
  g73
  (
    n161,
    n75
  );


  buf
  g74
  (
    n172,
    n63
  );


  buf
  g75
  (
    n248,
    n76
  );


  buf
  g76
  (
    n233,
    n52
  );


  not
  g77
  (
    KeyWire_0_44,
    n61
  );


  not
  g78
  (
    n219,
    n54
  );


  not
  g79
  (
    n268,
    n41
  );


  buf
  g80
  (
    n140,
    n46
  );


  buf
  g81
  (
    n115,
    n56
  );


  buf
  g82
  (
    n98,
    n42
  );


  not
  g83
  (
    n230,
    n61
  );


  buf
  g84
  (
    n267,
    n38
  );


  buf
  g85
  (
    n227,
    n72
  );


  not
  g86
  (
    n271,
    n47
  );


  buf
  g87
  (
    n191,
    n43
  );


  not
  g88
  (
    n221,
    n77
  );


  buf
  g89
  (
    KeyWire_0_22,
    n72
  );


  buf
  g90
  (
    n262,
    n34
  );


  buf
  g91
  (
    KeyWire_0_16,
    n34
  );


  buf
  g92
  (
    n137,
    n76
  );


  buf
  g93
  (
    n214,
    n51
  );


  not
  g94
  (
    n218,
    n64
  );


  not
  g95
  (
    n266,
    n64
  );


  not
  g96
  (
    n171,
    n40
  );


  not
  g97
  (
    n158,
    n54
  );


  not
  g98
  (
    n111,
    n64
  );


  not
  g99
  (
    n141,
    n73
  );


  buf
  g100
  (
    n265,
    n61
  );


  not
  g101
  (
    KeyWire_0_6,
    n33
  );


  not
  g102
  (
    n208,
    n71
  );


  buf
  g103
  (
    n136,
    n36
  );


  buf
  g104
  (
    n132,
    n45
  );


  buf
  g105
  (
    n256,
    n41
  );


  not
  g106
  (
    KeyWire_0_32,
    n69
  );


  buf
  g107
  (
    n176,
    n52
  );


  buf
  g108
  (
    n103,
    n44
  );


  buf
  g109
  (
    n112,
    n63
  );


  buf
  g110
  (
    KeyWire_0_29,
    n52
  );


  buf
  g111
  (
    n255,
    n66
  );


  not
  g112
  (
    n181,
    n67
  );


  not
  g113
  (
    n144,
    n37
  );


  not
  g114
  (
    n225,
    n60
  );


  buf
  g115
  (
    n156,
    n77
  );


  buf
  g116
  (
    n153,
    n45
  );


  not
  g117
  (
    n224,
    n50
  );


  buf
  g118
  (
    n107,
    n68
  );


  buf
  g119
  (
    n142,
    n70
  );


  buf
  g120
  (
    KeyWire_0_11,
    n35
  );


  buf
  g121
  (
    n257,
    n56
  );


  buf
  g122
  (
    n247,
    n46
  );


  buf
  g123
  (
    n226,
    n65
  );


  not
  g124
  (
    n253,
    n53
  );


  not
  g125
  (
    n155,
    n76
  );


  buf
  g126
  (
    n239,
    n62
  );


  buf
  g127
  (
    n196,
    n69
  );


  buf
  g128
  (
    n201,
    n39
  );


  not
  g129
  (
    n231,
    n36
  );


  buf
  g130
  (
    n237,
    n49
  );


  buf
  g131
  (
    n215,
    n59
  );


  buf
  g132
  (
    n164,
    n78
  );


  not
  g133
  (
    n198,
    n67
  );


  buf
  g134
  (
    n110,
    n65
  );


  buf
  g135
  (
    n254,
    n54
  );


  buf
  g136
  (
    n236,
    n40
  );


  buf
  g137
  (
    n212,
    n57
  );


  not
  g138
  (
    n92,
    n57
  );


  not
  g139
  (
    n124,
    n48
  );


  buf
  g140
  (
    n206,
    n59
  );


  buf
  g141
  (
    n147,
    n43
  );


  not
  g142
  (
    n91,
    n43
  );


  buf
  g143
  (
    n246,
    n39
  );


  not
  g144
  (
    n95,
    n37
  );


  buf
  g145
  (
    n89,
    n66
  );


  not
  g146
  (
    n177,
    n44
  );


  not
  g147
  (
    n186,
    n63
  );


  not
  g148
  (
    n194,
    n65
  );


  not
  g149
  (
    n163,
    n73
  );


  buf
  g150
  (
    n129,
    n70
  );


  not
  g151
  (
    n252,
    n34
  );


  buf
  g152
  (
    n211,
    n75
  );


  buf
  g153
  (
    n96,
    n65
  );


  not
  g154
  (
    n204,
    n33
  );


  not
  g155
  (
    n240,
    n48
  );


  not
  g156
  (
    n199,
    n55
  );


  not
  g157
  (
    n106,
    n35
  );


  not
  g158
  (
    n258,
    n62
  );


  buf
  g159
  (
    n125,
    n58
  );


  buf
  g160
  (
    n229,
    n79
  );


  not
  g161
  (
    n169,
    n75
  );


  buf
  g162
  (
    n134,
    n48
  );


  buf
  g163
  (
    n184,
    n50
  );


  not
  g164
  (
    n193,
    n78
  );


  buf
  g165
  (
    KeyWire_0_3,
    n74
  );


  buf
  g166
  (
    n167,
    n74
  );


  buf
  g167
  (
    n108,
    n78
  );


  not
  g168
  (
    n272,
    n39
  );


  buf
  g169
  (
    n128,
    n53
  );


  not
  g170
  (
    KeyWire_0_27,
    n39
  );


  not
  g171
  (
    KeyWire_0_54,
    n36
  );


  not
  g172
  (
    n220,
    n45
  );


  not
  g173
  (
    n146,
    n40
  );


  not
  g174
  (
    n228,
    n73
  );


  not
  g175
  (
    n138,
    n55
  );


  buf
  g176
  (
    n205,
    n60
  );


  not
  g177
  (
    n242,
    n75
  );


  not
  g178
  (
    n145,
    n35
  );


  not
  g179
  (
    n245,
    n69
  );


  not
  g180
  (
    n165,
    n74
  );


  not
  g181
  (
    KeyWire_0_38,
    n34
  );


  buf
  g182
  (
    n150,
    n66
  );


  buf
  g183
  (
    n179,
    n47
  );


  buf
  g184
  (
    n94,
    n76
  );


  not
  g185
  (
    n270,
    n38
  );


  not
  g186
  (
    KeyWire_0_20,
    n70
  );


  buf
  g187
  (
    n202,
    n77
  );


  buf
  g188
  (
    n152,
    n73
  );


  not
  g189
  (
    n114,
    n63
  );


  not
  g190
  (
    n241,
    n72
  );


  buf
  g191
  (
    n148,
    n58
  );


  not
  g192
  (
    n232,
    n41
  );


  not
  g193
  (
    n210,
    n62
  );


  buf
  g194
  (
    n139,
    n40
  );


  buf
  g195
  (
    n113,
    n64
  );


  buf
  g196
  (
    n261,
    n37
  );


  not
  g197
  (
    n104,
    n51
  );


  buf
  g198
  (
    n126,
    n59
  );


  not
  g199
  (
    n178,
    n37
  );


  buf
  g200
  (
    n185,
    n50
  );


  not
  g201
  (
    n180,
    n45
  );


  not
  g202
  (
    n263,
    n71
  );


  buf
  g203
  (
    n100,
    n67
  );


  not
  g204
  (
    n189,
    n51
  );


  buf
  g205
  (
    n235,
    n41
  );


  buf
  g206
  (
    n264,
    n52
  );


  not
  g207
  (
    n200,
    n61
  );


  not
  g208
  (
    n131,
    n53
  );


  buf
  g209
  (
    n203,
    n62
  );


  buf
  g210
  (
    n182,
    n42
  );


  not
  g211
  (
    n162,
    n57
  );


  buf
  g212
  (
    n118,
    n57
  );


  not
  g213
  (
    n195,
    n68
  );


  not
  g214
  (
    n154,
    n71
  );


  not
  g215
  (
    n251,
    n47
  );


  not
  g216
  (
    n99,
    n43
  );


  not
  g217
  (
    n222,
    n68
  );


  not
  g218
  (
    KeyWire_0_55,
    n48
  );


  not
  g219
  (
    n151,
    n55
  );


  buf
  g220
  (
    n190,
    n33
  );


  buf
  g221
  (
    n123,
    n49
  );


  not
  g222
  (
    n269,
    n56
  );


  not
  g223
  (
    n101,
    n53
  );


  not
  g224
  (
    KeyWire_0_19,
    n78
  );


  not
  g225
  (
    n170,
    n51
  );


  buf
  g226
  (
    n160,
    n58
  );


  buf
  g227
  (
    n260,
    n74
  );


  buf
  g228
  (
    n207,
    n60
  );


  buf
  g229
  (
    n109,
    n49
  );


  buf
  g230
  (
    n102,
    n58
  );


  not
  g231
  (
    n183,
    n66
  );


  buf
  g232
  (
    n223,
    n46
  );


  buf
  g233
  (
    n213,
    n56
  );


  not
  g234
  (
    n209,
    n55
  );


  buf
  g235
  (
    n90,
    n42
  );


  buf
  g236
  (
    n173,
    n44
  );


  buf
  g237
  (
    KeyWire_0_35,
    n59
  );


  buf
  g238
  (
    n197,
    n42
  );


  not
  g239
  (
    n133,
    n38
  );


  not
  g240
  (
    n243,
    n54
  );


  buf
  g241
  (
    n274,
    n117
  );


  buf
  g242
  (
    n459,
    n92
  );


  not
  g243
  (
    n351,
    n161
  );


  buf
  g244
  (
    n362,
    n97
  );


  buf
  g245
  (
    n458,
    n128
  );


  buf
  g246
  (
    n468,
    n135
  );


  buf
  g247
  (
    n331,
    n170
  );


  not
  g248
  (
    n310,
    n94
  );


  not
  g249
  (
    n430,
    n95
  );


  buf
  g250
  (
    n332,
    n155
  );


  buf
  g251
  (
    n431,
    n132
  );


  buf
  g252
  (
    n318,
    n83
  );


  not
  g253
  (
    n360,
    n128
  );


  buf
  g254
  (
    n438,
    n113
  );


  buf
  g255
  (
    n382,
    n173
  );


  not
  g256
  (
    n314,
    n99
  );


  not
  g257
  (
    n413,
    n146
  );


  not
  g258
  (
    n330,
    n99
  );


  not
  g259
  (
    n423,
    n104
  );


  not
  g260
  (
    n427,
    n90
  );


  not
  g261
  (
    n343,
    n112
  );


  not
  g262
  (
    n444,
    n178
  );


  buf
  g263
  (
    n387,
    n123
  );


  buf
  g264
  (
    n346,
    n140
  );


  buf
  g265
  (
    n355,
    n141
  );


  not
  g266
  (
    n469,
    n159
  );


  not
  g267
  (
    n422,
    n175
  );


  buf
  g268
  (
    n398,
    n83
  );


  not
  g269
  (
    n340,
    n86
  );


  not
  g270
  (
    n363,
    n114
  );


  not
  g271
  (
    n471,
    n79
  );


  buf
  g272
  (
    n386,
    n115
  );


  not
  g273
  (
    n424,
    n90
  );


  not
  g274
  (
    n349,
    n160
  );


  not
  g275
  (
    n335,
    n139
  );


  not
  g276
  (
    n359,
    n147
  );


  not
  g277
  (
    n383,
    n146
  );


  not
  g278
  (
    n396,
    n135
  );


  buf
  g279
  (
    n462,
    n136
  );


  buf
  g280
  (
    n436,
    n98
  );


  buf
  g281
  (
    n277,
    n98
  );


  not
  g282
  (
    n411,
    n160
  );


  buf
  g283
  (
    n367,
    n169
  );


  buf
  g284
  (
    n279,
    n162
  );


  not
  g285
  (
    n389,
    n109
  );


  not
  g286
  (
    KeyWire_0_10,
    n175
  );


  buf
  g287
  (
    n385,
    n79
  );


  not
  g288
  (
    n364,
    n166
  );


  not
  g289
  (
    n442,
    n89
  );


  buf
  g290
  (
    n434,
    n101
  );


  buf
  g291
  (
    n309,
    n170
  );


  buf
  g292
  (
    n305,
    n107
  );


  not
  g293
  (
    n410,
    n115
  );


  buf
  g294
  (
    n446,
    n108
  );


  buf
  g295
  (
    n454,
    n81
  );


  buf
  g296
  (
    n376,
    n93
  );


  not
  g297
  (
    n302,
    n176
  );


  buf
  g298
  (
    n393,
    n96
  );


  buf
  g299
  (
    n317,
    n166
  );


  not
  g300
  (
    n447,
    n161
  );


  not
  g301
  (
    n347,
    n100
  );


  not
  g302
  (
    n381,
    n123
  );


  not
  g303
  (
    n306,
    n126
  );


  not
  g304
  (
    n403,
    n147
  );


  not
  g305
  (
    n361,
    n174
  );


  buf
  g306
  (
    n407,
    n154
  );


  buf
  g307
  (
    n370,
    n157
  );


  not
  g308
  (
    n416,
    n98
  );


  not
  g309
  (
    n320,
    n122
  );


  not
  g310
  (
    n448,
    n151
  );


  not
  g311
  (
    n365,
    n100
  );


  not
  g312
  (
    n378,
    n133
  );


  buf
  g313
  (
    n428,
    n163
  );


  not
  g314
  (
    n429,
    n101
  );


  not
  g315
  (
    n409,
    n152
  );


  buf
  g316
  (
    n420,
    n180
  );


  buf
  g317
  (
    n298,
    n108
  );


  not
  g318
  (
    n445,
    n153
  );


  buf
  g319
  (
    n329,
    n161
  );


  buf
  g320
  (
    n399,
    n166
  );


  not
  g321
  (
    n278,
    n137
  );


  buf
  g322
  (
    n450,
    n94
  );


  not
  g323
  (
    n457,
    n162
  );


  not
  g324
  (
    KeyWire_0_50,
    n161
  );


  buf
  g325
  (
    n350,
    n172
  );


  not
  g326
  (
    n415,
    n111
  );


  buf
  g327
  (
    n345,
    n131
  );


  buf
  g328
  (
    n290,
    n152
  );


  not
  g329
  (
    n325,
    n107
  );


  buf
  g330
  (
    n281,
    n134
  );


  buf
  g331
  (
    n327,
    n100
  );


  not
  g332
  (
    n275,
    n160
  );


  not
  g333
  (
    KeyWire_0_39,
    n123
  );


  not
  g334
  (
    n467,
    n98
  );


  not
  g335
  (
    n282,
    n150
  );


  buf
  g336
  (
    n377,
    n121
  );


  not
  g337
  (
    n342,
    n137
  );


  buf
  g338
  (
    n449,
    n84
  );


  not
  g339
  (
    n297,
    n175
  );


  buf
  g340
  (
    n285,
    n82
  );


  not
  g341
  (
    n316,
    n126
  );


  not
  g342
  (
    n313,
    n135
  );


  not
  g343
  (
    KeyWire_0_14,
    n82
  );


  not
  g344
  (
    n283,
    n152
  );


  not
  g345
  (
    n394,
    n92
  );


  buf
  g346
  (
    n443,
    n176
  );


  buf
  g347
  (
    n456,
    n153
  );


  not
  g348
  (
    n280,
    n85
  );


  buf
  g349
  (
    n287,
    n179
  );


  not
  g350
  (
    KeyWire_0_45,
    n109
  );


  buf
  g351
  (
    n291,
    n90
  );


  not
  g352
  (
    n372,
    n141
  );


  buf
  g353
  (
    n452,
    n170
  );


  not
  g354
  (
    n304,
    n119
  );


  not
  g355
  (
    KeyWire_0_60,
    n87
  );


  buf
  g356
  (
    n440,
    n121
  );


  not
  g357
  (
    n461,
    n174
  );


  buf
  g358
  (
    n293,
    n111
  );


  not
  g359
  (
    n402,
    n153
  );


  not
  g360
  (
    n336,
    n125
  );


  buf
  g361
  (
    n397,
    n176
  );


  buf
  g362
  (
    n315,
    n89
  );


  buf
  g363
  (
    n324,
    n151
  );


  buf
  g364
  (
    n466,
    n92
  );


  buf
  g365
  (
    n414,
    n117
  );


  buf
  g366
  (
    n333,
    n136
  );


  not
  g367
  (
    n354,
    n84
  );


  not
  g368
  (
    n375,
    n137
  );


  buf
  g369
  (
    n391,
    n101
  );


  not
  g370
  (
    n432,
    n101
  );


  buf
  g371
  (
    n453,
    n144
  );


  not
  g372
  (
    n288,
    n118
  );


  not
  g373
  (
    n388,
    n119
  );


  or
  g374
  (
    n353,
    n177,
    n142,
    n111
  );


  xnor
  g375
  (
    n451,
    n144,
    n145,
    n134,
    n97
  );


  or
  g376
  (
    n419,
    n165,
    n169,
    n136,
    n163
  );


  xnor
  g377
  (
    n356,
    n99,
    n116,
    n129,
    n140
  );


  xnor
  g378
  (
    n426,
    n154,
    n86,
    n131,
    n166
  );


  nor
  g379
  (
    n301,
    n149,
    n145,
    n163,
    n95
  );


  nand
  g380
  (
    n292,
    n107,
    n154,
    n124,
    n104
  );


  or
  g381
  (
    n463,
    n126,
    n180,
    n112,
    n160
  );


  nor
  g382
  (
    n379,
    n180,
    n155,
    n142,
    n117
  );


  nand
  g383
  (
    n406,
    n128,
    n122,
    n130,
    n126
  );


  xnor
  g384
  (
    n294,
    n135,
    n105,
    n138,
    n97
  );


  and
  g385
  (
    n401,
    n110,
    n149,
    n172
  );


  xor
  g386
  (
    n395,
    n179,
    n151,
    n150,
    n142
  );


  xor
  g387
  (
    KeyWire_0_56,
    n132,
    n142,
    n120,
    n82
  );


  nand
  g388
  (
    n439,
    n153,
    n157,
    n149,
    n177
  );


  and
  g389
  (
    n384,
    n119,
    n140,
    n141,
    n171
  );


  xor
  g390
  (
    n421,
    n118,
    n106,
    n112,
    n176
  );


  nand
  g391
  (
    n308,
    n173,
    n134,
    n156,
    n146
  );


  nand
  g392
  (
    n344,
    n157,
    n124,
    n105,
    n95
  );


  nor
  g393
  (
    n358,
    n167,
    n94,
    n130,
    n125
  );


  or
  g394
  (
    n404,
    n156,
    n162,
    n90,
    n118
  );


  and
  g395
  (
    n455,
    n164,
    n147,
    n84,
    n91
  );


  and
  g396
  (
    n312,
    n103,
    n110,
    n129,
    n86
  );


  xnor
  g397
  (
    n374,
    n154,
    n165,
    n141,
    n139
  );


  xnor
  g398
  (
    KeyWire_0_31,
    n148,
    n82,
    n94,
    n174
  );


  xor
  g399
  (
    n418,
    n145,
    n116,
    n102,
    n131
  );


  or
  g400
  (
    n417,
    n159,
    n107,
    n146,
    n114
  );


  and
  g401
  (
    n357,
    n103,
    n100,
    n89,
    n175
  );


  xnor
  g402
  (
    n307,
    n143,
    n127,
    n109,
    n114
  );


  nand
  g403
  (
    n366,
    n83,
    n96,
    n120,
    n139
  );


  nand
  g404
  (
    n284,
    n110,
    n164,
    n144,
    n158
  );


  xnor
  g405
  (
    n311,
    n121,
    n105,
    n162,
    n81
  );


  nand
  g406
  (
    n369,
    n179,
    n159,
    n151,
    n96
  );


  nor
  g407
  (
    n352,
    n96,
    n163,
    n177,
    n133
  );


  nand
  g408
  (
    n465,
    n165,
    n158,
    n106,
    n112
  );


  nor
  g409
  (
    n392,
    n178,
    n158,
    n93,
    n138
  );


  and
  g410
  (
    n334,
    n133,
    n167,
    n116,
    n149
  );


  xor
  g411
  (
    n441,
    n99,
    n108,
    n81,
    n106
  );


  nand
  g412
  (
    n321,
    n172,
    n122,
    n128,
    n147
  );


  nor
  g413
  (
    n435,
    n170,
    n113,
    n171,
    n139
  );


  xor
  g414
  (
    n470,
    n156,
    n81,
    n102,
    n134
  );


  xnor
  g415
  (
    n300,
    n143,
    n85,
    n102
  );


  nand
  g416
  (
    n322,
    n143,
    n150,
    n127,
    n123
  );


  xnor
  g417
  (
    n368,
    n125,
    n173,
    n155,
    n168
  );


  or
  g418
  (
    n437,
    n121,
    n132,
    n111,
    n155
  );


  nor
  g419
  (
    n460,
    n117,
    n115,
    n103,
    n127
  );


  xor
  g420
  (
    n473,
    n80,
    n165,
    n93,
    n113
  );


  or
  g421
  (
    n328,
    n168,
    n157,
    n97,
    n138
  );


  and
  g422
  (
    n464,
    n118,
    n125,
    n168,
    n103
  );


  nand
  g423
  (
    KeyWire_0_28,
    n136,
    n116,
    n124
  );


  or
  g424
  (
    KeyWire_0_46,
    n171,
    n130,
    n129,
    n91
  );


  xor
  g425
  (
    n289,
    n150,
    n148,
    n115,
    n91
  );


  or
  g426
  (
    n326,
    n169,
    n92,
    n168,
    n105
  );


  nor
  g427
  (
    n433,
    n148,
    n114,
    n120,
    n85
  );


  nor
  g428
  (
    n299,
    n130,
    n129,
    n110,
    n80
  );


  nand
  g429
  (
    n295,
    n79,
    n127,
    n152,
    n167
  );


  nor
  g430
  (
    n405,
    n102,
    n95,
    n164,
    n143
  );


  nand
  g431
  (
    n371,
    n86,
    n159,
    n156,
    n104
  );


  and
  g432
  (
    n303,
    n106,
    n87,
    n179,
    n104
  );


  nand
  g433
  (
    n296,
    n138,
    n177,
    n80,
    n174
  );


  xnor
  g434
  (
    n341,
    n93,
    n108,
    n120,
    n132
  );


  or
  g435
  (
    n408,
    n89,
    n171,
    n140,
    n178
  );


  xor
  g436
  (
    n390,
    n133,
    n83,
    n178,
    n167
  );


  xnor
  g437
  (
    n400,
    n148,
    n122,
    n158,
    n80
  );


  and
  g438
  (
    n425,
    n169,
    n131,
    n119,
    n137
  );


  nor
  g439
  (
    n348,
    n113,
    n84,
    n173,
    n164
  );


  nor
  g440
  (
    n339,
    n145,
    n109,
    n91,
    n144
  );


  not
  g441
  (
    n615,
    n241
  );


  buf
  g442
  (
    n539,
    n377
  );


  not
  g443
  (
    n552,
    n245
  );


  not
  g444
  (
    n493,
    n240
  );


  not
  g445
  (
    n559,
    n233
  );


  not
  g446
  (
    n517,
    n184
  );


  not
  g447
  (
    n635,
    n395
  );


  buf
  g448
  (
    n495,
    n212
  );


  buf
  g449
  (
    n543,
    n270
  );


  not
  g450
  (
    n488,
    n259
  );


  buf
  g451
  (
    n581,
    n310
  );


  buf
  g452
  (
    n551,
    n367
  );


  buf
  g453
  (
    KeyWire_0_5,
    n228
  );


  not
  g454
  (
    n499,
    n250
  );


  buf
  g455
  (
    n501,
    n422
  );


  not
  g456
  (
    n476,
    n384
  );


  buf
  g457
  (
    n516,
    n205
  );


  buf
  g458
  (
    n546,
    n237
  );


  not
  g459
  (
    KeyWire_0_30,
    n189
  );


  not
  g460
  (
    n491,
    n205
  );


  buf
  g461
  (
    n528,
    n323
  );


  buf
  g462
  (
    n512,
    n366
  );


  not
  g463
  (
    n497,
    n184
  );


  buf
  g464
  (
    n579,
    n215
  );


  not
  g465
  (
    n569,
    n187
  );


  buf
  g466
  (
    n554,
    n227
  );


  not
  g467
  (
    n498,
    n231
  );


  buf
  g468
  (
    n519,
    n226
  );


  not
  g469
  (
    n636,
    n359
  );


  not
  g470
  (
    n607,
    n220
  );


  not
  g471
  (
    n475,
    n219
  );


  buf
  g472
  (
    n563,
    n224
  );


  buf
  g473
  (
    n606,
    n321
  );


  not
  g474
  (
    n614,
    n266
  );


  buf
  g475
  (
    n507,
    n249
  );


  buf
  g476
  (
    KeyWire_0_4,
    n244
  );


  not
  g477
  (
    n595,
    n421
  );


  buf
  g478
  (
    n537,
    n233
  );


  not
  g479
  (
    n618,
    n373
  );


  not
  g480
  (
    n490,
    n196
  );


  buf
  g481
  (
    n556,
    n238
  );


  buf
  g482
  (
    KeyWire_0_23,
    n197
  );


  buf
  g483
  (
    n483,
    n215
  );


  not
  g484
  (
    n631,
    n278
  );


  or
  g485
  (
    n584,
    n225,
    n185,
    n248
  );


  nor
  g486
  (
    n496,
    n191,
    n236,
    n192,
    n255
  );


  nand
  g487
  (
    n515,
    n260,
    n194,
    n195,
    n222
  );


  xor
  g488
  (
    n624,
    n200,
    n193,
    n192,
    n218
  );


  nor
  g489
  (
    n587,
    n255,
    n261,
    n250,
    n197
  );


  nor
  g490
  (
    n638,
    n237,
    n341,
    n198,
    n426
  );


  nand
  g491
  (
    n575,
    n230,
    n241,
    n398,
    n265
  );


  and
  g492
  (
    n542,
    n226,
    n216,
    n240,
    n268
  );


  nor
  g493
  (
    n536,
    n316,
    n426,
    n194,
    n285
  );


  and
  g494
  (
    n576,
    n232,
    n212,
    n249,
    n258
  );


  nand
  g495
  (
    n592,
    n224,
    n214,
    n187,
    n222
  );


  and
  g496
  (
    n520,
    n407,
    n206,
    n304,
    n218
  );


  xnor
  g497
  (
    n599,
    n302,
    n355,
    n275,
    n263
  );


  or
  g498
  (
    n530,
    n250,
    n263,
    n252,
    n203
  );


  nand
  g499
  (
    n583,
    n269,
    n257,
    n191,
    n252
  );


  xor
  g500
  (
    n524,
    n192,
    n268,
    n428,
    n208
  );


  or
  g501
  (
    n600,
    n213,
    n225,
    n265,
    n389
  );


  nor
  g502
  (
    n526,
    n201,
    n239,
    n295,
    n391
  );


  nand
  g503
  (
    n521,
    n257,
    n303,
    n267,
    n203
  );


  nand
  g504
  (
    n523,
    n343,
    n217,
    n210,
    n252
  );


  xnor
  g505
  (
    n608,
    n269,
    n260,
    n277,
    n338
  );


  and
  g506
  (
    n605,
    n426,
    n353,
    n234,
    n385
  );


  and
  g507
  (
    n590,
    n192,
    n187,
    n280,
    n320
  );


  or
  g508
  (
    n588,
    n183,
    n270,
    n246,
    n223
  );


  nand
  g509
  (
    n562,
    n235,
    n182,
    n219,
    n188
  );


  or
  g510
  (
    n482,
    n217,
    n257,
    n261,
    n208
  );


  xnor
  g511
  (
    n601,
    n247,
    n229,
    n248,
    n348
  );


  xor
  g512
  (
    n564,
    n202,
    n311,
    n264,
    n245
  );


  xnor
  g513
  (
    n508,
    n256,
    n204,
    n403,
    n227
  );


  nand
  g514
  (
    KeyWire_0_62,
    n260,
    n418,
    n186,
    n349
  );


  xor
  g515
  (
    n479,
    n284,
    n262,
    n228,
    n181
  );


  xnor
  g516
  (
    n548,
    n269,
    n427,
    n229,
    n354
  );


  xnor
  g517
  (
    n506,
    n419,
    n339,
    n221,
    n224
  );


  nor
  g518
  (
    n620,
    n404,
    n345,
    n257,
    n242
  );


  and
  g519
  (
    n541,
    n314,
    n219,
    n394,
    n232
  );


  and
  g520
  (
    n609,
    n202,
    n416,
    n209,
    n322
  );


  xor
  g521
  (
    n544,
    n234,
    n397,
    n258,
    n390
  );


  nand
  g522
  (
    KeyWire_0_2,
    n267,
    n211,
    n427,
    n221
  );


  and
  g523
  (
    n547,
    n235,
    n412,
    n414,
    n261
  );


  or
  g524
  (
    n582,
    n283,
    n324,
    n374,
    n211
  );


  xor
  g525
  (
    n586,
    n350,
    n294,
    n265,
    n335
  );


  nand
  g526
  (
    n555,
    n423,
    n263,
    n370,
    n251
  );


  and
  g527
  (
    KeyWire_0_25,
    n301,
    n193,
    n220,
    n229
  );


  or
  g528
  (
    KeyWire_0_21,
    n246,
    n382,
    n238,
    n251
  );


  nor
  g529
  (
    n550,
    n182,
    n427,
    n259,
    n245
  );


  xor
  g530
  (
    n572,
    n207,
    n368,
    n342,
    n240
  );


  xnor
  g531
  (
    n513,
    n227,
    n249,
    n372,
    n230
  );


  and
  g532
  (
    n589,
    n319,
    n182,
    n198,
    n186
  );


  or
  g533
  (
    KeyWire_0_61,
    n336,
    n361,
    n215,
    n264
  );


  and
  g534
  (
    n558,
    n282,
    n402,
    n228,
    n246
  );


  nor
  g535
  (
    n486,
    n234,
    n270,
    n190,
    n219
  );


  nand
  g536
  (
    n478,
    n190,
    n236,
    n363,
    n213
  );


  nor
  g537
  (
    n484,
    n194,
    n191,
    n378,
    n427
  );


  nor
  g538
  (
    n527,
    n400,
    n202,
    n223,
    n351
  );


  and
  g539
  (
    n492,
    n248,
    n279,
    n268,
    n189
  );


  or
  g540
  (
    n617,
    n194,
    n410,
    n241,
    n231
  );


  xor
  g541
  (
    n574,
    n239,
    n196,
    n199,
    n243
  );


  or
  g542
  (
    n594,
    n247,
    n369,
    n250,
    n364
  );


  nand
  g543
  (
    n621,
    n216,
    n288,
    n274,
    n212
  );


  nor
  g544
  (
    n634,
    n293,
    n276,
    n297,
    n189
  );


  xnor
  g545
  (
    n494,
    n259,
    n239,
    n428,
    n331
  );


  nor
  g546
  (
    n613,
    n281,
    n210,
    n188,
    n185
  );


  or
  g547
  (
    n502,
    n232,
    n228,
    n287,
    n207
  );


  nor
  g548
  (
    n623,
    n200,
    n216,
    n408,
    n286
  );


  xor
  g549
  (
    n626,
    n264,
    n203,
    n296,
    n291
  );


  xnor
  g550
  (
    n510,
    n263,
    n213,
    n199,
    n233
  );


  nand
  g551
  (
    n509,
    n217,
    n269,
    n208,
    n386
  );


  and
  g552
  (
    n532,
    n332,
    n218,
    n204,
    n326
  );


  and
  g553
  (
    n632,
    n191,
    n379,
    n241,
    n337
  );


  and
  g554
  (
    n598,
    n251,
    n198,
    n242,
    n267
  );


  nor
  g555
  (
    n570,
    n204,
    n222,
    n211,
    n392
  );


  nand
  g556
  (
    n568,
    n195,
    n388,
    n212,
    n357
  );


  and
  g557
  (
    n629,
    n266,
    n195,
    n214,
    n254
  );


  xnor
  g558
  (
    n578,
    n318,
    n193,
    n426,
    n333
  );


  xor
  g559
  (
    n511,
    n204,
    n387,
    n259,
    n218
  );


  xor
  g560
  (
    n560,
    n189,
    n181,
    n223,
    n305
  );


  xnor
  g561
  (
    n610,
    n184,
    n185,
    n265,
    n222
  );


  nor
  g562
  (
    n487,
    n185,
    n196,
    n425,
    n190
  );


  nor
  g563
  (
    n481,
    n417,
    n201,
    n254,
    n267
  );


  or
  g564
  (
    n565,
    n188,
    n356,
    n328,
    n182
  );


  nand
  g565
  (
    n616,
    n327,
    n220,
    n183,
    n334
  );


  xnor
  g566
  (
    KeyWire_0_58,
    n196,
    n245,
    n198,
    n239
  );


  xnor
  g567
  (
    n529,
    n290,
    n230,
    n225,
    n205
  );


  xor
  g568
  (
    n611,
    n217,
    n214,
    n413,
    n210
  );


  xnor
  g569
  (
    n597,
    n200,
    n298,
    n424,
    n238
  );


  or
  g570
  (
    n549,
    n188,
    n184,
    n200,
    n292
  );


  xor
  g571
  (
    n514,
    n247,
    n225,
    n365,
    n362
  );


  xor
  g572
  (
    n522,
    n202,
    n262,
    n243
  );


  and
  g573
  (
    n553,
    n313,
    n258,
    n183,
    n307
  );


  and
  g574
  (
    n557,
    n264,
    n230,
    n209,
    n396
  );


  xnor
  g575
  (
    n573,
    n266,
    n375,
    n243,
    n236
  );


  and
  g576
  (
    n580,
    n253,
    n399,
    n308,
    n199
  );


  nand
  g577
  (
    n625,
    n206,
    n201,
    n330,
    n220
  );


  xor
  g578
  (
    n622,
    n195,
    n221,
    n216,
    n381
  );


  xor
  g579
  (
    KeyWire_0_8,
    n262,
    n244,
    n344,
    n223
  );


  xor
  g580
  (
    n477,
    n231,
    n317,
    n197,
    n289
  );


  nor
  g581
  (
    n518,
    n240,
    n358,
    n235,
    n411
  );


  or
  g582
  (
    n604,
    n306,
    n181,
    n315,
    n258
  );


  and
  g583
  (
    n533,
    n300,
    n254,
    n207,
    n201
  );


  nor
  g584
  (
    n585,
    n233,
    n347,
    n213,
    n380
  );


  or
  g585
  (
    n500,
    n203,
    n208,
    n346,
    n237
  );


  xnor
  g586
  (
    n485,
    n207,
    n424,
    n193,
    n260
  );


  or
  g587
  (
    n577,
    n209,
    n236,
    n234,
    n340
  );


  xor
  g588
  (
    n540,
    n190,
    n253,
    n405,
    n211
  );


  nor
  g589
  (
    n503,
    n242,
    n325,
    n401,
    n425
  );


  nor
  g590
  (
    n630,
    n209,
    n197,
    n299,
    n252
  );


  nor
  g591
  (
    n596,
    n235,
    n237,
    n205,
    n253
  );


  nand
  g592
  (
    n567,
    n180,
    n221,
    n266,
    n262
  );


  xor
  g593
  (
    n637,
    n246,
    n186,
    n210,
    n270
  );


  and
  g594
  (
    n561,
    n181,
    n271,
    n309,
    n360
  );


  nand
  g595
  (
    n480,
    n183,
    n255,
    n242,
    n244
  );


  or
  g596
  (
    n612,
    n253,
    n256,
    n393,
    n238
  );


  xor
  g597
  (
    n603,
    n186,
    n415,
    n206,
    n226
  );


  xor
  g598
  (
    n619,
    n261,
    n312,
    n247,
    n215
  );


  and
  g599
  (
    n531,
    n206,
    n244,
    n329,
    n254
  );


  or
  g600
  (
    n504,
    n199,
    n268,
    n352,
    n428
  );


  nor
  g601
  (
    n627,
    n226,
    n406,
    n251,
    n371
  );


  xor
  g602
  (
    n602,
    n187,
    n376,
    n255,
    n224
  );


  and
  g603
  (
    KeyWire_0_36,
    n256,
    n227,
    n420,
    n249
  );


  nor
  g604
  (
    n545,
    n383,
    n409,
    n214,
    n229
  );


  xnor
  g605
  (
    n535,
    n232,
    n256,
    n248,
    n231
  );


  or
  g606
  (
    n652,
    n430,
    n478
  );


  xnor
  g607
  (
    n649,
    n455,
    n447,
    n499,
    n431
  );


  nand
  g608
  (
    n670,
    n454,
    n489,
    n443,
    n440
  );


  nor
  g609
  (
    n655,
    n452,
    n475,
    n437,
    n497
  );


  xnor
  g610
  (
    n658,
    n429,
    n510,
    n455,
    n442
  );


  xnor
  g611
  (
    n646,
    n433,
    n430,
    n441,
    n458
  );


  nand
  g612
  (
    n654,
    n451,
    n450,
    n456,
    n458
  );


  nand
  g613
  (
    KeyWire_0_15,
    n445,
    n450,
    n431,
    n447
  );


  xnor
  g614
  (
    n651,
    n459,
    n447,
    n504,
    n438
  );


  nor
  g615
  (
    n640,
    n438,
    n432,
    n516
  );


  nor
  g616
  (
    n650,
    n460,
    n456,
    n496,
    n431
  );


  or
  g617
  (
    n678,
    n455,
    n457,
    n435,
    n451
  );


  nor
  g618
  (
    n660,
    n444,
    n455,
    n458,
    n433
  );


  and
  g619
  (
    KeyWire_0_53,
    n432,
    n507,
    n437
  );


  xor
  g620
  (
    n648,
    n434,
    n517,
    n433,
    n482
  );


  nor
  g621
  (
    n671,
    n454,
    n453,
    n452,
    n436
  );


  xnor
  g622
  (
    n667,
    n435,
    n441,
    n485,
    n487
  );


  or
  g623
  (
    n676,
    n459,
    n454,
    n450,
    n480
  );


  xor
  g624
  (
    n664,
    n434,
    n445,
    n429,
    n446
  );


  xnor
  g625
  (
    n669,
    n498,
    n445,
    n451,
    n448
  );


  nor
  g626
  (
    n662,
    n439,
    n491,
    n438,
    n484
  );


  or
  g627
  (
    n673,
    n442,
    n435,
    n474,
    n440
  );


  or
  g628
  (
    KeyWire_0_13,
    n495,
    n451,
    n437,
    n457
  );


  xnor
  g629
  (
    n675,
    n436,
    n456,
    n481,
    n503
  );


  nor
  g630
  (
    n661,
    n448,
    n439,
    n444,
    n442
  );


  and
  g631
  (
    KeyWire_0_42,
    n460,
    n515,
    n505,
    n458
  );


  nor
  g632
  (
    n672,
    n443,
    n452,
    n440,
    n429
  );


  or
  g633
  (
    n679,
    n441,
    n460,
    n443,
    n486
  );


  nand
  g634
  (
    n663,
    n449,
    n479,
    n436,
    n461
  );


  and
  g635
  (
    n657,
    n501,
    n449,
    n444,
    n441
  );


  and
  g636
  (
    n643,
    n509,
    n444,
    n454,
    n453
  );


  xnor
  g637
  (
    n665,
    n431,
    n446,
    n506,
    n447
  );


  nand
  g638
  (
    n682,
    n460,
    n446,
    n453,
    n476
  );


  or
  g639
  (
    n641,
    n434,
    n459,
    n492,
    n477
  );


  xor
  g640
  (
    n668,
    n512,
    n449,
    n433,
    n453
  );


  or
  g641
  (
    n681,
    n438,
    n430,
    n450,
    n436
  );


  nand
  g642
  (
    KeyWire_0_34,
    n439,
    n448,
    n456,
    n500
  );


  nand
  g643
  (
    n642,
    n439,
    n430,
    n443,
    n442
  );


  xor
  g644
  (
    n674,
    n428,
    n508,
    n445,
    n440
  );


  xor
  g645
  (
    n659,
    n446,
    n494,
    n449,
    n483
  );


  nor
  g646
  (
    n677,
    n429,
    n514,
    n488,
    n459
  );


  and
  g647
  (
    n647,
    n448,
    n435,
    n502,
    n490
  );


  or
  g648
  (
    n666,
    n513,
    n457,
    n434,
    n511
  );


  nor
  g649
  (
    n645,
    n432,
    n493,
    n452,
    n457
  );


  xor
  g650
  (
    n723,
    n625,
    n535,
    n577,
    n588
  );


  and
  g651
  (
    n702,
    n623,
    n605,
    n650,
    n644
  );


  or
  g652
  (
    n750,
    n561,
    n653,
    n570
  );


  or
  g653
  (
    n757,
    n526,
    n563,
    n581,
    n647
  );


  or
  g654
  (
    n748,
    n611,
    n639,
    n525,
    n606
  );


  or
  g655
  (
    n686,
    n640,
    n627,
    n578,
    n612
  );


  nor
  g656
  (
    n739,
    n576,
    n560,
    n645,
    n639
  );


  xnor
  g657
  (
    n698,
    n528,
    n560,
    n625,
    n631
  );


  nand
  g658
  (
    n684,
    n623,
    n659,
    n640,
    n604
  );


  xor
  g659
  (
    n764,
    n577,
    n554,
    n590,
    n656
  );


  and
  g660
  (
    n695,
    n569,
    n639,
    n622,
    n586
  );


  xor
  g661
  (
    n760,
    n574,
    n574,
    n597,
    n648
  );


  or
  g662
  (
    n732,
    n610,
    n660,
    n571,
    n620
  );


  xnor
  g663
  (
    n749,
    n596,
    n612,
    n630,
    n609
  );


  xnor
  g664
  (
    n711,
    n626,
    n580,
    n647,
    n630
  );


  nor
  g665
  (
    n768,
    n598,
    n646,
    n613,
    n622
  );


  or
  g666
  (
    n759,
    n616,
    n608,
    n634,
    n606
  );


  xor
  g667
  (
    n755,
    n566,
    n538,
    n632,
    n642
  );


  and
  g668
  (
    n713,
    n645,
    n618,
    n608,
    n615
  );


  and
  g669
  (
    n719,
    n630,
    n594,
    n653,
    n584
  );


  nand
  g670
  (
    n693,
    n547,
    n630,
    n631,
    n617
  );


  or
  g671
  (
    n687,
    n520,
    n631,
    n649,
    n635
  );


  xnor
  g672
  (
    n700,
    n603,
    n611,
    n559,
    n605
  );


  and
  g673
  (
    n712,
    n579,
    n566,
    n645,
    n584
  );


  or
  g674
  (
    n741,
    n650,
    n580,
    n583,
    n620
  );


  or
  g675
  (
    n722,
    n606,
    n657,
    n650,
    n558
  );


  nor
  g676
  (
    n716,
    n644,
    n558,
    n616,
    n572
  );


  and
  g677
  (
    n726,
    n591,
    n655,
    n629,
    n643
  );


  and
  g678
  (
    n756,
    n628,
    n621,
    n564,
    n565
  );


  nand
  g679
  (
    n699,
    n658,
    n620,
    n568
  );


  nor
  g680
  (
    n697,
    n641,
    n657,
    n565
  );


  and
  g681
  (
    n761,
    n575,
    n619,
    n631,
    n593
  );


  and
  g682
  (
    n769,
    n562,
    n593,
    n658,
    n552
  );


  or
  g683
  (
    n689,
    n615,
    n625,
    n633,
    n567
  );


  or
  g684
  (
    n767,
    n654,
    n642,
    n644,
    n651
  );


  xnor
  g685
  (
    n730,
    n602,
    n626,
    n627,
    n659
  );


  nor
  g686
  (
    n692,
    n555,
    n621,
    n649,
    n647
  );


  nor
  g687
  (
    n737,
    n572,
    n607,
    n660
  );


  nand
  g688
  (
    n685,
    n607,
    n616,
    n650,
    n530
  );


  xnor
  g689
  (
    n733,
    n600,
    n643,
    n573,
    n653
  );


  xor
  g690
  (
    n727,
    n656,
    n622,
    n578,
    n628
  );


  nor
  g691
  (
    n706,
    n614,
    n591,
    n563,
    n627
  );


  xnor
  g692
  (
    n683,
    n562,
    n613,
    n634,
    n575
  );


  or
  g693
  (
    n740,
    n587,
    n629,
    n592,
    n615
  );


  xnor
  g694
  (
    n744,
    n621,
    n628,
    n594,
    n541
  );


  xor
  g695
  (
    n766,
    n648,
    n553,
    n570,
    n523
  );


  xor
  g696
  (
    n717,
    n610,
    n606,
    n640,
    n651
  );


  and
  g697
  (
    n731,
    n641,
    n618,
    n536,
    n592
  );


  nand
  g698
  (
    n728,
    n583,
    n648,
    n617
  );


  nor
  g699
  (
    n688,
    n581,
    n534,
    n597,
    n654
  );


  xor
  g700
  (
    n762,
    n548,
    n620,
    n660,
    n586
  );


  nor
  g701
  (
    n747,
    n564,
    n622,
    n557,
    n646
  );


  nor
  g702
  (
    n734,
    n599,
    n550,
    n614,
    n655
  );


  nor
  g703
  (
    n746,
    n540,
    n602,
    n652,
    n614
  );


  xor
  g704
  (
    n751,
    n604,
    n641,
    n655,
    n539
  );


  nor
  g705
  (
    n708,
    n652,
    n624,
    n582,
    n555
  );


  and
  g706
  (
    n701,
    n626,
    n576,
    n643,
    n654
  );


  and
  g707
  (
    n754,
    n609,
    n613,
    n611,
    n623
  );


  nand
  g708
  (
    n714,
    n642,
    n646,
    n573,
    n656
  );


  or
  g709
  (
    KeyWire_0_41,
    n543,
    n644,
    n527,
    n619
  );


  xor
  g710
  (
    n691,
    n571,
    n604,
    n612,
    n633
  );


  or
  g711
  (
    n721,
    n652,
    n569,
    n561,
    n589
  );


  nor
  g712
  (
    n738,
    n628,
    n596,
    n518,
    n579
  );


  or
  g713
  (
    n715,
    n646,
    n521,
    n542,
    n598
  );


  nor
  g714
  (
    n724,
    n601,
    n595,
    n546,
    n633
  );


  and
  g715
  (
    n763,
    n588,
    n608,
    n519,
    n651
  );


  xnor
  g716
  (
    n707,
    n626,
    n634,
    n589,
    n654
  );


  nor
  g717
  (
    KeyWire_0_12,
    n624,
    n615,
    n595,
    n609
  );


  xnor
  g718
  (
    n709,
    n551,
    n585,
    n624,
    n655
  );


  nor
  g719
  (
    n736,
    n640,
    n554,
    n643,
    n600
  );


  or
  g720
  (
    n752,
    n649,
    n651,
    n618,
    n614
  );


  nor
  g721
  (
    n729,
    n599,
    n617,
    n610,
    n607
  );


  nor
  g722
  (
    n703,
    n549,
    n632,
    n639,
    n647
  );


  and
  g723
  (
    n704,
    n618,
    n621,
    n629,
    n617
  );


  nor
  g724
  (
    KeyWire_0_7,
    n601,
    n619,
    n623,
    n559
  );


  nor
  g725
  (
    n753,
    n627,
    n556,
    n633
  );


  nand
  g726
  (
    n765,
    n616,
    n642,
    n659,
    n582
  );


  xnor
  g727
  (
    n735,
    n533,
    n652,
    n641,
    n529
  );


  and
  g728
  (
    n742,
    n605,
    n613,
    n658,
    n537
  );


  and
  g729
  (
    n690,
    n657,
    n544,
    n619,
    n632
  );


  xnor
  g730
  (
    n710,
    n524,
    n590,
    n567,
    n604
  );


  xor
  g731
  (
    n705,
    n645,
    n608,
    n605,
    n649
  );


  xor
  g732
  (
    n694,
    n545,
    n611,
    n587,
    n557
  );


  xor
  g733
  (
    n745,
    n629,
    n656,
    n625,
    n609
  );


  xnor
  g734
  (
    n696,
    n610,
    n522,
    n658,
    n585
  );


  xnor
  g735
  (
    n758,
    n659,
    n632,
    n531,
    n612
  );


  xnor
  g736
  (
    n743,
    n634,
    n532,
    n624,
    n603
  );


  xor
  g737
  (
    KeyWire_0_17,
    n665,
    n664,
    n689,
    n672
  );


  xor
  g738
  (
    n784,
    n697,
    n695,
    n661,
    n670
  );


  xnor
  g739
  (
    n780,
    n663,
    n672,
    n665,
    n666
  );


  nor
  g740
  (
    n781,
    n670,
    n661,
    n664,
    n671
  );


  nor
  g741
  (
    n772,
    n666,
    n665,
    n685,
    n693
  );


  and
  g742
  (
    n774,
    n694,
    n661,
    n667,
    n665
  );


  xor
  g743
  (
    n783,
    n672,
    n667,
    n662,
    n668
  );


  xnor
  g744
  (
    KeyWire_0_47,
    n688,
    n692,
    n671,
    n662
  );


  or
  g745
  (
    n785,
    n669,
    n669,
    n690,
    n663
  );


  xnor
  g746
  (
    n782,
    n664,
    n670,
    n668
  );


  nor
  g747
  (
    n770,
    n669,
    n691,
    n687,
    n668
  );


  xor
  g748
  (
    n778,
    n671,
    n684,
    n669,
    n660
  );


  nor
  g749
  (
    n776,
    n663,
    n667,
    n671,
    n686
  );


  or
  g750
  (
    n779,
    n698,
    n662,
    n666
  );


  nor
  g751
  (
    n775,
    n663,
    n664,
    n668,
    n662
  );


  xnor
  g752
  (
    n773,
    n667,
    n696,
    n683,
    n661
  );


  nor
  g753
  (
    n788,
    n773,
    n770,
    n771,
    n701
  );


  xor
  g754
  (
    n789,
    n707,
    n710,
    n700,
    n709
  );


  xnor
  g755
  (
    n786,
    n706,
    n699,
    n702,
    n705
  );


  xor
  g756
  (
    n787,
    n708,
    n704,
    n703,
    n772
  );


  xor
  g757
  (
    n795,
    n677,
    n787,
    n721,
    n675
  );


  nand
  g758
  (
    n800,
    n674,
    n717,
    n673,
    n672
  );


  nor
  g759
  (
    n792,
    n673,
    n673,
    n676,
    n713
  );


  nor
  g760
  (
    n790,
    n788,
    n674,
    n728,
    n675
  );


  nor
  g761
  (
    n794,
    n675,
    n788,
    n786,
    n727
  );


  nand
  g762
  (
    n796,
    n724,
    n726,
    n719,
    n676
  );


  or
  g763
  (
    n798,
    n673,
    n786,
    n674
  );


  xnor
  g764
  (
    n799,
    n789,
    n675,
    n788,
    n786
  );


  nor
  g765
  (
    n791,
    n715,
    n711,
    n720,
    n718
  );


  xor
  g766
  (
    n793,
    n788,
    n722,
    n786,
    n787
  );


  and
  g767
  (
    n797,
    n787,
    n677,
    n676
  );


  xnor
  g768
  (
    n801,
    n676,
    n787,
    n712,
    n716
  );


  nor
  g769
  (
    n802,
    n729,
    n725,
    n714,
    n723
  );


  not
  g770
  (
    n822,
    n797
  );


  not
  g771
  (
    n804,
    n793
  );


  buf
  g772
  (
    n807,
    n794
  );


  not
  g773
  (
    n825,
    n798
  );


  not
  g774
  (
    n812,
    n677
  );


  buf
  g775
  (
    n824,
    n800
  );


  buf
  g776
  (
    n806,
    n797
  );


  buf
  g777
  (
    n810,
    n730
  );


  buf
  g778
  (
    n819,
    n461
  );


  buf
  g779
  (
    n809,
    n790
  );


  buf
  g780
  (
    n815,
    n798
  );


  buf
  g781
  (
    n821,
    n796
  );


  buf
  g782
  (
    n803,
    n799
  );


  buf
  g783
  (
    n818,
    n798
  );


  not
  g784
  (
    n811,
    n800
  );


  not
  g785
  (
    n808,
    n797
  );


  buf
  g786
  (
    n820,
    n799
  );


  not
  g787
  (
    n826,
    n789
  );


  buf
  g788
  (
    n816,
    n795
  );


  not
  g789
  (
    n813,
    n799
  );


  not
  g790
  (
    n814,
    n789
  );


  xnor
  g791
  (
    n823,
    n789,
    n798,
    n800,
    n797
  );


  xor
  g792
  (
    n817,
    n795,
    n796,
    n461,
    n792
  );


  xnor
  g793
  (
    n805,
    n462,
    n461,
    n799,
    n791
  );


  xor
  g794
  (
    n828,
    n803,
    n801
  );


  nand
  g795
  (
    n827,
    n801,
    n802,
    n800,
    n803
  );


  nor
  g796
  (
    n829,
    n803,
    n827
  );


  buf
  g797
  (
    n832,
    n804
  );


  nand
  g798
  (
    n831,
    n829,
    n805
  );


  and
  g799
  (
    n833,
    n804,
    n829
  );


  nor
  g800
  (
    n830,
    n829,
    n829,
    n804,
    n803
  );


  not
  g801
  (
    n837,
    n831
  );


  buf
  g802
  (
    n842,
    n833
  );


  buf
  g803
  (
    n836,
    n832
  );


  not
  g804
  (
    n845,
    n831
  );


  buf
  g805
  (
    KeyWire_0_63,
    n805
  );


  buf
  g806
  (
    n847,
    n832
  );


  not
  g807
  (
    n844,
    n831
  );


  not
  g808
  (
    n841,
    n830
  );


  buf
  g809
  (
    n843,
    n833
  );


  buf
  g810
  (
    n835,
    n830
  );


  buf
  g811
  (
    n846,
    n805
  );


  buf
  g812
  (
    n839,
    n833
  );


  xor
  g813
  (
    n838,
    n830,
    n832
  );


  and
  g814
  (
    n848,
    n805,
    n832
  );


  nor
  g815
  (
    n834,
    n830,
    n831
  );


  nand
  g816
  (
    n866,
    n465,
    n816,
    n271
  );


  and
  g817
  (
    n867,
    n816,
    n835,
    n784
  );


  and
  g818
  (
    n877,
    n812,
    n844,
    n748
  );


  and
  g819
  (
    n881,
    n840,
    n808,
    n745
  );


  and
  g820
  (
    n885,
    n844,
    n464,
    n838
  );


  and
  g821
  (
    n849,
    n839,
    n809,
    n678
  );


  or
  g822
  (
    n894,
    n835,
    n814,
    n839
  );


  nor
  g823
  (
    KeyWire_0_52,
    n731,
    n843,
    n678
  );


  or
  g824
  (
    n893,
    n813,
    n811,
    n465
  );


  nor
  g825
  (
    n861,
    n811,
    n818,
    n271
  );


  or
  g826
  (
    n859,
    n740,
    n746,
    n813
  );


  xor
  g827
  (
    n853,
    n844,
    n816,
    n835
  );


  or
  g828
  (
    n890,
    n810,
    n833,
    n742
  );


  nor
  g829
  (
    n883,
    n734,
    n732,
    n842
  );


  xor
  g830
  (
    n863,
    n785,
    n735,
    n783
  );


  nor
  g831
  (
    n857,
    n272,
    n750,
    n814
  );


  xor
  g832
  (
    n872,
    n806,
    n844,
    n820,
    n842
  );


  nor
  g833
  (
    n887,
    n744,
    n828,
    n817,
    n272
  );


  or
  g834
  (
    n852,
    n837,
    n733,
    n807,
    n815
  );


  nand
  g835
  (
    n871,
    n815,
    n812,
    n813,
    n838
  );


  or
  g836
  (
    n850,
    n836,
    n842,
    n464,
    n813
  );


  nor
  g837
  (
    n870,
    n840,
    n816,
    n841
  );


  or
  g838
  (
    n865,
    n818,
    n811,
    n834,
    n802
  );


  xnor
  g839
  (
    n874,
    n838,
    n837,
    n743,
    n781
  );


  or
  g840
  (
    n886,
    n819,
    n838,
    n463,
    n779
  );


  xnor
  g841
  (
    n879,
    n839,
    n807,
    n464,
    n778
  );


  and
  g842
  (
    n860,
    n814,
    n775,
    n840,
    n466
  );


  nand
  g843
  (
    n873,
    n817,
    n806,
    n810,
    n820
  );


  nand
  g844
  (
    n895,
    n741,
    n776,
    n809,
    n841
  );


  or
  g845
  (
    n889,
    n679,
    n777,
    n845,
    n811
  );


  nand
  g846
  (
    n876,
    n819,
    n842,
    n806,
    n815
  );


  nand
  g847
  (
    n882,
    n817,
    n463,
    n780,
    n845
  );


  nand
  g848
  (
    n856,
    n463,
    n466,
    n812,
    n678
  );


  nand
  g849
  (
    n891,
    n841,
    n807,
    n635,
    n738
  );


  nor
  g850
  (
    n864,
    n739,
    n814,
    n782,
    n465
  );


  xnor
  g851
  (
    n875,
    n464,
    n812,
    n806,
    n808
  );


  nand
  g852
  (
    n851,
    n679,
    n837,
    n678,
    n465
  );


  nand
  g853
  (
    n888,
    n839,
    n737,
    n271,
    n818
  );


  xor
  g854
  (
    n868,
    n462,
    n462,
    n463,
    n808
  );


  xor
  g855
  (
    n869,
    n635,
    n819,
    n774,
    n845
  );


  xor
  g856
  (
    n858,
    n679,
    n817,
    n810
  );


  xor
  g857
  (
    n862,
    n808,
    n834,
    n807
  );


  nor
  g858
  (
    n884,
    n843,
    n819,
    n837,
    n736
  );


  and
  g859
  (
    n880,
    n843,
    n749,
    n679,
    n462
  );


  and
  g860
  (
    n878,
    n834,
    n843,
    n747,
    n809
  );


  nand
  g861
  (
    n892,
    n836,
    n815,
    n809,
    n818
  );


  nand
  g862
  (
    n854,
    n835,
    n840,
    n836
  );


  buf
  g863
  (
    n896,
    n850
  );


  buf
  g864
  (
    n897,
    n466
  );


  not
  g865
  (
    n898,
    n851
  );


  or
  g866
  (
    n899,
    n852,
    n849,
    n466
  );


  or
  g867
  (
    n909,
    n898,
    n858,
    n17,
    n896
  );


  nand
  g868
  (
    n906,
    n863,
    n18,
    n15,
    n897
  );


  and
  g869
  (
    n900,
    n18,
    n866,
    n16
  );


  nor
  g870
  (
    n903,
    n861,
    n898,
    n896
  );


  nand
  g871
  (
    n902,
    n18,
    n897,
    n860,
    n864
  );


  and
  g872
  (
    n910,
    n16,
    n898,
    n272,
    n865
  );


  and
  g873
  (
    n901,
    n857,
    n15,
    n272,
    n17
  );


  xor
  g874
  (
    n907,
    n854,
    n855,
    n273,
    n896
  );


  and
  g875
  (
    n905,
    n866,
    n863,
    n853,
    n897
  );


  and
  g876
  (
    n911,
    n865,
    n15,
    n862,
    n17
  );


  xnor
  g877
  (
    n904,
    n859,
    n15,
    n897,
    n864
  );


  nand
  g878
  (
    n908,
    n896,
    n17,
    n856,
    n16
  );


  not
  g879
  (
    n912,
    n907
  );


  xnor
  g880
  (
    n915,
    n87,
    n88
  );


  xnor
  g881
  (
    n914,
    n909,
    n88
  );


  nor
  g882
  (
    n913,
    n910,
    n908,
    n87
  );


  buf
  g883
  (
    n916,
    n912
  );


  buf
  g884
  (
    KeyWire_0_51,
    n913
  );


  nand
  g885
  (
    n918,
    n753,
    n916,
    n470
  );


  and
  g886
  (
    n919,
    n917,
    n917,
    n467,
    n468
  );


  and
  g887
  (
    n923,
    n469,
    n916,
    n752,
    n470
  );


  nand
  g888
  (
    n920,
    n469,
    n467,
    n468
  );


  nand
  g889
  (
    n921,
    n469,
    n916,
    n468
  );


  xnor
  g890
  (
    n922,
    n469,
    n467,
    n470,
    n751
  );


  or
  g891
  (
    n927,
    n636,
    n636,
    n638,
    n921
  );


  nand
  g892
  (
    n924,
    n637,
    n637,
    n638,
    n636
  );


  xor
  g893
  (
    n925,
    n636,
    n637,
    n920
  );


  nor
  g894
  (
    n926,
    n638,
    n919,
    n922,
    n635
  );


  xor
  g895
  (
    n928,
    n927,
    n470,
    n680,
    n471
  );


  or
  g896
  (
    KeyWire_0_26,
    n758,
    n759,
    n757,
    n928
  );


  nor
  g897
  (
    n929,
    n928,
    n756,
    n754,
    n755
  );


  nor
  g898
  (
    n931,
    n929,
    n680
  );


  nor
  g899
  (
    n933,
    n762,
    n471,
    n931
  );


  nand
  g900
  (
    n935,
    n931,
    n761,
    n471,
    n760
  );


  and
  g901
  (
    n932,
    n765,
    n472,
    n931,
    n764
  );


  xnor
  g902
  (
    n934,
    n930,
    n471,
    n763,
    n472
  );


  xor
  g903
  (
    n937,
    n473,
    n472,
    n933
  );


  nand
  g904
  (
    n936,
    n934,
    n473
  );


  nand
  g905
  (
    n938,
    n937,
    n820
  );


  buf
  g906
  (
    n939,
    n938
  );


  nand
  g907
  (
    n940,
    n802,
    n938,
    n935
  );


  xnor
  g908
  (
    n943,
    n940,
    n823,
    n824,
    n681
  );


  nand
  g909
  (
    n946,
    n823,
    n823,
    n939,
    n681
  );


  nand
  g910
  (
    n942,
    n823,
    n824,
    n940
  );


  or
  g911
  (
    n944,
    n940,
    n824,
    n766,
    n821
  );


  or
  g912
  (
    n948,
    n939,
    n822,
    n821,
    n681
  );


  xnor
  g913
  (
    n945,
    n939,
    n767,
    n821,
    n940
  );


  nand
  g914
  (
    n947,
    n681,
    n822,
    n939,
    n825
  );


  and
  g915
  (
    KeyWire_0_37,
    n821,
    n820,
    n822
  );


  nor
  g916
  (
    n951,
    n768,
    n682,
    n941
  );


  xor
  g917
  (
    KeyWire_0_0,
    n941,
    n682
  );


  xnor
  g918
  (
    n950,
    n638,
    n941,
    n769,
    n682
  );


  xor
  g919
  (
    n963,
    n847,
    n941,
    n946,
    n951
  );


  xor
  g920
  (
    n962,
    n943,
    n942,
    n845,
    n847
  );


  xnor
  g921
  (
    n956,
    n847,
    n943,
    n945,
    n950
  );


  nand
  g922
  (
    n954,
    n950,
    n944,
    n949
  );


  and
  g923
  (
    n955,
    n944,
    n946,
    n951
  );


  xnor
  g924
  (
    n958,
    n846,
    n847,
    n945,
    n943
  );


  xor
  g925
  (
    n961,
    n947,
    n949,
    n846
  );


  and
  g926
  (
    n960,
    n846,
    n947,
    n950,
    n944
  );


  and
  g927
  (
    n959,
    n942,
    n942,
    n947,
    n951
  );


  and
  g928
  (
    n953,
    n950,
    n942,
    n949,
    n945
  );


  xnor
  g929
  (
    n952,
    n945,
    n846,
    n848,
    n943
  );


  or
  g930
  (
    n957,
    n848,
    n946,
    n951,
    n947
  );


  nor
  g931
  (
    n967,
    n886,
    n952,
    n957,
    n880
  );


  nor
  g932
  (
    n990,
    n885,
    n869,
    n879,
    n877
  );


  nand
  g933
  (
    n973,
    n874,
    n962,
    n867,
    n881
  );


  nand
  g934
  (
    n975,
    n961,
    n890,
    n959,
    n878
  );


  and
  g935
  (
    n970,
    n891,
    n880,
    n884,
    n883
  );


  and
  g936
  (
    n988,
    n954,
    n884,
    n893,
    n876
  );


  xor
  g937
  (
    n980,
    n963,
    n961,
    n885,
    n887
  );


  or
  g938
  (
    n984,
    n877,
    n877,
    n959,
    n953
  );


  nor
  g939
  (
    n995,
    n875,
    n956,
    n886,
    n871
  );


  or
  g940
  (
    n966,
    n872,
    n888,
    n955,
    n962
  );


  or
  g941
  (
    KeyWire_0_59,
    n959,
    n882,
    n890,
    n868
  );


  or
  g942
  (
    n971,
    n874,
    n880,
    n873,
    n960
  );


  xor
  g943
  (
    n974,
    n873,
    n873,
    n883,
    n878
  );


  nor
  g944
  (
    n991,
    n891,
    n868,
    n890,
    n881
  );


  or
  g945
  (
    n993,
    n961,
    n891,
    n876,
    n892
  );


  nand
  g946
  (
    n989,
    n960,
    n958,
    n883,
    n891
  );


  nand
  g947
  (
    n964,
    n885,
    n889,
    n872,
    n963
  );


  xnor
  g948
  (
    n979,
    n893,
    n890,
    n879,
    n960
  );


  xnor
  g949
  (
    n981,
    n892,
    n875,
    n886,
    n882
  );


  xnor
  g950
  (
    n987,
    n892,
    n884,
    n954,
    n878
  );


  xor
  g951
  (
    n968,
    n874,
    n874,
    n893,
    n883
  );


  and
  g952
  (
    n986,
    n887,
    n962,
    n888,
    n882
  );


  xor
  g953
  (
    n978,
    n956,
    n961,
    n875,
    n892
  );


  or
  g954
  (
    n977,
    n875,
    n886,
    n881,
    n869
  );


  and
  g955
  (
    KeyWire_0_40,
    n873,
    n870,
    n889,
    n879
  );


  nor
  g956
  (
    n982,
    n878,
    n889,
    n962,
    n876
  );


  xnor
  g957
  (
    n992,
    n881,
    n884,
    n888,
    n879
  );


  nor
  g958
  (
    n965,
    n882,
    n952,
    n889,
    n877
  );


  xnor
  g959
  (
    n994,
    n887,
    n885,
    n959,
    n953
  );


  or
  g960
  (
    n983,
    n893,
    n871,
    n955,
    n887
  );


  xor
  g961
  (
    n972,
    n957,
    n888,
    n867,
    n880
  );


  nand
  g962
  (
    n976,
    n870,
    n876,
    n958,
    n960
  );


  or
  g963
  (
    n1007,
    n967,
    n993,
    n965,
    n915
  );


  and
  g964
  (
    n1010,
    n994,
    n895,
    n980,
    n894
  );


  nand
  g965
  (
    n1003,
    n894,
    n894,
    n971,
    n895
  );


  and
  g966
  (
    n1002,
    n826,
    n826,
    n848,
    n825
  );


  nor
  g967
  (
    n1009,
    n894,
    n826,
    n273,
    n991
  );


  nand
  g968
  (
    n1011,
    n915,
    n992,
    n948,
    n989
  );


  or
  g969
  (
    n998,
    n899,
    n914,
    n979,
    n981
  );


  nor
  g970
  (
    n1013,
    n964,
    n975,
    n963,
    n970
  );


  nand
  g971
  (
    n1012,
    n972,
    n848,
    n273,
    n915
  );


  xor
  g972
  (
    n1001,
    n968,
    n899,
    n917,
    n948
  );


  and
  g973
  (
    n1008,
    n990,
    n895,
    n915,
    n986
  );


  nor
  g974
  (
    n1004,
    n969,
    n988,
    n825
  );


  or
  g975
  (
    n1006,
    n987,
    n948,
    n802,
    n899
  );


  nand
  g976
  (
    n999,
    n995,
    n976,
    n826,
    n917
  );


  and
  g977
  (
    n997,
    n895,
    n963,
    n973,
    n948
  );


  xor
  g978
  (
    n1000,
    n899,
    n273,
    n911,
    n974
  );


  nor
  g979
  (
    n996,
    n984,
    n923,
    n983,
    n977
  );


  and
  g980
  (
    n1005,
    n985,
    n966,
    n978,
    n982
  );


  or
  g981
  (
    n1017,
    n1006,
    n23,
    n1003,
    n32
  );


  or
  g982
  (
    n1015,
    n28,
    n1005,
    n32,
    n1013
  );


  or
  g983
  (
    n1024,
    n1004,
    n30,
    n25,
    n19
  );


  and
  g984
  (
    n1032,
    n20,
    n29,
    n22,
    n21
  );


  xnor
  g985
  (
    n1031,
    n998,
    n26,
    n997,
    n23
  );


  nand
  g986
  (
    n1022,
    n1008,
    n22,
    n20,
    n23
  );


  xor
  g987
  (
    n1025,
    n19,
    n31,
    n1011
  );


  nand
  g988
  (
    n1021,
    n1002,
    n1000,
    n27,
    n29
  );


  and
  g989
  (
    n1016,
    n19,
    n1010,
    n25,
    n27
  );


  nor
  g990
  (
    n1027,
    n24,
    n27,
    n31,
    n28
  );


  or
  g991
  (
    n1026,
    n18,
    n22,
    n996,
    n1013
  );


  nand
  g992
  (
    n1018,
    n1012,
    n32,
    n22,
    n29
  );


  or
  g993
  (
    n1029,
    n26,
    n24,
    n20
  );


  xor
  g994
  (
    n1028,
    n30,
    n28
  );


  nand
  g995
  (
    n1030,
    n25,
    n32,
    n20,
    n30
  );


  nor
  g996
  (
    KeyWire_0_49,
    n1009,
    n21,
    n999
  );


  nand
  g997
  (
    n1023,
    n26,
    n29,
    n19,
    n1007
  );


  and
  g998
  (
    n1019,
    n25,
    n31,
    n24,
    n26
  );


  or
  g999
  (
    KeyWire_0_48,
    n27,
    n1001,
    n23,
    n21
  );


  xnor
  KeyGate_0_0
  (
    n949,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n93,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n628,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n273,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n489,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n474,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n159,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n718,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n505,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n36,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n380,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n188,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n720,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n639,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n323,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n680,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n105,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n777,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n57,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n174,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n117,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n525,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n244,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n534,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n249,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n571,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n930,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n216,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n337,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n250,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n593,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n412,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n127,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n187,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n644,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n168,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n591,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n941,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n122,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n472,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n969,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n725,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n653,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n83,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n217,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n338,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n373,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n771,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n1014,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n1020,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n276,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n917,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n855,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n656,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n135,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n238,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n319,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n69,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n566,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n985,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n286,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n538,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n633,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n840,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

