

module Stat_2675_57_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n94,
  n256,
  n636,
  n627,
  n609,
  n626,
  n848,
  n858,
  n1036,
  n1826,
  n1941,
  n1948,
  n1940,
  n1947,
  n1942,
  n1943,
  n1946,
  n1938,
  n1936,
  n1944,
  n2699,
  n2691,
  n2687,
  n2688,
  n2692,
  n2693,
  n2689,
  n2685,
  n2700,
  n2681,
  n2697,
  n2690,
  n2683,
  n2701,
  n2684,
  n2696,
  n2694,
  n2686,
  n2695,
  n2682,
  n2698,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n94;
  output n256;
  output n636;
  output n627;
  output n609;
  output n626;
  output n848;
  output n858;
  output n1036;
  output n1826;
  output n1941;
  output n1948;
  output n1940;
  output n1947;
  output n1942;
  output n1943;
  output n1946;
  output n1938;
  output n1936;
  output n1944;
  output n2699;
  output n2691;
  output n2687;
  output n2688;
  output n2692;
  output n2693;
  output n2689;
  output n2685;
  output n2700;
  output n2681;
  output n2697;
  output n2690;
  output n2683;
  output n2701;
  output n2684;
  output n2696;
  output n2694;
  output n2686;
  output n2695;
  output n2682;
  output n2698;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1937;
  wire n1939;
  wire n1945;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n59,
    n11
  );


  not
  g1
  (
    n90,
    n11
  );


  not
  g2
  (
    n106,
    n7
  );


  buf
  g3
  (
    n112,
    n5
  );


  not
  g4
  (
    n48,
    n16
  );


  not
  g5
  (
    n77,
    n9
  );


  buf
  g6
  (
    n37,
    n20
  );


  buf
  g7
  (
    n52,
    n18
  );


  buf
  g8
  (
    n44,
    n22
  );


  not
  g9
  (
    n69,
    n16
  );


  buf
  g10
  (
    n100,
    n18
  );


  not
  g11
  (
    n41,
    n11
  );


  buf
  g12
  (
    n98,
    n20
  );


  not
  g13
  (
    n72,
    n14
  );


  buf
  g14
  (
    n40,
    n13
  );


  not
  g15
  (
    n118,
    n23
  );


  not
  g16
  (
    n34,
    n15
  );


  buf
  g17
  (
    n57,
    n4
  );


  not
  g18
  (
    n45,
    n3
  );


  buf
  g19
  (
    n61,
    n1
  );


  buf
  g20
  (
    n38,
    n17
  );


  not
  g21
  (
    n39,
    n21
  );


  buf
  g22
  (
    n32,
    n5
  );


  not
  g23
  (
    n46,
    n10
  );


  not
  g24
  (
    n64,
    n15
  );


  not
  g25
  (
    n55,
    n4
  );


  not
  g26
  (
    n49,
    n1
  );


  not
  g27
  (
    n42,
    n14
  );


  buf
  g28
  (
    n89,
    n17
  );


  buf
  g29
  (
    n43,
    n12
  );


  buf
  g30
  (
    n115,
    n15
  );


  not
  g31
  (
    n104,
    n22
  );


  buf
  g32
  (
    n78,
    n19
  );


  buf
  g33
  (
    n58,
    n3
  );


  buf
  g34
  (
    n96,
    n21
  );


  buf
  g35
  (
    n84,
    n21
  );


  not
  g36
  (
    n27,
    n14
  );


  not
  g37
  (
    n107,
    n13
  );


  not
  g38
  (
    n94,
    n9
  );


  not
  g39
  (
    n105,
    n20
  );


  not
  g40
  (
    n74,
    n8
  );


  buf
  g41
  (
    n117,
    n8
  );


  not
  g42
  (
    n75,
    n17
  );


  buf
  g43
  (
    n109,
    n16
  );


  buf
  g44
  (
    n65,
    n6
  );


  not
  g45
  (
    n36,
    n21
  );


  not
  g46
  (
    n73,
    n5
  );


  buf
  g47
  (
    n71,
    n23
  );


  buf
  g48
  (
    n63,
    n19
  );


  not
  g49
  (
    n54,
    n19
  );


  not
  g50
  (
    n29,
    n10
  );


  not
  g51
  (
    n67,
    n18
  );


  buf
  g52
  (
    n70,
    n10
  );


  not
  g53
  (
    n92,
    n6
  );


  buf
  g54
  (
    n111,
    n13
  );


  not
  g55
  (
    KeyWire_0_51,
    n6
  );


  buf
  g56
  (
    n51,
    n7
  );


  not
  g57
  (
    n88,
    n4
  );


  buf
  g58
  (
    n62,
    n20
  );


  buf
  g59
  (
    n116,
    n18
  );


  buf
  g60
  (
    n60,
    n8
  );


  not
  g61
  (
    n103,
    n1
  );


  buf
  g62
  (
    n99,
    n22
  );


  not
  g63
  (
    n113,
    n13
  );


  buf
  g64
  (
    n56,
    n10
  );


  buf
  g65
  (
    n93,
    n14
  );


  not
  g66
  (
    n53,
    n2
  );


  buf
  g67
  (
    n102,
    n19
  );


  not
  g68
  (
    n85,
    n8
  );


  buf
  g69
  (
    n76,
    n6
  );


  not
  g70
  (
    n108,
    n9
  );


  buf
  g71
  (
    n91,
    n2
  );


  buf
  g72
  (
    n68,
    n7
  );


  not
  g73
  (
    n82,
    n3
  );


  buf
  g74
  (
    n80,
    n23
  );


  not
  g75
  (
    n114,
    n17
  );


  buf
  g76
  (
    n95,
    n7
  );


  not
  g77
  (
    n87,
    n11
  );


  not
  g78
  (
    n50,
    n12
  );


  not
  g79
  (
    n83,
    n2
  );


  not
  g80
  (
    n86,
    n15
  );


  buf
  g81
  (
    n28,
    n22
  );


  not
  g82
  (
    n30,
    n1
  );


  not
  g83
  (
    n81,
    n12
  );


  not
  g84
  (
    n97,
    n23
  );


  not
  g85
  (
    n66,
    n3
  );


  buf
  g86
  (
    n79,
    n9
  );


  not
  g87
  (
    n31,
    n4
  );


  not
  g88
  (
    n47,
    n16
  );


  not
  g89
  (
    n35,
    n2
  );


  not
  g90
  (
    n110,
    n5
  );


  buf
  g91
  (
    KeyWire_0_18,
    n12
  );


  buf
  g92
  (
    n163,
    n28
  );


  not
  g93
  (
    n128,
    n51
  );


  not
  g94
  (
    n119,
    n46
  );


  buf
  g95
  (
    n120,
    n51
  );


  buf
  g96
  (
    n158,
    n39
  );


  buf
  g97
  (
    n135,
    n33
  );


  not
  g98
  (
    n148,
    n48
  );


  buf
  g99
  (
    n134,
    n52
  );


  not
  g100
  (
    n138,
    n40
  );


  buf
  g101
  (
    n136,
    n36
  );


  not
  g102
  (
    n131,
    n43
  );


  buf
  g103
  (
    n124,
    n32
  );


  not
  g104
  (
    n167,
    n42
  );


  buf
  g105
  (
    n145,
    n45
  );


  buf
  g106
  (
    n146,
    n31
  );


  buf
  g107
  (
    n144,
    n27
  );


  buf
  g108
  (
    n154,
    n50
  );


  not
  g109
  (
    n137,
    n30
  );


  buf
  g110
  (
    n123,
    n33
  );


  not
  g111
  (
    n153,
    n36
  );


  buf
  g112
  (
    n156,
    n46
  );


  not
  g113
  (
    n141,
    n42
  );


  buf
  g114
  (
    n142,
    n38
  );


  buf
  g115
  (
    n161,
    n49
  );


  buf
  g116
  (
    n132,
    n38
  );


  buf
  g117
  (
    n133,
    n43
  );


  not
  g118
  (
    n164,
    n32
  );


  not
  g119
  (
    n121,
    n31
  );


  not
  g120
  (
    n129,
    n40
  );


  not
  g121
  (
    n147,
    n44
  );


  buf
  g122
  (
    n151,
    n51
  );


  buf
  g123
  (
    n165,
    n32
  );


  not
  g124
  (
    n166,
    n34
  );


  buf
  g125
  (
    n126,
    n28
  );


  xor
  g126
  (
    n152,
    n35,
    n39,
    n41,
    n48
  );


  or
  g127
  (
    n157,
    n43,
    n46,
    n37
  );


  or
  g128
  (
    n139,
    n33,
    n36,
    n50
  );


  and
  g129
  (
    n168,
    n40,
    n48,
    n52,
    n41
  );


  xor
  g130
  (
    n125,
    n34,
    n48,
    n44,
    n42
  );


  nand
  g131
  (
    n150,
    n37,
    n29,
    n28
  );


  nor
  g132
  (
    n127,
    n52,
    n46,
    n47,
    n31
  );


  and
  g133
  (
    n160,
    n40,
    n33,
    n27,
    n39
  );


  or
  g134
  (
    n140,
    n47,
    n28,
    n41,
    n30
  );


  or
  g135
  (
    n155,
    n49,
    n30,
    n34,
    n39
  );


  nand
  g136
  (
    n162,
    n42,
    n49,
    n35,
    n44
  );


  nand
  g137
  (
    n122,
    n52,
    n50,
    n30,
    n43
  );


  nor
  g138
  (
    KeyWire_0_49,
    n36,
    n47,
    n41,
    n44
  );


  nor
  g139
  (
    n159,
    n45,
    n34,
    n35,
    n29
  );


  nor
  g140
  (
    n149,
    n49,
    n38,
    n47,
    n37
  );


  and
  g141
  (
    n130,
    n45,
    n38,
    n51,
    n32
  );


  xor
  g142
  (
    n169,
    n31,
    n45,
    n29,
    n35
  );


  not
  g143
  (
    n270,
    n129
  );


  buf
  g144
  (
    n186,
    n164
  );


  not
  g145
  (
    n263,
    n148
  );


  not
  g146
  (
    n238,
    n161
  );


  buf
  g147
  (
    n252,
    n146
  );


  not
  g148
  (
    n175,
    n149
  );


  not
  g149
  (
    n283,
    n144
  );


  buf
  g150
  (
    n174,
    n159
  );


  not
  g151
  (
    n281,
    n166
  );


  not
  g152
  (
    n272,
    n165
  );


  not
  g153
  (
    n284,
    n164
  );


  not
  g154
  (
    n199,
    n153
  );


  buf
  g155
  (
    n188,
    n152
  );


  not
  g156
  (
    n209,
    n167
  );


  buf
  g157
  (
    n268,
    n123
  );


  buf
  g158
  (
    KeyWire_0_35,
    n131
  );


  buf
  g159
  (
    n227,
    n161
  );


  not
  g160
  (
    n266,
    n140
  );


  not
  g161
  (
    n249,
    n135
  );


  not
  g162
  (
    n286,
    n127
  );


  buf
  g163
  (
    n242,
    n124
  );


  buf
  g164
  (
    n192,
    n162
  );


  buf
  g165
  (
    n196,
    n137
  );


  buf
  g166
  (
    n194,
    n158
  );


  buf
  g167
  (
    n285,
    n126
  );


  buf
  g168
  (
    n229,
    n142
  );


  not
  g169
  (
    n226,
    n162
  );


  not
  g170
  (
    n172,
    n134
  );


  not
  g171
  (
    n289,
    n123
  );


  not
  g172
  (
    n290,
    n145
  );


  buf
  g173
  (
    n248,
    n119
  );


  buf
  g174
  (
    n235,
    n132
  );


  not
  g175
  (
    n234,
    n153
  );


  not
  g176
  (
    n178,
    n163
  );


  buf
  g177
  (
    n221,
    n169
  );


  not
  g178
  (
    n177,
    n134
  );


  buf
  g179
  (
    n222,
    n163
  );


  buf
  g180
  (
    n171,
    n147
  );


  buf
  g181
  (
    n244,
    n138
  );


  not
  g182
  (
    n182,
    n122
  );


  buf
  g183
  (
    n205,
    n155
  );


  buf
  g184
  (
    n273,
    n151
  );


  buf
  g185
  (
    n212,
    n156
  );


  not
  g186
  (
    n190,
    n136
  );


  buf
  g187
  (
    n203,
    n129
  );


  buf
  g188
  (
    n223,
    n137
  );


  buf
  g189
  (
    n202,
    n166
  );


  buf
  g190
  (
    n233,
    n150
  );


  not
  g191
  (
    n237,
    n131
  );


  buf
  g192
  (
    n277,
    n120
  );


  buf
  g193
  (
    n267,
    n163
  );


  buf
  g194
  (
    n220,
    n149
  );


  buf
  g195
  (
    n184,
    n130
  );


  buf
  g196
  (
    n271,
    n152
  );


  buf
  g197
  (
    n213,
    n124
  );


  buf
  g198
  (
    n288,
    n128
  );


  buf
  g199
  (
    n262,
    n165
  );


  buf
  g200
  (
    n258,
    n140
  );


  buf
  g201
  (
    n204,
    n169
  );


  buf
  g202
  (
    n239,
    n150
  );


  buf
  g203
  (
    n280,
    n146
  );


  buf
  g204
  (
    n173,
    n167
  );


  not
  g205
  (
    n232,
    n125
  );


  not
  g206
  (
    n274,
    n163
  );


  buf
  g207
  (
    n219,
    n168
  );


  buf
  g208
  (
    n257,
    n141
  );


  not
  g209
  (
    n198,
    n162
  );


  buf
  g210
  (
    n243,
    n154
  );


  not
  g211
  (
    n247,
    n139
  );


  not
  g212
  (
    n250,
    n133
  );


  not
  g213
  (
    n253,
    n151
  );


  buf
  g214
  (
    n187,
    n130
  );


  buf
  g215
  (
    n245,
    n147
  );


  not
  g216
  (
    n211,
    n122
  );


  buf
  g217
  (
    n197,
    n160
  );


  not
  g218
  (
    n214,
    n164
  );


  not
  g219
  (
    n193,
    n128
  );


  not
  g220
  (
    n225,
    n160
  );


  buf
  g221
  (
    n228,
    n136
  );


  buf
  g222
  (
    n279,
    n165
  );


  buf
  g223
  (
    n287,
    n164
  );


  not
  g224
  (
    n278,
    n167
  );


  not
  g225
  (
    n207,
    n127
  );


  not
  g226
  (
    n236,
    n121
  );


  buf
  g227
  (
    n251,
    n148
  );


  buf
  g228
  (
    n179,
    n143
  );


  not
  g229
  (
    n206,
    n158
  );


  buf
  g230
  (
    n218,
    n133
  );


  buf
  g231
  (
    n215,
    n161
  );


  not
  g232
  (
    n208,
    n155
  );


  not
  g233
  (
    n231,
    n162
  );


  not
  g234
  (
    n246,
    n157
  );


  buf
  g235
  (
    n180,
    n168
  );


  not
  g236
  (
    n183,
    n126
  );


  buf
  g237
  (
    KeyWire_0_2,
    n167
  );


  not
  g238
  (
    n269,
    n156
  );


  buf
  g239
  (
    n189,
    n168
  );


  buf
  g240
  (
    n224,
    n161
  );


  not
  g241
  (
    n255,
    n168
  );


  buf
  g242
  (
    n210,
    n160
  );


  not
  g243
  (
    n240,
    n138
  );


  not
  g244
  (
    n259,
    n142
  );


  buf
  g245
  (
    n241,
    n120
  );


  buf
  g246
  (
    n230,
    n141
  );


  not
  g247
  (
    n201,
    n159
  );


  buf
  g248
  (
    n191,
    n154
  );


  not
  g249
  (
    n260,
    n166
  );


  buf
  g250
  (
    n265,
    n144
  );


  buf
  g251
  (
    n264,
    n169
  );


  not
  g252
  (
    n185,
    n125
  );


  buf
  g253
  (
    n200,
    n166
  );


  buf
  g254
  (
    n254,
    n169
  );


  buf
  g255
  (
    n216,
    n121
  );


  buf
  g256
  (
    n181,
    n119
  );


  not
  g257
  (
    n275,
    n132
  );


  not
  g258
  (
    n276,
    n157
  );


  buf
  g259
  (
    n217,
    n145
  );


  buf
  g260
  (
    n282,
    n165
  );


  buf
  g261
  (
    n256,
    n143
  );


  buf
  g262
  (
    n176,
    n139
  );


  not
  g263
  (
    n261,
    n135
  );


  buf
  g264
  (
    n351,
    n170
  );


  buf
  g265
  (
    n328,
    n179
  );


  buf
  g266
  (
    n379,
    n183
  );


  not
  g267
  (
    n333,
    n184
  );


  buf
  g268
  (
    n388,
    n192
  );


  not
  g269
  (
    n365,
    n173
  );


  not
  g270
  (
    n394,
    n183
  );


  not
  g271
  (
    n310,
    n173
  );


  buf
  g272
  (
    n385,
    n188
  );


  buf
  g273
  (
    n295,
    n184
  );


  not
  g274
  (
    n338,
    n182
  );


  not
  g275
  (
    n312,
    n195
  );


  buf
  g276
  (
    n350,
    n179
  );


  not
  g277
  (
    n393,
    n174
  );


  buf
  g278
  (
    n324,
    n171
  );


  not
  g279
  (
    n369,
    n53
  );


  not
  g280
  (
    n326,
    n188
  );


  buf
  g281
  (
    n358,
    n191
  );


  buf
  g282
  (
    n313,
    n172
  );


  not
  g283
  (
    n361,
    n180
  );


  buf
  g284
  (
    n378,
    n190
  );


  buf
  g285
  (
    n390,
    n180
  );


  not
  g286
  (
    n356,
    n194
  );


  not
  g287
  (
    KeyWire_0_27,
    n174
  );


  not
  g288
  (
    n331,
    n171
  );


  buf
  g289
  (
    n367,
    n186
  );


  buf
  g290
  (
    n294,
    n192
  );


  buf
  g291
  (
    n364,
    n185
  );


  not
  g292
  (
    n337,
    n195
  );


  buf
  g293
  (
    n382,
    n188
  );


  buf
  g294
  (
    n380,
    n171
  );


  buf
  g295
  (
    n321,
    n174
  );


  buf
  g296
  (
    n302,
    n191
  );


  buf
  g297
  (
    n372,
    n174
  );


  buf
  g298
  (
    n305,
    n190
  );


  buf
  g299
  (
    n348,
    n195
  );


  buf
  g300
  (
    n343,
    n186
  );


  not
  g301
  (
    n387,
    n190
  );


  not
  g302
  (
    n339,
    n185
  );


  buf
  g303
  (
    n301,
    n170
  );


  buf
  g304
  (
    n357,
    n181
  );


  buf
  g305
  (
    KeyWire_0_4,
    n189
  );


  not
  g306
  (
    n325,
    n179
  );


  not
  g307
  (
    n330,
    n177
  );


  buf
  g308
  (
    n314,
    n177
  );


  buf
  g309
  (
    n291,
    n187
  );


  not
  g310
  (
    n342,
    n175
  );


  buf
  g311
  (
    n355,
    n193
  );


  not
  g312
  (
    n340,
    n192
  );


  not
  g313
  (
    n299,
    n173
  );


  buf
  g314
  (
    n383,
    n177
  );


  buf
  g315
  (
    n368,
    n189
  );


  buf
  g316
  (
    n353,
    n189
  );


  buf
  g317
  (
    n376,
    n187
  );


  not
  g318
  (
    n381,
    n175
  );


  buf
  g319
  (
    n360,
    n194
  );


  not
  g320
  (
    n347,
    n190
  );


  not
  g321
  (
    n304,
    n182
  );


  not
  g322
  (
    n318,
    n186
  );


  not
  g323
  (
    n322,
    n171
  );


  buf
  g324
  (
    n384,
    n195
  );


  not
  g325
  (
    n344,
    n178
  );


  buf
  g326
  (
    n308,
    n176
  );


  not
  g327
  (
    n377,
    n178
  );


  buf
  g328
  (
    n303,
    n181
  );


  buf
  g329
  (
    n297,
    n180
  );


  not
  g330
  (
    n336,
    n175
  );


  not
  g331
  (
    n307,
    n194
  );


  buf
  g332
  (
    n300,
    n192
  );


  not
  g333
  (
    n373,
    n176
  );


  buf
  g334
  (
    n371,
    n193
  );


  not
  g335
  (
    n309,
    n183
  );


  not
  g336
  (
    n292,
    n170
  );


  buf
  g337
  (
    n335,
    n194
  );


  buf
  g338
  (
    n354,
    n182
  );


  not
  g339
  (
    n323,
    n184
  );


  not
  g340
  (
    n311,
    n193
  );


  buf
  g341
  (
    n349,
    n191
  );


  not
  g342
  (
    n362,
    n185
  );


  buf
  g343
  (
    n374,
    n188
  );


  buf
  g344
  (
    n375,
    n176
  );


  not
  g345
  (
    n392,
    n183
  );


  not
  g346
  (
    n316,
    n186
  );


  buf
  g347
  (
    n391,
    n179
  );


  buf
  g348
  (
    n341,
    n180
  );


  not
  g349
  (
    n327,
    n172
  );


  buf
  g350
  (
    n386,
    n196
  );


  not
  g351
  (
    n319,
    n172
  );


  buf
  g352
  (
    n334,
    n187
  );


  not
  g353
  (
    n352,
    n178
  );


  not
  g354
  (
    n320,
    n176
  );


  buf
  g355
  (
    n359,
    n182
  );


  not
  g356
  (
    n315,
    n175
  );


  buf
  g357
  (
    n363,
    n191
  );


  buf
  g358
  (
    n366,
    n181
  );


  not
  g359
  (
    n389,
    n185
  );


  not
  g360
  (
    n332,
    n173
  );


  not
  g361
  (
    n329,
    n172
  );


  buf
  g362
  (
    n306,
    n193
  );


  buf
  g363
  (
    n298,
    n177
  );


  not
  g364
  (
    n345,
    n181
  );


  not
  g365
  (
    n293,
    n184
  );


  buf
  g366
  (
    n296,
    n178
  );


  or
  g367
  (
    n370,
    n189,
    n187
  );


  not
  g368
  (
    n485,
    n260
  );


  not
  g369
  (
    n506,
    n268
  );


  xnor
  g370
  (
    n450,
    n275,
    n227,
    n208,
    n252
  );


  nand
  g371
  (
    n512,
    n275,
    n246,
    n208,
    n207
  );


  xnor
  g372
  (
    n473,
    n235,
    n254,
    n273,
    n274
  );


  xor
  g373
  (
    n472,
    n196,
    n276,
    n263,
    n267
  );


  or
  g374
  (
    KeyWire_0_23,
    n263,
    n257,
    n254,
    n358
  );


  and
  g375
  (
    n492,
    n237,
    n287,
    n256,
    n244
  );


  nor
  g376
  (
    n484,
    n269,
    n389,
    n268,
    n365
  );


  and
  g377
  (
    n493,
    n283,
    n274,
    n272,
    n261
  );


  and
  g378
  (
    n432,
    n353,
    n199,
    n261,
    n268
  );


  or
  g379
  (
    n517,
    n271,
    n258,
    n281,
    n238
  );


  xor
  g380
  (
    n519,
    n361,
    n233,
    n275,
    n260
  );


  nand
  g381
  (
    n428,
    n236,
    n218,
    n221,
    n223
  );


  nor
  g382
  (
    n470,
    n216,
    n274,
    n252,
    n198
  );


  nor
  g383
  (
    n509,
    n281,
    n228,
    n241,
    n332
  );


  nor
  g384
  (
    n494,
    n202,
    n242,
    n201,
    n256
  );


  nor
  g385
  (
    n443,
    n255,
    n211,
    n333,
    n374
  );


  xor
  g386
  (
    n399,
    n277,
    n214,
    n251,
    n213
  );


  xor
  g387
  (
    n458,
    n284,
    n232,
    n214,
    n197
  );


  nand
  g388
  (
    n507,
    n217,
    n387,
    n390,
    n330
  );


  nor
  g389
  (
    n395,
    n198,
    n356,
    n222,
    n209
  );


  and
  g390
  (
    n410,
    n352,
    n384,
    n215,
    n197
  );


  xnor
  g391
  (
    n477,
    n196,
    n364,
    n250,
    n256
  );


  nor
  g392
  (
    n421,
    n248,
    n204,
    n224,
    n336
  );


  nor
  g393
  (
    n418,
    n280,
    n334,
    n282,
    n375
  );


  or
  g394
  (
    n463,
    n262,
    n309,
    n236,
    n207
  );


  nand
  g395
  (
    n436,
    n251,
    n340,
    n327,
    n202
  );


  or
  g396
  (
    n430,
    n252,
    n337,
    n247,
    n265
  );


  or
  g397
  (
    n467,
    n314,
    n247,
    n267,
    n239
  );


  and
  g398
  (
    n462,
    n393,
    n273,
    n229,
    n227
  );


  xor
  g399
  (
    n455,
    n253,
    n247,
    n209,
    n371
  );


  xor
  g400
  (
    n454,
    n349,
    n386,
    n205
  );


  and
  g401
  (
    n461,
    n285,
    n229,
    n283,
    n372
  );


  nor
  g402
  (
    n515,
    n213,
    n216,
    n391
  );


  or
  g403
  (
    n491,
    n250,
    n202,
    n339,
    n221
  );


  xnor
  g404
  (
    n502,
    n272,
    n273,
    n231,
    n259
  );


  nand
  g405
  (
    n396,
    n363,
    n392,
    n283,
    n241
  );


  or
  g406
  (
    n434,
    n297,
    n215,
    n278,
    n206
  );


  or
  g407
  (
    n398,
    n273,
    n280,
    n263,
    n272
  );


  nand
  g408
  (
    n488,
    n212,
    n286,
    n264,
    n229
  );


  xor
  g409
  (
    n415,
    n279,
    n300,
    n354,
    n199
  );


  and
  g410
  (
    n404,
    n282,
    n210,
    n204,
    n380
  );


  and
  g411
  (
    n486,
    n272,
    n266,
    n282,
    n382
  );


  nand
  g412
  (
    KeyWire_0_3,
    n338,
    n202,
    n381,
    n270
  );


  nand
  g413
  (
    n407,
    n322,
    n318,
    n224,
    n221
  );


  nor
  g414
  (
    n449,
    n203,
    n335,
    n381,
    n384
  );


  nor
  g415
  (
    n420,
    n351,
    n209,
    n311,
    n261
  );


  and
  g416
  (
    n500,
    n243,
    n305,
    n285,
    n246
  );


  or
  g417
  (
    n401,
    n219,
    n203,
    n223,
    n279
  );


  xnor
  g418
  (
    n427,
    n232,
    n357,
    n203,
    n285
  );


  nand
  g419
  (
    KeyWire_0_12,
    n230,
    n350,
    n270,
    n341
  );


  xor
  g420
  (
    n478,
    n215,
    n230,
    n294,
    n284
  );


  nand
  g421
  (
    n504,
    n386,
    n265,
    n240,
    n263
  );


  nor
  g422
  (
    n417,
    n367,
    n234,
    n271,
    n320
  );


  xnor
  g423
  (
    n416,
    n245,
    n220,
    n312,
    n315
  );


  xnor
  g424
  (
    n496,
    n226,
    n208,
    n246,
    n390
  );


  nand
  g425
  (
    n503,
    n231,
    n258,
    n219,
    n282
  );


  xnor
  g426
  (
    n513,
    n205,
    n299,
    n213,
    n288
  );


  and
  g427
  (
    n413,
    n362,
    n227,
    n242,
    n248
  );


  nor
  g428
  (
    n426,
    n262,
    n237,
    n306,
    n198
  );


  or
  g429
  (
    n440,
    n385,
    n264,
    n287,
    n212
  );


  or
  g430
  (
    n412,
    n211,
    n383,
    n252,
    n319
  );


  xor
  g431
  (
    n431,
    n379,
    n253,
    n301,
    n212
  );


  nor
  g432
  (
    n422,
    n265,
    n207,
    n360,
    n236
  );


  nor
  g433
  (
    n497,
    n228,
    n383,
    n388,
    n284
  );


  or
  g434
  (
    n508,
    n269,
    n271,
    n287,
    n235
  );


  and
  g435
  (
    n442,
    n372,
    n317,
    n281,
    n260
  );


  or
  g436
  (
    n409,
    n387,
    n347,
    n262,
    n259
  );


  and
  g437
  (
    n402,
    n266,
    n243,
    n218,
    n257
  );


  and
  g438
  (
    n481,
    n277,
    n254,
    n214,
    n225
  );


  and
  g439
  (
    n439,
    n215,
    n201,
    n310,
    n242
  );


  and
  g440
  (
    n474,
    n216,
    n255,
    n375,
    n331
  );


  nor
  g441
  (
    n469,
    n250,
    n224,
    n244,
    n368
  );


  or
  g442
  (
    n433,
    n223,
    n246,
    n265,
    n204
  );


  and
  g443
  (
    n483,
    n276,
    n359,
    n236,
    n241
  );


  nor
  g444
  (
    n414,
    n268,
    n380,
    n378,
    n240
  );


  nand
  g445
  (
    n482,
    n208,
    n233,
    n266,
    n248
  );


  and
  g446
  (
    n456,
    n373,
    n239,
    n392,
    n245
  );


  xnor
  g447
  (
    n510,
    n225,
    n229,
    n277,
    n355
  );


  nor
  g448
  (
    n505,
    n222,
    n223,
    n379,
    n217
  );


  and
  g449
  (
    n475,
    n243,
    n235,
    n276,
    n197
  );


  nor
  g450
  (
    n447,
    n303,
    n259,
    n376,
    n247
  );


  and
  g451
  (
    n419,
    n235,
    n205,
    n298,
    n260
  );


  nand
  g452
  (
    n452,
    n230,
    n220,
    n280,
    n237
  );


  nand
  g453
  (
    n457,
    n226,
    n211,
    n258,
    n234
  );


  and
  g454
  (
    n476,
    n206,
    n233,
    n232,
    n283
  );


  xnor
  g455
  (
    n453,
    n271,
    n199,
    n220,
    n324
  );


  or
  g456
  (
    n501,
    n321,
    n308,
    n276,
    n234
  );


  and
  g457
  (
    n444,
    n296,
    n284,
    n201,
    n316
  );


  and
  g458
  (
    n445,
    n220,
    n200,
    n251,
    n249
  );


  xnor
  g459
  (
    n498,
    n245,
    n262,
    n342,
    n217
  );


  or
  g460
  (
    n465,
    n288,
    n293,
    n278,
    n302
  );


  xor
  g461
  (
    n406,
    n219,
    n280,
    n348,
    n231
  );


  and
  g462
  (
    n514,
    n287,
    n389,
    n258,
    n218
  );


  nor
  g463
  (
    n425,
    n250,
    n382,
    n231,
    n206
  );


  or
  g464
  (
    n423,
    n270,
    n345,
    n212,
    n388
  );


  or
  g465
  (
    n490,
    n240,
    n228,
    n261,
    n207
  );


  or
  g466
  (
    n429,
    n374,
    n269,
    n274,
    n277
  );


  xnor
  g467
  (
    n511,
    n343,
    n371,
    n377,
    n264
  );


  nor
  g468
  (
    n438,
    n233,
    n292,
    n224,
    n249
  );


  xnor
  g469
  (
    n408,
    n203,
    n328,
    n217,
    n267
  );


  nor
  g470
  (
    n516,
    n245,
    n251,
    n213,
    n377
  );


  and
  g471
  (
    n499,
    n295,
    n237,
    n291,
    n286
  );


  or
  g472
  (
    n411,
    n198,
    n256,
    n228,
    n248
  );


  nand
  g473
  (
    n448,
    n254,
    n249,
    n238
  );


  xor
  g474
  (
    n400,
    n323,
    n225,
    n216,
    n255
  );


  xor
  g475
  (
    n451,
    n239,
    n244,
    n210,
    n376
  );


  or
  g476
  (
    n424,
    n196,
    n373,
    n197,
    n218
  );


  and
  g477
  (
    n441,
    n313,
    n200,
    n286,
    n304
  );


  xor
  g478
  (
    KeyWire_0_38,
    n226,
    n199,
    n279,
    n259
  );


  or
  g479
  (
    n489,
    n242,
    n253,
    n204,
    n244
  );


  or
  g480
  (
    n479,
    n329,
    n232,
    n378,
    n255
  );


  nand
  g481
  (
    n466,
    n201,
    n278,
    n266,
    n209
  );


  nand
  g482
  (
    n397,
    n281,
    n222,
    n238,
    n239
  );


  and
  g483
  (
    n518,
    n278,
    n286,
    n264,
    n225
  );


  and
  g484
  (
    n437,
    n307,
    n234,
    n214,
    n210
  );


  and
  g485
  (
    n460,
    n221,
    n285,
    n219,
    n369
  );


  nand
  g486
  (
    n487,
    n226,
    n200,
    n249,
    n325
  );


  nor
  g487
  (
    n464,
    n200,
    n326,
    n227,
    n346
  );


  nor
  g488
  (
    n446,
    n240,
    n241,
    n230,
    n206
  );


  nor
  g489
  (
    n495,
    n370,
    n270,
    n210,
    n366
  );


  and
  g490
  (
    n435,
    n275,
    n257,
    n279
  );


  xor
  g491
  (
    n471,
    n269,
    n243,
    n385,
    n267
  );


  xnor
  g492
  (
    n403,
    n253,
    n344,
    n211,
    n222
  );


  nand
  g493
  (
    n543,
    n400,
    n63,
    n70,
    n73
  );


  nor
  g494
  (
    KeyWire_0_61,
    n76,
    n53,
    n74,
    n62
  );


  nand
  g495
  (
    n526,
    n66,
    n62,
    n73,
    n64
  );


  nand
  g496
  (
    n535,
    n66,
    n56,
    n57,
    n74
  );


  xnor
  g497
  (
    n554,
    n77,
    n401,
    n62,
    n82
  );


  xor
  g498
  (
    n530,
    n56,
    n429,
    n410,
    n79
  );


  nor
  g499
  (
    n545,
    n79,
    n76,
    n80,
    n63
  );


  xor
  g500
  (
    n521,
    n74,
    n395,
    n73,
    n57
  );


  xnor
  g501
  (
    n533,
    n402,
    n409,
    n67,
    n421
  );


  and
  g502
  (
    n544,
    n61,
    n412,
    n55
  );


  or
  g503
  (
    n546,
    n75,
    n66,
    n59,
    n78
  );


  and
  g504
  (
    n541,
    n62,
    n64,
    n56,
    n432
  );


  nand
  g505
  (
    KeyWire_0_8,
    n65,
    n59,
    n399,
    n78
  );


  nor
  g506
  (
    n548,
    n72,
    n80,
    n63,
    n64
  );


  nand
  g507
  (
    n520,
    n425,
    n80,
    n58,
    n71
  );


  xor
  g508
  (
    n550,
    n427,
    n61,
    n428
  );


  xnor
  g509
  (
    n557,
    n423,
    n406,
    n79,
    n81
  );


  xnor
  g510
  (
    n528,
    n418,
    n54,
    n70,
    n69
  );


  and
  g511
  (
    n552,
    n398,
    n413,
    n408,
    n78
  );


  nor
  g512
  (
    n525,
    n426,
    n65,
    n67,
    n288
  );


  and
  g513
  (
    n536,
    n68,
    n422,
    n61,
    n424
  );


  nor
  g514
  (
    n529,
    n58,
    n403,
    n56,
    n76
  );


  or
  g515
  (
    n558,
    n396,
    n71,
    n55,
    n60
  );


  and
  g516
  (
    n542,
    n60,
    n72,
    n71
  );


  xnor
  g517
  (
    n549,
    n54,
    n414,
    n70,
    n76
  );


  or
  g518
  (
    n539,
    n430,
    n419,
    n53,
    n68
  );


  xnor
  g519
  (
    n532,
    n53,
    n67,
    n75,
    n77
  );


  xor
  g520
  (
    n527,
    n57,
    n415,
    n433,
    n71
  );


  nand
  g521
  (
    n540,
    n411,
    n80,
    n68,
    n54
  );


  or
  g522
  (
    n547,
    n59,
    n64,
    n69,
    n78
  );


  or
  g523
  (
    n553,
    n405,
    n72,
    n431,
    n79
  );


  nor
  g524
  (
    n524,
    n397,
    n58,
    n60,
    n65
  );


  or
  g525
  (
    n534,
    n67,
    n75,
    n57,
    n58
  );


  nand
  g526
  (
    n555,
    n55,
    n60,
    n416,
    n81
  );


  and
  g527
  (
    n531,
    n59,
    n69,
    n65,
    n77
  );


  and
  g528
  (
    n522,
    n63,
    n407,
    n75,
    n420
  );


  or
  g529
  (
    n551,
    n70,
    n66,
    n417,
    n69
  );


  nand
  g530
  (
    n523,
    n81,
    n54,
    n73,
    n404
  );


  xor
  g531
  (
    n556,
    n74,
    n68,
    n81,
    n77
  );


  buf
  g532
  (
    KeyWire_0_33,
    n520
  );


  not
  g533
  (
    n561,
    n521
  );


  not
  g534
  (
    n563,
    n522
  );


  buf
  g535
  (
    n565,
    n520
  );


  buf
  g536
  (
    n564,
    n520
  );


  not
  g537
  (
    n566,
    n521
  );


  not
  g538
  (
    n569,
    n520
  );


  buf
  g539
  (
    n567,
    n521
  );


  buf
  g540
  (
    n562,
    n522
  );


  not
  g541
  (
    n559,
    n522
  );


  not
  g542
  (
    n568,
    n521
  );


  buf
  g543
  (
    n599,
    n559
  );


  buf
  g544
  (
    n573,
    n564
  );


  buf
  g545
  (
    n580,
    n561
  );


  not
  g546
  (
    n585,
    n562
  );


  not
  g547
  (
    n570,
    n560
  );


  buf
  g548
  (
    n594,
    n563
  );


  buf
  g549
  (
    n586,
    n565
  );


  not
  g550
  (
    n595,
    n563
  );


  not
  g551
  (
    n574,
    n566
  );


  not
  g552
  (
    n571,
    n562
  );


  not
  g553
  (
    n587,
    n566
  );


  not
  g554
  (
    n593,
    n559
  );


  buf
  g555
  (
    n596,
    n564
  );


  buf
  g556
  (
    n598,
    n563
  );


  buf
  g557
  (
    n579,
    n561
  );


  buf
  g558
  (
    n578,
    n565
  );


  buf
  g559
  (
    n572,
    n565
  );


  buf
  g560
  (
    n575,
    n559
  );


  not
  g561
  (
    KeyWire_0_21,
    n563
  );


  not
  g562
  (
    n581,
    n564
  );


  not
  g563
  (
    n584,
    n561
  );


  buf
  g564
  (
    n576,
    n560
  );


  not
  g565
  (
    n590,
    n561
  );


  buf
  g566
  (
    n597,
    n562
  );


  not
  g567
  (
    n577,
    n565
  );


  buf
  g568
  (
    n591,
    n562
  );


  not
  g569
  (
    n592,
    n559
  );


  buf
  g570
  (
    n588,
    n564
  );


  buf
  g571
  (
    n583,
    n560
  );


  not
  g572
  (
    n582,
    n560
  );


  xnor
  g573
  (
    n633,
    n571,
    n453,
    n483,
    n478
  );


  xnor
  g574
  (
    n606,
    n500,
    n497,
    n570,
    n575
  );


  nor
  g575
  (
    n635,
    n507,
    n454,
    n578,
    n442
  );


  xnor
  g576
  (
    n604,
    n577,
    n447,
    n504,
    n570
  );


  xor
  g577
  (
    n631,
    n483,
    n439,
    n490,
    n576
  );


  or
  g578
  (
    n612,
    n480,
    n572,
    n574
  );


  or
  g579
  (
    n618,
    n495,
    n472,
    n575,
    n573
  );


  xnor
  g580
  (
    n611,
    n498,
    n489,
    n472,
    n492
  );


  or
  g581
  (
    n600,
    n500,
    n479,
    n570,
    n576
  );


  xor
  g582
  (
    n624,
    n465,
    n478,
    n574,
    n576
  );


  xnor
  g583
  (
    n610,
    n482,
    n571,
    n503,
    n471
  );


  nand
  g584
  (
    n636,
    n497,
    n575,
    n476,
    n506
  );


  or
  g585
  (
    n607,
    n494,
    n493,
    n474,
    n435
  );


  nand
  g586
  (
    n617,
    n577,
    n477,
    n448,
    n451
  );


  xnor
  g587
  (
    KeyWire_0_44,
    n444,
    n456,
    n578,
    n457
  );


  or
  g588
  (
    n628,
    n506,
    n436,
    n434,
    n485
  );


  xnor
  g589
  (
    n625,
    n574,
    n572,
    n481,
    n578
  );


  xor
  g590
  (
    n601,
    n452,
    n501,
    n443,
    n491
  );


  nand
  g591
  (
    n608,
    n503,
    n504,
    n471,
    n440
  );


  nor
  g592
  (
    n620,
    n502,
    n571,
    n486,
    n464
  );


  or
  g593
  (
    n613,
    n570,
    n473,
    n577,
    n469
  );


  nand
  g594
  (
    n605,
    n494,
    n460,
    n437,
    n480
  );


  xnor
  g595
  (
    n616,
    n477,
    n496,
    n473,
    n487
  );


  nor
  g596
  (
    n621,
    n488,
    n462,
    n450,
    n505
  );


  or
  g597
  (
    n626,
    n484,
    n498,
    n499,
    n492
  );


  xnor
  g598
  (
    n602,
    n481,
    n475,
    n474,
    n479
  );


  xnor
  g599
  (
    n629,
    n482,
    n488,
    n461,
    n573
  );


  and
  g600
  (
    n619,
    n463,
    n486,
    n489,
    n438
  );


  and
  g601
  (
    n623,
    n445,
    n491,
    n499,
    n484
  );


  nor
  g602
  (
    n634,
    n476,
    n468,
    n577,
    n573
  );


  and
  g603
  (
    n614,
    n455,
    n490,
    n573,
    n470
  );


  or
  g604
  (
    n622,
    n495,
    n579,
    n475,
    n496
  );


  nor
  g605
  (
    n603,
    n449,
    n446,
    n470,
    n502
  );


  nor
  g606
  (
    n609,
    n501,
    n459,
    n571,
    n576
  );


  nand
  g607
  (
    n632,
    n441,
    n487,
    n485,
    n578
  );


  or
  g608
  (
    n630,
    n575,
    n466,
    n458,
    n467
  );


  xnor
  g609
  (
    n627,
    n574,
    n572,
    n505,
    n493
  );


  not
  g610
  (
    n658,
    n618
  );


  buf
  g611
  (
    n639,
    n621
  );


  buf
  g612
  (
    n655,
    n625
  );


  buf
  g613
  (
    n656,
    n606
  );


  not
  g614
  (
    n647,
    n620
  );


  not
  g615
  (
    n654,
    n622
  );


  buf
  g616
  (
    n646,
    n613
  );


  not
  g617
  (
    n644,
    n607
  );


  buf
  g618
  (
    n637,
    n612
  );


  buf
  g619
  (
    n650,
    n616
  );


  not
  g620
  (
    n642,
    n619
  );


  not
  g621
  (
    n638,
    n611
  );


  buf
  g622
  (
    n657,
    n604
  );


  not
  g623
  (
    n648,
    n605
  );


  not
  g624
  (
    n649,
    n623
  );


  buf
  g625
  (
    n653,
    n615
  );


  not
  g626
  (
    n651,
    n608
  );


  buf
  g627
  (
    n640,
    n617
  );


  buf
  g628
  (
    n652,
    n614
  );


  buf
  g629
  (
    n643,
    n609
  );


  buf
  g630
  (
    n645,
    n610
  );


  buf
  g631
  (
    n641,
    n624
  );


  not
  g632
  (
    n693,
    n594
  );


  buf
  g633
  (
    n666,
    n650
  );


  not
  g634
  (
    n709,
    n639
  );


  buf
  g635
  (
    n679,
    n642
  );


  buf
  g636
  (
    n713,
    n544
  );


  buf
  g637
  (
    n703,
    n528
  );


  or
  g638
  (
    n667,
    n545,
    n532
  );


  nor
  g639
  (
    n700,
    n638,
    n640,
    n523
  );


  and
  g640
  (
    n670,
    n651,
    n648,
    n637,
    n587
  );


  and
  g641
  (
    n717,
    n645,
    n530,
    n548,
    n556
  );


  nor
  g642
  (
    n699,
    n536,
    n537,
    n543,
    n648
  );


  or
  g643
  (
    n688,
    n551,
    n538,
    n532,
    n548
  );


  or
  g644
  (
    n726,
    n591,
    n644,
    n531,
    n539
  );


  xnor
  g645
  (
    n715,
    n533,
    n538,
    n594,
    n591
  );


  nand
  g646
  (
    n721,
    n582,
    n544,
    n641,
    n550
  );


  xnor
  g647
  (
    n698,
    n554,
    n580,
    n540,
    n535
  );


  nand
  g648
  (
    n720,
    n524,
    n522,
    n583,
    n536
  );


  xnor
  g649
  (
    n677,
    n533,
    n553,
    n654,
    n532
  );


  xnor
  g650
  (
    n665,
    n541,
    n556,
    n523,
    n525
  );


  xor
  g651
  (
    n696,
    n650,
    n580,
    n655,
    n539
  );


  xnor
  g652
  (
    n675,
    n531,
    n647,
    n580,
    n555
  );


  or
  g653
  (
    n687,
    n637,
    n535,
    n643,
    n546
  );


  xnor
  g654
  (
    n724,
    n539,
    n529,
    n533,
    n650
  );


  xnor
  g655
  (
    n695,
    n542,
    n586,
    n530,
    n639
  );


  xor
  g656
  (
    n723,
    n556,
    n541,
    n543,
    n581
  );


  and
  g657
  (
    n668,
    n591,
    n534,
    n645,
    n641
  );


  nand
  g658
  (
    n690,
    n528,
    n653,
    n581,
    n540
  );


  and
  g659
  (
    n692,
    n590,
    n638,
    n532,
    n537
  );


  or
  g660
  (
    n680,
    n651,
    n588,
    n524,
    n582
  );


  or
  g661
  (
    n718,
    n641,
    n590,
    n584,
    n530
  );


  or
  g662
  (
    n730,
    n529,
    n549,
    n586,
    n646
  );


  xnor
  g663
  (
    n722,
    n653,
    n541,
    n588,
    n543
  );


  xnor
  g664
  (
    n669,
    n647,
    n548,
    n594,
    n539
  );


  xor
  g665
  (
    n681,
    n553,
    n643,
    n588,
    n651
  );


  and
  g666
  (
    n707,
    n582,
    n643,
    n528,
    n654
  );


  xor
  g667
  (
    n694,
    n550,
    n593,
    n646,
    n538
  );


  nor
  g668
  (
    n682,
    n590,
    n649,
    n542,
    n652
  );


  xnor
  g669
  (
    n706,
    n579,
    n652,
    n589
  );


  nor
  g670
  (
    n662,
    n642,
    n587,
    n542,
    n641
  );


  nand
  g671
  (
    n672,
    n651,
    n643,
    n589
  );


  xor
  g672
  (
    n701,
    n582,
    n585,
    n534,
    n640
  );


  xnor
  g673
  (
    n702,
    n586,
    n648,
    n551
  );


  nand
  g674
  (
    n684,
    n654,
    n592,
    n546,
    n536
  );


  nand
  g675
  (
    n712,
    n537,
    n646,
    n542,
    n549
  );


  or
  g676
  (
    n705,
    n645,
    n556,
    n535,
    n642
  );


  xnor
  g677
  (
    n697,
    n554,
    n554,
    n642,
    n580
  );


  xnor
  g678
  (
    n676,
    n637,
    n587,
    n523,
    n553
  );


  nand
  g679
  (
    n689,
    n585,
    n528,
    n544,
    n653
  );


  xnor
  g680
  (
    n710,
    n526,
    n549,
    n553,
    n552
  );


  and
  g681
  (
    n711,
    n585,
    n590,
    n649
  );


  xnor
  g682
  (
    n683,
    n644,
    n654,
    n592,
    n550
  );


  xnor
  g683
  (
    n708,
    n586,
    n584,
    n526
  );


  or
  g684
  (
    n674,
    n551,
    n527,
    n549,
    n540
  );


  xor
  g685
  (
    n728,
    n546,
    n545,
    n581,
    n593
  );


  xnor
  g686
  (
    n729,
    n588,
    n545,
    n555,
    n579
  );


  or
  g687
  (
    n671,
    n583,
    n531,
    n585,
    n527
  );


  xor
  g688
  (
    n725,
    n547,
    n640,
    n534,
    n593
  );


  xor
  g689
  (
    n704,
    n526,
    n552,
    n545,
    n527
  );


  or
  g690
  (
    n727,
    n547,
    n644,
    n531,
    n592
  );


  nor
  g691
  (
    n731,
    n639,
    n547,
    n592,
    n581
  );


  or
  g692
  (
    n716,
    n587,
    n552,
    n646,
    n554
  );


  or
  g693
  (
    n719,
    n589,
    n529,
    n550,
    n637
  );


  xor
  g694
  (
    n660,
    n538,
    n543,
    n639,
    n525
  );


  xor
  g695
  (
    n661,
    n638,
    n530,
    n584,
    n548
  );


  nand
  g696
  (
    n663,
    n650,
    n524,
    n525,
    n579
  );


  nand
  g697
  (
    n691,
    n555,
    n584,
    n647,
    n529
  );


  or
  g698
  (
    n686,
    n547,
    n533,
    n541,
    n540
  );


  nand
  g699
  (
    n678,
    n555,
    n525,
    n536,
    n534
  );


  xnor
  g700
  (
    n714,
    n647,
    n644,
    n524,
    n583
  );


  xor
  g701
  (
    n685,
    n653,
    n591,
    n552,
    n640
  );


  xor
  g702
  (
    n664,
    n648,
    n527,
    n645,
    n535
  );


  xnor
  g703
  (
    n659,
    n537,
    n544,
    n546,
    n593
  );


  nor
  g704
  (
    n673,
    n652,
    n649,
    n583,
    n638
  );


  not
  g705
  (
    n743,
    n663
  );


  buf
  g706
  (
    n738,
    n685
  );


  not
  g707
  (
    n765,
    n686
  );


  buf
  g708
  (
    n751,
    n673
  );


  not
  g709
  (
    n766,
    n668
  );


  buf
  g710
  (
    n760,
    n662
  );


  not
  g711
  (
    n757,
    n690
  );


  buf
  g712
  (
    n737,
    n675
  );


  not
  g713
  (
    n759,
    n684
  );


  buf
  g714
  (
    n736,
    n667
  );


  buf
  g715
  (
    n763,
    n678
  );


  not
  g716
  (
    n732,
    n661
  );


  buf
  g717
  (
    n761,
    n676
  );


  not
  g718
  (
    n762,
    n672
  );


  not
  g719
  (
    n748,
    n677
  );


  buf
  g720
  (
    n749,
    n692
  );


  buf
  g721
  (
    n741,
    n682
  );


  not
  g722
  (
    n735,
    n681
  );


  not
  g723
  (
    n733,
    n680
  );


  buf
  g724
  (
    n742,
    n670
  );


  not
  g725
  (
    n753,
    n665
  );


  buf
  g726
  (
    n744,
    n669
  );


  buf
  g727
  (
    n767,
    n683
  );


  not
  g728
  (
    n745,
    n689
  );


  not
  g729
  (
    n754,
    n659
  );


  not
  g730
  (
    n764,
    n679
  );


  not
  g731
  (
    n750,
    n666
  );


  buf
  g732
  (
    n747,
    n688
  );


  buf
  g733
  (
    n739,
    n693
  );


  buf
  g734
  (
    n755,
    n664
  );


  not
  g735
  (
    n740,
    n671
  );


  buf
  g736
  (
    n734,
    n687
  );


  not
  g737
  (
    n752,
    n694
  );


  not
  g738
  (
    n756,
    n660
  );


  buf
  g739
  (
    n746,
    n691
  );


  not
  g740
  (
    n758,
    n674
  );


  buf
  g741
  (
    n783,
    n599
  );


  buf
  g742
  (
    n770,
    n732
  );


  buf
  g743
  (
    n773,
    n597
  );


  buf
  g744
  (
    n786,
    n596
  );


  not
  g745
  (
    n779,
    n734
  );


  not
  g746
  (
    n771,
    n599
  );


  buf
  g747
  (
    n776,
    n596
  );


  not
  g748
  (
    n775,
    n596
  );


  not
  g749
  (
    n772,
    n598
  );


  not
  g750
  (
    n774,
    n595
  );


  not
  g751
  (
    n781,
    n734
  );


  buf
  g752
  (
    n777,
    n735
  );


  buf
  g753
  (
    n787,
    n736
  );


  xnor
  g754
  (
    n780,
    n594,
    n734,
    n595
  );


  xnor
  g755
  (
    n785,
    n733,
    n733,
    n734,
    n595
  );


  xnor
  g756
  (
    n784,
    n733,
    n736,
    n732,
    n599
  );


  nand
  g757
  (
    n778,
    n597,
    n735,
    n598
  );


  xor
  g758
  (
    n782,
    n733,
    n736,
    n597,
    n598
  );


  xnor
  g759
  (
    n768,
    n598,
    n732,
    n736
  );


  and
  g760
  (
    n769,
    n596,
    n597,
    n735,
    n595
  );


  buf
  g761
  (
    n798,
    n771
  );


  buf
  g762
  (
    n814,
    n745
  );


  not
  g763
  (
    n799,
    n770
  );


  not
  g764
  (
    n806,
    n746
  );


  buf
  g765
  (
    n807,
    n741
  );


  buf
  g766
  (
    n804,
    n743
  );


  xor
  g767
  (
    n813,
    n769,
    n748,
    n768,
    n749
  );


  nand
  g768
  (
    n801,
    n739,
    n740,
    n567
  );


  nor
  g769
  (
    n797,
    n740,
    n744,
    n631,
    n629
  );


  and
  g770
  (
    n791,
    n741,
    n567,
    n742,
    n737
  );


  xor
  g771
  (
    n795,
    n655,
    n747,
    n773,
    n634
  );


  xnor
  g772
  (
    n788,
    n743,
    n770,
    n747,
    n744
  );


  and
  g773
  (
    n790,
    n630,
    n738,
    n626,
    n769
  );


  and
  g774
  (
    n796,
    n741,
    n773,
    n566,
    n636
  );


  and
  g775
  (
    KeyWire_0_7,
    n746,
    n772,
    n749,
    n743
  );


  xor
  g776
  (
    n803,
    n740,
    n627,
    n748,
    n745
  );


  or
  g777
  (
    n810,
    n768,
    n744,
    n772,
    n771
  );


  nand
  g778
  (
    KeyWire_0_62,
    n739,
    n772,
    n744,
    n742
  );


  or
  g779
  (
    KeyWire_0_0,
    n746,
    n769,
    n738,
    n773
  );


  nand
  g780
  (
    n792,
    n773,
    n771,
    n655
  );


  nor
  g781
  (
    n816,
    n750,
    n740,
    n632,
    n739
  );


  and
  g782
  (
    n817,
    n774,
    n770,
    n745,
    n747
  );


  xnor
  g783
  (
    n789,
    n633,
    n749,
    n748,
    n567
  );


  nor
  g784
  (
    n809,
    n774,
    n742,
    n738,
    n566
  );


  and
  g785
  (
    n805,
    n775,
    n742,
    n774,
    n749
  );


  or
  g786
  (
    n808,
    n769,
    n775,
    n628,
    n770
  );


  xor
  g787
  (
    n815,
    n747,
    n768,
    n739
  );


  xor
  g788
  (
    n793,
    n745,
    n737,
    n748
  );


  xor
  g789
  (
    n794,
    n737,
    n746,
    n743,
    n772
  );


  xor
  g790
  (
    n802,
    n741,
    n774,
    n635,
    n738
  );


  and
  g791
  (
    n830,
    n805,
    n807,
    n809
  );


  and
  g792
  (
    n841,
    n797,
    n789,
    n788
  );


  nand
  g793
  (
    n822,
    n798,
    n801,
    n804
  );


  and
  g794
  (
    n844,
    n809,
    n794,
    n810
  );


  and
  g795
  (
    n821,
    n809,
    n793,
    n814
  );


  nor
  g796
  (
    n833,
    n808,
    n802,
    n792
  );


  nor
  g797
  (
    n835,
    n793,
    n801,
    n805
  );


  and
  g798
  (
    n834,
    n797,
    n798,
    n813,
    n808
  );


  nand
  g799
  (
    n832,
    n800,
    n799,
    n790,
    n797
  );


  and
  g800
  (
    n819,
    n801,
    n805,
    n796,
    n790
  );


  or
  g801
  (
    n838,
    n804,
    n813,
    n800,
    n791
  );


  nand
  g802
  (
    n831,
    n794,
    n810,
    n797,
    n790
  );


  or
  g803
  (
    n825,
    n812,
    n796,
    n803,
    n805
  );


  or
  g804
  (
    n840,
    n793,
    n814,
    n795,
    n813
  );


  nand
  g805
  (
    n828,
    n795,
    n811,
    n803,
    n807
  );


  xnor
  g806
  (
    n836,
    n812,
    n794,
    n788,
    n799
  );


  xnor
  g807
  (
    n829,
    n798,
    n796,
    n807,
    n808
  );


  and
  g808
  (
    n839,
    n812,
    n806,
    n803,
    n792
  );


  xor
  g809
  (
    n818,
    n808,
    n788,
    n799
  );


  and
  g810
  (
    n845,
    n806,
    n807,
    n789,
    n810
  );


  nor
  g811
  (
    n827,
    n802,
    n791,
    n804,
    n796
  );


  nand
  g812
  (
    n823,
    n800,
    n806,
    n812,
    n799
  );


  nor
  g813
  (
    n842,
    n790,
    n795,
    n811,
    n800
  );


  or
  g814
  (
    n843,
    n791,
    n806,
    n809,
    n810
  );


  and
  g815
  (
    n824,
    n793,
    n802,
    n804
  );


  xnor
  g816
  (
    n820,
    n792,
    n798,
    n811,
    n789
  );


  nor
  g817
  (
    n837,
    n803,
    n792,
    n795,
    n811
  );


  or
  g818
  (
    n826,
    n791,
    n789,
    n813,
    n794
  );


  not
  g819
  (
    n849,
    n818
  );


  not
  g820
  (
    n846,
    n819
  );


  not
  g821
  (
    n850,
    n818
  );


  not
  g822
  (
    n848,
    n819
  );


  not
  g823
  (
    n847,
    n818
  );


  not
  g824
  (
    n851,
    n818
  );


  buf
  g825
  (
    n856,
    n850
  );


  buf
  g826
  (
    n853,
    n851
  );


  not
  g827
  (
    n852,
    n851
  );


  not
  g828
  (
    n854,
    n850
  );


  buf
  g829
  (
    n855,
    n849
  );


  buf
  g830
  (
    n857,
    n852
  );


  nor
  g831
  (
    n859,
    n819,
    n820
  );


  or
  g832
  (
    n858,
    n857,
    n857,
    n819,
    n820
  );


  buf
  g833
  (
    n860,
    n859
  );


  not
  g834
  (
    n862,
    n858
  );


  buf
  g835
  (
    n861,
    n859
  );


  buf
  g836
  (
    n863,
    n860
  );


  not
  g837
  (
    n864,
    n863
  );


  buf
  g838
  (
    n865,
    n863
  );


  nor
  g839
  (
    n867,
    n865,
    n85
  );


  xor
  g840
  (
    n871,
    n82,
    n864
  );


  nor
  g841
  (
    n866,
    n85,
    n865
  );


  xnor
  g842
  (
    n870,
    n83,
    n85
  );


  or
  g843
  (
    n869,
    n864,
    n865
  );


  xor
  g844
  (
    KeyWire_0_16,
    n82,
    n84
  );


  xnor
  g845
  (
    n872,
    n865,
    n84,
    n83
  );


  or
  g846
  (
    n873,
    n83,
    n864,
    n84
  );


  buf
  g847
  (
    n885,
    n867
  );


  not
  g848
  (
    n879,
    n751
  );


  buf
  g849
  (
    n903,
    n873
  );


  buf
  g850
  (
    n890,
    n871
  );


  buf
  g851
  (
    n886,
    n753
  );


  not
  g852
  (
    n900,
    n87
  );


  buf
  g853
  (
    KeyWire_0_34,
    n873
  );


  buf
  g854
  (
    n878,
    n394
  );


  buf
  g855
  (
    n883,
    n86
  );


  not
  g856
  (
    n877,
    n871
  );


  buf
  g857
  (
    n899,
    n867
  );


  not
  g858
  (
    n896,
    n754
  );


  buf
  g859
  (
    n894,
    n868
  );


  buf
  g860
  (
    n875,
    n750
  );


  not
  g861
  (
    n895,
    n822
  );


  buf
  g862
  (
    n874,
    n753
  );


  or
  g863
  (
    n884,
    n821,
    n87,
    n873,
    n751
  );


  xor
  g864
  (
    n898,
    n822,
    n754,
    n752,
    n867
  );


  nand
  g865
  (
    n897,
    n752,
    n751,
    n872,
    n869
  );


  or
  g866
  (
    n904,
    n870,
    n393,
    n872,
    n871
  );


  xor
  g867
  (
    n888,
    n862,
    n86,
    n867,
    n87
  );


  nand
  g868
  (
    n901,
    n752,
    n87,
    n822,
    n754
  );


  xnor
  g869
  (
    n902,
    n750,
    n823,
    n821,
    n866
  );


  xor
  g870
  (
    n891,
    n823,
    n866,
    n85,
    n753
  );


  and
  g871
  (
    n892,
    n750,
    n868,
    n872
  );


  xnor
  g872
  (
    n893,
    n869,
    n870,
    n821
  );


  xnor
  g873
  (
    n887,
    n871,
    n751,
    n823,
    n821
  );


  and
  g874
  (
    n881,
    n86,
    n823,
    n394,
    n868
  );


  and
  g875
  (
    n882,
    n861,
    n754,
    n866,
    n872
  );


  or
  g876
  (
    n889,
    n752,
    n869,
    n753
  );


  or
  g877
  (
    n880,
    n870,
    n86,
    n866,
    n822
  );


  buf
  g878
  (
    n905,
    n874
  );


  not
  g879
  (
    n907,
    n905
  );


  buf
  g880
  (
    n906,
    n905
  );


  buf
  g881
  (
    n911,
    n907
  );


  buf
  g882
  (
    n910,
    n906
  );


  not
  g883
  (
    n909,
    n906
  );


  buf
  g884
  (
    n908,
    n907
  );


  nor
  g885
  (
    n918,
    n89,
    n93,
    n91
  );


  or
  g886
  (
    n920,
    n92,
    n911,
    n94,
    n826
  );


  xor
  g887
  (
    n926,
    n827,
    n908,
    n910,
    n94
  );


  xnor
  g888
  (
    n917,
    n909,
    n91,
    n828
  );


  or
  g889
  (
    n927,
    n93,
    n827,
    n824
  );


  or
  g890
  (
    n923,
    n95,
    n90,
    n826,
    n910
  );


  xnor
  g891
  (
    n925,
    n90,
    n909,
    n89,
    n826
  );


  nor
  g892
  (
    n913,
    n88,
    n911,
    n825,
    n92
  );


  nor
  g893
  (
    n914,
    n911,
    n908,
    n92,
    n909
  );


  nand
  g894
  (
    n924,
    n825,
    n88,
    n911,
    n824
  );


  xor
  g895
  (
    n919,
    n93,
    n94,
    n90,
    n88
  );


  or
  g896
  (
    n912,
    n824,
    n908,
    n91,
    n94
  );


  xor
  g897
  (
    n915,
    n827,
    n826,
    n89,
    n825
  );


  nor
  g898
  (
    n921,
    n910,
    n873,
    n93,
    n908
  );


  xnor
  g899
  (
    n922,
    n824,
    n88,
    n909,
    n90
  );


  or
  g900
  (
    n916,
    n825,
    n89,
    n92,
    n910
  );


  nor
  g901
  (
    n976,
    n914,
    n913
  );


  nand
  g902
  (
    n946,
    n599,
    n855
  );


  nand
  g903
  (
    n975,
    n886,
    n901
  );


  xnor
  g904
  (
    n990,
    n894,
    n877
  );


  nand
  g905
  (
    n933,
    n856,
    n853,
    n922
  );


  xor
  g906
  (
    n978,
    n898,
    n899,
    n921
  );


  nand
  g907
  (
    n965,
    n919,
    n899,
    n896
  );


  xnor
  g908
  (
    n967,
    n912,
    n880,
    n885
  );


  or
  g909
  (
    n987,
    n894,
    n904,
    n917
  );


  nand
  g910
  (
    n970,
    n896,
    n920,
    n568
  );


  and
  g911
  (
    n968,
    n902,
    n886,
    n879
  );


  or
  g912
  (
    n989,
    n926,
    n877,
    n919
  );


  and
  g913
  (
    n961,
    n920,
    n889,
    n856
  );


  and
  g914
  (
    n964,
    n886,
    n927
  );


  nor
  g915
  (
    n972,
    n921,
    n855,
    n914
  );


  nor
  g916
  (
    n981,
    n894,
    n884,
    n888
  );


  xnor
  g917
  (
    n985,
    n856,
    n897,
    n568
  );


  and
  g918
  (
    n938,
    n918,
    n893,
    n874
  );


  or
  g919
  (
    n931,
    n893,
    n876,
    n891
  );


  nand
  g920
  (
    n935,
    n892,
    n874,
    n922
  );


  nor
  g921
  (
    n948,
    n912,
    n904,
    n879
  );


  nand
  g922
  (
    n953,
    n902,
    n916,
    n903
  );


  xnor
  g923
  (
    n945,
    n902,
    n569,
    n877
  );


  nor
  g924
  (
    n977,
    n816,
    n903,
    n817
  );


  nor
  g925
  (
    n980,
    n883,
    n883,
    n901,
    n889
  );


  xnor
  g926
  (
    n939,
    n854,
    n891,
    n876,
    n902
  );


  nand
  g927
  (
    n954,
    n904,
    n874,
    n914,
    n891
  );


  and
  g928
  (
    n959,
    n916,
    n925,
    n882,
    n923
  );


  or
  g929
  (
    n973,
    n925,
    n288,
    n876,
    n926
  );


  xor
  g930
  (
    n947,
    n885,
    n853,
    n913,
    n816
  );


  nand
  g931
  (
    n962,
    n888,
    n856,
    n854,
    n881
  );


  nand
  g932
  (
    n955,
    n885,
    n888,
    n898,
    n817
  );


  nor
  g933
  (
    n984,
    n903,
    n886,
    n882,
    n904
  );


  or
  g934
  (
    n937,
    n927,
    n815,
    n852,
    n901
  );


  xor
  g935
  (
    n949,
    n897,
    n923,
    n568,
    n817
  );


  xor
  g936
  (
    n982,
    n917,
    n915,
    n900,
    n916
  );


  and
  g937
  (
    n956,
    n881,
    n894,
    n887,
    n889
  );


  nand
  g938
  (
    n974,
    n879,
    n892,
    n875
  );


  or
  g939
  (
    n986,
    n925,
    n895,
    n890,
    n917
  );


  nor
  g940
  (
    n941,
    n887,
    n569,
    n915,
    n912
  );


  nor
  g941
  (
    n934,
    n920,
    n883,
    n896,
    n901
  );


  or
  g942
  (
    n983,
    n898,
    n917,
    n897,
    n889
  );


  xor
  g943
  (
    n936,
    n854,
    n815,
    n921,
    n913
  );


  nand
  g944
  (
    n951,
    n852,
    n855,
    n878,
    n875
  );


  and
  g945
  (
    n963,
    n923,
    n877,
    n883,
    n900
  );


  or
  g946
  (
    n929,
    n892,
    n890,
    n880,
    n924
  );


  or
  g947
  (
    n950,
    n919,
    n816,
    n895,
    n924
  );


  or
  g948
  (
    n979,
    n852,
    n899,
    n893,
    n895
  );


  nand
  g949
  (
    n966,
    n900,
    n897,
    n915,
    n814
  );


  xor
  g950
  (
    n932,
    n919,
    n884,
    n903,
    n922
  );


  nand
  g951
  (
    n942,
    n885,
    n568,
    n914,
    n921
  );


  and
  g952
  (
    n971,
    n853,
    n918,
    n880,
    n887
  );


  nand
  g953
  (
    n928,
    n920,
    n878,
    n899
  );


  and
  g954
  (
    n988,
    n888,
    n912,
    n815,
    n887
  );


  nand
  g955
  (
    n944,
    n916,
    n891,
    n927,
    n896
  );


  nand
  g956
  (
    n943,
    n853,
    n817,
    n923,
    n855
  );


  nor
  g957
  (
    KeyWire_0_24,
    n881,
    n884,
    n924,
    n926
  );


  and
  g958
  (
    n969,
    n854,
    n895,
    n875,
    n918
  );


  or
  g959
  (
    n952,
    n926,
    n881,
    n890,
    n882
  );


  and
  g960
  (
    n930,
    n816,
    n879,
    n876,
    n878
  );


  nor
  g961
  (
    n960,
    n922,
    n815,
    n880,
    n892
  );


  nor
  g962
  (
    n957,
    n924,
    n884,
    n900,
    n893
  );


  or
  g963
  (
    n958,
    n890,
    n814,
    n898,
    n915
  );


  xor
  g964
  (
    n991,
    n925,
    n918,
    n913,
    n882
  );


  not
  g965
  (
    n1000,
    n928
  );


  not
  g966
  (
    n994,
    n929
  );


  not
  g967
  (
    n1001,
    n930
  );


  not
  g968
  (
    n995,
    n929
  );


  not
  g969
  (
    n998,
    n928
  );


  buf
  g970
  (
    n997,
    n929
  );


  not
  g971
  (
    n999,
    n928
  );


  buf
  g972
  (
    n996,
    n929
  );


  not
  g973
  (
    n993,
    n928
  );


  buf
  g974
  (
    n992,
    n930
  );


  or
  g975
  (
    n1033,
    n932,
    n939
  );


  xnor
  g976
  (
    n1041,
    n938,
    n828
  );


  nand
  g977
  (
    n1030,
    n996,
    n998
  );


  xor
  g978
  (
    n1028,
    n931,
    n930
  );


  xnor
  g979
  (
    n1008,
    n933,
    n999
  );


  buf
  g980
  (
    n1029,
    n934
  );


  xor
  g981
  (
    n1016,
    n996,
    n930
  );


  buf
  g982
  (
    n1002,
    n995
  );


  and
  g983
  (
    n1015,
    n996,
    n936
  );


  buf
  g984
  (
    n1013,
    n1000
  );


  nand
  g985
  (
    n1032,
    n1001,
    n994
  );


  or
  g986
  (
    n1026,
    n939,
    n937
  );


  xnor
  g987
  (
    n1010,
    n996,
    n993
  );


  nand
  g988
  (
    n1037,
    n992,
    n997
  );


  xor
  g989
  (
    n1038,
    n934,
    n938
  );


  nor
  g990
  (
    n1039,
    n931,
    n992
  );


  and
  g991
  (
    n1014,
    n999,
    n993
  );


  nand
  g992
  (
    n1040,
    n289,
    n936
  );


  or
  g993
  (
    n1007,
    n997,
    n933
  );


  nor
  g994
  (
    n1006,
    n933,
    n931
  );


  xor
  g995
  (
    n1024,
    n1001,
    n936
  );


  xor
  g996
  (
    n1012,
    n935,
    n937
  );


  or
  g997
  (
    n1022,
    n994,
    n992
  );


  or
  g998
  (
    KeyWire_0_57,
    n935,
    n932
  );


  or
  g999
  (
    n1017,
    n999,
    n993
  );


  or
  g1000
  (
    n1031,
    n992,
    n998
  );


  nand
  g1001
  (
    n1035,
    n932,
    n997
  );


  xnor
  g1002
  (
    n1019,
    n936,
    n995
  );


  or
  g1003
  (
    n1023,
    n933,
    n1000
  );


  and
  g1004
  (
    n1027,
    n932,
    n569
  );


  xnor
  g1005
  (
    n1034,
    n997,
    n998
  );


  and
  g1006
  (
    n1021,
    n934,
    n998
  );


  and
  g1007
  (
    n1004,
    n935,
    n1001
  );


  and
  g1008
  (
    n1003,
    n937,
    n289
  );


  nor
  g1009
  (
    n1018,
    n995,
    n931
  );


  or
  g1010
  (
    n1025,
    n1001,
    n938
  );


  nor
  g1011
  (
    n1011,
    n937,
    n999
  );


  nand
  g1012
  (
    n1020,
    n935,
    n938
  );


  xnor
  g1013
  (
    n1009,
    n994,
    n1000
  );


  xor
  g1014
  (
    n1036,
    n993,
    n994
  );


  not
  g1015
  (
    n1136,
    n1021
  );


  buf
  g1016
  (
    n1127,
    n1006
  );


  not
  g1017
  (
    n1146,
    n95
  );


  buf
  g1018
  (
    n1092,
    n1028
  );


  not
  g1019
  (
    n1089,
    n109
  );


  buf
  g1020
  (
    n1121,
    n1035
  );


  buf
  g1021
  (
    n1144,
    n1008
  );


  not
  g1022
  (
    n1164,
    n101
  );


  buf
  g1023
  (
    n1180,
    n1024
  );


  not
  g1024
  (
    n1069,
    n759
  );


  not
  g1025
  (
    n1159,
    n764
  );


  buf
  g1026
  (
    n1129,
    n1012
  );


  buf
  g1027
  (
    n1179,
    n1025
  );


  not
  g1028
  (
    n1198,
    n1018
  );


  buf
  g1029
  (
    n1168,
    n108
  );


  buf
  g1030
  (
    n1177,
    n1025
  );


  not
  g1031
  (
    n1183,
    n1027
  );


  not
  g1032
  (
    n1110,
    n1022
  );


  buf
  g1033
  (
    n1175,
    n113
  );


  buf
  g1034
  (
    n1196,
    n764
  );


  not
  g1035
  (
    n1126,
    n508
  );


  buf
  g1036
  (
    n1085,
    n1027
  );


  buf
  g1037
  (
    n1079,
    n1027
  );


  buf
  g1038
  (
    n1197,
    n1036
  );


  buf
  g1039
  (
    n1170,
    n1025
  );


  not
  g1040
  (
    n1054,
    n111
  );


  not
  g1041
  (
    n1070,
    n112
  );


  not
  g1042
  (
    n1082,
    n762
  );


  not
  g1043
  (
    n1200,
    n760
  );


  not
  g1044
  (
    n1154,
    n107
  );


  not
  g1045
  (
    KeyWire_0_53,
    n108
  );


  not
  g1046
  (
    n1072,
    n1038
  );


  buf
  g1047
  (
    n1119,
    n1019
  );


  not
  g1048
  (
    n1161,
    n103
  );


  buf
  g1049
  (
    n1147,
    n1010
  );


  not
  g1050
  (
    n1077,
    n1005
  );


  not
  g1051
  (
    n1058,
    n103
  );


  not
  g1052
  (
    n1102,
    n113
  );


  not
  g1053
  (
    n1106,
    n1005
  );


  not
  g1054
  (
    n1149,
    n508
  );


  buf
  g1055
  (
    n1128,
    n104
  );


  not
  g1056
  (
    n1067,
    n758
  );


  buf
  g1057
  (
    n1145,
    n507
  );


  not
  g1058
  (
    n1162,
    n109
  );


  buf
  g1059
  (
    n1105,
    n1007
  );


  not
  g1060
  (
    n1169,
    n763
  );


  buf
  g1061
  (
    n1131,
    n765
  );


  not
  g1062
  (
    n1140,
    n764
  );


  buf
  g1063
  (
    n1093,
    n1028
  );


  buf
  g1064
  (
    KeyWire_0_22,
    n1037
  );


  buf
  g1065
  (
    n1053,
    n510
  );


  buf
  g1066
  (
    n1108,
    n115
  );


  buf
  g1067
  (
    n1194,
    n1015
  );


  not
  g1068
  (
    n1096,
    n1002
  );


  not
  g1069
  (
    n1171,
    n762
  );


  not
  g1070
  (
    n1163,
    n1004
  );


  buf
  g1071
  (
    n1125,
    n1030
  );


  buf
  g1072
  (
    n1078,
    n939
  );


  buf
  g1073
  (
    n1176,
    n1040
  );


  not
  g1074
  (
    n1073,
    n102
  );


  not
  g1075
  (
    n1055,
    n101
  );


  buf
  g1076
  (
    n1044,
    n101
  );


  buf
  g1077
  (
    n1167,
    n1020
  );


  not
  g1078
  (
    n1049,
    n1041
  );


  not
  g1079
  (
    n1181,
    n1029
  );


  not
  g1080
  (
    KeyWire_0_48,
    n1006
  );


  buf
  g1081
  (
    n1080,
    n1014
  );


  not
  g1082
  (
    n1123,
    n107
  );


  buf
  g1083
  (
    n1081,
    n101
  );


  buf
  g1084
  (
    n1142,
    n763
  );


  buf
  g1085
  (
    n1050,
    n761
  );


  not
  g1086
  (
    n1158,
    n96
  );


  not
  g1087
  (
    n1104,
    n1022
  );


  not
  g1088
  (
    n1111,
    n1026
  );


  not
  g1089
  (
    n1042,
    n111
  );


  buf
  g1090
  (
    n1043,
    n762
  );


  buf
  g1091
  (
    n1088,
    n756
  );


  buf
  g1092
  (
    n1090,
    n106
  );


  not
  g1093
  (
    n1094,
    n1010
  );


  not
  g1094
  (
    n1165,
    n1039
  );


  buf
  g1095
  (
    n1134,
    n766
  );


  buf
  g1096
  (
    n1139,
    n109
  );


  buf
  g1097
  (
    n1095,
    n510
  );


  not
  g1098
  (
    n1091,
    n1014
  );


  not
  g1099
  (
    n1156,
    n1034
  );


  not
  g1100
  (
    n1157,
    n1033
  );


  buf
  g1101
  (
    n1133,
    n1041
  );


  buf
  g1102
  (
    n1184,
    n102
  );


  buf
  g1103
  (
    n1174,
    n1006
  );


  buf
  g1104
  (
    n1135,
    n1013
  );


  buf
  g1105
  (
    n1193,
    n1011
  );


  not
  g1106
  (
    n1084,
    n761
  );


  not
  g1107
  (
    n1114,
    n1038
  );


  not
  g1108
  (
    n1124,
    n1029
  );


  buf
  g1109
  (
    n1189,
    n1020
  );


  buf
  g1110
  (
    n1192,
    n1023
  );


  not
  g1111
  (
    n1118,
    n1022
  );


  buf
  g1112
  (
    n1191,
    n755
  );


  not
  g1113
  (
    n1195,
    n766
  );


  buf
  g1114
  (
    n1122,
    n1009
  );


  not
  g1115
  (
    n1112,
    n764
  );


  not
  g1116
  (
    n1138,
    n95
  );


  buf
  g1117
  (
    n1107,
    n759
  );


  buf
  g1118
  (
    n1117,
    n115
  );


  buf
  g1119
  (
    n1062,
    n116
  );


  buf
  g1120
  (
    n1086,
    n1030
  );


  buf
  g1121
  (
    n1052,
    n1017
  );


  not
  g1122
  (
    n1172,
    n109
  );


  not
  g1123
  (
    n1137,
    n1024
  );


  xnor
  g1124
  (
    n1120,
    n1023,
    n763,
    n100,
    n1035
  );


  xor
  g1125
  (
    n1182,
    n98,
    n1008,
    n106,
    n100
  );


  nand
  g1126
  (
    n1076,
    n1014,
    n102,
    n1020,
    n1038
  );


  nand
  g1127
  (
    n1061,
    n1041,
    n106,
    n1013,
    n509
  );


  nand
  g1128
  (
    n1199,
    n939,
    n1034,
    n1024,
    n1023
  );


  nor
  g1129
  (
    n1143,
    n1011,
    n1033,
    n1031,
    n96
  );


  xnor
  g1130
  (
    n1101,
    n1039,
    n1004,
    n114,
    n98
  );


  nor
  g1131
  (
    n1155,
    n1028,
    n110,
    n1036,
    n758
  );


  xor
  g1132
  (
    n1151,
    n1002,
    n760,
    n1024,
    n759
  );


  nand
  g1133
  (
    n1056,
    n1014,
    n1008,
    n1016,
    n100
  );


  nand
  g1134
  (
    n1071,
    n755,
    n1018,
    n99,
    n1041
  );


  and
  g1135
  (
    n1141,
    n1021,
    n110,
    n761,
    n1032
  );


  nand
  g1136
  (
    n1097,
    n763,
    n1029,
    n1017,
    n1031
  );


  xor
  g1137
  (
    n1160,
    n97,
    n1020,
    n1037,
    n105
  );


  or
  g1138
  (
    n1185,
    n98,
    n1023,
    n115
  );


  or
  g1139
  (
    n1173,
    n1027,
    n105,
    n1037,
    n1034
  );


  xnor
  g1140
  (
    n1047,
    n512,
    n761,
    n96,
    n1032
  );


  nand
  g1141
  (
    n1116,
    n760,
    n765,
    n1010,
    n1040
  );


  and
  g1142
  (
    n1187,
    n1032,
    n1033,
    n1003,
    n765
  );


  nor
  g1143
  (
    n1045,
    n104,
    n111,
    n107,
    n756
  );


  or
  g1144
  (
    n1046,
    n98,
    n104,
    n1007,
    n1025
  );


  or
  g1145
  (
    n1059,
    n762,
    n96,
    n1009,
    n757
  );


  xor
  g1146
  (
    n1152,
    n757,
    n1004,
    n1026,
    n1036
  );


  nor
  g1147
  (
    n1148,
    n1039,
    n767,
    n766,
    n1005
  );


  and
  g1148
  (
    n1113,
    n1012,
    n1039,
    n1013,
    n1034
  );


  nor
  g1149
  (
    n1068,
    n1026,
    n103,
    n1021,
    n110
  );


  nand
  g1150
  (
    n1178,
    n97,
    n99,
    n940,
    n1018
  );


  or
  g1151
  (
    n1065,
    n99,
    n97,
    n1017
  );


  xor
  g1152
  (
    n1066,
    n1036,
    n757,
    n1016,
    n758
  );


  xor
  g1153
  (
    n1100,
    n102,
    n511,
    n1031,
    n1011
  );


  xnor
  g1154
  (
    n1098,
    n1009,
    n1022,
    n1028,
    n765
  );


  and
  g1155
  (
    n1166,
    n111,
    n756,
    n1026,
    n755
  );


  and
  g1156
  (
    n1115,
    n511,
    n1019,
    n1029
  );


  or
  g1157
  (
    KeyWire_0_28,
    n113,
    n97,
    n755,
    n758
  );


  xnor
  g1158
  (
    n1083,
    n1040,
    n1007,
    n766,
    n107
  );


  xor
  g1159
  (
    n1064,
    n1007,
    n1037,
    n1031,
    n1013
  );


  xnor
  g1160
  (
    n1057,
    n1032,
    n1016,
    n1021,
    n1011
  );


  nand
  g1161
  (
    n1099,
    n509,
    n1033,
    n103,
    n757
  );


  and
  g1162
  (
    n1060,
    n112,
    n100,
    n108,
    n1003
  );


  nor
  g1163
  (
    n1051,
    n112,
    n105,
    n767
  );


  xor
  g1164
  (
    n1153,
    n114,
    n756,
    n1030,
    n95
  );


  xor
  g1165
  (
    n1132,
    n1035,
    n113,
    n99,
    n1040
  );


  xnor
  g1166
  (
    n1074,
    n1003,
    n512,
    n1035,
    n759
  );


  nor
  g1167
  (
    n1048,
    n1015,
    n1003,
    n114,
    n760
  );


  xor
  g1168
  (
    n1186,
    n1005,
    n104,
    n114,
    n1009
  );


  and
  g1169
  (
    n1103,
    n1016,
    n1006,
    n767,
    n1019
  );


  or
  g1170
  (
    n1063,
    n112,
    n1038,
    n1010,
    n1008
  );


  or
  g1171
  (
    n1130,
    n1018,
    n1015,
    n1012
  );


  or
  g1172
  (
    n1188,
    n106,
    n105,
    n1002,
    n1004
  );


  and
  g1173
  (
    n1150,
    n1030,
    n110,
    n108,
    n1012
  );


  nor
  g1174
  (
    n1364,
    n1137,
    n724
  );


  nor
  g1175
  (
    n1273,
    n1056,
    n1134
  );


  or
  g1176
  (
    n1410,
    n784,
    n1167
  );


  xnor
  g1177
  (
    n1332,
    n981,
    n1176
  );


  and
  g1178
  (
    n1503,
    n1181,
    n1092
  );


  nor
  g1179
  (
    n1378,
    n1091,
    n717
  );


  nand
  g1180
  (
    n1326,
    n557,
    n1144
  );


  xor
  g1181
  (
    n1271,
    n1181,
    n721
  );


  or
  g1182
  (
    n1461,
    n1158,
    n966
  );


  or
  g1183
  (
    n1495,
    n1158,
    n1098
  );


  xor
  g1184
  (
    n1430,
    n979,
    n1182
  );


  xnor
  g1185
  (
    n1368,
    n988,
    n1176
  );


  xor
  g1186
  (
    n1449,
    n956,
    n967
  );


  and
  g1187
  (
    n1452,
    n1085,
    n962
  );


  nand
  g1188
  (
    n1291,
    n978,
    n1185
  );


  nand
  g1189
  (
    n1279,
    n1165,
    n777
  );


  nor
  g1190
  (
    KeyWire_0_13,
    n1200,
    n1171
  );


  or
  g1191
  (
    n1236,
    n1059,
    n1194
  );


  and
  g1192
  (
    n1239,
    n1057,
    n1143
  );


  xnor
  g1193
  (
    n1497,
    n1046,
    n981
  );


  or
  g1194
  (
    n1274,
    n1107,
    n779
  );


  or
  g1195
  (
    n1386,
    n1111,
    n775
  );


  nor
  g1196
  (
    n1505,
    n1108,
    n945
  );


  xnor
  g1197
  (
    n1463,
    n1146,
    n986
  );


  or
  g1198
  (
    n1301,
    n1147,
    n1097
  );


  nand
  g1199
  (
    n1212,
    n704,
    n1093
  );


  and
  g1200
  (
    KeyWire_0_9,
    n1088,
    n1103
  );


  nand
  g1201
  (
    n1474,
    n1054,
    n1175
  );


  or
  g1202
  (
    n1339,
    n1076,
    n1170
  );


  or
  g1203
  (
    n1290,
    n1175,
    n787
  );


  nor
  g1204
  (
    n1507,
    n1060,
    n1165
  );


  nand
  g1205
  (
    KeyWire_0_52,
    n1137,
    n1113
  );


  xnor
  g1206
  (
    n1229,
    n1061,
    n1144
  );


  and
  g1207
  (
    n1499,
    n1053,
    n1166
  );


  and
  g1208
  (
    n1389,
    n984,
    n1104
  );


  and
  g1209
  (
    n1422,
    n1111,
    n1072
  );


  and
  g1210
  (
    n1335,
    n1051,
    n1099
  );


  or
  g1211
  (
    n1382,
    n1179,
    n1059
  );


  xor
  g1212
  (
    n1299,
    n960,
    n1073
  );


  or
  g1213
  (
    n1446,
    n1092,
    n1188
  );


  xnor
  g1214
  (
    n1275,
    n1132,
    n1146
  );


  nand
  g1215
  (
    n1402,
    n942,
    n941
  );


  and
  g1216
  (
    n1456,
    n720,
    n708
  );


  nand
  g1217
  (
    n1296,
    n1152,
    n947
  );


  or
  g1218
  (
    n1216,
    n956,
    n780
  );


  xnor
  g1219
  (
    n1202,
    n1057,
    n1088
  );


  or
  g1220
  (
    n1224,
    n977,
    n1183
  );


  or
  g1221
  (
    n1464,
    n1088,
    n1075
  );


  xnor
  g1222
  (
    n1476,
    n1096,
    n1080
  );


  and
  g1223
  (
    n1489,
    n776,
    n976
  );


  or
  g1224
  (
    n1300,
    n1169,
    n1057
  );


  and
  g1225
  (
    n1460,
    n955,
    n1184
  );


  nor
  g1226
  (
    n1214,
    n779,
    n1102
  );


  or
  g1227
  (
    n1331,
    n1111,
    n1150
  );


  nand
  g1228
  (
    n1520,
    n1110,
    n965
  );


  nor
  g1229
  (
    n1518,
    n1164,
    n983
  );


  nor
  g1230
  (
    n1268,
    n1087,
    n1143
  );


  and
  g1231
  (
    n1306,
    n1060,
    n1174
  );


  xnor
  g1232
  (
    n1350,
    n1073,
    n1126
  );


  and
  g1233
  (
    n1303,
    n1130,
    n1101
  );


  and
  g1234
  (
    n1523,
    n558,
    n954
  );


  xor
  g1235
  (
    n1221,
    n1066,
    n1161
  );


  nor
  g1236
  (
    n1321,
    n1077,
    n1108
  );


  nor
  g1237
  (
    n1286,
    n707,
    n1056
  );


  xnor
  g1238
  (
    n1228,
    n985,
    n1135
  );


  and
  g1239
  (
    n1457,
    n965,
    n1180
  );


  nand
  g1240
  (
    n1515,
    n723,
    n1089
  );


  nor
  g1241
  (
    n1270,
    n1117,
    n1124
  );


  nor
  g1242
  (
    n1390,
    n1043,
    n948
  );


  xnor
  g1243
  (
    n1218,
    n1135,
    n1082
  );


  nor
  g1244
  (
    n1213,
    n1054,
    n1081
  );


  or
  g1245
  (
    n1431,
    n1047,
    n1157
  );


  xnor
  g1246
  (
    n1387,
    n1089,
    n1195
  );


  xor
  g1247
  (
    n1437,
    n1165,
    n943
  );


  xnor
  g1248
  (
    n1512,
    n1145,
    n941
  );


  not
  g1249
  (
    n1365,
    n954
  );


  xor
  g1250
  (
    n1360,
    n1163,
    n1087
  );


  nor
  g1251
  (
    n1217,
    n1109,
    n1063
  );


  nand
  g1252
  (
    n1435,
    n962,
    n969
  );


  and
  g1253
  (
    n1408,
    n1129,
    n1067
  );


  nor
  g1254
  (
    n1338,
    n975,
    n1072
  );


  and
  g1255
  (
    n1278,
    n780,
    n1049
  );


  xnor
  g1256
  (
    n1281,
    n1072,
    n954
  );


  and
  g1257
  (
    n1334,
    n1118,
    n775
  );


  xnor
  g1258
  (
    n1486,
    n1185,
    n989
  );


  and
  g1259
  (
    n1406,
    n1141,
    n1092
  );


  xor
  g1260
  (
    n1429,
    n1170,
    n1161
  );


  or
  g1261
  (
    n1438,
    n1132,
    n946
  );


  and
  g1262
  (
    n1372,
    n1183,
    n969
  );


  and
  g1263
  (
    n1348,
    n1129,
    n1052
  );


  nand
  g1264
  (
    n1468,
    n1144,
    n1175
  );


  or
  g1265
  (
    n1374,
    n1077,
    n1081
  );


  xnor
  g1266
  (
    n1333,
    n944,
    n1081
  );


  nand
  g1267
  (
    n1307,
    n964,
    n1055
  );


  xnor
  g1268
  (
    n1447,
    n1045,
    n1053
  );


  and
  g1269
  (
    n1442,
    n1118,
    n1191
  );


  and
  g1270
  (
    n1425,
    n1058,
    n1177
  );


  xor
  g1271
  (
    n1357,
    n1140,
    n1079
  );


  nand
  g1272
  (
    n1478,
    n1070,
    n1101
  );


  xnor
  g1273
  (
    n1353,
    n989,
    n983
  );


  and
  g1274
  (
    n1248,
    n712,
    n1162
  );


  and
  g1275
  (
    n1342,
    n982,
    n1162
  );


  or
  g1276
  (
    n1491,
    n1132,
    n1178
  );


  and
  g1277
  (
    n1396,
    n1126,
    n956
  );


  xnor
  g1278
  (
    n1209,
    n1044,
    n1142
  );


  and
  g1279
  (
    n1472,
    n1159,
    n951
  );


  xor
  g1280
  (
    n1488,
    n1145,
    n1115
  );


  or
  g1281
  (
    n1211,
    n1095,
    n1196
  );


  nor
  g1282
  (
    n1205,
    n1109,
    n1127
  );


  or
  g1283
  (
    n1380,
    n1165,
    n1095
  );


  xor
  g1284
  (
    n1511,
    n956,
    n1151
  );


  xor
  g1285
  (
    n1525,
    n1125,
    n945
  );


  and
  g1286
  (
    n1250,
    n716,
    n1197
  );


  or
  g1287
  (
    n1385,
    n1090,
    n782
  );


  xnor
  g1288
  (
    n1277,
    n1164,
    n1130
  );


  and
  g1289
  (
    n1289,
    n1087,
    n701
  );


  nand
  g1290
  (
    n1423,
    n962,
    n1196
  );


  nor
  g1291
  (
    n1448,
    n1084,
    n1152
  );


  nor
  g1292
  (
    n1346,
    n1139,
    n1115
  );


  nand
  g1293
  (
    n1359,
    n978,
    n955
  );


  xor
  g1294
  (
    n1256,
    n702,
    n728
  );


  xnor
  g1295
  (
    n1369,
    n1045,
    n1157
  );


  or
  g1296
  (
    n1496,
    n1121,
    n1133
  );


  nor
  g1297
  (
    KeyWire_0_50,
    n960,
    n1079
  );


  or
  g1298
  (
    n1356,
    n973,
    n725
  );


  xor
  g1299
  (
    n1417,
    n975,
    n1050
  );


  xor
  g1300
  (
    n1226,
    n1180,
    n1076
  );


  nand
  g1301
  (
    n1407,
    n1143,
    n1090
  );


  or
  g1302
  (
    n1394,
    n1091,
    n1189
  );


  xnor
  g1303
  (
    n1475,
    n957,
    n1190
  );


  nand
  g1304
  (
    n1376,
    n1199,
    n1064
  );


  and
  g1305
  (
    n1305,
    n1097,
    n959
  );


  xnor
  g1306
  (
    n1421,
    n1114,
    n1174
  );


  or
  g1307
  (
    n1498,
    n1189,
    n1150
  );


  or
  g1308
  (
    n1258,
    n1129,
    n781
  );


  or
  g1309
  (
    n1254,
    n1093,
    n1149
  );


  nor
  g1310
  (
    n1293,
    n1076,
    n1139
  );


  and
  g1311
  (
    n1409,
    n1154,
    n1044
  );


  xnor
  g1312
  (
    n1383,
    n1058,
    n1159
  );


  nor
  g1313
  (
    n1233,
    n1117,
    n1161
  );


  xnor
  g1314
  (
    n1480,
    n780,
    n1116
  );


  nor
  g1315
  (
    n1343,
    n1139,
    n557
  );


  nand
  g1316
  (
    n1500,
    n709,
    n1153
  );


  and
  g1317
  (
    n1427,
    n1070,
    n1042
  );


  xor
  g1318
  (
    n1312,
    n977,
    n1138
  );


  and
  g1319
  (
    n1398,
    n1105,
    n1162
  );


  and
  g1320
  (
    n1384,
    n778,
    n1146
  );


  nor
  g1321
  (
    n1424,
    n949,
    n1115
  );


  nor
  g1322
  (
    n1314,
    n1128,
    n977
  );


  xor
  g1323
  (
    n1481,
    n907,
    n1061
  );


  and
  g1324
  (
    n1487,
    n967,
    n726
  );


  xnor
  g1325
  (
    n1375,
    n1197,
    n1168
  );


  xnor
  g1326
  (
    n1249,
    n777,
    n1095
  );


  nor
  g1327
  (
    n1280,
    n1194,
    n1172
  );


  xnor
  g1328
  (
    n1237,
    n785,
    n1061
  );


  xnor
  g1329
  (
    n1276,
    n1110,
    n966
  );


  or
  g1330
  (
    n1473,
    n1125,
    n1080
  );


  xnor
  g1331
  (
    n1227,
    n1048,
    n1104
  );


  nand
  g1332
  (
    n1434,
    n717,
    n1043
  );


  or
  g1333
  (
    n1392,
    n1198,
    n557
  );


  or
  g1334
  (
    KeyWire_0_36,
    n1106,
    n1084
  );


  xor
  g1335
  (
    n1320,
    n1158,
    n946
  );


  or
  g1336
  (
    n1311,
    n959,
    n1085
  );


  or
  g1337
  (
    n1230,
    n1178,
    n1173
  );


  nand
  g1338
  (
    n1315,
    n1154,
    n946
  );


  nor
  g1339
  (
    n1304,
    n949,
    n991
  );


  xor
  g1340
  (
    n1415,
    n1145,
    n715
  );


  nor
  g1341
  (
    n1257,
    n1085,
    n787
  );


  nand
  g1342
  (
    n1400,
    n1146,
    n1142
  );


  and
  g1343
  (
    n1285,
    n1116,
    n974
  );


  xnor
  g1344
  (
    n1469,
    n974,
    n1101
  );


  or
  g1345
  (
    n1308,
    n951,
    n1117
  );


  nand
  g1346
  (
    n1506,
    n1176,
    n943
  );


  and
  g1347
  (
    n1458,
    n1069,
    n1116
  );


  xnor
  g1348
  (
    n1349,
    n955,
    n1166
  );


  or
  g1349
  (
    n1318,
    n1169,
    n1159
  );


  nand
  g1350
  (
    n1208,
    n1085,
    n1142
  );


  nor
  g1351
  (
    n1440,
    n1110,
    n1160,
    n958,
    n1073
  );


  and
  g1352
  (
    n1215,
    n970,
    n990,
    n1159,
    n1102
  );


  xor
  g1353
  (
    n1483,
    n982,
    n1153,
    n1113,
    n1074
  );


  nor
  g1354
  (
    n1344,
    n1105,
    n1125,
    n1062,
    n990
  );


  or
  g1355
  (
    n1242,
    n968,
    n1199,
    n1107,
    n1134
  );


  and
  g1356
  (
    n1521,
    n729,
    n967,
    n1136,
    n1194
  );


  nor
  g1357
  (
    n1524,
    n1187,
    n1118,
    n782,
    n1197
  );


  or
  g1358
  (
    n1340,
    n1066,
    n1148,
    n1112,
    n1141
  );


  or
  g1359
  (
    n1465,
    n1081,
    n1119,
    n786,
    n1157
  );


  and
  g1360
  (
    n1207,
    n1198,
    n1080,
    n971,
    n1149
  );


  xor
  g1361
  (
    KeyWire_0_43,
    n955,
    n1172,
    n1099,
    n784
  );


  nor
  g1362
  (
    n1492,
    n1063,
    n1156,
    n558,
    n1180
  );


  xor
  g1363
  (
    n1244,
    n1114,
    n964,
    n940,
    n1128
  );


  or
  g1364
  (
    n1414,
    n946,
    n1112,
    n1138,
    n948
  );


  nand
  g1365
  (
    n1405,
    n988,
    n984,
    n1142,
    n778
  );


  or
  g1366
  (
    n1235,
    n948,
    n724,
    n1152,
    n1122
  );


  xnor
  g1367
  (
    n1381,
    n1103,
    n1107,
    n1046,
    n783
  );


  nand
  g1368
  (
    n1401,
    n1141,
    n787,
    n940,
    n943
  );


  nand
  g1369
  (
    n1467,
    n1100,
    n1193,
    n1063,
    n1169
  );


  xnor
  g1370
  (
    n1513,
    n1048,
    n980,
    n1190,
    n1181
  );


  or
  g1371
  (
    n1328,
    n1086,
    n1163,
    n1192,
    n1190
  );


  xnor
  g1372
  (
    n1514,
    n1128,
    n960,
    n949,
    n1193
  );


  xnor
  g1373
  (
    n1420,
    n727,
    n1170,
    n1188,
    n1069
  );


  nand
  g1374
  (
    n1526,
    n777,
    n969,
    n981,
    n944
  );


  nand
  g1375
  (
    n1522,
    n1179,
    n1192,
    n1108,
    n953
  );


  xor
  g1376
  (
    n1220,
    n952,
    n1067,
    n1154,
    n1124
  );


  and
  g1377
  (
    n1288,
    n940,
    n785,
    n1084,
    n1193
  );


  nand
  g1378
  (
    n1238,
    n1133,
    n1149,
    n958,
    n1052
  );


  nand
  g1379
  (
    KeyWire_0_10,
    n1178,
    n1099,
    n977,
    n1121
  );


  xor
  g1380
  (
    n1240,
    n776,
    n1127,
    n1105,
    n1136
  );


  nor
  g1381
  (
    n1466,
    n714,
    n1084,
    n972,
    n1122
  );


  and
  g1382
  (
    n1527,
    n1195,
    n982,
    n1104,
    n1059
  );


  nor
  g1383
  (
    n1419,
    n1155,
    n1097,
    n976,
    n1106
  );


  xor
  g1384
  (
    n1426,
    n1048,
    n1096,
    n949,
    n1199
  );


  and
  g1385
  (
    n1260,
    n970,
    n947,
    n1057,
    n1160
  );


  and
  g1386
  (
    n1453,
    n1062,
    n1133,
    n1055,
    n721
  );


  xnor
  g1387
  (
    n1319,
    n1056,
    n1133,
    n947,
    n1172
  );


  and
  g1388
  (
    n1445,
    n1050,
    n1123,
    n776,
    n1144
  );


  xor
  g1389
  (
    n1266,
    n786,
    n1156,
    n1155,
    n944
  );


  and
  g1390
  (
    n1509,
    n1058,
    n987,
    n1172,
    n1200
  );


  or
  g1391
  (
    n1245,
    n985,
    n1065,
    n1157,
    n711
  );


  nand
  g1392
  (
    n1310,
    n1088,
    n1195,
    n1171,
    n991
  );


  xor
  g1393
  (
    n1223,
    n784,
    n972,
    n1061,
    n978
  );


  or
  g1394
  (
    n1259,
    n719,
    n558,
    n967,
    n1099
  );


  and
  g1395
  (
    n1361,
    n1188,
    n730,
    n960,
    n1168
  );


  nand
  g1396
  (
    n1265,
    n970,
    n1046,
    n1082,
    n1097
  );


  xnor
  g1397
  (
    n1367,
    n1089,
    n1140,
    n968,
    n1134
  );


  and
  g1398
  (
    n1388,
    n722,
    n783,
    n990,
    n1194
  );


  xnor
  g1399
  (
    n1263,
    n959,
    n1124,
    n968,
    n1138
  );


  nor
  g1400
  (
    n1206,
    n1166,
    n1042,
    n1055,
    n720
  );


  xnor
  g1401
  (
    n1341,
    n1093,
    n957,
    n1072,
    n976
  );


  or
  g1402
  (
    n1234,
    n986,
    n1073,
    n718,
    n1103
  );


  xor
  g1403
  (
    n1444,
    n1122,
    n981,
    n957,
    n1066
  );


  nor
  g1404
  (
    n1201,
    n1173,
    n696,
    n1068,
    n1120
  );


  xor
  g1405
  (
    n1329,
    n1049,
    n1075,
    n1199,
    n991
  );


  or
  g1406
  (
    n1391,
    n966,
    n1151,
    n1054,
    n941
  );


  or
  g1407
  (
    n1284,
    n1114,
    n1079,
    n1121,
    n1094
  );


  and
  g1408
  (
    n1327,
    n1196,
    n1186,
    n1071,
    n1083
  );


  xor
  g1409
  (
    n1345,
    n961,
    n718,
    n983,
    n1107
  );


  xnor
  g1410
  (
    n1519,
    n1067,
    n1189,
    n986,
    n984
  );


  xor
  g1411
  (
    n1436,
    n1051,
    n1068,
    n979,
    n1050
  );


  and
  g1412
  (
    n1399,
    n1145,
    n781,
    n1198,
    n1186
  );


  xor
  g1413
  (
    n1282,
    n1175,
    n1068,
    n962,
    n1078
  );


  and
  g1414
  (
    n1295,
    n965,
    n1174,
    n1191,
    n1055
  );


  or
  g1415
  (
    n1439,
    n1069,
    n964,
    n705,
    n1131
  );


  xnor
  g1416
  (
    n1316,
    n1166,
    n1047,
    n1113,
    n1135
  );


  and
  g1417
  (
    n1484,
    n1082,
    n1164,
    n781,
    n1174
  );


  xor
  g1418
  (
    n1412,
    n1191,
    n786,
    n1042,
    n1083
  );


  or
  g1419
  (
    n1325,
    n1148,
    n1151,
    n965,
    n948
  );


  or
  g1420
  (
    n1377,
    n1191,
    n1075,
    n1070,
    n569
  );


  xnor
  g1421
  (
    n1262,
    n1120,
    n1079,
    n1187,
    n1098
  );


  or
  g1422
  (
    n1309,
    n1127,
    n1108,
    n1164,
    n1065
  );


  and
  g1423
  (
    n1454,
    n966,
    n1187,
    n1152,
    n1131
  );


  and
  g1424
  (
    n1508,
    n729,
    n1058,
    n1149,
    n1049
  );


  or
  g1425
  (
    n1322,
    n979,
    n973,
    n1180,
    n1052
  );


  nand
  g1426
  (
    n1267,
    n1193,
    n1120,
    n1130,
    n1197
  );


  or
  g1427
  (
    n1355,
    n557,
    n1069,
    n1184
  );


  or
  g1428
  (
    n1459,
    n1119,
    n1117,
    n1178,
    n1051
  );


  or
  g1429
  (
    n1441,
    n1102,
    n974,
    n778,
    n971
  );


  xor
  g1430
  (
    n1370,
    n1137,
    n1125,
    n950,
    n1183
  );


  nor
  g1431
  (
    n1247,
    n1177,
    n723,
    n988,
    n698
  );


  nor
  g1432
  (
    n1471,
    n1074,
    n1154,
    n700,
    n947
  );


  xnor
  g1433
  (
    n1443,
    n970,
    n950,
    n1116,
    n1179
  );


  or
  g1434
  (
    n1413,
    n980,
    n783,
    n1160
  );


  nand
  g1435
  (
    n1482,
    n1045,
    n1163,
    n1101
  );


  and
  g1436
  (
    n1347,
    n945,
    n1100,
    n1113,
    n1143
  );


  nand
  g1437
  (
    n1297,
    n1066,
    n1111,
    n1062,
    n963
  );


  or
  g1438
  (
    n1451,
    n1074,
    n1047,
    n710,
    n1119
  );


  nand
  g1439
  (
    n1504,
    n697,
    n706,
    n944,
    n1140
  );


  and
  g1440
  (
    n1337,
    n1185,
    n1086,
    n1071,
    n959
  );


  and
  g1441
  (
    n1462,
    n1168,
    n1076,
    n1128,
    n1137
  );


  and
  g1442
  (
    KeyWire_0_40,
    n1053,
    n1183,
    n1182,
    n1100
  );


  nand
  g1443
  (
    n1336,
    n1044,
    n988,
    n1126,
    n1043
  );


  and
  g1444
  (
    n1231,
    n1120,
    n1060,
    n1150,
    n1155
  );


  or
  g1445
  (
    n1502,
    n716,
    n1132,
    n1112,
    n778
  );


  or
  g1446
  (
    n1450,
    n726,
    n1141,
    n1123,
    n1167
  );


  or
  g1447
  (
    n1225,
    n942,
    n1075,
    n1104,
    n1095
  );


  xnor
  g1448
  (
    n1373,
    n978,
    n703,
    n982,
    n1090
  );


  nor
  g1449
  (
    n1416,
    n782,
    n968,
    n1062,
    n727
  );


  nand
  g1450
  (
    n1433,
    n1105,
    n1078,
    n980,
    n975
  );


  nand
  g1451
  (
    n1261,
    n1156,
    n1060,
    n725,
    n728
  );


  xnor
  g1452
  (
    n1203,
    n1077,
    n1086,
    n1091,
    n781
  );


  nand
  g1453
  (
    n1418,
    n785,
    n1167,
    n991,
    n1126
  );


  xnor
  g1454
  (
    n1255,
    n984,
    n1109,
    n952,
    n787
  );


  xor
  g1455
  (
    n1358,
    n1177,
    n961,
    n777,
    n953
  );


  and
  g1456
  (
    n1411,
    n1063,
    n1042,
    n951,
    n1195
  );


  xnor
  g1457
  (
    n1494,
    n1064,
    n1112,
    n1200,
    n1059
  );


  nor
  g1458
  (
    n1292,
    n1184,
    n1070,
    n722,
    n1078
  );


  xnor
  g1459
  (
    n1432,
    n1147,
    n963,
    n1044,
    n558
  );


  nand
  g1460
  (
    n1354,
    n1182,
    n1080,
    n1043,
    n1065
  );


  nand
  g1461
  (
    n1404,
    n952,
    n1110,
    n1092,
    n1171
  );


  or
  g1462
  (
    n1330,
    n1083,
    n786,
    n945,
    n1123
  );


  xnor
  g1463
  (
    n1269,
    n1167,
    n1054,
    n951,
    n1139
  );


  or
  g1464
  (
    n1470,
    n1056,
    n1130,
    n1118,
    n961
  );


  and
  g1465
  (
    n1204,
    n1155,
    n1186,
    n1078,
    n942
  );


  or
  g1466
  (
    n1317,
    n699,
    n1090,
    n1170,
    n1179
  );


  xnor
  g1467
  (
    n1393,
    n1161,
    n957,
    n695,
    n1135
  );


  xor
  g1468
  (
    n1485,
    n1148,
    n974,
    n1151,
    n1071
  );


  xnor
  g1469
  (
    n1253,
    n971,
    n989,
    n1109,
    n1071
  );


  nand
  g1470
  (
    n1490,
    n973,
    n942,
    n1091,
    n1169
  );


  nand
  g1471
  (
    n1251,
    n1129,
    n1114,
    n1094,
    n1171
  );


  xnor
  g1472
  (
    n1428,
    n980,
    n1138,
    n953,
    n1173
  );


  and
  g1473
  (
    n1379,
    n1188,
    n952,
    n964,
    n1083
  );


  xnor
  g1474
  (
    n1232,
    n1124,
    n1098,
    n1050,
    n1182
  );


  xor
  g1475
  (
    n1352,
    n784,
    n1045,
    n975,
    n1123
  );


  and
  g1476
  (
    n1210,
    n1158,
    n1121,
    n780,
    n976
  );


  nand
  g1477
  (
    n1493,
    n1196,
    n1122,
    n1087,
    n1147
  );


  and
  g1478
  (
    n1366,
    n1115,
    n1119,
    n776,
    n1094
  );


  nand
  g1479
  (
    n1302,
    n1168,
    n1150,
    n1100,
    n1134
  );


  nand
  g1480
  (
    n1403,
    n1127,
    n1093,
    n1106,
    n950
  );


  nand
  g1481
  (
    n1455,
    n1153,
    n1185,
    n1047,
    n987
  );


  nand
  g1482
  (
    n1363,
    n1046,
    n1200,
    n1136,
    n987
  );


  or
  g1483
  (
    n1517,
    n1131,
    n1136,
    n1048,
    n950
  );


  nand
  g1484
  (
    KeyWire_0_63,
    n1065,
    n958,
    n1086,
    n719
  );


  nand
  g1485
  (
    n1395,
    n1187,
    n1051,
    n1094,
    n783
  );


  nand
  g1486
  (
    n1313,
    n1148,
    n983,
    n963,
    n989
  );


  and
  g1487
  (
    n1294,
    n1067,
    n1192,
    n1173,
    n969
  );


  and
  g1488
  (
    n1516,
    n1162,
    n1106,
    n985,
    n1147
  );


  nand
  g1489
  (
    n1371,
    n1190,
    n1068,
    n1089,
    n1052
  );


  and
  g1490
  (
    n1501,
    n1074,
    n1176,
    n779,
    n1198
  );


  or
  g1491
  (
    n1222,
    n1177,
    n1186,
    n713,
    n1096
  );


  and
  g1492
  (
    n1252,
    n1156,
    n987,
    n1192,
    n779
  );


  nand
  g1493
  (
    n1351,
    n1098,
    n963,
    n1064,
    n953
  );


  nand
  g1494
  (
    n1219,
    n972,
    n1189,
    n1049,
    n943
  );


  and
  g1495
  (
    n1241,
    n961,
    n986,
    n1064,
    n1096
  );


  and
  g1496
  (
    KeyWire_0_11,
    n1053,
    n1102,
    n979,
    n730
  );


  xnor
  g1497
  (
    n1287,
    n1103,
    n990,
    n985,
    n1082
  );


  xnor
  g1498
  (
    n1510,
    n782,
    n971,
    n1181,
    n785
  );


  xnor
  g1499
  (
    n1479,
    n973,
    n972,
    n941,
    n1077
  );


  and
  g1500
  (
    n1283,
    n1131,
    n958,
    n1153,
    n1140
  );


  xnor
  g1501
  (
    n1646,
    n1356,
    n1455,
    n1266,
    n1465
  );


  xnor
  g1502
  (
    n1622,
    n1220,
    n1402,
    n1217,
    n1307
  );


  xor
  g1503
  (
    n1587,
    n1327,
    n1455,
    n1374,
    n1387
  );


  and
  g1504
  (
    n1599,
    n1302,
    n1272,
    n1392,
    n1259
  );


  nand
  g1505
  (
    n1565,
    n1210,
    n1440,
    n1246,
    n1415
  );


  xor
  g1506
  (
    n1769,
    n1334,
    n1307,
    n1363,
    n1262
  );


  xnor
  g1507
  (
    n1585,
    n1451,
    n1305,
    n1315,
    n1340
  );


  nor
  g1508
  (
    n1594,
    n1314,
    n1347,
    n1386,
    n1326
  );


  xnor
  g1509
  (
    n1637,
    n1274,
    n1278,
    n1432,
    n1456
  );


  or
  g1510
  (
    n1579,
    n1319,
    n1459,
    n1256,
    n1477
  );


  xnor
  g1511
  (
    n1702,
    n1378,
    n1264,
    n1207,
    n1423
  );


  xnor
  g1512
  (
    n1548,
    n1271,
    n1287,
    n1386,
    n1347
  );


  nor
  g1513
  (
    n1606,
    n1321,
    n1299,
    n1277,
    n1393
  );


  and
  g1514
  (
    n1649,
    n1216,
    n1375,
    n1287,
    n1476
  );


  nor
  g1515
  (
    n1669,
    n1439,
    n1273,
    n1254,
    n1420
  );


  nor
  g1516
  (
    n1614,
    n1390,
    n1445,
    n1330,
    n1426
  );


  nor
  g1517
  (
    n1597,
    n1341,
    n1234,
    n1212,
    n1313
  );


  nor
  g1518
  (
    n1608,
    n1446,
    n1295,
    n1238,
    n1210
  );


  and
  g1519
  (
    n1712,
    n1275,
    n1334,
    n1265,
    n1431
  );


  nor
  g1520
  (
    n1791,
    n1297,
    n1218,
    n1379,
    n1222
  );


  and
  g1521
  (
    n1535,
    n1288,
    n1368,
    n1409,
    n1327
  );


  xor
  g1522
  (
    n1638,
    n1448,
    n1447,
    n1445,
    n1204
  );


  or
  g1523
  (
    n1567,
    n1411,
    n1288,
    n1469,
    n1427
  );


  xnor
  g1524
  (
    n1659,
    n1237,
    n1234,
    n1447,
    n1350
  );


  nor
  g1525
  (
    n1656,
    n1479,
    n1419,
    n1407,
    n1317
  );


  nor
  g1526
  (
    n1549,
    n1374,
    n1436,
    n1257,
    n1254
  );


  nand
  g1527
  (
    n1759,
    n1400,
    n1418,
    n1279,
    n1201
  );


  nand
  g1528
  (
    n1803,
    n1229,
    n1350,
    n1392,
    n1473
  );


  xor
  g1529
  (
    n1551,
    n1283,
    n1260,
    n1352,
    n1293
  );


  xnor
  g1530
  (
    n1741,
    n1403,
    n1435,
    n1314,
    n1212
  );


  xor
  g1531
  (
    KeyWire_0_25,
    n1258,
    n1429,
    n1219,
    n1406
  );


  nand
  g1532
  (
    n1568,
    n1448,
    n1222,
    n1249,
    n1418
  );


  nor
  g1533
  (
    n1623,
    n1373,
    n1281,
    n1456,
    n1377
  );


  xor
  g1534
  (
    n1732,
    n1286,
    n1397,
    n1301,
    n1292
  );


  and
  g1535
  (
    n1711,
    n1287,
    n1372,
    n1201,
    n1401
  );


  xor
  g1536
  (
    n1770,
    n1463,
    n1255,
    n1252,
    n1375
  );


  nor
  g1537
  (
    n1738,
    n1296,
    n1460,
    n1432,
    n1414
  );


  or
  g1538
  (
    n1717,
    n1390,
    n1310,
    n1366,
    n1244
  );


  nor
  g1539
  (
    n1678,
    n1376,
    n1393,
    n1348,
    n1429
  );


  xnor
  g1540
  (
    n1716,
    n1427,
    n1335,
    n1325,
    n1213
  );


  nand
  g1541
  (
    n1633,
    n1205,
    n1333,
    n1384,
    n1434
  );


  and
  g1542
  (
    n1616,
    n1397,
    n1353,
    n1297,
    n1315
  );


  or
  g1543
  (
    n1763,
    n1413,
    n1421,
    n1239,
    n1312
  );


  nand
  g1544
  (
    n1677,
    n1387,
    n1362,
    n1453,
    n1420
  );


  xnor
  g1545
  (
    n1675,
    n1431,
    n1356,
    n1223,
    n1403
  );


  xnor
  g1546
  (
    n1650,
    n1324,
    n1358,
    n1478,
    n1342
  );


  and
  g1547
  (
    n1529,
    n1469,
    n1214,
    n1333,
    n1261
  );


  xor
  g1548
  (
    n1593,
    n1291,
    n1464,
    n1320,
    n1419
  );


  or
  g1549
  (
    n1636,
    n1328,
    n1430,
    n1330,
    n1362
  );


  and
  g1550
  (
    n1706,
    n1452,
    n1435,
    n1224,
    n1407
  );


  xnor
  g1551
  (
    n1583,
    n1361,
    n1444,
    n1362,
    n1395
  );


  nor
  g1552
  (
    n1612,
    n1372,
    n1229,
    n1391,
    n1346
  );


  xor
  g1553
  (
    n1784,
    n1236,
    n1284,
    n1354,
    n1276
  );


  or
  g1554
  (
    n1542,
    n1282,
    n1281,
    n1404,
    n1411
  );


  or
  g1555
  (
    n1540,
    n1458,
    n1450,
    n1221,
    n1392
  );


  nor
  g1556
  (
    n1619,
    n1290,
    n1410,
    n1223,
    n1325
  );


  or
  g1557
  (
    n1600,
    n1238,
    n1376,
    n1421,
    n1396
  );


  nand
  g1558
  (
    n1737,
    n1351,
    n1366,
    n1232,
    n1469
  );


  xor
  g1559
  (
    n1557,
    n1361,
    n1364,
    n1345,
    n1329
  );


  and
  g1560
  (
    n1584,
    n1324,
    n1260,
    n1284,
    n1446
  );


  nor
  g1561
  (
    n1642,
    n1301,
    n1230,
    n1332,
    n1323
  );


  xor
  g1562
  (
    n1682,
    n1415,
    n1295,
    n1206,
    n1331
  );


  nor
  g1563
  (
    n1624,
    n1340,
    n1212,
    n1337,
    n1425
  );


  nand
  g1564
  (
    n1546,
    n1240,
    n1343,
    n1394,
    n1438
  );


  or
  g1565
  (
    n1797,
    n1320,
    n1329,
    n1442,
    n1275
  );


  xnor
  g1566
  (
    n1699,
    n1363,
    n1306,
    n1384,
    n1221
  );


  or
  g1567
  (
    n1734,
    n1278,
    n1371,
    n1388,
    n1418
  );


  xnor
  g1568
  (
    n1545,
    n1217,
    n1345,
    n1474,
    n1415
  );


  or
  g1569
  (
    n1625,
    n1406,
    n1299,
    n1476,
    n1251
  );


  or
  g1570
  (
    n1730,
    n1338,
    n1433,
    n1329,
    n1233
  );


  or
  g1571
  (
    n1644,
    n1441,
    n1253,
    n1317,
    n1405
  );


  xor
  g1572
  (
    n1604,
    n1363,
    n1302,
    n1266,
    n1264
  );


  xnor
  g1573
  (
    n1787,
    n1227,
    n1249,
    n1430,
    n1254
  );


  nor
  g1574
  (
    n1762,
    n1390,
    n1389,
    n1357,
    n1319
  );


  xor
  g1575
  (
    n1708,
    n1245,
    n1427,
    n1224,
    n1358
  );


  nor
  g1576
  (
    n1532,
    n1344,
    n1332,
    n1253,
    n1243
  );


  xnor
  g1577
  (
    n1657,
    n1416,
    n1256,
    n1242,
    n1316
  );


  nor
  g1578
  (
    n1686,
    n1404,
    n1214,
    n1215,
    n1378
  );


  xor
  g1579
  (
    n1660,
    n1410,
    n1369,
    n1349,
    n1477
  );


  or
  g1580
  (
    n1561,
    n1208,
    n1237,
    n1419,
    n1340
  );


  and
  g1581
  (
    n1704,
    n1479,
    n1437,
    n1208,
    n1369
  );


  nor
  g1582
  (
    n1740,
    n1348,
    n1341,
    n1432,
    n1255
  );


  and
  g1583
  (
    n1689,
    n1347,
    n1218,
    n1457,
    n1473
  );


  and
  g1584
  (
    n1774,
    n1460,
    n1465,
    n1259,
    n1298
  );


  nand
  g1585
  (
    n1707,
    n1380,
    n1453,
    n1389,
    n1296
  );


  nand
  g1586
  (
    n1785,
    n1248,
    n1250,
    n1236,
    n1457
  );


  xor
  g1587
  (
    n1658,
    n1442,
    n1400,
    n1316,
    n1339
  );


  xor
  g1588
  (
    n1592,
    n1294,
    n1285,
    n1291,
    n1448
  );


  nand
  g1589
  (
    n1778,
    n1397,
    n1323,
    n1399,
    n1328
  );


  nor
  g1590
  (
    KeyWire_0_14,
    n1325,
    n1251,
    n1274,
    n1423
  );


  and
  g1591
  (
    n1747,
    n1454,
    n1453,
    n116,
    n1401
  );


  and
  g1592
  (
    n1793,
    n1452,
    n1334,
    n1267,
    n1467
  );


  or
  g1593
  (
    n1692,
    n1213,
    n1315,
    n1302,
    n1257
  );


  nand
  g1594
  (
    n1701,
    n1356,
    n1370,
    n1437,
    n1470
  );


  xor
  g1595
  (
    n1742,
    n1339,
    n1206,
    n1458
  );


  xor
  g1596
  (
    n1647,
    n1416,
    n1303,
    n1333,
    n1267
  );


  or
  g1597
  (
    n1581,
    n1342,
    n1226,
    n1253,
    n1365
  );


  xor
  g1598
  (
    n1615,
    n1252,
    n1414,
    n1229,
    n1240
  );


  or
  g1599
  (
    n1773,
    n1338,
    n1209,
    n1457,
    n1288
  );


  or
  g1600
  (
    n1795,
    n1311,
    n1383,
    n1309,
    n1305
  );


  and
  g1601
  (
    n1630,
    n1397,
    n1277,
    n1450,
    n1259
  );


  and
  g1602
  (
    n1569,
    n1311,
    n1365,
    n1341,
    n1416
  );


  or
  g1603
  (
    n1552,
    n1361,
    n1422,
    n1476,
    n1424
  );


  nand
  g1604
  (
    n1672,
    n1351,
    n1331,
    n1308,
    n1309
  );


  xnor
  g1605
  (
    n1687,
    n1321,
    n1235,
    n1311,
    n1471
  );


  nand
  g1606
  (
    n1556,
    n1352,
    n1460,
    n1438,
    n1286
  );


  xor
  g1607
  (
    n1541,
    n1408,
    n1446,
    n1438,
    n1261
  );


  and
  g1608
  (
    n1543,
    n1230,
    n1443,
    n1273,
    n1308
  );


  or
  g1609
  (
    n1671,
    n1424,
    n1370,
    n1381,
    n1407
  );


  nand
  g1610
  (
    n1536,
    n1300,
    n1417,
    n1350,
    n1426
  );


  xnor
  g1611
  (
    n1804,
    n1312,
    n1236,
    n1348,
    n1325
  );


  and
  g1612
  (
    n1643,
    n1204,
    n1441,
    n1235,
    n1276
  );


  and
  g1613
  (
    n1794,
    n1217,
    n1346,
    n1350,
    n1211
  );


  xnor
  g1614
  (
    n1586,
    n1336,
    n1386,
    n1406,
    n1480
  );


  nand
  g1615
  (
    n1605,
    n1354,
    n1233,
    n1368,
    n1237
  );


  nand
  g1616
  (
    n1553,
    n1203,
    n1354,
    n1232,
    n1410
  );


  xor
  g1617
  (
    n1697,
    n1372,
    n1300,
    n1223,
    n1462
  );


  nand
  g1618
  (
    KeyWire_0_32,
    n1408,
    n1412,
    n1472,
    n1364
  );


  nand
  g1619
  (
    n1598,
    n1209,
    n1281,
    n1241,
    n1401
  );


  xor
  g1620
  (
    n1753,
    n1411,
    n1357,
    n1210,
    n1380
  );


  nor
  g1621
  (
    n1634,
    n1339,
    n1319,
    n1270,
    n1308
  );


  xnor
  g1622
  (
    n1801,
    n1225,
    n1461,
    n1405,
    n1240
  );


  and
  g1623
  (
    n1746,
    n1207,
    n1422,
    n1437,
    n1452
  );


  or
  g1624
  (
    n1698,
    n1222,
    n1298,
    n1220,
    n1320
  );


  and
  g1625
  (
    n1772,
    n1215,
    n1435,
    n1260,
    n1399
  );


  xnor
  g1626
  (
    n1531,
    n1412,
    n1218,
    n1364,
    n1396
  );


  or
  g1627
  (
    n1544,
    n1478,
    n1363,
    n1431,
    n1216
  );


  and
  g1628
  (
    n1566,
    n1429,
    n1304,
    n1289,
    n1265
  );


  xor
  g1629
  (
    n1739,
    n1222,
    n1344,
    n1349,
    n1439
  );


  and
  g1630
  (
    n1806,
    n1270,
    n1310,
    n1466,
    n1352
  );


  or
  g1631
  (
    n1653,
    n1318,
    n1239,
    n1474,
    n1205
  );


  or
  g1632
  (
    n1798,
    n1428,
    n1293,
    n1464,
    n1251
  );


  and
  g1633
  (
    n1700,
    n1284,
    n1326,
    n1274,
    n1214
  );


  nand
  g1634
  (
    n1691,
    n1421,
    n1354,
    n1274,
    n1391
  );


  nand
  g1635
  (
    n1617,
    n1331,
    n1290,
    n1336,
    n1309
  );


  nor
  g1636
  (
    n1722,
    n1459,
    n1399,
    n1297,
    n1208
  );


  xor
  g1637
  (
    n1758,
    n1279,
    n1208,
    n1270,
    n1336
  );


  xor
  g1638
  (
    n1618,
    n1473,
    n1242,
    n1403,
    n1229
  );


  nor
  g1639
  (
    n1752,
    n1262,
    n1353,
    n1245,
    n1449
  );


  and
  g1640
  (
    n1628,
    n1314,
    n1384,
    n1398,
    n1327
  );


  or
  g1641
  (
    n1670,
    n1252,
    n1394,
    n1265,
    n1283
  );


  nand
  g1642
  (
    n1539,
    n1472,
    n1441,
    n1440,
    n1334
  );


  nor
  g1643
  (
    n1729,
    n1278,
    n1477,
    n1302,
    n1247
  );


  nand
  g1644
  (
    n1673,
    n1285,
    n1210,
    n1295,
    n1417
  );


  nor
  g1645
  (
    n1663,
    n1346,
    n1362,
    n1455,
    n1328
  );


  xor
  g1646
  (
    n1648,
    n1358,
    n1398,
    n1297,
    n1299
  );


  xnor
  g1647
  (
    n1765,
    n1322,
    n1241,
    n1306,
    n1353
  );


  or
  g1648
  (
    n1595,
    n1373,
    n1272,
    n1349,
    n1443
  );


  or
  g1649
  (
    n1627,
    n1445,
    n1291,
    n1261,
    n1205
  );


  and
  g1650
  (
    n1693,
    n1353,
    n1331,
    n1220,
    n1318
  );


  or
  g1651
  (
    n1574,
    n1468,
    n1371,
    n1269,
    n1227
  );


  and
  g1652
  (
    n1610,
    n1313,
    n1430,
    n1323,
    n1466
  );


  or
  g1653
  (
    n1547,
    n1426,
    n1212,
    n1359,
    n1219
  );


  xor
  g1654
  (
    n1635,
    n1226,
    n1271,
    n1368,
    n1417
  );


  nand
  g1655
  (
    n1555,
    n1234,
    n1405,
    n1243,
    n1382
  );


  or
  g1656
  (
    n1766,
    n1206,
    n1244,
    n1235,
    n1406
  );


  xor
  g1657
  (
    n1575,
    n1378,
    n1423,
    n1449,
    n1462
  );


  nand
  g1658
  (
    n1767,
    n1273,
    n1396,
    n1361,
    n1268
  );


  xnor
  g1659
  (
    n1710,
    n1249,
    n1338,
    n1336,
    n1220
  );


  nor
  g1660
  (
    n1668,
    n1370,
    n1204,
    n1301,
    n1247
  );


  nand
  g1661
  (
    n1777,
    n1228,
    n1303,
    n1340,
    n1464
  );


  or
  g1662
  (
    n1718,
    n1463,
    n1207,
    n1223,
    n1314
  );


  or
  g1663
  (
    n1775,
    n1330,
    n1217,
    n1407,
    n1460
  );


  xnor
  g1664
  (
    n1602,
    n1254,
    n1423,
    n1458,
    n1475
  );


  or
  g1665
  (
    n1723,
    n1424,
    n1468,
    n1322,
    n1352
  );


  and
  g1666
  (
    n1530,
    n1379,
    n1367,
    n1474,
    n1281
  );


  or
  g1667
  (
    n1538,
    n1335,
    n1365,
    n1429,
    n1395
  );


  and
  g1668
  (
    n1573,
    n1280,
    n1242,
    n1464,
    n1401
  );


  and
  g1669
  (
    n1577,
    n1342,
    n1365,
    n1475,
    n1293
  );


  xnor
  g1670
  (
    n1727,
    n1382,
    n1385,
    n1360,
    n1287
  );


  xnor
  g1671
  (
    n1667,
    n1271,
    n1323,
    n1256,
    n1273
  );


  xnor
  g1672
  (
    n1684,
    n1310,
    n1313,
    n1421,
    n1275
  );


  nor
  g1673
  (
    n1776,
    n1224,
    n1467,
    n1291,
    n1389
  );


  xnor
  g1674
  (
    n1786,
    n1277,
    n1231,
    n1266,
    n1230
  );


  nand
  g1675
  (
    n1613,
    n1244,
    n1303,
    n1300,
    n1398
  );


  or
  g1676
  (
    n1744,
    n1470,
    n1425,
    n1472,
    n1437
  );


  nand
  g1677
  (
    n1750,
    n1256,
    n1225,
    n1355,
    n1440
  );


  nand
  g1678
  (
    n1632,
    n1304,
    n1463,
    n1269,
    n1471
  );


  or
  g1679
  (
    n1728,
    n1321,
    n1289,
    n1468,
    n1282
  );


  and
  g1680
  (
    n1664,
    n1444,
    n1298,
    n1459,
    n1386
  );


  and
  g1681
  (
    n1764,
    n1387,
    n1230,
    n1371,
    n1218
  );


  and
  g1682
  (
    n1683,
    n1213,
    n1358,
    n1245,
    n1459
  );


  nor
  g1683
  (
    n1676,
    n1461,
    n1415,
    n1206,
    n1250
  );


  and
  g1684
  (
    n1783,
    n1260,
    n1319,
    n1266,
    n1360
  );


  xnor
  g1685
  (
    n1799,
    n1349,
    n1215,
    n1290,
    n1322
  );


  and
  g1686
  (
    n1715,
    n1388,
    n1367,
    n1231,
    n1405
  );


  xor
  g1687
  (
    n1564,
    n1313,
    n1318,
    n1442,
    n1360
  );


  nand
  g1688
  (
    n1796,
    n117,
    n1369,
    n1408,
    n1255
  );


  xnor
  g1689
  (
    n1679,
    n1240,
    n1454,
    n1451,
    n1211
  );


  xnor
  g1690
  (
    n1780,
    n1346,
    n1409,
    n1427,
    n1337
  );


  xor
  g1691
  (
    n1537,
    n1299,
    n1213,
    n1245,
    n1269
  );


  xnor
  g1692
  (
    n1768,
    n1463,
    n1466,
    n1227,
    n1422
  );


  nor
  g1693
  (
    n1749,
    n1376,
    n1383,
    n1377,
    n1351
  );


  xnor
  g1694
  (
    n1681,
    n1440,
    n1271,
    n1435,
    n1219
  );


  nor
  g1695
  (
    n1570,
    n1461,
    n1451,
    n1379,
    n1376
  );


  xnor
  g1696
  (
    n1588,
    n1434,
    n1399,
    n1479,
    n1216
  );


  xor
  g1697
  (
    n1641,
    n1292,
    n1202,
    n1284,
    n1373
  );


  xnor
  g1698
  (
    n1736,
    n1478,
    n1374,
    n1395,
    n1338
  );


  xnor
  g1699
  (
    n1607,
    n1439,
    n1417,
    n1393,
    n1391
  );


  xnor
  g1700
  (
    n1731,
    n1296,
    n1337,
    n1324,
    n1436
  );


  and
  g1701
  (
    n1603,
    n1263,
    n1250,
    n1380,
    n1419
  );


  or
  g1702
  (
    n1609,
    n1400,
    n1288,
    n1413,
    n1219
  );


  and
  g1703
  (
    n1709,
    n1359,
    n1316,
    n1265,
    n1317
  );


  nor
  g1704
  (
    n1748,
    n1367,
    n1428,
    n1447,
    n1303
  );


  or
  g1705
  (
    n1688,
    n1442,
    n1241,
    n1418,
    n1471
  );


  and
  g1706
  (
    n1654,
    n1431,
    n1300,
    n1263,
    n1375
  );


  nor
  g1707
  (
    n1788,
    n1307,
    n1278,
    n1412,
    n1456
  );


  nor
  g1708
  (
    n1620,
    n1369,
    n1473,
    n1263,
    n1388
  );


  xnor
  g1709
  (
    n1719,
    n1304,
    n1207,
    n1301,
    n1286
  );


  nor
  g1710
  (
    n1721,
    n1296,
    n1374,
    n1247,
    n1357
  );


  xor
  g1711
  (
    n1589,
    n1293,
    n1355,
    n1320,
    n1311
  );


  and
  g1712
  (
    n1757,
    n1448,
    n1309,
    n1379,
    n1246
  );


  xnor
  g1713
  (
    n1534,
    n1324,
    n1333,
    n1378,
    n1298
  );


  or
  g1714
  (
    n1560,
    n1403,
    n1347,
    n1211,
    n1202
  );


  nand
  g1715
  (
    n1703,
    n1285,
    n1392,
    n1409,
    n1382
  );


  nand
  g1716
  (
    n1725,
    n1269,
    n1275,
    n1414,
    n1202
  );


  nor
  g1717
  (
    n1743,
    n1450,
    n1235,
    n1304,
    n1259
  );


  xnor
  g1718
  (
    n1571,
    n1462,
    n1247,
    n1394,
    n1250
  );


  nor
  g1719
  (
    n1800,
    n1471,
    n1380,
    n1225,
    n1326
  );


  and
  g1720
  (
    n1572,
    n1381,
    n1444,
    n1251,
    n1326
  );


  or
  g1721
  (
    n1533,
    n1420,
    n1439,
    n1355,
    n1328
  );


  nand
  g1722
  (
    n1666,
    n1465,
    n1430,
    n1345,
    n1317
  );


  nand
  g1723
  (
    n1626,
    n1383,
    n1337,
    n1402,
    n1410
  );


  and
  g1724
  (
    n1559,
    n1316,
    n1232,
    n1404,
    n1305
  );


  xnor
  g1725
  (
    n1661,
    n1472,
    n1211,
    n1228,
    n1226
  );


  or
  g1726
  (
    n1754,
    n1467,
    n1264,
    n1267,
    n1312
  );


  xnor
  g1727
  (
    n1629,
    n1225,
    n1276,
    n1424,
    n1307
  );


  xnor
  g1728
  (
    n1578,
    n1310,
    n1400,
    n1454,
    n1453
  );


  nor
  g1729
  (
    n1802,
    n1359,
    n1402,
    n1390,
    n1449
  );


  xor
  g1730
  (
    n1601,
    n1443,
    n1209,
    n1248,
    n1268
  );


  nor
  g1731
  (
    n1726,
    n1446,
    n1329,
    n1201,
    n1282
  );


  nand
  g1732
  (
    n1696,
    n1332,
    n1209,
    n1467,
    n1425
  );


  and
  g1733
  (
    n1655,
    n1294,
    n1457,
    n1465,
    n1356
  );


  nor
  g1734
  (
    n1713,
    n1332,
    n1243,
    n1366,
    n1234
  );


  or
  g1735
  (
    n1745,
    n1475,
    n1258,
    n1428,
    n1375
  );


  nor
  g1736
  (
    n1596,
    n1395,
    n1294,
    n1432,
    n1470
  );


  and
  g1737
  (
    n1805,
    n1382,
    n1231,
    n116,
    n1345
  );


  or
  g1738
  (
    n1685,
    n1377,
    n1461,
    n1404,
    n1456
  );


  nand
  g1739
  (
    n1735,
    n1285,
    n1221,
    n1263,
    n1335
  );


  xnor
  g1740
  (
    n1720,
    n1306,
    n1444,
    n1227,
    n1295
  );


  nand
  g1741
  (
    n1590,
    n1280,
    n1364,
    n1294,
    n1343
  );


  or
  g1742
  (
    n1563,
    n1339,
    n1436,
    n1322,
    n1469
  );


  nand
  g1743
  (
    n1705,
    n1394,
    n1359,
    n1203,
    n1455
  );


  or
  g1744
  (
    n1782,
    n1289,
    n1253,
    n1221,
    n1388
  );


  nand
  g1745
  (
    n1645,
    n1216,
    n1443,
    n1477,
    n1434
  );


  nand
  g1746
  (
    n1662,
    n1224,
    n1387,
    n1228,
    n1283
  );


  nand
  g1747
  (
    n1771,
    n1383,
    n1226,
    n1434,
    n1438
  );


  nand
  g1748
  (
    n1751,
    n1262,
    n1282,
    n1468,
    n1279
  );


  nand
  g1749
  (
    n1651,
    n1412,
    n1478,
    n1357,
    n1355
  );


  xnor
  g1750
  (
    n1554,
    n1454,
    n1408,
    n1367,
    n1277
  );


  nor
  g1751
  (
    n1733,
    n1258,
    n1241,
    n1343,
    n1228
  );


  or
  g1752
  (
    n1724,
    n1445,
    n1385,
    n1272,
    n1233
  );


  xnor
  g1753
  (
    n1558,
    n1261,
    n1239,
    n1381,
    n1452
  );


  xnor
  g1754
  (
    n1591,
    n1286,
    n1420,
    n1433,
    n1268
  );


  or
  g1755
  (
    n1789,
    n1279,
    n1413,
    n1414,
    n1348
  );


  or
  g1756
  (
    n1761,
    n1385,
    n1416,
    n1396,
    n1292
  );


  nand
  g1757
  (
    n1562,
    n1476,
    n1318,
    n1344,
    n1272
  );


  nor
  g1758
  (
    n1611,
    n1371,
    n1258,
    n1262,
    n1398
  );


  or
  g1759
  (
    n1781,
    n1474,
    n1232,
    n1268,
    n1248
  );


  xnor
  g1760
  (
    n1779,
    n1451,
    n1385,
    n1292,
    n1373
  );


  xor
  g1761
  (
    n1714,
    n116,
    n1249,
    n1283,
    n1252
  );


  xor
  g1762
  (
    n1690,
    n1255,
    n1436,
    n1246,
    n1344
  );


  xnor
  g1763
  (
    n1760,
    n1306,
    n1242,
    n1370,
    n1422
  );


  and
  g1764
  (
    n1580,
    n1341,
    n1391,
    n1360,
    n1246
  );


  nand
  g1765
  (
    n1756,
    n1203,
    n1267,
    n1450,
    n1393
  );


  xnor
  g1766
  (
    n1680,
    n1308,
    n1290,
    n1384,
    n1215
  );


  and
  g1767
  (
    n1652,
    n1343,
    n1368,
    n1270,
    n1449
  );


  and
  g1768
  (
    n1695,
    n1327,
    n1470,
    n1413,
    n1238
  );


  and
  g1769
  (
    n1674,
    n1280,
    n1409,
    n1433,
    n1305
  );


  xor
  g1770
  (
    n1528,
    n1233,
    n1428,
    n1426,
    n1425
  );


  nor
  g1771
  (
    n1790,
    n1238,
    n1257,
    n1321
  );


  nor
  g1772
  (
    n1665,
    n1248,
    n1315,
    n1447,
    n1433
  );


  nand
  g1773
  (
    n1621,
    n1411,
    n1289,
    n1479,
    n1231
  );


  nor
  g1774
  (
    n1640,
    n1402,
    n1330,
    n1475,
    n1244
  );


  or
  g1775
  (
    n1755,
    n1214,
    n1264,
    n1366,
    n1335
  );


  xor
  g1776
  (
    n1792,
    n1243,
    n1276,
    n1441,
    n1280
  );


  or
  g1777
  (
    n1582,
    n1462,
    n1351,
    n1377,
    n1312
  );


  xor
  g1778
  (
    n1631,
    n1372,
    n1239,
    n1236,
    n1342
  );


  xor
  g1779
  (
    n1576,
    n1237,
    n1381,
    n1389,
    n1466
  );


  not
  g1780
  (
    n1813,
    n1531
  );


  not
  g1781
  (
    n1810,
    n1528
  );


  not
  g1782
  (
    n1808,
    n1528
  );


  buf
  g1783
  (
    n1814,
    n1529
  );


  buf
  g1784
  (
    n1809,
    n1530
  );


  buf
  g1785
  (
    n1811,
    n1531
  );


  buf
  g1786
  (
    n1812,
    n1529
  );


  buf
  g1787
  (
    n1807,
    n1530
  );


  buf
  g1788
  (
    n1821,
    n1532
  );


  buf
  g1789
  (
    n1815,
    n1532
  );


  buf
  g1790
  (
    n1818,
    n1537
  );


  buf
  g1791
  (
    n1816,
    n1536
  );


  not
  g1792
  (
    n1817,
    n1533
  );


  not
  g1793
  (
    n1824,
    n1533
  );


  or
  g1794
  (
    n1822,
    n1534,
    n1535,
    n1809,
    n1807
  );


  and
  g1795
  (
    n1819,
    n1811,
    n1810,
    n1809,
    n1537
  );


  xnor
  g1796
  (
    n1823,
    n1808,
    n1535,
    n1536,
    n1811
  );


  or
  g1797
  (
    n1820,
    n1810,
    n1808,
    n1807,
    n1534
  );


  xnor
  g1798
  (
    n1825,
    n1815,
    n1538
  );


  xnor
  g1799
  (
    n1827,
    n1816,
    n1816,
    n1825,
    n1817
  );


  nor
  g1800
  (
    n1826,
    n1815,
    n1816,
    n1825
  );


  not
  g1801
  (
    n1828,
    n1827
  );


  and
  g1802
  (
    n1829,
    n1818,
    n1828,
    n1819,
    n1817
  );


  nand
  g1803
  (
    n1830,
    n1819,
    n1828,
    n1818
  );


  xnor
  g1804
  (
    n1831,
    n1818,
    n1817
  );


  buf
  g1805
  (
    n1832,
    n1829
  );


  xor
  g1806
  (
    n1833,
    n1812,
    n1832
  );


  nor
  g1807
  (
    KeyWire_0_17,
    n1833,
    n1820
  );


  nor
  g1808
  (
    n1836,
    n1819,
    n1820
  );


  nand
  g1809
  (
    n1835,
    n1833,
    n1833,
    n1820,
    n1819
  );


  nor
  g1810
  (
    n1846,
    n656,
    n656,
    n1830,
    n657
  );


  xor
  g1811
  (
    n1843,
    n657,
    n658,
    n1831
  );


  nor
  g1812
  (
    n1837,
    n1834,
    n1835,
    n1821,
    n828
  );


  or
  g1813
  (
    n1844,
    n829,
    n657,
    n1829,
    n1835
  );


  xnor
  g1814
  (
    n1839,
    n656,
    n1830,
    n1836
  );


  xnor
  g1815
  (
    n1838,
    n1821,
    n1836,
    n1829
  );


  and
  g1816
  (
    n1841,
    n829,
    n1821,
    n1836,
    n1832
  );


  xor
  g1817
  (
    n1845,
    n829,
    n1835,
    n1831,
    n657
  );


  nor
  g1818
  (
    n1847,
    n1835,
    n658,
    n828
  );


  nand
  g1819
  (
    n1848,
    n656,
    n655,
    n1834,
    n1828
  );


  or
  g1820
  (
    n1842,
    n1831,
    n1830,
    n658,
    n1833
  );


  xnor
  g1821
  (
    n1840,
    n1821,
    n1834,
    n1836
  );


  and
  g1822
  (
    n1850,
    n1483,
    n1846,
    n1837,
    n1482
  );


  nor
  g1823
  (
    n1874,
    n1481,
    n1540,
    n1484,
    n1823
  );


  xor
  g1824
  (
    n1857,
    n1822,
    n1543,
    n290,
    n1841
  );


  nor
  g1825
  (
    n1870,
    n1483,
    n1839,
    n289,
    n1847
  );


  xnor
  g1826
  (
    n1873,
    n1541,
    n1848,
    n1837,
    n1823
  );


  or
  g1827
  (
    n1860,
    n1484,
    n1548,
    n1487,
    n1485
  );


  or
  g1828
  (
    n1863,
    n1848,
    n1846,
    n1841,
    n1484
  );


  nor
  g1829
  (
    n1865,
    n1539,
    n1546,
    n289
  );


  nand
  g1830
  (
    n1861,
    n1549,
    n1480,
    n1841,
    n1844
  );


  nor
  g1831
  (
    n1849,
    n1545,
    n1837,
    n1543,
    n1542
  );


  and
  g1832
  (
    n1868,
    n1842,
    n1547,
    n1551,
    n1550
  );


  nand
  g1833
  (
    n1866,
    n1842,
    n1838,
    n1488,
    n1549
  );


  or
  g1834
  (
    n1851,
    n1845,
    n1823,
    n1839,
    n1837
  );


  and
  g1835
  (
    n1864,
    n1843,
    n1822,
    n1487,
    n1842
  );


  or
  g1836
  (
    n1877,
    n1841,
    n731,
    n1481,
    n1823
  );


  nor
  g1837
  (
    n1852,
    n1485,
    n1485,
    n1540,
    n1483
  );


  and
  g1838
  (
    n1867,
    n1488,
    n1544,
    n1844,
    n1838
  );


  nor
  g1839
  (
    n1858,
    n1482,
    n290,
    n1486,
    n1484
  );


  or
  g1840
  (
    n1862,
    n1848,
    n290,
    n1845,
    n1840
  );


  nand
  g1841
  (
    n1854,
    n1482,
    n1822,
    n1838,
    n1548
  );


  nor
  g1842
  (
    n1855,
    n290,
    n1840,
    n1486
  );


  xnor
  g1843
  (
    n1872,
    n1487,
    n1845,
    n1488,
    n1485
  );


  nand
  g1844
  (
    n1876,
    n1542,
    n1847,
    n1844,
    n1487
  );


  or
  g1845
  (
    n1856,
    n1839,
    n1838,
    n1822,
    n1846
  );


  nor
  g1846
  (
    n1869,
    n1842,
    n1481,
    n1845,
    n1843
  );


  or
  g1847
  (
    n1878,
    n1847,
    n731,
    n1547,
    n1839
  );


  or
  g1848
  (
    n1879,
    n1846,
    n1483,
    n1545,
    n1486
  );


  xnor
  g1849
  (
    n1875,
    n1541,
    n1486,
    n1480,
    n1550
  );


  nor
  g1850
  (
    n1871,
    n1848,
    n1843,
    n1544
  );


  xnor
  g1851
  (
    n1859,
    n1539,
    n1488,
    n1480,
    n1844
  );


  and
  g1852
  (
    n1853,
    n1482,
    n1840,
    n1481,
    n1847
  );


  not
  g1853
  (
    n1888,
    n1849
  );


  buf
  g1854
  (
    n1884,
    n1851
  );


  not
  g1855
  (
    n1880,
    n1850
  );


  buf
  g1856
  (
    n1886,
    n1851
  );


  buf
  g1857
  (
    n1889,
    n1849
  );


  not
  g1858
  (
    n1882,
    n1849
  );


  buf
  g1859
  (
    n1887,
    n1850
  );


  not
  g1860
  (
    n1885,
    n1849
  );


  not
  g1861
  (
    n1881,
    n1850
  );


  not
  g1862
  (
    n1883,
    n1850
  );


  xor
  g1863
  (
    KeyWire_0_60,
    n1869,
    n1881,
    n1887,
    n1888
  );


  xnor
  g1864
  (
    n1913,
    n1855,
    n1880,
    n1859,
    n1861
  );


  xnor
  g1865
  (
    n1920,
    n1876,
    n1856,
    n1858,
    n1860
  );


  xor
  g1866
  (
    n1929,
    n1878,
    n1851,
    n1854,
    n1889
  );


  nor
  g1867
  (
    n1890,
    n1883,
    n1863,
    n1856,
    n1866
  );


  nor
  g1868
  (
    n1895,
    n1862,
    n1886,
    n1866,
    n1876
  );


  or
  g1869
  (
    n1919,
    n1884,
    n1887,
    n1874,
    n1859
  );


  xnor
  g1870
  (
    n1909,
    n1861,
    n1889,
    n1885,
    n1870
  );


  xnor
  g1871
  (
    n1899,
    n1877,
    n1872,
    n1812,
    n1882
  );


  or
  g1872
  (
    n1898,
    n1870,
    n1861,
    n1871
  );


  and
  g1873
  (
    n1902,
    n1877,
    n1869,
    n1884,
    n1866
  );


  nor
  g1874
  (
    n1910,
    n1858,
    n1880,
    n1886,
    n1862
  );


  nor
  g1875
  (
    n1925,
    n1860,
    n1888,
    n1879,
    n1873
  );


  xnor
  g1876
  (
    n1891,
    n1881,
    n1882,
    n1853,
    n1813
  );


  xor
  g1877
  (
    n1915,
    n1865,
    n1872,
    n1855,
    n1879
  );


  or
  g1878
  (
    n1911,
    n1875,
    n1885,
    n1863,
    n1883
  );


  xor
  g1879
  (
    n1893,
    n1867,
    n1869,
    n1870,
    n1857
  );


  xnor
  g1880
  (
    n1922,
    n1852,
    n1852,
    n1878,
    n1882
  );


  xor
  g1881
  (
    n1918,
    n1871,
    n1884,
    n1814,
    n1873
  );


  xnor
  g1882
  (
    n1921,
    n1881,
    n1880,
    n1864,
    n1859
  );


  and
  g1883
  (
    n1914,
    n1865,
    n1881,
    n1863,
    n1874
  );


  nand
  g1884
  (
    n1907,
    n1855,
    n1857,
    n1851,
    n1885
  );


  nand
  g1885
  (
    n1905,
    n1871,
    n1860,
    n1867,
    n1888
  );


  or
  g1886
  (
    n1927,
    n1858,
    n1852,
    n1889,
    n1860
  );


  xnor
  g1887
  (
    n1928,
    n1875,
    n1876,
    n1867,
    n1853
  );


  xnor
  g1888
  (
    n1904,
    n1884,
    n1883,
    n1877,
    n1814
  );


  or
  g1889
  (
    n1906,
    n1857,
    n1878,
    n1853,
    n1814
  );


  xnor
  g1890
  (
    n1897,
    n1885,
    n1854
  );


  and
  g1891
  (
    n1926,
    n1874,
    n1856,
    n1883,
    n1875
  );


  nand
  g1892
  (
    n1923,
    n1868,
    n1864,
    n1870,
    n1872
  );


  and
  g1893
  (
    n1894,
    n1865,
    n1878,
    n1886,
    n1880
  );


  nand
  g1894
  (
    n1917,
    n1867,
    n1873,
    n1858,
    n1871
  );


  or
  g1895
  (
    n1896,
    n1853,
    n1877,
    n1879
  );


  nand
  g1896
  (
    n1892,
    n1875,
    n1855,
    n1874,
    n1873
  );


  xnor
  g1897
  (
    n1924,
    n1868,
    n1888,
    n1876,
    n1857
  );


  xnor
  g1898
  (
    n1900,
    n1864,
    n1866,
    n1859,
    n1872
  );


  xnor
  g1899
  (
    n1903,
    n1864,
    n1882,
    n1862,
    n1868
  );


  xnor
  g1900
  (
    n1901,
    n1852,
    n1886,
    n1856,
    n1863
  );


  nand
  g1901
  (
    n1916,
    n1889,
    n1865,
    n1862,
    n1868
  );


  and
  g1902
  (
    n1908,
    n1813,
    n1887,
    n1869
  );


  xor
  g1903
  (
    n1930,
    n1890,
    n1824
  );


  and
  g1904
  (
    n1932,
    n1891,
    n1930,
    n1892
  );


  nand
  g1905
  (
    n1934,
    n1890,
    n1892,
    n1895
  );


  and
  g1906
  (
    n1933,
    n1894,
    n1930,
    n1893,
    n1896
  );


  nor
  g1907
  (
    n1931,
    n1891,
    n1893,
    n1930,
    n1894
  );


  and
  g1908
  (
    n1945,
    n832,
    n1933,
    n1910
  );


  nand
  g1909
  (
    n1937,
    n1898,
    n1911,
    n1908,
    n1902
  );


  nor
  g1910
  (
    n1939,
    n1933,
    n1899,
    n1931,
    n1905
  );


  or
  g1911
  (
    KeyWire_0_30,
    n1932,
    n1933,
    n1909,
    n831
  );


  and
  g1912
  (
    n1935,
    n1910,
    n1904,
    n1934,
    n1901
  );


  nor
  g1913
  (
    n1948,
    n1900,
    n1896,
    n832,
    n830
  );


  or
  g1914
  (
    n1947,
    n833,
    n1931,
    n1905
  );


  nor
  g1915
  (
    n1946,
    n1901,
    n1932,
    n1898,
    n1906
  );


  xor
  g1916
  (
    n1949,
    n832,
    n830,
    n1906
  );


  nand
  g1917
  (
    n1941,
    n832,
    n1911,
    n831,
    n1909
  );


  nor
  g1918
  (
    n1942,
    n1932,
    n1902,
    n1907,
    n1897
  );


  or
  g1919
  (
    n1938,
    n831,
    n1907,
    n1934,
    n1931
  );


  xor
  g1920
  (
    n1943,
    n831,
    n1934,
    n1908,
    n1899
  );


  nor
  g1921
  (
    n1940,
    n1932,
    n1903,
    n1904,
    n1900
  );


  nand
  g1922
  (
    n1936,
    n1897,
    n829,
    n830,
    n1903
  );


  not
  g1923
  (
    n1953,
    n1948
  );


  buf
  g1924
  (
    n1954,
    n1947
  );


  buf
  g1925
  (
    n1952,
    n1949
  );


  buf
  g1926
  (
    n1951,
    n1949
  );


  not
  g1927
  (
    n1950,
    n1948
  );


  nand
  g1928
  (
    n1961,
    n1924,
    n1951,
    n1950,
    n1927
  );


  xor
  g1929
  (
    n1969,
    n1921,
    n1953,
    n1912
  );


  and
  g1930
  (
    n1964,
    n1914,
    n1954,
    n1918,
    n1922
  );


  and
  g1931
  (
    n1956,
    n1921,
    n1950,
    n1915,
    n1926
  );


  and
  g1932
  (
    n1962,
    n1952,
    n1929,
    n1928,
    n1925
  );


  and
  g1933
  (
    n1958,
    n1916,
    n1921,
    n1923
  );


  xor
  g1934
  (
    n1968,
    n1951,
    n1919,
    n1920
  );


  and
  g1935
  (
    n1959,
    n1924,
    n1929,
    n1950
  );


  xor
  g1936
  (
    n1957,
    n1954,
    n1927,
    n1917,
    n1952
  );


  and
  g1937
  (
    n1970,
    n1925,
    n1924,
    n1952,
    n1926
  );


  xnor
  g1938
  (
    n1971,
    n1923,
    n1915,
    n1928,
    n1913
  );


  and
  g1939
  (
    n1955,
    n1926,
    n1914,
    n1919,
    n1928
  );


  and
  g1940
  (
    n1974,
    n1927,
    n1928,
    n1923,
    n1916
  );


  xor
  g1941
  (
    KeyWire_0_6,
    n1954,
    n1922,
    n1952,
    n1953
  );


  nor
  g1942
  (
    n1960,
    n1950,
    n1913,
    n1924,
    n1951
  );


  nor
  g1943
  (
    n1966,
    n1920,
    n1927,
    n1918
  );


  nand
  g1944
  (
    n1972,
    n1919,
    n1953,
    n1925,
    n1926
  );


  nor
  g1945
  (
    n1963,
    n1929,
    n1951,
    n1923,
    n1920
  );


  xor
  g1946
  (
    n1965,
    n1918,
    n1922,
    n1954
  );


  and
  g1947
  (
    n1967,
    n1925,
    n1917,
    n1920,
    n1912
  );


  nand
  g1948
  (
    n1985,
    n1973,
    n1517,
    n1513,
    n1491
  );


  nand
  g1949
  (
    n2043,
    n834,
    n1508,
    n1496,
    n1500
  );


  nor
  g1950
  (
    n1984,
    n841,
    n1526,
    n1969,
    n1492
  );


  xnor
  g1951
  (
    n2027,
    n843,
    n1493,
    n845,
    n1934
  );


  or
  g1952
  (
    n2035,
    n1505,
    n843,
    n1559,
    n1557
  );


  nor
  g1953
  (
    n2039,
    n1492,
    n833,
    n1556,
    n1968
  );


  and
  g1954
  (
    n1996,
    n1516,
    n1489,
    n845,
    n1955
  );


  nor
  g1955
  (
    n2013,
    n1503,
    n1969,
    n843,
    n1525
  );


  xor
  g1956
  (
    KeyWire_0_39,
    n1493,
    n1971,
    n1512,
    n842
  );


  xnor
  g1957
  (
    n2022,
    n1520,
    n1521,
    n1492,
    n1502
  );


  xor
  g1958
  (
    n2005,
    n836,
    n1516,
    n1523,
    n1965
  );


  xor
  g1959
  (
    n2008,
    n1968,
    n1960,
    n1519,
    n1521
  );


  or
  g1960
  (
    n1981,
    n1489,
    n513,
    n840,
    n1967
  );


  and
  g1961
  (
    n1991,
    n843,
    n1526,
    n837,
    n1517
  );


  nor
  g1962
  (
    n1986,
    n1961,
    n1960,
    n1524,
    n844
  );


  xor
  g1963
  (
    n2025,
    n1509,
    n1493,
    n518,
    n1494
  );


  xnor
  g1964
  (
    n2033,
    n1963,
    n1514,
    n1526,
    n1512
  );


  and
  g1965
  (
    n2003,
    n513,
    n1501,
    n1512,
    n1522
  );


  nor
  g1966
  (
    n2047,
    n1553,
    n517,
    n1554,
    n1555
  );


  nand
  g1967
  (
    n2015,
    n1959,
    n1518,
    n1558,
    n1500
  );


  nor
  g1968
  (
    n2052,
    n1508,
    n1968,
    n835,
    n1516
  );


  nor
  g1969
  (
    n2029,
    n834,
    n1503,
    n1499
  );


  nand
  g1970
  (
    n2010,
    n1512,
    n1495,
    n1504,
    n1499
  );


  nand
  g1971
  (
    n2012,
    n1498,
    n1519,
    n833,
    n1964
  );


  or
  g1972
  (
    n2046,
    n1506,
    n1527,
    n1956,
    n1518
  );


  xor
  g1973
  (
    n1998,
    n1525,
    n1959,
    n1497,
    n1504
  );


  or
  g1974
  (
    n1979,
    n1515,
    n836,
    n1525,
    n1974
  );


  nor
  g1975
  (
    n2006,
    n1517,
    n842,
    n1552,
    n1504
  );


  or
  g1976
  (
    n2040,
    n1496,
    n1519,
    n1507,
    n1513
  );


  xnor
  g1977
  (
    n1999,
    n1970,
    n1510,
    n835,
    n1522
  );


  and
  g1978
  (
    n2031,
    n841,
    n514,
    n834,
    n1958
  );


  nor
  g1979
  (
    n1975,
    n841,
    n1511,
    n1502
  );


  nor
  g1980
  (
    n1997,
    n837,
    n1522,
    n840,
    n1970
  );


  nor
  g1981
  (
    n2034,
    n1959,
    n835,
    n1495,
    n1824
  );


  and
  g1982
  (
    n2049,
    n517,
    n1521,
    n1507,
    n1962
  );


  xnor
  g1983
  (
    n2016,
    n1514,
    n1498,
    n1518,
    n515
  );


  nor
  g1984
  (
    n1990,
    n1520,
    n839,
    n1963,
    n1956
  );


  and
  g1985
  (
    n2023,
    n838,
    n845,
    n1489,
    n1554
  );


  nor
  g1986
  (
    n2011,
    n1495,
    n1972,
    n1965,
    n844
  );


  xnor
  g1987
  (
    n2001,
    n1961,
    n1955,
    n1967,
    n1969
  );


  xnor
  g1988
  (
    n2000,
    n1510,
    n1502,
    n838,
    n519
  );


  nor
  g1989
  (
    n1988,
    n1520,
    n1973,
    n1523,
    n1522
  );


  nand
  g1990
  (
    n2032,
    n1499,
    n1973,
    n1524,
    n1491
  );


  xnor
  g1991
  (
    n1976,
    n1966,
    n1497,
    n1515,
    n1491
  );


  nor
  g1992
  (
    n2017,
    n1504,
    n1490,
    n1500,
    n1514
  );


  or
  g1993
  (
    n1993,
    n1524,
    n1959,
    n1964,
    n1527
  );


  nor
  g1994
  (
    n2041,
    n1490,
    n1496,
    n1973,
    n1516
  );


  nand
  g1995
  (
    n2038,
    n1507,
    n1557,
    n1508,
    n1490
  );


  and
  g1996
  (
    n1982,
    n1964,
    n1972,
    n514,
    n1957
  );


  nand
  g1997
  (
    n2019,
    n1972,
    n840,
    n1974,
    n836
  );


  xor
  g1998
  (
    n1995,
    n1501,
    n844,
    n1513,
    n1494
  );


  xnor
  g1999
  (
    n2004,
    n1505,
    n1510,
    n1559,
    n1511
  );


  nand
  g2000
  (
    n2002,
    n1958,
    n1958,
    n1966,
    n518
  );


  or
  g2001
  (
    n2042,
    n1490,
    n1524,
    n1501,
    n1527
  );


  and
  g2002
  (
    n2045,
    n1957,
    n1971,
    n1513,
    n1511
  );


  or
  g2003
  (
    n1977,
    n1960,
    n1968,
    n845,
    n1527
  );


  xnor
  g2004
  (
    n1983,
    n1963,
    n1553,
    n1961,
    n838
  );


  nand
  g2005
  (
    n1994,
    n1515,
    n1493,
    n833,
    n1496
  );


  xnor
  g2006
  (
    n2036,
    n837,
    n1967,
    n1957,
    n840
  );


  nand
  g2007
  (
    n2051,
    n1970,
    n1523,
    n1518,
    n1965
  );


  xor
  g2008
  (
    n2024,
    n1511,
    n1498,
    n1515,
    n1507
  );


  xor
  g2009
  (
    n1987,
    n837,
    n1506,
    n1520,
    n1971
  );


  or
  g2010
  (
    n2021,
    n1974,
    n1514,
    n1556,
    n1500
  );


  nor
  g2011
  (
    n2020,
    n834,
    n515,
    n1489,
    n1505
  );


  xnor
  g2012
  (
    KeyWire_0_55,
    n1961,
    n1555,
    n1505,
    n836
  );


  xnor
  g2013
  (
    n1980,
    n1956,
    n1508,
    n1497,
    n1966
  );


  nand
  g2014
  (
    n2030,
    n1519,
    n1509,
    n1491,
    n842
  );


  nor
  g2015
  (
    n2037,
    n839,
    n841,
    n1962,
    n516
  );


  nand
  g2016
  (
    n2050,
    n1492,
    n839,
    n1498,
    n1957
  );


  and
  g2017
  (
    n2026,
    n1962,
    n1521,
    n1964,
    n1525
  );


  or
  g2018
  (
    n2014,
    n1501,
    n1509,
    n1494,
    n1497
  );


  or
  g2019
  (
    n2054,
    n842,
    n1509,
    n1506,
    n1503
  );


  and
  g2020
  (
    n2009,
    n1970,
    n1971,
    n1962,
    n1960
  );


  nand
  g2021
  (
    n1989,
    n1494,
    n839,
    n519,
    n1499
  );


  nor
  g2022
  (
    n1978,
    n1558,
    n1963,
    n844,
    n1967
  );


  nor
  g2023
  (
    n1992,
    n1956,
    n835,
    n1969,
    n1552
  );


  nor
  g2024
  (
    KeyWire_0_5,
    n1965,
    n1526,
    n1955
  );


  and
  g2025
  (
    n2007,
    n1510,
    n1551,
    n1966,
    n1506
  );


  or
  g2026
  (
    n2048,
    n838,
    n1523,
    n1974,
    n1972
  );


  or
  g2027
  (
    n2028,
    n1958,
    n1517,
    n516,
    n1495
  );


  and
  g2028
  (
    n2164,
    n1633,
    n1737,
    n1791,
    n1990
  );


  or
  g2029
  (
    n2187,
    n1578,
    n2016,
    n1591,
    n1796
  );


  nand
  g2030
  (
    KeyWire_0_31,
    n2014,
    n2050,
    n1575,
    n1584
  );


  and
  g2031
  (
    n2266,
    n2022,
    n2047,
    n2034,
    n1699
  );


  xor
  g2032
  (
    n2319,
    n1625,
    n2009,
    n1594,
    n1700
  );


  xnor
  g2033
  (
    n2085,
    n1640,
    n1607,
    n1604,
    n1660
  );


  nand
  g2034
  (
    n2242,
    n1687,
    n1666,
    n2042,
    n1592
  );


  nor
  g2035
  (
    n2120,
    n1741,
    n2039,
    n1984,
    n1690
  );


  nand
  g2036
  (
    n2357,
    n1607,
    n1606,
    n2044,
    n1713
  );


  and
  g2037
  (
    n2354,
    n1800,
    n1991,
    n2024,
    n1706
  );


  xor
  g2038
  (
    n2059,
    n1699,
    n1688,
    n1787,
    n2032
  );


  nor
  g2039
  (
    n2244,
    n1623,
    n1734,
    n1560,
    n1780
  );


  xnor
  g2040
  (
    n2190,
    n1781,
    n1993,
    n1711,
    n1563
  );


  or
  g2041
  (
    n2307,
    n1739,
    n2016,
    n1989,
    n1673
  );


  and
  g2042
  (
    n2073,
    n1695,
    n1711,
    n1798,
    n1665
  );


  xnor
  g2043
  (
    n2122,
    n1626,
    n1617,
    n1794,
    n1618
  );


  and
  g2044
  (
    n2070,
    n1805,
    n1736,
    n1740,
    n1634
  );


  nor
  g2045
  (
    n2333,
    n1762,
    n1770,
    n1730,
    n2019
  );


  nand
  g2046
  (
    n2151,
    n1641,
    n2015,
    n2036,
    n2026
  );


  and
  g2047
  (
    n2168,
    n2053,
    n1762,
    n1682,
    n1668
  );


  or
  g2048
  (
    n2135,
    n1657,
    n2030,
    n1987,
    n1624
  );


  xor
  g2049
  (
    n2111,
    n1647,
    n1591,
    n1688,
    n1999
  );


  or
  g2050
  (
    n2094,
    n1781,
    n1646,
    n1569,
    n1977
  );


  and
  g2051
  (
    n2277,
    n2002,
    n2028,
    n1650,
    n1667
  );


  xnor
  g2052
  (
    n2121,
    n2026,
    n1801,
    n1603,
    n1755
  );


  xor
  g2053
  (
    n2271,
    n1748,
    n1802,
    n1978,
    n1570
  );


  xor
  g2054
  (
    n2199,
    n1992,
    n1999,
    n1565,
    n2049
  );


  and
  g2055
  (
    n2213,
    n1988,
    n2011,
    n1785,
    n1716
  );


  xor
  g2056
  (
    n2347,
    n1726,
    n1562,
    n1787,
    n1977
  );


  or
  g2057
  (
    n2336,
    n1567,
    n1672,
    n1985,
    n1713
  );


  xnor
  g2058
  (
    n2256,
    n2006,
    n1983,
    n1705,
    n2025
  );


  xnor
  g2059
  (
    n2063,
    n1686,
    n1995,
    n1631,
    n1671
  );


  nand
  g2060
  (
    n2203,
    n1764,
    n1779,
    n1655,
    n1606
  );


  and
  g2061
  (
    n2143,
    n1564,
    n1609,
    n1651,
    n2007
  );


  nand
  g2062
  (
    n2218,
    n1752,
    n1797,
    n1668,
    n1645
  );


  xnor
  g2063
  (
    n2175,
    n2019,
    n1648,
    n1986
  );


  xnor
  g2064
  (
    n2329,
    n1745,
    n1679,
    n1800,
    n1576
  );


  xor
  g2065
  (
    n2237,
    n1711,
    n1795,
    n1585,
    n1641
  );


  and
  g2066
  (
    n2189,
    n1777,
    n1771,
    n1980,
    n1698
  );


  xnor
  g2067
  (
    n2344,
    n1983,
    n1741,
    n1752,
    n1761
  );


  nor
  g2068
  (
    n2207,
    n1593,
    n1606,
    n1785,
    n1759
  );


  nand
  g2069
  (
    n2263,
    n1662,
    n1645,
    n2054,
    n1588
  );


  nor
  g2070
  (
    n2351,
    n1582,
    n1610,
    n1770,
    n1712
  );


  xnor
  g2071
  (
    n2126,
    n1782,
    n1565,
    n1764,
    n1576
  );


  nor
  g2072
  (
    n2300,
    n1993,
    n1717,
    n1609,
    n2039
  );


  or
  g2073
  (
    n2148,
    n2036,
    n1766,
    n1753,
    n1733
  );


  and
  g2074
  (
    n2310,
    n2027,
    n1804,
    n2033,
    n1722
  );


  xor
  g2075
  (
    n2119,
    n1583,
    n1639,
    n1732,
    n2017
  );


  and
  g2076
  (
    n2255,
    n1747,
    n1604,
    n1599,
    n1616
  );


  nand
  g2077
  (
    n2340,
    n1701,
    n1694,
    n1999,
    n1564
  );


  and
  g2078
  (
    n2231,
    n1569,
    n1633,
    n2004,
    n2041
  );


  nand
  g2079
  (
    n2246,
    n1667,
    n1632,
    n1670,
    n1985
  );


  nor
  g2080
  (
    n2069,
    n1792,
    n2033,
    n1684,
    n1715
  );


  nor
  g2081
  (
    n2259,
    n1607,
    n1695,
    n1601,
    n1629
  );


  nand
  g2082
  (
    n2243,
    n1566,
    n1602,
    n1684,
    n1750
  );


  nand
  g2083
  (
    n2249,
    n1791,
    n1634,
    n2001,
    n1596
  );


  xnor
  g2084
  (
    n2299,
    n2040,
    n1577,
    n1990,
    n1749
  );


  xnor
  g2085
  (
    n2303,
    n1642,
    n1744,
    n2049,
    n1975
  );


  or
  g2086
  (
    n2147,
    n1561,
    n1997,
    n1782,
    n1767
  );


  nor
  g2087
  (
    n2154,
    n1585,
    n2039,
    n1699,
    n1705
  );


  or
  g2088
  (
    n2087,
    n1981,
    n1565,
    n1705,
    n1646
  );


  nor
  g2089
  (
    n2077,
    n1731,
    n1649,
    n2017,
    n1635
  );


  nand
  g2090
  (
    n2309,
    n1790,
    n1651,
    n2051,
    n1782
  );


  or
  g2091
  (
    n2356,
    n1805,
    n1567,
    n2034,
    n1683
  );


  or
  g2092
  (
    n2176,
    n1707,
    n1564,
    n1681,
    n2011
  );


  or
  g2093
  (
    n2366,
    n1772,
    n1652,
    n2042,
    n1727
  );


  xnor
  g2094
  (
    n2233,
    n1671,
    n1751,
    n1613,
    n1786
  );


  nor
  g2095
  (
    n2269,
    n1773,
    n1687,
    n1578,
    n2046
  );


  or
  g2096
  (
    n2224,
    n1571,
    n1686,
    n1640,
    n1743
  );


  nor
  g2097
  (
    n2323,
    n1641,
    n1789,
    n2002,
    n1629
  );


  xnor
  g2098
  (
    KeyWire_0_29,
    n1673,
    n2020,
    n1805,
    n1663
  );


  nand
  g2099
  (
    n2359,
    n1990,
    n1637,
    n1629,
    n1577
  );


  xor
  g2100
  (
    n2208,
    n1715,
    n1602,
    n2002,
    n1749
  );


  and
  g2101
  (
    n2225,
    n1745,
    n2043,
    n2003,
    n2025
  );


  nor
  g2102
  (
    n2273,
    n1717,
    n1798,
    n1758,
    n1984
  );


  nor
  g2103
  (
    n2338,
    n1672,
    n1560,
    n1734,
    n1987
  );


  and
  g2104
  (
    n2315,
    n1751,
    n2050,
    n1698,
    n1756
  );


  and
  g2105
  (
    n2130,
    n1603,
    n2021,
    n1794
  );


  nor
  g2106
  (
    n2239,
    n1999,
    n1795,
    n1588,
    n1574
  );


  xor
  g2107
  (
    n2312,
    n1587,
    n1667,
    n1621,
    n2018
  );


  nor
  g2108
  (
    n2082,
    n1744,
    n1620,
    n1611,
    n1709
  );


  or
  g2109
  (
    n2262,
    n1749,
    n1776,
    n1788,
    n2001
  );


  nor
  g2110
  (
    n2220,
    n2053,
    n1738,
    n2023,
    n1599
  );


  and
  g2111
  (
    n2332,
    n1758,
    n2011,
    n1776,
    n2019
  );


  and
  g2112
  (
    n2355,
    n1976,
    n1648,
    n2012,
    n1656
  );


  nor
  g2113
  (
    n2095,
    n1682,
    n1721,
    n1594,
    n1988
  );


  nor
  g2114
  (
    n2250,
    n1775,
    n1713,
    n1601,
    n1610
  );


  nand
  g2115
  (
    n2295,
    n1720,
    n1722,
    n1753,
    n1771
  );


  nand
  g2116
  (
    n2251,
    n1589,
    n1997,
    n1725,
    n1790
  );


  or
  g2117
  (
    n2308,
    n1772,
    n1610,
    n1628,
    n1581
  );


  xnor
  g2118
  (
    n2058,
    n1994,
    n1662,
    n1675,
    n2020
  );


  and
  g2119
  (
    n2289,
    n2019,
    n1561,
    n2050,
    n1640
  );


  or
  g2120
  (
    n2293,
    n1717,
    n1685,
    n1705,
    n1629
  );


  nand
  g2121
  (
    n2223,
    n1633,
    n1684,
    n2001,
    n1634
  );


  xnor
  g2122
  (
    n2304,
    n1673,
    n1727,
    n1691,
    n1589
  );


  and
  g2123
  (
    n2186,
    n1979,
    n1738,
    n1571,
    n1770
  );


  and
  g2124
  (
    n2125,
    n2008,
    n1758,
    n2042,
    n1568
  );


  nor
  g2125
  (
    n2089,
    n1773,
    n1607,
    n1696,
    n1726
  );


  and
  g2126
  (
    n2112,
    n1651,
    n1778,
    n1975,
    n2011
  );


  xnor
  g2127
  (
    n2342,
    n1615,
    n1640,
    n1636,
    n2006
  );


  nand
  g2128
  (
    n2162,
    n1590,
    n1777,
    n1649,
    n1587
  );


  xnor
  g2129
  (
    n2345,
    n1706,
    n1744,
    n1774,
    n1769
  );


  xor
  g2130
  (
    n2292,
    n2037,
    n1701,
    n1674,
    n1586
  );


  nor
  g2131
  (
    n2173,
    n1706,
    n1718,
    n2045,
    n2009
  );


  or
  g2132
  (
    n2104,
    n1681,
    n1665,
    n1998,
    n1746
  );


  xnor
  g2133
  (
    n2171,
    n1979,
    n1756,
    n1994,
    n1594
  );


  or
  g2134
  (
    n2064,
    n1581,
    n2036,
    n2024,
    n1732
  );


  xor
  g2135
  (
    n2296,
    n1782,
    n1694,
    n1721,
    n1644
  );


  and
  g2136
  (
    n2353,
    n1676,
    n1708,
    n1707,
    n1572
  );


  xnor
  g2137
  (
    n2330,
    n1661,
    n1996,
    n1739,
    n1757
  );


  xor
  g2138
  (
    n2214,
    n1624,
    n1996,
    n1602,
    n1643
  );


  xor
  g2139
  (
    n2201,
    n1755,
    n1697,
    n2031,
    n1792
  );


  or
  g2140
  (
    n2280,
    n1563,
    n1700,
    n1989,
    n1775
  );


  or
  g2141
  (
    n2097,
    n1605,
    n1574,
    n1737,
    n1717
  );


  and
  g2142
  (
    n2313,
    n1724,
    n2038,
    n1560,
    n2004
  );


  xnor
  g2143
  (
    n2114,
    n1626,
    n1765,
    n2032,
    n1977
  );


  xnor
  g2144
  (
    n2221,
    n2044,
    n1799,
    n1780,
    n1597
  );


  nor
  g2145
  (
    n2177,
    n1731,
    n1735,
    n1748,
    n1995
  );


  and
  g2146
  (
    n2285,
    n2031,
    n1765,
    n1628,
    n1653
  );


  or
  g2147
  (
    n2193,
    n1644,
    n1689,
    n1635,
    n1725
  );


  xnor
  g2148
  (
    n2202,
    n2015,
    n1738,
    n1692,
    n1728
  );


  xnor
  g2149
  (
    n2352,
    n1662,
    n1659,
    n1613,
    n1597
  );


  nor
  g2150
  (
    n2341,
    n2028,
    n1801,
    n1746,
    n1769
  );


  or
  g2151
  (
    n2258,
    n2052,
    n2025,
    n1563,
    n1736
  );


  nand
  g2152
  (
    n2105,
    n1775,
    n1741,
    n1663,
    n1796
  );


  nand
  g2153
  (
    n2363,
    n1631,
    n1994,
    n1658,
    n1691
  );


  xnor
  g2154
  (
    n2179,
    n1784,
    n2020,
    n2009,
    n2053
  );


  nor
  g2155
  (
    n2294,
    n1619,
    n1675,
    n1788,
    n1753
  );


  nor
  g2156
  (
    n2174,
    n2045,
    n1621,
    n1656,
    n2024
  );


  nor
  g2157
  (
    n2099,
    n2052,
    n1784,
    n2047,
    n1777
  );


  xnor
  g2158
  (
    n2320,
    n1573,
    n1797,
    n1608,
    n1659
  );


  or
  g2159
  (
    n2182,
    n2030,
    n1718,
    n1730,
    n1997
  );


  and
  g2160
  (
    n2109,
    n1793,
    n1710,
    n1689,
    n2035
  );


  nand
  g2161
  (
    n2267,
    n1784,
    n1980,
    n1768,
    n1756
  );


  and
  g2162
  (
    n2056,
    n2027,
    n1733,
    n1651,
    n1708
  );


  xor
  g2163
  (
    n2282,
    n2004,
    n1987,
    n1698,
    n1754
  );


  or
  g2164
  (
    n2209,
    n1731,
    n1600,
    n1976,
    n1646
  );


  and
  g2165
  (
    n2358,
    n2022,
    n1792,
    n1636,
    n2026
  );


  nor
  g2166
  (
    n2248,
    n1723,
    n1766,
    n2037,
    n2006
  );


  xor
  g2167
  (
    n2160,
    n2010,
    n2004,
    n2040,
    n1595
  );


  nor
  g2168
  (
    n2149,
    n1781,
    n1620,
    n1590,
    n1746
  );


  xnor
  g2169
  (
    n2362,
    n1632,
    n1692,
    n1763,
    n2054
  );


  and
  g2170
  (
    n2346,
    n1690,
    n2050,
    n1587,
    n2000
  );


  xnor
  g2171
  (
    n2150,
    n1674,
    n1979,
    n2002,
    n1645
  );


  and
  g2172
  (
    n2116,
    n2048,
    n2018,
    n1780,
    n1676
  );


  nand
  g2173
  (
    n2178,
    n1643,
    n1984,
    n1608,
    n1790
  );


  xor
  g2174
  (
    n2327,
    n1750,
    n1625,
    n2046,
    n1789
  );


  xor
  g2175
  (
    n2159,
    n1645,
    n1804,
    n1981,
    n1991
  );


  or
  g2176
  (
    n2337,
    n2027,
    n1642,
    n2008,
    n1727
  );


  and
  g2177
  (
    n2291,
    n2005,
    n1572,
    n2052,
    n1685
  );


  nand
  g2178
  (
    n2311,
    n1991,
    n1664,
    n2020
  );


  xor
  g2179
  (
    n2194,
    n1623,
    n1617,
    n2022,
    n1803
  );


  nand
  g2180
  (
    n2368,
    n1673,
    n1609,
    n1686,
    n1630
  );


  and
  g2181
  (
    n2305,
    n1762,
    n1684,
    n2005,
    n1672
  );


  and
  g2182
  (
    KeyWire_0_54,
    n1638,
    n1584,
    n1704,
    n1740
  );


  and
  g2183
  (
    n2170,
    n1665,
    n1773,
    n1703,
    n1783
  );


  nand
  g2184
  (
    n2195,
    n2013,
    n2030,
    n1668,
    n1679
  );


  nand
  g2185
  (
    n2367,
    n2023,
    n1784,
    n1990,
    n1725
  );


  xnor
  g2186
  (
    n2086,
    n1605,
    n1706,
    n1562,
    n2049
  );


  nand
  g2187
  (
    n2166,
    n1787,
    n1710,
    n1593,
    n1737
  );


  or
  g2188
  (
    n2079,
    n2012,
    n1644,
    n1683,
    n1767
  );


  xor
  g2189
  (
    n2096,
    n1709,
    n2041,
    n1781,
    n1644
  );


  or
  g2190
  (
    n2228,
    n1986,
    n1693,
    n1590,
    n1622
  );


  and
  g2191
  (
    n2211,
    n1752,
    n1616,
    n1666,
    n1592
  );


  or
  g2192
  (
    KeyWire_0_56,
    n1982,
    n2032,
    n1617,
    n2003
  );


  or
  g2193
  (
    n2146,
    n1997,
    n1724,
    n2000,
    n1753
  );


  nand
  g2194
  (
    n2227,
    n1790,
    n1976,
    n1744,
    n1666
  );


  nand
  g2195
  (
    n2072,
    n1700,
    n1709,
    n1586,
    n1802
  );


  nand
  g2196
  (
    n2372,
    n1627,
    n1759,
    n1630,
    n1568
  );


  nor
  g2197
  (
    n2068,
    n1799,
    n1598,
    n2007,
    n1681
  );


  and
  g2198
  (
    n2314,
    n1632,
    n1592,
    n1669,
    n1614
  );


  and
  g2199
  (
    n2106,
    n1697,
    n1586,
    n1617,
    n1587
  );


  xor
  g2200
  (
    n2286,
    n1714,
    n1635,
    n1789,
    n1621
  );


  or
  g2201
  (
    n2091,
    n2024,
    n1729,
    n2017,
    n1797
  );


  xor
  g2202
  (
    n2092,
    n1748,
    n1652,
    n1778,
    n1768
  );


  and
  g2203
  (
    n2210,
    n1609,
    n1654,
    n1596,
    n1710
  );


  or
  g2204
  (
    n2074,
    n1598,
    n2000,
    n1716,
    n1559
  );


  nor
  g2205
  (
    n2191,
    n1566,
    n1996,
    n1992,
    n1574
  );


  and
  g2206
  (
    n2057,
    n2022,
    n1765,
    n1754,
    n1599
  );


  nand
  g2207
  (
    n2373,
    n1678,
    n1662,
    n1622,
    n1589
  );


  nand
  g2208
  (
    n2110,
    n1690,
    n2006,
    n1760,
    n1601
  );


  and
  g2209
  (
    n2371,
    n1799,
    n1680,
    n1754,
    n2021
  );


  xor
  g2210
  (
    n2075,
    n1571,
    n1583,
    n1783,
    n1652
  );


  and
  g2211
  (
    n2158,
    n1688,
    n2035,
    n2005,
    n2015
  );


  xnor
  g2212
  (
    n2076,
    n1622,
    n1795,
    n1708,
    n1734
  );


  nor
  g2213
  (
    n2055,
    n1674,
    n1988,
    n1579,
    n1760
  );


  xnor
  g2214
  (
    n2276,
    n1780,
    n1978,
    n1566,
    n1995
  );


  xor
  g2215
  (
    n2226,
    n1653,
    n2000,
    n1675,
    n1772
  );


  or
  g2216
  (
    n2155,
    n2045,
    n1616,
    n1750,
    n2046
  );


  or
  g2217
  (
    n2138,
    n1614,
    n1605,
    n1738,
    n1726
  );


  nor
  g2218
  (
    n2197,
    n1663,
    n1712,
    n2031,
    n1610
  );


  and
  g2219
  (
    n2298,
    n1691,
    n1660,
    n1742,
    n1639
  );


  nor
  g2220
  (
    n2115,
    n1677,
    n1998,
    n1755,
    n1695
  );


  nor
  g2221
  (
    n2254,
    n1723,
    n1580,
    n1601,
    n1791
  );


  xnor
  g2222
  (
    n2163,
    n1719,
    n2027,
    n1639,
    n1656
  );


  xnor
  g2223
  (
    n2134,
    n1741,
    n1659,
    n1746,
    n1779
  );


  xnor
  g2224
  (
    n2245,
    n1793,
    n1631,
    n1657,
    n1772
  );


  xnor
  g2225
  (
    n2360,
    n1721,
    n1800,
    n2035,
    n1660
  );


  xor
  g2226
  (
    n2369,
    n1730,
    n1590,
    n1794,
    n1650
  );


  and
  g2227
  (
    n2137,
    n1768,
    n2040,
    n1723,
    n1732
  );


  xor
  g2228
  (
    n2067,
    n1591,
    n1618,
    n1981,
    n1977
  );


  xnor
  g2229
  (
    n2257,
    n1740,
    n1766,
    n1612,
    n1575
  );


  or
  g2230
  (
    n2290,
    n2038,
    n1693,
    n1718,
    n1747
  );


  xnor
  g2231
  (
    n2275,
    n1690,
    n1716,
    n2043,
    n1728
  );


  xor
  g2232
  (
    n2062,
    n1761,
    n1742,
    n1600,
    n1624
  );


  xor
  g2233
  (
    n2350,
    n1760,
    n1745,
    n2041,
    n1655
  );


  nor
  g2234
  (
    n2157,
    n1649,
    n2036,
    n1658,
    n1612
  );


  nand
  g2235
  (
    n2325,
    n1763,
    n1693,
    n1983,
    n1646
  );


  nand
  g2236
  (
    KeyWire_0_47,
    n1774,
    n1619,
    n1647,
    n2033
  );


  xnor
  g2237
  (
    n2088,
    n1678,
    n2008,
    n1655,
    n1597
  );


  and
  g2238
  (
    n2136,
    n1663,
    n1632,
    n1597,
    n2049
  );


  or
  g2239
  (
    n2212,
    n2040,
    n1803,
    n1775,
    n2044
  );


  xnor
  g2240
  (
    n2264,
    n1715,
    n1742,
    n2016,
    n1639
  );


  xor
  g2241
  (
    n2102,
    n1804,
    n1615,
    n1619,
    n1623
  );


  xnor
  g2242
  (
    n2216,
    n1777,
    n1714,
    n1643,
    n2026
  );


  nor
  g2243
  (
    n2205,
    n2025,
    n1570,
    n1759,
    n2029
  );


  xnor
  g2244
  (
    n2272,
    n1731,
    n1743,
    n1608,
    n1704
  );


  or
  g2245
  (
    n2078,
    n1650,
    n2029,
    n1769,
    n1728
  );


  nand
  g2246
  (
    n2124,
    n2035,
    n1612,
    n1685,
    n1701
  );


  and
  g2247
  (
    n2284,
    n1710,
    n1603,
    n2023,
    n1618
  );


  and
  g2248
  (
    n2321,
    n1698,
    n1707,
    n1763,
    n1982
  );


  and
  g2249
  (
    n2181,
    n1704,
    n1719,
    n1680,
    n1702
  );


  or
  g2250
  (
    n2229,
    n1570,
    n1779,
    n1613,
    n1611
  );


  nand
  g2251
  (
    n2061,
    n2010,
    n1762,
    n1573,
    n2029
  );


  nor
  g2252
  (
    n2217,
    n1642,
    n1567,
    n1711,
    n2028
  );


  xor
  g2253
  (
    n2331,
    n1748,
    n1694,
    n1671,
    n1771
  );


  nor
  g2254
  (
    n2169,
    n1757,
    n1585,
    n1682,
    n2034
  );


  nor
  g2255
  (
    n2180,
    n1724,
    n1692,
    n1761,
    n2048
  );


  xor
  g2256
  (
    KeyWire_0_20,
    n1653,
    n1672,
    n1647,
    n1670
  );


  and
  g2257
  (
    n2100,
    n2053,
    n1802,
    n1670,
    n1759
  );


  or
  g2258
  (
    n2297,
    n2033,
    n2047,
    n1712,
    n1665
  );


  xor
  g2259
  (
    n2071,
    n1580,
    n1995,
    n2015,
    n1616
  );


  or
  g2260
  (
    n2117,
    n1985,
    n2037,
    n1692,
    n1735
  );


  or
  g2261
  (
    n2172,
    n2038,
    n1703,
    n2031,
    n1789
  );


  or
  g2262
  (
    n2339,
    n1720,
    n1767,
    n1975,
    n2017
  );


  or
  g2263
  (
    n2238,
    n2007,
    n1726,
    n1643,
    n1729
  );


  and
  g2264
  (
    n2265,
    n1700,
    n1798,
    n1796,
    n1989
  );


  xor
  g2265
  (
    n2335,
    n1728,
    n1624,
    n1761,
    n1724
  );


  nor
  g2266
  (
    n2240,
    n1577,
    n1614,
    n2045,
    n1788
  );


  xnor
  g2267
  (
    KeyWire_0_26,
    n1579,
    n2038,
    n2054,
    n1769
  );


  nand
  g2268
  (
    n2196,
    n1621,
    n1976,
    n1750,
    n1679
  );


  xnor
  g2269
  (
    n2167,
    n1581,
    n2052,
    n1667,
    n1569
  );


  nand
  g2270
  (
    n2198,
    n2037,
    n1732,
    n1801,
    n1800
  );


  nand
  g2271
  (
    n2328,
    n1661,
    n1647,
    n1776,
    n1658
  );


  nor
  g2272
  (
    n2145,
    n1699,
    n1803,
    n1614,
    n1593
  );


  xnor
  g2273
  (
    n2270,
    n1701,
    n1794,
    n1804,
    n2012
  );


  and
  g2274
  (
    n2129,
    n1656,
    n1625,
    n1757,
    n1991
  );


  and
  g2275
  (
    n2317,
    n2034,
    n2018,
    n1733,
    n1757
  );


  nor
  g2276
  (
    n2361,
    n1707,
    n2054,
    n1604,
    n1600
  );


  nand
  g2277
  (
    n2184,
    n1573,
    n1975,
    n1737,
    n1603
  );


  nand
  g2278
  (
    n2316,
    n1677,
    n1982,
    n1987,
    n1745
  );


  or
  g2279
  (
    n2302,
    n1792,
    n1716,
    n1730,
    n1595
  );


  or
  g2280
  (
    n2334,
    n1626,
    n1697,
    n1668,
    n2043
  );


  and
  g2281
  (
    n2215,
    n1619,
    n1685,
    n1584,
    n1704
  );


  and
  g2282
  (
    n2185,
    n2051,
    n1760,
    n1580,
    n2039
  );


  xor
  g2283
  (
    n2192,
    n1702,
    n1758,
    n1627,
    n1747
  );


  and
  g2284
  (
    n2241,
    n1998,
    n1721,
    n1715,
    n1671
  );


  and
  g2285
  (
    n2128,
    n1615,
    n1756,
    n1678,
    n1586
  );


  nand
  g2286
  (
    n2165,
    n1779,
    n1747,
    n1638,
    n1768
  );


  or
  g2287
  (
    n2348,
    n1681,
    n1689,
    n1996,
    n1992
  );


  nor
  g2288
  (
    n2326,
    n2003,
    n2029,
    n1791,
    n1579
  );


  or
  g2289
  (
    n2144,
    n1594,
    n1654,
    n2018,
    n1626
  );


  xor
  g2290
  (
    n2232,
    n1786,
    n1766,
    n1686,
    n1709
  );


  xor
  g2291
  (
    n2131,
    n1691,
    n1993,
    n1778,
    n1983
  );


  xnor
  g2292
  (
    n2080,
    n1736,
    n1994,
    n1637,
    n2014
  );


  nand
  g2293
  (
    n2084,
    n1742,
    n1751,
    n2032,
    n1783
  );


  xnor
  g2294
  (
    n2301,
    n1591,
    n1799,
    n1578,
    n2013
  );


  xnor
  g2295
  (
    n2206,
    n1613,
    n1695,
    n1605,
    n1720
  );


  nor
  g2296
  (
    n2060,
    n1630,
    n1670,
    n1679,
    n1714
  );


  xor
  g2297
  (
    n2222,
    n1654,
    n1992,
    n2042,
    n1702
  );


  or
  g2298
  (
    n2247,
    n1712,
    n2009,
    n1675,
    n1676
  );


  and
  g2299
  (
    n2204,
    n1764,
    n1582,
    n1755,
    n1593
  );


  nand
  g2300
  (
    KeyWire_0_45,
    n2021,
    n2030,
    n2023,
    n1635
  );


  xnor
  g2301
  (
    n2142,
    n1661,
    n1687,
    n1678,
    n1620
  );


  nor
  g2302
  (
    n2200,
    n1793,
    n1638,
    n1798,
    n1979
  );


  and
  g2303
  (
    n2324,
    n2016,
    n1669,
    n1676,
    n1637
  );


  nor
  g2304
  (
    n2123,
    n2051,
    n1689,
    n1718,
    n1719
  );


  nand
  g2305
  (
    KeyWire_0_42,
    n1598,
    n1729,
    n1722,
    n1764
  );


  xnor
  g2306
  (
    n2156,
    n1739,
    n1776,
    n1683,
    n1608
  );


  nand
  g2307
  (
    n2253,
    n1696,
    n1561,
    n1988,
    n2008
  );


  nand
  g2308
  (
    n2153,
    n1596,
    n1664,
    n1806,
    n1652
  );


  xnor
  g2309
  (
    n2081,
    n1655,
    n1785,
    n1568,
    n1611
  );


  xor
  g2310
  (
    KeyWire_0_15,
    n2013,
    n1743,
    n1658,
    n1666
  );


  and
  g2311
  (
    n2279,
    n1598,
    n1572,
    n2051,
    n2047
  );


  nor
  g2312
  (
    n2236,
    n1714,
    n1575,
    n2013,
    n1725
  );


  nor
  g2313
  (
    n2349,
    n2010,
    n1733,
    n2046,
    n1774
  );


  nand
  g2314
  (
    n2268,
    n1797,
    n1669,
    n1618,
    n2048
  );


  xor
  g2315
  (
    n2235,
    n1683,
    n1722,
    n2028,
    n1734
  );


  or
  g2316
  (
    n2230,
    n1978,
    n1802,
    n1773,
    n1653
  );


  and
  g2317
  (
    n2188,
    n1615,
    n1736,
    n1978,
    n1767
  );


  xnor
  g2318
  (
    n2108,
    n1648,
    n2001,
    n1650,
    n1739
  );


  or
  g2319
  (
    n2107,
    n1628,
    n1636,
    n1752,
    n2014
  );


  xor
  g2320
  (
    n2281,
    n1596,
    n1778,
    n2014,
    n1763
  );


  xor
  g2321
  (
    n2098,
    n1795,
    n1688,
    n1592,
    n1633
  );


  xnor
  g2322
  (
    n2090,
    n1599,
    n1788,
    n1751,
    n1588
  );


  nand
  g2323
  (
    n2364,
    n1783,
    n1664,
    n1765,
    n1582
  );


  nor
  g2324
  (
    n2288,
    n1682,
    n1602,
    n1687,
    n2041
  );


  and
  g2325
  (
    n2133,
    n1743,
    n1719,
    n1986,
    n1677
  );


  or
  g2326
  (
    n2118,
    n1576,
    n2005,
    n1735,
    n1680
  );


  nand
  g2327
  (
    n2093,
    n1674,
    n1985,
    n1771,
    n1680
  );


  xor
  g2328
  (
    n2101,
    n1754,
    n1604,
    n1989,
    n1786
  );


  xnor
  g2329
  (
    n2318,
    n1696,
    n1627,
    n2003,
    n1770
  );


  xor
  g2330
  (
    n2139,
    n1740,
    n1696,
    n1620,
    n1628
  );


  xor
  g2331
  (
    n2066,
    n2043,
    n1729,
    n1583,
    n1659
  );


  xor
  g2332
  (
    n2234,
    n2044,
    n1625,
    n1693,
    n1803
  );


  xor
  g2333
  (
    n2260,
    n1785,
    n2048,
    n1649,
    n1998
  );


  nor
  g2334
  (
    n2283,
    n1986,
    n1630,
    n1727,
    n1720
  );


  and
  g2335
  (
    n2127,
    n1708,
    n1787,
    n1634,
    n1774
  );


  nand
  g2336
  (
    n2287,
    n1612,
    n1980,
    n1622,
    n1589
  );


  nor
  g2337
  (
    n2374,
    n2007,
    n1660,
    n1713,
    n1637
  );


  nor
  g2338
  (
    n2140,
    n1606,
    n1642,
    n1641,
    n1702
  );


  nor
  g2339
  (
    n2161,
    n1657,
    n1636,
    n1627,
    n1981
  );


  or
  g2340
  (
    n2278,
    n1982,
    n1805,
    n1677,
    n1703
  );


  or
  g2341
  (
    n2141,
    n1984,
    n1654,
    n1749,
    n1631
  );


  and
  g2342
  (
    n2322,
    n1980,
    n1595,
    n2010,
    n2012
  );


  nand
  g2343
  (
    n2365,
    n1801,
    n1697,
    n1595,
    n1669
  );


  nor
  g2344
  (
    n2113,
    n1588,
    n1638,
    n1694,
    n1657
  );


  xor
  g2345
  (
    n2343,
    n1723,
    n1735,
    n1623,
    n1993
  );


  and
  g2346
  (
    n2132,
    n1661,
    n1611,
    n1562,
    n1600
  );


  xnor
  g2347
  (
    n2083,
    n1796,
    n1793,
    n1703,
    n1786
  );


  or
  g2348
  (
    n2499,
    n2307,
    n2123,
    n2284,
    n2357
  );


  and
  g2349
  (
    n2414,
    n2354,
    n2199,
    n2125,
    n2351
  );


  and
  g2350
  (
    n2426,
    n2335,
    n2339,
    n2169,
    n2267
  );


  and
  g2351
  (
    n2584,
    n2290,
    n2360,
    n2192,
    n2109
  );


  and
  g2352
  (
    n2506,
    n2315,
    n2187,
    n2321,
    n2133
  );


  or
  g2353
  (
    n2585,
    n2079,
    n2167,
    n2297,
    n2368
  );


  xnor
  g2354
  (
    n2539,
    n2158,
    n2369,
    n2348,
    n2344
  );


  nand
  g2355
  (
    n2487,
    n2168,
    n26,
    n2344,
    n2193
  );


  xnor
  g2356
  (
    n2516,
    n2103,
    n2345,
    n2246,
    n2362
  );


  nand
  g2357
  (
    n2489,
    n2303,
    n2248,
    n2113,
    n2070
  );


  nand
  g2358
  (
    n2559,
    n2276,
    n2371,
    n2296,
    n2352
  );


  xnor
  g2359
  (
    n2511,
    n2217,
    n2370,
    n2145,
    n2281
  );


  nor
  g2360
  (
    n2530,
    n2116,
    n2299,
    n2164,
    n2349
  );


  nor
  g2361
  (
    n2532,
    n2221,
    n2130,
    n2085,
    n2280
  );


  nand
  g2362
  (
    n2382,
    n2196,
    n2279,
    n2300,
    n2075
  );


  nor
  g2363
  (
    n2454,
    n2273,
    n2342,
    n2337,
    n2132
  );


  nor
  g2364
  (
    n2500,
    n2302,
    n2262,
    n2367,
    n2366
  );


  xnor
  g2365
  (
    n2450,
    n2231,
    n2117,
    n2141,
    n2223
  );


  and
  g2366
  (
    n2550,
    n2363,
    n2120,
    n2293,
    n2282
  );


  or
  g2367
  (
    n2419,
    n2250,
    n2194,
    n2153,
    n2112
  );


  and
  g2368
  (
    n2518,
    n2277,
    n2233,
    n1806,
    n2349
  );


  nor
  g2369
  (
    n2557,
    n2316,
    n2284,
    n2308,
    n2217
  );


  nor
  g2370
  (
    n2411,
    n2231,
    n2246,
    n2292,
    n2163
  );


  and
  g2371
  (
    n2482,
    n2287,
    n2132,
    n2358,
    n2273
  );


  and
  g2372
  (
    n2400,
    n2369,
    n2118,
    n2144,
    n2082
  );


  and
  g2373
  (
    n2407,
    n2222,
    n2343,
    n2247,
    n26
  );


  or
  g2374
  (
    n2442,
    n2306,
    n2251,
    n2328,
    n2356
  );


  nor
  g2375
  (
    n2394,
    n2275,
    n2183,
    n2292,
    n2370
  );


  or
  g2376
  (
    n2387,
    n2166,
    n2290,
    n118,
    n2057
  );


  xor
  g2377
  (
    n2467,
    n2091,
    n2308,
    n2225,
    n2331
  );


  and
  g2378
  (
    n2441,
    n2135,
    n2154,
    n2361,
    n2370
  );


  or
  g2379
  (
    n2455,
    n2215,
    n2342,
    n2241,
    n2238
  );


  xnor
  g2380
  (
    n2383,
    n2092,
    n2314,
    n2359,
    n2357
  );


  nor
  g2381
  (
    n2527,
    n2318,
    n2353,
    n2090,
    n2365
  );


  nand
  g2382
  (
    n2390,
    n2245,
    n2314,
    n2283,
    n2348
  );


  nor
  g2383
  (
    n2471,
    n2159,
    n2333,
    n2234,
    n2367
  );


  nand
  g2384
  (
    n2401,
    n2373,
    n2098,
    n2288,
    n2238
  );


  nand
  g2385
  (
    n2582,
    n2323,
    n2285,
    n2278,
    n2331
  );


  or
  g2386
  (
    n2542,
    n2165,
    n2269,
    n2297,
    n2328
  );


  and
  g2387
  (
    n2447,
    n2269,
    n2311,
    n2374,
    n2299
  );


  nor
  g2388
  (
    n2586,
    n2336,
    n2334,
    n2076,
    n2322
  );


  nor
  g2389
  (
    n2449,
    n2223,
    n2373,
    n2266,
    n2099
  );


  xnor
  g2390
  (
    n2592,
    n2311,
    n2122,
    n2358,
    n2298
  );


  nand
  g2391
  (
    n2521,
    n2198,
    n2334,
    n2174,
    n2063
  );


  xor
  g2392
  (
    n2463,
    n2355,
    n2118,
    n2264,
    n2347
  );


  xnor
  g2393
  (
    n2476,
    n2142,
    n2321,
    n2359,
    n2312
  );


  xor
  g2394
  (
    n2552,
    n2279,
    n2293,
    n2266,
    n2106
  );


  and
  g2395
  (
    n2497,
    n2111,
    n2207,
    n2344,
    n2358
  );


  nand
  g2396
  (
    n2398,
    n2156,
    n2303,
    n2326,
    n2374
  );


  and
  g2397
  (
    n2510,
    n2304,
    n2333,
    n2259,
    n2088
  );


  or
  g2398
  (
    n2503,
    n2280,
    n2371,
    n2267,
    n2285
  );


  nor
  g2399
  (
    KeyWire_0_58,
    n2268,
    n2268,
    n2308,
    n2265
  );


  nand
  g2400
  (
    n2474,
    n2272,
    n2178,
    n2240,
    n2168
  );


  or
  g2401
  (
    n2464,
    n2188,
    n2137,
    n2212,
    n2312
  );


  xnor
  g2402
  (
    n2409,
    n2283,
    n2332,
    n2312
  );


  xor
  g2403
  (
    n2547,
    n2286,
    n2319,
    n2341,
    n2073
  );


  xor
  g2404
  (
    n2457,
    n2286,
    n2229,
    n2349,
    n2086
  );


  nor
  g2405
  (
    n2458,
    n2346,
    n2319,
    n2314,
    n2355
  );


  and
  g2406
  (
    n2579,
    n2260,
    n2363,
    n2092,
    n2275
  );


  or
  g2407
  (
    n2393,
    n2288,
    n2360,
    n2268,
    n2245
  );


  xor
  g2408
  (
    n2576,
    n2371,
    n2078,
    n2081,
    n2067
  );


  nand
  g2409
  (
    n2490,
    n2242,
    n2096,
    n2307,
    n2249
  );


  and
  g2410
  (
    n2477,
    n2083,
    n2214,
    n2172,
    n2066
  );


  nand
  g2411
  (
    KeyWire_0_59,
    n2251,
    n2158,
    n2127,
    n2327
  );


  nor
  g2412
  (
    n2508,
    n2345,
    n2346,
    n2253,
    n2279
  );


  nand
  g2413
  (
    n2375,
    n2101,
    n2310,
    n2096,
    n2151
  );


  or
  g2414
  (
    n2438,
    n2373,
    n2327,
    n2349,
    n2278
  );


  and
  g2415
  (
    KeyWire_0_37,
    n2366,
    n2290,
    n2300,
    n2156
  );


  xor
  g2416
  (
    n2488,
    n2325,
    n2317,
    n26,
    n2374
  );


  xor
  g2417
  (
    n2406,
    n2105,
    n2150,
    n2311,
    n2318
  );


  nand
  g2418
  (
    n2502,
    n2294,
    n2263,
    n2165,
    n2093
  );


  nor
  g2419
  (
    n2572,
    n2291,
    n2220,
    n2080,
    n2279
  );


  nand
  g2420
  (
    n2556,
    n2095,
    n2093,
    n2182,
    n2315
  );


  and
  g2421
  (
    n2415,
    n2301,
    n2195,
    n2330,
    n2071
  );


  and
  g2422
  (
    n2563,
    n2147,
    n2176,
    n2350,
    n2099
  );


  nand
  g2423
  (
    n2445,
    n2285,
    n2182,
    n2298,
    n2155
  );


  xor
  g2424
  (
    n2595,
    n2146,
    n2259,
    n2124,
    n2324
  );


  nand
  g2425
  (
    n2405,
    n2250,
    n2200,
    n2285,
    n2301
  );


  or
  g2426
  (
    n2468,
    n2360,
    n2347,
    n2324,
    n2256
  );


  nor
  g2427
  (
    n2587,
    n2288,
    n2235,
    n2278,
    n2329
  );


  and
  g2428
  (
    n2523,
    n2362,
    n2225,
    n2313,
    n2261
  );


  xnor
  g2429
  (
    n2562,
    n2271,
    n2304,
    n2249,
    n2367
  );


  xnor
  g2430
  (
    n2492,
    n2193,
    n2345,
    n2318,
    n2262
  );


  nor
  g2431
  (
    n2388,
    n2210,
    n2323,
    n2216,
    n2140
  );


  nor
  g2432
  (
    n2420,
    n2289,
    n2261,
    n2243,
    n2102
  );


  nor
  g2433
  (
    n2531,
    n2330,
    n2148,
    n2192,
    n2202
  );


  and
  g2434
  (
    n2514,
    n2195,
    n2112,
    n2125,
    n2166
  );


  and
  g2435
  (
    n2470,
    n2198,
    n2336,
    n2322,
    n2265
  );


  nand
  g2436
  (
    n2491,
    n2061,
    n2167,
    n2339,
    n2179
  );


  xnor
  g2437
  (
    n2408,
    n2346,
    n2128,
    n2257,
    n2064
  );


  nand
  g2438
  (
    n2486,
    n2084,
    n2219,
    n2316,
    n2272
  );


  xnor
  g2439
  (
    n2386,
    n2151,
    n2184,
    n2147,
    n2292
  );


  xnor
  g2440
  (
    n2428,
    n2065,
    n2320,
    n2180,
    n2269
  );


  or
  g2441
  (
    n2432,
    n2110,
    n2162,
    n2342,
    n2244
  );


  xnor
  g2442
  (
    n2573,
    n2140,
    n2353,
    n2074,
    n2244
  );


  nor
  g2443
  (
    n2403,
    n2270,
    n2350,
    n2100,
    n2219
  );


  xor
  g2444
  (
    n2484,
    n2138,
    n2338,
    n2227,
    n2061
  );


  and
  g2445
  (
    n2448,
    n2131,
    n2191,
    n2333,
    n2309
  );


  nor
  g2446
  (
    n2541,
    n2272,
    n2203,
    n2320,
    n2236
  );


  nor
  g2447
  (
    n2574,
    n2135,
    n2243,
    n2103,
    n2319
  );


  nor
  g2448
  (
    n2493,
    n2201,
    n2282,
    n2373,
    n2355
  );


  and
  g2449
  (
    n2588,
    n2282,
    n2351,
    n2055,
    n2089
  );


  nor
  g2450
  (
    n2427,
    n2056,
    n2364,
    n2309,
    n2293
  );


  xnor
  g2451
  (
    n2568,
    n2161,
    n2359,
    n2186,
    n2076
  );


  nand
  g2452
  (
    n2554,
    n2073,
    n2324,
    n2173,
    n2175
  );


  nand
  g2453
  (
    n2412,
    n2296,
    n2063,
    n2197,
    n2233
  );


  xor
  g2454
  (
    n2564,
    n2320,
    n2097,
    n2331,
    n2308
  );


  and
  g2455
  (
    n2569,
    n2316,
    n2083,
    n2337,
    n2263
  );


  nor
  g2456
  (
    n2551,
    n2304,
    n2365,
    n2300,
    n2211
  );


  nor
  g2457
  (
    n2480,
    n2085,
    n2109,
    n2264,
    n2139
  );


  and
  g2458
  (
    n2446,
    n2062,
    n2354,
    n2077,
    n2106
  );


  and
  g2459
  (
    n2593,
    n2281,
    n2149,
    n2097,
    n2143
  );


  xor
  g2460
  (
    n2513,
    n2129,
    n2312,
    n2257,
    n2253
  );


  and
  g2461
  (
    n2379,
    n2327,
    n2181,
    n2313,
    n2228
  );


  nand
  g2462
  (
    n2560,
    n2372,
    n2184,
    n117,
    n2295
  );


  nand
  g2463
  (
    n2377,
    n2254,
    n2107,
    n2267,
    n26
  );


  xnor
  g2464
  (
    n2496,
    n2256,
    n2298,
    n2154,
    n25
  );


  xnor
  g2465
  (
    n2591,
    n2159,
    n2153,
    n2364,
    n2072
  );


  nor
  g2466
  (
    n2429,
    n2368,
    n2260,
    n2095,
    n2065
  );


  xnor
  g2467
  (
    n2501,
    n2321,
    n2352,
    n2280,
    n2296
  );


  xnor
  g2468
  (
    n2596,
    n2368,
    n25,
    n2330,
    n2255
  );


  xnor
  g2469
  (
    n2567,
    n2177,
    n2203,
    n2296,
    n2286
  );


  nand
  g2470
  (
    n2529,
    n2241,
    n25,
    n2293,
    n2059
  );


  xnor
  g2471
  (
    n2418,
    n2336,
    n2077,
    n2113,
    n117
  );


  xnor
  g2472
  (
    n2395,
    n2190,
    n2196,
    n2098,
    n2262
  );


  or
  g2473
  (
    n2473,
    n2286,
    n2080,
    n2155,
    n2262
  );


  and
  g2474
  (
    n2431,
    n2273,
    n2127,
    n2347,
    n2356
  );


  or
  g2475
  (
    n2504,
    n2359,
    n2372,
    n2171,
    n2353
  );


  or
  g2476
  (
    n2456,
    n2338,
    n2297,
    n2101,
    n2211
  );


  nor
  g2477
  (
    n2570,
    n2229,
    n2365,
    n2100,
    n2372
  );


  xor
  g2478
  (
    n2453,
    n2144,
    n2091,
    n2289,
    n2288
  );


  nand
  g2479
  (
    n2440,
    n2248,
    n2175,
    n2367,
    n2315
  );


  and
  g2480
  (
    n2481,
    n2163,
    n2066,
    n2294,
    n2354
  );


  xnor
  g2481
  (
    n2545,
    n2309,
    n2104,
    n2222,
    n2228
  );


  and
  g2482
  (
    n2433,
    n2268,
    n2357,
    n2302,
    n2139
  );


  or
  g2483
  (
    n2577,
    n2289,
    n2289,
    n2117,
    n2197
  );


  nor
  g2484
  (
    n2452,
    n2277,
    n2340,
    n2209,
    n2087
  );


  xnor
  g2485
  (
    n2590,
    n2275,
    n2074,
    n2346,
    n2089
  );


  and
  g2486
  (
    n2392,
    n2317,
    n2341,
    n2305,
    n118
  );


  xor
  g2487
  (
    KeyWire_0_1,
    n2291,
    n2152,
    n2102,
    n2301
  );


  xnor
  g2488
  (
    n2543,
    n2176,
    n2278,
    n2205,
    n2081
  );


  xnor
  g2489
  (
    n2528,
    n2075,
    n1806,
    n2187,
    n2227
  );


  xor
  g2490
  (
    n2540,
    n2208,
    n2291,
    n2295,
    n2274
  );


  or
  g2491
  (
    KeyWire_0_19,
    n2321,
    n2255,
    n2120,
    n2298
  );


  xor
  g2492
  (
    n2466,
    n2269,
    n2301,
    n2364,
    n2305
  );


  nor
  g2493
  (
    n2397,
    n2072,
    n2141,
    n2194,
    n2306
  );


  xnor
  g2494
  (
    n2526,
    n2145,
    n2361,
    n2055,
    n2311
  );


  xor
  g2495
  (
    n2469,
    n2084,
    n2208,
    n2116,
    n118
  );


  xnor
  g2496
  (
    n2378,
    n2304,
    n2291,
    n2287,
    n2206
  );


  xor
  g2497
  (
    n2561,
    n2318,
    n2283,
    n2371,
    n2355
  );


  nor
  g2498
  (
    n2451,
    n2338,
    n2230,
    n2133,
    n2287
  );


  xnor
  g2499
  (
    n2384,
    n2274,
    n2328,
    n2221,
    n2218
  );


  nor
  g2500
  (
    n2413,
    n2322,
    n1806,
    n2351,
    n2235
  );


  nand
  g2501
  (
    n2424,
    n2272,
    n2363,
    n2366,
    n2332
  );


  nand
  g2502
  (
    n2434,
    n2071,
    n2068,
    n2079,
    n2258
  );


  and
  g2503
  (
    n2461,
    n2058,
    n2340,
    n2237,
    n2110
  );


  or
  g2504
  (
    n2444,
    n2108,
    n2212,
    n2276,
    n2216
  );


  nand
  g2505
  (
    n2422,
    n2240,
    n2325,
    n2340,
    n2281
  );


  xor
  g2506
  (
    n2525,
    n2171,
    n2361,
    n2310,
    n2354
  );


  or
  g2507
  (
    n2380,
    n2356,
    n2224,
    n2057,
    n2258
  );


  xor
  g2508
  (
    n2479,
    n2134,
    n2340,
    n2111,
    n2191
  );


  nand
  g2509
  (
    n2421,
    n2173,
    n2339,
    n2114,
    n2108
  );


  xor
  g2510
  (
    n2583,
    n2115,
    n2341,
    n2070,
    n24
  );


  or
  g2511
  (
    n2460,
    n2126,
    n2148,
    n2366,
    n2236
  );


  and
  g2512
  (
    n2410,
    n2343,
    n2335,
    n2334,
    n2157
  );


  and
  g2513
  (
    n2381,
    n2201,
    n2267,
    n2274,
    n2213
  );


  nand
  g2514
  (
    n2565,
    n2252,
    n2160,
    n2368,
    n2310
  );


  and
  g2515
  (
    n2495,
    n2232,
    n2315,
    n2290,
    n2088
  );


  or
  g2516
  (
    KeyWire_0_46,
    n2190,
    n2164,
    n2337,
    n2305
  );


  nor
  g2517
  (
    n2430,
    n2239,
    n2129,
    n24,
    n2169
  );


  nor
  g2518
  (
    n2515,
    n2107,
    n2360,
    n2121,
    n2185
  );


  and
  g2519
  (
    n2512,
    n2363,
    n2270,
    n2143,
    n2094
  );


  xnor
  g2520
  (
    n2578,
    n2300,
    n2326,
    n2142,
    n2275
  );


  nand
  g2521
  (
    n2555,
    n2185,
    n2336,
    n2317,
    n2162
  );


  nor
  g2522
  (
    n2391,
    n2183,
    n2369,
    n2138,
    n2206
  );


  or
  g2523
  (
    n2553,
    n2350,
    n2094,
    n2302,
    n2294
  );


  nand
  g2524
  (
    n2571,
    n2161,
    n2352,
    n2131,
    n2218
  );


  nand
  g2525
  (
    n2580,
    n2320,
    n2329,
    n2263,
    n2330
  );


  xnor
  g2526
  (
    n2399,
    n2266,
    n2207,
    n2306,
    n2357
  );


  xor
  g2527
  (
    n2396,
    n2362,
    n2149,
    n2214,
    n2264
  );


  xor
  g2528
  (
    n2475,
    n2263,
    n2090,
    n2265,
    n2264
  );


  nand
  g2529
  (
    n2498,
    n2329,
    n2348,
    n2130,
    n2332
  );


  or
  g2530
  (
    n2483,
    n2351,
    n2281,
    n2220,
    n2306
  );


  or
  g2531
  (
    n2459,
    n2343,
    n2180,
    n2280,
    n2239
  );


  or
  g2532
  (
    n2425,
    n2358,
    n2242,
    n2345,
    n2104
  );


  nand
  g2533
  (
    n2566,
    n2316,
    n2294,
    n2331,
    n2334
  );


  nor
  g2534
  (
    n2537,
    n2128,
    n2067,
    n2189,
    n2271
  );


  and
  g2535
  (
    n2416,
    n2210,
    n2078,
    n2209,
    n2252
  );


  or
  g2536
  (
    n2548,
    n24,
    n2232,
    n2115,
    n2364
  );


  nor
  g2537
  (
    n2594,
    n2314,
    n2297,
    n2317,
    n2369
  );


  nand
  g2538
  (
    n2538,
    n2299,
    n2350,
    n2284,
    n2170
  );


  xor
  g2539
  (
    n2485,
    n2177,
    n2137,
    n2344,
    n118
  );


  and
  g2540
  (
    n2376,
    n2056,
    n2200,
    n2295,
    n2347
  );


  xor
  g2541
  (
    n2544,
    n2205,
    n2266,
    n24,
    n2337
  );


  nand
  g2542
  (
    n2423,
    n2189,
    n2188,
    n2058,
    n2356
  );


  nand
  g2543
  (
    n2505,
    n2069,
    n2069,
    n2122,
    n117
  );


  or
  g2544
  (
    n2546,
    n2307,
    n2305,
    n2309,
    n2325
  );


  and
  g2545
  (
    n2520,
    n2339,
    n25,
    n2059,
    n2276
  );


  and
  g2546
  (
    n2435,
    n2202,
    n2295,
    n2303,
    n2179
  );


  nand
  g2547
  (
    n2402,
    n2157,
    n2365,
    n2325,
    n2299
  );


  nand
  g2548
  (
    n2437,
    n2247,
    n2215,
    n2124,
    n2064
  );


  nor
  g2549
  (
    n2524,
    n2302,
    n2068,
    n2276,
    n2282
  );


  nor
  g2550
  (
    n2478,
    n2270,
    n2174,
    n2341,
    n2119
  );


  or
  g2551
  (
    n2507,
    n2086,
    n2060,
    n2136,
    n2292
  );


  xor
  g2552
  (
    n2581,
    n2082,
    n2352,
    n2274,
    n2323
  );


  xnor
  g2553
  (
    n2522,
    n2333,
    n2372,
    n2307,
    n2327
  );


  nand
  g2554
  (
    n2534,
    n2277,
    n2172,
    n2126,
    n2310
  );


  nor
  g2555
  (
    n2385,
    n2199,
    n2362,
    n2335,
    n2178
  );


  and
  g2556
  (
    n2417,
    n2313,
    n2342,
    n2230,
    n2270
  );


  and
  g2557
  (
    n2535,
    n2303,
    n2114,
    n2060,
    n2273
  );


  or
  g2558
  (
    n2439,
    n2136,
    n2226,
    n2234,
    n2152
  );


  nor
  g2559
  (
    n2472,
    n2277,
    n2123,
    n2271,
    n2265
  );


  xnor
  g2560
  (
    n2519,
    n2324,
    n2313,
    n2237,
    n2181
  );


  or
  g2561
  (
    n2436,
    n2121,
    n2328,
    n2119,
    n2150
  );


  or
  g2562
  (
    n2494,
    n2224,
    n2319,
    n2254,
    n2283
  );


  xor
  g2563
  (
    n2549,
    n2335,
    n2226,
    n2062,
    n2213
  );


  xor
  g2564
  (
    n2443,
    n2326,
    n2323,
    n2146,
    n2134
  );


  xor
  g2565
  (
    n2536,
    n2348,
    n2204,
    n2361,
    n2287
  );


  xor
  g2566
  (
    n2589,
    n2322,
    n2284,
    n2326,
    n2374
  );


  xnor
  g2567
  (
    n2465,
    n2186,
    n2353,
    n2087,
    n2343
  );


  xor
  g2568
  (
    n2509,
    n2204,
    n2105,
    n2329,
    n2370
  );


  and
  g2569
  (
    n2533,
    n2170,
    n2271,
    n2338,
    n2160
  );


  nand
  g2570
  (
    n2622,
    n2410,
    n2484,
    n2465,
    n2546
  );


  and
  g2571
  (
    n2617,
    n2541,
    n2488,
    n2469,
    n2550
  );


  nand
  g2572
  (
    n2597,
    n2522,
    n2487,
    n2376,
    n2488
  );


  nand
  g2573
  (
    n2670,
    n2425,
    n2512,
    n2504,
    n2513
  );


  and
  g2574
  (
    n2642,
    n2584,
    n2494,
    n2515,
    n2567
  );


  xor
  g2575
  (
    n2652,
    n2572,
    n2562,
    n2472,
    n2478
  );


  and
  g2576
  (
    n2650,
    n2497,
    n2418,
    n2391,
    n2450
  );


  nor
  g2577
  (
    n2655,
    n2589,
    n2521,
    n2412,
    n2424
  );


  or
  g2578
  (
    n2613,
    n2579,
    n2455,
    n2575,
    n2459
  );


  xor
  g2579
  (
    n2623,
    n2551,
    n2386,
    n2545,
    n2511
  );


  nand
  g2580
  (
    n2657,
    n2502,
    n2451,
    n2547,
    n2398
  );


  xnor
  g2581
  (
    n2631,
    n2379,
    n2573,
    n2580,
    n2596
  );


  xnor
  g2582
  (
    n2614,
    n2542,
    n2452,
    n2399,
    n2409
  );


  nor
  g2583
  (
    n2665,
    n2477,
    n2416,
    n2485,
    n2435
  );


  and
  g2584
  (
    n2639,
    n2534,
    n2419,
    n2573,
    n2564
  );


  xnor
  g2585
  (
    n2608,
    n2458,
    n2524,
    n2434,
    n2537
  );


  nand
  g2586
  (
    n2680,
    n2548,
    n2540,
    n2387,
    n2556
  );


  xor
  g2587
  (
    n2618,
    n2403,
    n2490,
    n2591,
    n2421
  );


  xnor
  g2588
  (
    n2653,
    n2510,
    n2540,
    n2583,
    n2496
  );


  or
  g2589
  (
    n2647,
    n2578,
    n2500,
    n2462,
    n2547
  );


  or
  g2590
  (
    n2666,
    n2557,
    n2595,
    n2475,
    n2392
  );


  or
  g2591
  (
    n2605,
    n2588,
    n2548,
    n2491,
    n2571
  );


  nor
  g2592
  (
    n2633,
    n2440,
    n2480,
    n2476,
    n2554
  );


  xor
  g2593
  (
    n2643,
    n2569,
    n2567,
    n2447,
    n2430
  );


  xnor
  g2594
  (
    n2677,
    n2562,
    n2394,
    n2571,
    n2431
  );


  xor
  g2595
  (
    n2660,
    n2503,
    n2483,
    n2498,
    n2524
  );


  xor
  g2596
  (
    n2671,
    n2474,
    n2589,
    n2592,
    n2552
  );


  or
  g2597
  (
    n2616,
    n2570,
    n2555,
    n2530,
    n2526
  );


  or
  g2598
  (
    n2611,
    n2549,
    n2449,
    n2436,
    n2445
  );


  and
  g2599
  (
    n2646,
    n2574,
    n2413,
    n2499,
    n2507
  );


  nor
  g2600
  (
    n2676,
    n2563,
    n2587,
    n2532,
    n2560
  );


  and
  g2601
  (
    n2607,
    n2539,
    n2519,
    n2443,
    n2520
  );


  or
  g2602
  (
    n2598,
    n2534,
    n2522,
    n2481,
    n2494
  );


  xor
  g2603
  (
    n2662,
    n2565,
    n2518,
    n2508,
    n2545
  );


  nor
  g2604
  (
    n2672,
    n2543,
    n2583,
    n2414,
    n2595
  );


  or
  g2605
  (
    n2621,
    n2558,
    n2395,
    n2542,
    n2557
  );


  nand
  g2606
  (
    n2644,
    n2526,
    n2528,
    n2385,
    n2493
  );


  xnor
  g2607
  (
    n2599,
    n2384,
    n2565,
    n2487,
    n2553
  );


  nand
  g2608
  (
    n2636,
    n2561,
    n2579,
    n2486,
    n2439
  );


  xnor
  g2609
  (
    n2601,
    n2586,
    n2411,
    n2537,
    n2561
  );


  nor
  g2610
  (
    n2674,
    n2591,
    n2558,
    n2576,
    n2517
  );


  nor
  g2611
  (
    n2604,
    n2420,
    n2551,
    n2577,
    n2505
  );


  xor
  g2612
  (
    n2637,
    n2529,
    n2588,
    n2564,
    n2587
  );


  xor
  g2613
  (
    n2620,
    n2427,
    n2417,
    n2536,
    n2507
  );


  nand
  g2614
  (
    n2656,
    n2503,
    n2569,
    n2495,
    n2596
  );


  and
  g2615
  (
    n2659,
    n2492,
    n2501,
    n2377,
    n2592
  );


  nand
  g2616
  (
    n2628,
    n2433,
    n2489,
    n2514,
    n2584
  );


  nand
  g2617
  (
    n2669,
    n2553,
    n2559,
    n2593,
    n2543
  );


  xnor
  g2618
  (
    n2640,
    n2544,
    n2509,
    n2549,
    n2468
  );


  xnor
  g2619
  (
    n2615,
    n2461,
    n2544,
    n2502,
    n2532
  );


  nor
  g2620
  (
    n2641,
    n2375,
    n2536,
    n2446,
    n2457
  );


  xor
  g2621
  (
    n2658,
    n2438,
    n2501,
    n2516,
    n2566
  );


  nand
  g2622
  (
    n2609,
    n2552,
    n2460,
    n2590
  );


  nor
  g2623
  (
    n2625,
    n2415,
    n2531,
    n2484,
    n2577
  );


  or
  g2624
  (
    n2629,
    n2510,
    n2406,
    n2511,
    n2432
  );


  and
  g2625
  (
    n2663,
    n2466,
    n2594,
    n2422,
    n2533
  );


  xor
  g2626
  (
    n2626,
    n2383,
    n2525,
    n2550,
    n2504
  );


  xor
  g2627
  (
    n2634,
    n2560,
    n2400,
    n2470,
    n2581
  );


  nor
  g2628
  (
    n2675,
    n2528,
    n2527,
    n2498,
    n2508
  );


  nor
  g2629
  (
    n2600,
    n2378,
    n2444,
    n2541,
    n2388
  );


  xnor
  g2630
  (
    n2667,
    n2495,
    n2382,
    n2396,
    n2556
  );


  and
  g2631
  (
    KeyWire_0_41,
    n2491,
    n2380,
    n2402,
    n2485
  );


  xor
  g2632
  (
    n2651,
    n2521,
    n2585,
    n2529,
    n2453
  );


  or
  g2633
  (
    n2627,
    n2496,
    n2429,
    n2539,
    n2506
  );


  nand
  g2634
  (
    n2624,
    n2397,
    n2580,
    n2594,
    n2578
  );


  nor
  g2635
  (
    n2679,
    n2437,
    n2515,
    n2585,
    n2582
  );


  and
  g2636
  (
    n2602,
    n2581,
    n2497,
    n2486,
    n2519
  );


  or
  g2637
  (
    n2668,
    n2525,
    n2489,
    n2408,
    n2505
  );


  nor
  g2638
  (
    n2606,
    n2530,
    n2442,
    n2492,
    n2518
  );


  xnor
  g2639
  (
    n2603,
    n2593,
    n2517,
    n2514,
    n2574
  );


  xnor
  g2640
  (
    n2612,
    n2464,
    n2572,
    n2512,
    n2428
  );


  xnor
  g2641
  (
    n2630,
    n2389,
    n2576,
    n2523,
    n2506
  );


  nor
  g2642
  (
    n2661,
    n2559,
    n2554,
    n2483,
    n2538
  );


  xnor
  g2643
  (
    n2648,
    n2527,
    n2426,
    n2538,
    n2405
  );


  xnor
  g2644
  (
    n2654,
    n2390,
    n2381,
    n2568,
    n2479
  );


  and
  g2645
  (
    n2619,
    n2493,
    n2454,
    n2570,
    n2499
  );


  and
  g2646
  (
    n2664,
    n2393,
    n2490,
    n2568,
    n2531
  );


  or
  g2647
  (
    n2635,
    n2520,
    n2482,
    n2566,
    n2463
  );


  nor
  g2648
  (
    n2673,
    n2407,
    n2575,
    n2563,
    n2404
  );


  or
  g2649
  (
    n2645,
    n2467,
    n2586,
    n2441,
    n2523
  );


  nand
  g2650
  (
    n2638,
    n2516,
    n2456,
    n2535,
    n2473
  );


  and
  g2651
  (
    n2632,
    n2513,
    n2401,
    n2582,
    n2471
  );


  xnor
  g2652
  (
    n2610,
    n2533,
    n2546,
    n2509,
    n2423
  );


  nand
  g2653
  (
    n2678,
    n2500,
    n2535,
    n2555,
    n2448
  );


  xnor
  g2654
  (
    n2688,
    n2680,
    n2661,
    n2599,
    n2673
  );


  or
  g2655
  (
    n2686,
    n2632,
    n2648,
    n2674,
    n2640
  );


  or
  g2656
  (
    n2687,
    n2669,
    n2641,
    n2638,
    n2603
  );


  xor
  g2657
  (
    n2695,
    n2620,
    n2606,
    n2644,
    n2646
  );


  nand
  g2658
  (
    n2693,
    n2667,
    n2598,
    n2631,
    n2671
  );


  nor
  g2659
  (
    n2681,
    n2621,
    n2635,
    n2672,
    n2676
  );


  nor
  g2660
  (
    n2691,
    n2654,
    n2626,
    n2653,
    n2642
  );


  xnor
  g2661
  (
    n2689,
    n2651,
    n2622,
    n2668,
    n2605
  );


  nor
  g2662
  (
    n2694,
    n2675,
    n2608,
    n2633,
    n2678
  );


  xor
  g2663
  (
    n2685,
    n2645,
    n2666,
    n2609,
    n2610
  );


  and
  g2664
  (
    n2698,
    n2604,
    n2662,
    n2679,
    n2677
  );


  nor
  g2665
  (
    n2701,
    n2656,
    n2658,
    n2597,
    n2612
  );


  xor
  g2666
  (
    n2683,
    n2663,
    n2650,
    n2660,
    n2643
  );


  nand
  g2667
  (
    n2697,
    n2629,
    n2670,
    n2655,
    n2602
  );


  or
  g2668
  (
    n2700,
    n2625,
    n2607,
    n2627,
    n2636
  );


  or
  g2669
  (
    n2699,
    n2611,
    n2601,
    n2639,
    n2600
  );


  or
  g2670
  (
    n2684,
    n2659,
    n2637,
    n2665,
    n2623
  );


  xnor
  g2671
  (
    n2690,
    n2614,
    n2664,
    n2616,
    n2657
  );


  xnor
  g2672
  (
    n2696,
    n2628,
    n2634,
    n2617,
    n2647
  );


  or
  g2673
  (
    n2692,
    n2649,
    n2615,
    n2613,
    n2619
  );


  xor
  g2674
  (
    n2682,
    n2630,
    n2618,
    n2652,
    n2624
  );


  xnor
  KeyGate_0_0
  (
    n811,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n2558,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n195,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n468,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n346,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n2018,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1973,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n812,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n537,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1298,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1272,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1324,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n459,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1243,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1694,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n2219,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n868,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1834,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n101,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n2389,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n2261,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n589,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1109,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n405,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n940,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1639,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n2306,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n317,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1190,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n2274,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1944,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n2252,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n1550,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n560,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n876,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n170,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1264,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n2517,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n480,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n2044,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n1323,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n2649,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n2103,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n1362,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n615,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n2065,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n2575,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n2183,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n1087,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n143,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n1246,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n33,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n1397,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1075,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n2370,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n2053,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n2152,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n1005,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n2404,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n2462,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n1912,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n538,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n800,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n1477,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

