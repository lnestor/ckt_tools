

module Stat_1459_54_3
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n921,
  n922,
  n996,
  n988,
  n990,
  n998,
  n995,
  n1000,
  n985,
  n999,
  n997,
  n993,
  n991,
  n994,
  n983,
  n1053,
  n1085,
  n1086,
  n1080,
  n1084,
  n1081,
  n1078,
  n1082,
  n1077,
  n1136,
  n1134,
  n1131,
  n1132,
  n1135,
  n1137,
  n1133,
  n1495,
  n1496,
  n1497,
  n1493,
  n1494,
  n1491,
  n1490,
  n1492
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n921;output n922;output n996;output n988;output n990;output n998;output n995;output n1000;output n985;output n999;output n997;output n993;output n991;output n994;output n983;output n1053;output n1085;output n1086;output n1080;output n1084;output n1081;output n1078;output n1082;output n1077;output n1136;output n1134;output n1131;output n1132;output n1135;output n1137;output n1133;output n1495;output n1496;output n1497;output n1493;output n1494;output n1491;output n1490;output n1492;
  wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n984;wire n986;wire n987;wire n989;wire n992;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1079;wire n1083;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n106,
    n12
  );


  not
  g1
  (
    n109,
    n19
  );


  not
  g2
  (
    n91,
    n1
  );


  not
  g3
  (
    n96,
    n6
  );


  not
  g4
  (
    n48,
    n5
  );


  buf
  g5
  (
    n57,
    n21
  );


  buf
  g6
  (
    n41,
    n1
  );


  not
  g7
  (
    n101,
    n22
  );


  buf
  g8
  (
    n89,
    n8
  );


  buf
  g9
  (
    n116,
    n18
  );


  not
  g10
  (
    n66,
    n4
  );


  not
  g11
  (
    n62,
    n6
  );


  not
  g12
  (
    n58,
    n12
  );


  not
  g13
  (
    KeyWire_0_5,
    n11
  );


  not
  g14
  (
    n47,
    n3
  );


  not
  g15
  (
    n70,
    n8
  );


  not
  g16
  (
    n79,
    n16
  );


  not
  g17
  (
    n59,
    n15
  );


  buf
  g18
  (
    n90,
    n19
  );


  buf
  g19
  (
    n104,
    n5
  );


  buf
  g20
  (
    n40,
    n17
  );


  not
  g21
  (
    n61,
    n17
  );


  buf
  g22
  (
    n54,
    n15
  );


  buf
  g23
  (
    n78,
    n4
  );


  buf
  g24
  (
    n111,
    n19
  );


  buf
  g25
  (
    n105,
    n8
  );


  not
  g26
  (
    n100,
    n16
  );


  buf
  g27
  (
    n93,
    n6
  );


  buf
  g28
  (
    n94,
    n7
  );


  buf
  g29
  (
    n67,
    n17
  );


  buf
  g30
  (
    n42,
    n22
  );


  buf
  g31
  (
    n45,
    n20
  );


  not
  g32
  (
    n99,
    n11
  );


  not
  g33
  (
    n124,
    n4
  );


  buf
  g34
  (
    n55,
    n7
  );


  buf
  g35
  (
    n49,
    n10
  );


  not
  g36
  (
    n107,
    n6
  );


  buf
  g37
  (
    n110,
    n1
  );


  not
  g38
  (
    n64,
    n13
  );


  buf
  g39
  (
    n88,
    n10
  );


  buf
  g40
  (
    n121,
    n11
  );


  buf
  g41
  (
    n71,
    n20
  );


  buf
  g42
  (
    n43,
    n18
  );


  buf
  g43
  (
    n65,
    n14
  );


  buf
  g44
  (
    n76,
    n10
  );


  not
  g45
  (
    n44,
    n20
  );


  buf
  g46
  (
    n108,
    n15
  );


  buf
  g47
  (
    n84,
    n13
  );


  not
  g48
  (
    KeyWire_0_24,
    n5
  );


  not
  g49
  (
    n46,
    n9
  );


  buf
  g50
  (
    n95,
    n9
  );


  buf
  g51
  (
    n98,
    n13
  );


  buf
  g52
  (
    n81,
    n3
  );


  buf
  g53
  (
    n39,
    n8
  );


  buf
  g54
  (
    n63,
    n14
  );


  buf
  g55
  (
    n114,
    n21
  );


  not
  g56
  (
    n115,
    n9
  );


  buf
  g57
  (
    n102,
    n14
  );


  buf
  g58
  (
    n92,
    n19
  );


  not
  g59
  (
    n86,
    n18
  );


  not
  g60
  (
    n68,
    n2
  );


  buf
  g61
  (
    n122,
    n4
  );


  not
  g62
  (
    n56,
    n12
  );


  buf
  g63
  (
    n82,
    n3
  );


  not
  g64
  (
    n87,
    n21
  );


  buf
  g65
  (
    n77,
    n14
  );


  buf
  g66
  (
    n113,
    n21
  );


  buf
  g67
  (
    n85,
    n9
  );


  buf
  g68
  (
    n117,
    n13
  );


  buf
  g69
  (
    n75,
    n3
  );


  buf
  g70
  (
    n119,
    n1
  );


  buf
  g71
  (
    n60,
    n20
  );


  not
  g72
  (
    n103,
    n16
  );


  not
  g73
  (
    KeyWire_0_13,
    n5
  );


  not
  g74
  (
    n123,
    n2
  );


  buf
  g75
  (
    n53,
    n7
  );


  buf
  g76
  (
    n80,
    n16
  );


  not
  g77
  (
    n52,
    n10
  );


  not
  g78
  (
    n72,
    n17
  );


  not
  g79
  (
    n112,
    n18
  );


  buf
  g80
  (
    n69,
    n15
  );


  buf
  g81
  (
    n50,
    n7
  );


  buf
  g82
  (
    n73,
    n11
  );


  not
  g83
  (
    n97,
    n12
  );


  not
  g84
  (
    n74,
    n2
  );


  buf
  g85
  (
    n83,
    n2
  );


  not
  g86
  (
    n250,
    n43
  );


  buf
  g87
  (
    n197,
    n98
  );


  not
  g88
  (
    n327,
    n61
  );


  buf
  g89
  (
    n281,
    n96
  );


  not
  g90
  (
    n370,
    n52
  );


  not
  g91
  (
    n442,
    n70
  );


  buf
  g92
  (
    n264,
    n95
  );


  buf
  g93
  (
    n266,
    n81
  );


  not
  g94
  (
    n276,
    n114
  );


  buf
  g95
  (
    n210,
    n88
  );


  buf
  g96
  (
    n257,
    n105
  );


  buf
  g97
  (
    n341,
    n112
  );


  not
  g98
  (
    n126,
    n100
  );


  not
  g99
  (
    n223,
    n45
  );


  buf
  g100
  (
    n353,
    n94
  );


  not
  g101
  (
    n377,
    n78
  );


  buf
  g102
  (
    n166,
    n56
  );


  not
  g103
  (
    n300,
    n115
  );


  buf
  g104
  (
    n150,
    n112
  );


  not
  g105
  (
    n339,
    n114
  );


  buf
  g106
  (
    n418,
    n68
  );


  not
  g107
  (
    n129,
    n87
  );


  buf
  g108
  (
    n164,
    n50
  );


  buf
  g109
  (
    n406,
    n92
  );


  not
  g110
  (
    n272,
    n74
  );


  not
  g111
  (
    n224,
    n91
  );


  buf
  g112
  (
    n260,
    n94
  );


  not
  g113
  (
    n167,
    n92
  );


  not
  g114
  (
    n364,
    n116
  );


  buf
  g115
  (
    n261,
    n90
  );


  not
  g116
  (
    n410,
    n71
  );


  buf
  g117
  (
    n330,
    n54
  );


  buf
  g118
  (
    n422,
    n62
  );


  not
  g119
  (
    n438,
    n62
  );


  buf
  g120
  (
    n446,
    n80
  );


  buf
  g121
  (
    n193,
    n112
  );


  buf
  g122
  (
    n331,
    n106
  );


  not
  g123
  (
    n285,
    n114
  );


  buf
  g124
  (
    n348,
    n53
  );


  not
  g125
  (
    n192,
    n79
  );


  not
  g126
  (
    n371,
    n99
  );


  buf
  g127
  (
    n302,
    n121
  );


  buf
  g128
  (
    n297,
    n49
  );


  buf
  g129
  (
    n397,
    n115
  );


  buf
  g130
  (
    n369,
    n76
  );


  not
  g131
  (
    n296,
    n85
  );


  buf
  g132
  (
    n243,
    n76
  );


  buf
  g133
  (
    n130,
    n69
  );


  buf
  g134
  (
    n320,
    n43
  );


  not
  g135
  (
    n153,
    n65
  );


  buf
  g136
  (
    n242,
    n75
  );


  not
  g137
  (
    n148,
    n116
  );


  not
  g138
  (
    n235,
    n104
  );


  buf
  g139
  (
    n337,
    n60
  );


  buf
  g140
  (
    n165,
    n73
  );


  not
  g141
  (
    n267,
    n105
  );


  not
  g142
  (
    n209,
    n101
  );


  buf
  g143
  (
    n424,
    n90
  );


  not
  g144
  (
    n157,
    n119
  );


  buf
  g145
  (
    n200,
    n49
  );


  buf
  g146
  (
    n273,
    n60
  );


  not
  g147
  (
    n283,
    n69
  );


  buf
  g148
  (
    n398,
    n64
  );


  buf
  g149
  (
    n189,
    n60
  );


  not
  g150
  (
    n322,
    n95
  );


  buf
  g151
  (
    n402,
    n101
  );


  not
  g152
  (
    n433,
    n58
  );


  buf
  g153
  (
    n380,
    n85
  );


  buf
  g154
  (
    n408,
    n111
  );


  not
  g155
  (
    n247,
    n122
  );


  not
  g156
  (
    n163,
    n100
  );


  not
  g157
  (
    n182,
    n77
  );


  buf
  g158
  (
    n429,
    n74
  );


  not
  g159
  (
    n313,
    n47
  );


  not
  g160
  (
    n404,
    n95
  );


  not
  g161
  (
    n388,
    n96
  );


  not
  g162
  (
    n231,
    n69
  );


  not
  g163
  (
    n301,
    n118
  );


  buf
  g164
  (
    n376,
    n74
  );


  not
  g165
  (
    n354,
    n57
  );


  not
  g166
  (
    n439,
    n104
  );


  not
  g167
  (
    n318,
    n84
  );


  buf
  g168
  (
    n444,
    n63
  );


  not
  g169
  (
    n382,
    n59
  );


  buf
  g170
  (
    n183,
    n67
  );


  buf
  g171
  (
    n390,
    n68
  );


  not
  g172
  (
    n350,
    n82
  );


  not
  g173
  (
    n396,
    n75
  );


  buf
  g174
  (
    n191,
    n104
  );


  buf
  g175
  (
    n291,
    n77
  );


  not
  g176
  (
    n335,
    n81
  );


  buf
  g177
  (
    n425,
    n83
  );


  not
  g178
  (
    KeyWire_0_10,
    n110
  );


  not
  g179
  (
    n234,
    n44
  );


  not
  g180
  (
    n360,
    n120
  );


  not
  g181
  (
    n217,
    n85
  );


  not
  g182
  (
    n365,
    n108
  );


  not
  g183
  (
    n315,
    n54
  );


  buf
  g184
  (
    n212,
    n121
  );


  not
  g185
  (
    n405,
    n61
  );


  not
  g186
  (
    n171,
    n120
  );


  buf
  g187
  (
    n141,
    n72
  );


  buf
  g188
  (
    n345,
    n58
  );


  buf
  g189
  (
    n338,
    n77
  );


  buf
  g190
  (
    n393,
    n70
  );


  buf
  g191
  (
    n308,
    n72
  );


  buf
  g192
  (
    n415,
    n106
  );


  not
  g193
  (
    n132,
    n94
  );


  buf
  g194
  (
    n188,
    n91
  );


  not
  g195
  (
    n222,
    n78
  );


  buf
  g196
  (
    n340,
    n93
  );


  buf
  g197
  (
    n352,
    n117
  );


  not
  g198
  (
    n394,
    n73
  );


  buf
  g199
  (
    n201,
    n99
  );


  not
  g200
  (
    n254,
    n110
  );


  buf
  g201
  (
    n351,
    n72
  );


  not
  g202
  (
    n280,
    n107
  );


  not
  g203
  (
    n149,
    n92
  );


  not
  g204
  (
    n204,
    n115
  );


  buf
  g205
  (
    n147,
    n54
  );


  not
  g206
  (
    n328,
    n96
  );


  not
  g207
  (
    n431,
    n89
  );


  not
  g208
  (
    n437,
    n41
  );


  buf
  g209
  (
    n259,
    n83
  );


  not
  g210
  (
    n307,
    n40
  );


  not
  g211
  (
    n133,
    n52
  );


  not
  g212
  (
    n262,
    n61
  );


  buf
  g213
  (
    n258,
    n48
  );


  not
  g214
  (
    n135,
    n117
  );


  not
  g215
  (
    n187,
    n109
  );


  buf
  g216
  (
    n395,
    n86
  );


  not
  g217
  (
    n303,
    n116
  );


  not
  g218
  (
    n277,
    n63
  );


  not
  g219
  (
    n202,
    n101
  );


  buf
  g220
  (
    n289,
    n105
  );


  buf
  g221
  (
    KeyWire_0_29,
    n107
  );


  not
  g222
  (
    n420,
    n70
  );


  not
  g223
  (
    n215,
    n117
  );


  buf
  g224
  (
    n158,
    n117
  );


  not
  g225
  (
    n332,
    n94
  );


  not
  g226
  (
    n411,
    n39
  );


  buf
  g227
  (
    n391,
    n105
  );


  not
  g228
  (
    n241,
    n45
  );


  not
  g229
  (
    n387,
    n39
  );


  not
  g230
  (
    n220,
    n103
  );


  not
  g231
  (
    n237,
    n82
  );


  buf
  g232
  (
    n363,
    n99
  );


  not
  g233
  (
    n227,
    n40
  );


  not
  g234
  (
    n416,
    n102
  );


  buf
  g235
  (
    n426,
    n39
  );


  not
  g236
  (
    n373,
    n76
  );


  buf
  g237
  (
    n143,
    n116
  );


  buf
  g238
  (
    n137,
    n55
  );


  not
  g239
  (
    n274,
    n75
  );


  buf
  g240
  (
    n269,
    n101
  );


  buf
  g241
  (
    n190,
    n88
  );


  not
  g242
  (
    n435,
    n42
  );


  buf
  g243
  (
    n379,
    n48
  );


  not
  g244
  (
    n385,
    n79
  );


  buf
  g245
  (
    n314,
    n85
  );


  buf
  g246
  (
    n229,
    n100
  );


  not
  g247
  (
    n228,
    n50
  );


  buf
  g248
  (
    n145,
    n115
  );


  buf
  g249
  (
    n233,
    n122
  );


  buf
  g250
  (
    n134,
    n110
  );


  buf
  g251
  (
    n127,
    n89
  );


  buf
  g252
  (
    n427,
    n53
  );


  not
  g253
  (
    n305,
    n40
  );


  not
  g254
  (
    n419,
    n79
  );


  buf
  g255
  (
    n403,
    n60
  );


  not
  g256
  (
    n172,
    n78
  );


  buf
  g257
  (
    n181,
    n73
  );


  buf
  g258
  (
    n255,
    n49
  );


  not
  g259
  (
    n256,
    n82
  );


  buf
  g260
  (
    n432,
    n80
  );


  buf
  g261
  (
    n178,
    n46
  );


  buf
  g262
  (
    n434,
    n84
  );


  not
  g263
  (
    n361,
    n118
  );


  not
  g264
  (
    KeyWire_0_1,
    n64
  );


  not
  g265
  (
    n151,
    n58
  );


  buf
  g266
  (
    n177,
    n118
  );


  not
  g267
  (
    n428,
    n55
  );


  not
  g268
  (
    n218,
    n108
  );


  not
  g269
  (
    n139,
    n91
  );


  buf
  g270
  (
    n414,
    n55
  );


  buf
  g271
  (
    n381,
    n51
  );


  buf
  g272
  (
    n184,
    n67
  );


  not
  g273
  (
    n312,
    n50
  );


  buf
  g274
  (
    n236,
    n51
  );


  buf
  g275
  (
    n386,
    n86
  );


  not
  g276
  (
    n142,
    n71
  );


  not
  g277
  (
    n238,
    n48
  );


  not
  g278
  (
    n389,
    n66
  );


  not
  g279
  (
    n430,
    n113
  );


  buf
  g280
  (
    n329,
    n84
  );


  not
  g281
  (
    n248,
    n41
  );


  buf
  g282
  (
    n203,
    n93
  );


  buf
  g283
  (
    n282,
    n71
  );


  not
  g284
  (
    n349,
    n110
  );


  buf
  g285
  (
    n316,
    n121
  );


  not
  g286
  (
    n358,
    n98
  );


  buf
  g287
  (
    n162,
    n57
  );


  buf
  g288
  (
    n319,
    n90
  );


  not
  g289
  (
    n214,
    n43
  );


  buf
  g290
  (
    n356,
    n109
  );


  buf
  g291
  (
    n372,
    n42
  );


  not
  g292
  (
    n293,
    n42
  );


  not
  g293
  (
    n436,
    n120
  );


  buf
  g294
  (
    n186,
    n66
  );


  not
  g295
  (
    n230,
    n67
  );


  buf
  g296
  (
    n249,
    n87
  );


  buf
  g297
  (
    n213,
    n57
  );


  not
  g298
  (
    n265,
    n63
  );


  buf
  g299
  (
    n275,
    n113
  );


  not
  g300
  (
    n383,
    n58
  );


  buf
  g301
  (
    n138,
    n67
  );


  not
  g302
  (
    n384,
    n59
  );


  buf
  g303
  (
    n292,
    n51
  );


  buf
  g304
  (
    n195,
    n106
  );


  not
  g305
  (
    n154,
    n91
  );


  not
  g306
  (
    n136,
    n107
  );


  not
  g307
  (
    n357,
    n107
  );


  not
  g308
  (
    n325,
    n78
  );


  not
  g309
  (
    n263,
    n76
  );


  not
  g310
  (
    n421,
    n103
  );


  not
  g311
  (
    n342,
    n89
  );


  buf
  g312
  (
    n445,
    n81
  );


  buf
  g313
  (
    n176,
    n97
  );


  buf
  g314
  (
    n399,
    n103
  );


  buf
  g315
  (
    n226,
    n92
  );


  not
  g316
  (
    n413,
    n81
  );


  buf
  g317
  (
    n284,
    n46
  );


  not
  g318
  (
    n199,
    n74
  );


  not
  g319
  (
    n179,
    n77
  );


  not
  g320
  (
    n441,
    n122
  );


  buf
  g321
  (
    n288,
    n47
  );


  buf
  g322
  (
    n309,
    n119
  );


  not
  g323
  (
    n392,
    n123
  );


  not
  g324
  (
    n225,
    n97
  );


  buf
  g325
  (
    n245,
    n111
  );


  not
  g326
  (
    n175,
    n56
  );


  buf
  g327
  (
    n378,
    n90
  );


  not
  g328
  (
    n140,
    n88
  );


  not
  g329
  (
    n169,
    n83
  );


  not
  g330
  (
    n423,
    n89
  );


  buf
  g331
  (
    n294,
    n41
  );


  not
  g332
  (
    n270,
    n57
  );


  not
  g333
  (
    n152,
    n69
  );


  buf
  g334
  (
    n278,
    n56
  );


  not
  g335
  (
    n232,
    n80
  );


  buf
  g336
  (
    n180,
    n68
  );


  not
  g337
  (
    n271,
    n119
  );


  buf
  g338
  (
    n170,
    n66
  );


  buf
  g339
  (
    n295,
    n93
  );


  not
  g340
  (
    n362,
    n122
  );


  buf
  g341
  (
    n317,
    n68
  );


  buf
  g342
  (
    n207,
    n87
  );


  buf
  g343
  (
    n359,
    n53
  );


  buf
  g344
  (
    n174,
    n59
  );


  not
  g345
  (
    n251,
    n62
  );


  buf
  g346
  (
    n311,
    n120
  );


  buf
  g347
  (
    n173,
    n98
  );


  buf
  g348
  (
    n366,
    n121
  );


  buf
  g349
  (
    n198,
    n102
  );


  buf
  g350
  (
    n367,
    n62
  );


  not
  g351
  (
    n334,
    n104
  );


  buf
  g352
  (
    n219,
    n45
  );


  not
  g353
  (
    n168,
    n66
  );


  buf
  g354
  (
    n206,
    n108
  );


  buf
  g355
  (
    n159,
    n123
  );


  not
  g356
  (
    n125,
    n80
  );


  buf
  g357
  (
    n333,
    n46
  );


  buf
  g358
  (
    n185,
    n114
  );


  buf
  g359
  (
    n401,
    n102
  );


  not
  g360
  (
    n194,
    n97
  );


  not
  g361
  (
    n298,
    n86
  );


  not
  g362
  (
    n412,
    n79
  );


  not
  g363
  (
    KeyWire_0_21,
    n44
  );


  not
  g364
  (
    n409,
    n118
  );


  not
  g365
  (
    n346,
    n113
  );


  buf
  g366
  (
    n355,
    n100
  );


  not
  g367
  (
    n321,
    n70
  );


  not
  g368
  (
    n344,
    n55
  );


  buf
  g369
  (
    n221,
    n103
  );


  buf
  g370
  (
    n374,
    n83
  );


  not
  g371
  (
    n268,
    n71
  );


  buf
  g372
  (
    n323,
    n63
  );


  buf
  g373
  (
    n286,
    n64
  );


  buf
  g374
  (
    n304,
    n82
  );


  not
  g375
  (
    n290,
    n119
  );


  buf
  g376
  (
    n324,
    n109
  );


  buf
  g377
  (
    n407,
    n111
  );


  buf
  g378
  (
    n146,
    n52
  );


  not
  g379
  (
    n310,
    n95
  );


  not
  g380
  (
    n205,
    n93
  );


  buf
  g381
  (
    n131,
    n99
  );


  buf
  g382
  (
    n240,
    n65
  );


  buf
  g383
  (
    n400,
    n112
  );


  not
  g384
  (
    n336,
    n61
  );


  not
  g385
  (
    n156,
    n56
  );


  buf
  g386
  (
    n326,
    n84
  );


  not
  g387
  (
    KeyWire_0_4,
    n108
  );


  buf
  g388
  (
    n368,
    n87
  );


  buf
  g389
  (
    n375,
    n102
  );


  not
  g390
  (
    n440,
    n109
  );


  not
  g391
  (
    n246,
    n96
  );


  buf
  g392
  (
    n279,
    n111
  );


  buf
  g393
  (
    n347,
    n88
  );


  buf
  g394
  (
    n128,
    n59
  );


  not
  g395
  (
    n161,
    n106
  );


  not
  g396
  (
    n144,
    n44
  );


  buf
  g397
  (
    n417,
    n65
  );


  buf
  g398
  (
    n155,
    n73
  );


  not
  g399
  (
    n287,
    n64
  );


  buf
  g400
  (
    n211,
    n72
  );


  buf
  g401
  (
    n239,
    n113
  );


  buf
  g402
  (
    n253,
    n98
  );


  buf
  g403
  (
    n208,
    n97
  );


  buf
  g404
  (
    n306,
    n75
  );


  buf
  g405
  (
    n160,
    n65
  );


  not
  g406
  (
    n196,
    n47
  );


  not
  g407
  (
    n299,
    n86
  );


  xnor
  g408
  (
    n591,
    n308,
    n269,
    n322,
    n141
  );


  xor
  g409
  (
    n487,
    n234,
    n302,
    n210,
    n313
  );


  xor
  g410
  (
    n480,
    n157,
    n324,
    n224,
    n195
  );


  or
  g411
  (
    n481,
    n213,
    n148,
    n300,
    n128
  );


  and
  g412
  (
    n674,
    n223,
    n201,
    n221,
    n212
  );


  xnor
  g413
  (
    n455,
    n170,
    n238,
    n269,
    n279
  );


  xnor
  g414
  (
    n597,
    n146,
    n332,
    n168,
    n195
  );


  xnor
  g415
  (
    n657,
    n343,
    n144,
    n289,
    n262
  );


  nor
  g416
  (
    n449,
    n145,
    n127,
    n223,
    n137
  );


  and
  g417
  (
    n550,
    n280,
    n338,
    n319,
    n245
  );


  nand
  g418
  (
    n479,
    n346,
    n235,
    n243,
    n337
  );


  or
  g419
  (
    n466,
    n237,
    n310,
    n279,
    n184
  );


  xor
  g420
  (
    n620,
    n242,
    n305,
    n265,
    n206
  );


  nor
  g421
  (
    n531,
    n137,
    n271,
    n215,
    n161
  );


  nor
  g422
  (
    n561,
    n293,
    n328,
    n244,
    n158
  );


  nand
  g423
  (
    n634,
    n239,
    n292,
    n351,
    n149
  );


  nor
  g424
  (
    n488,
    n287,
    n213,
    n180,
    n177
  );


  or
  g425
  (
    n460,
    n205,
    n160,
    n129,
    n346
  );


  nand
  g426
  (
    n575,
    n229,
    n309,
    n163,
    n177
  );


  xor
  g427
  (
    n463,
    n178,
    n209,
    n334,
    n174
  );


  nand
  g428
  (
    n662,
    n293,
    n155,
    n191,
    n148
  );


  xnor
  g429
  (
    n483,
    n127,
    n195,
    n321,
    n349
  );


  xnor
  g430
  (
    n667,
    n132,
    n310,
    n230,
    n171
  );


  nand
  g431
  (
    n485,
    n242,
    n256,
    n301,
    n183
  );


  nand
  g432
  (
    n643,
    n150,
    n310,
    n222,
    n140
  );


  xnor
  g433
  (
    n453,
    n221,
    n169,
    n273,
    n298
  );


  nand
  g434
  (
    n607,
    n340,
    n345,
    n319,
    n173
  );


  or
  g435
  (
    n604,
    n350,
    n299,
    n333,
    n343
  );


  or
  g436
  (
    n489,
    n271,
    n304,
    n348,
    n215
  );


  xnor
  g437
  (
    n580,
    n341,
    n140,
    n332,
    n268
  );


  or
  g438
  (
    n652,
    n180,
    n129,
    n164,
    n179
  );


  and
  g439
  (
    n474,
    n186,
    n224,
    n211,
    n257
  );


  nand
  g440
  (
    n648,
    n171,
    n312,
    n319,
    n239
  );


  nor
  g441
  (
    n525,
    n294,
    n151,
    n309,
    n212
  );


  nand
  g442
  (
    KeyWire_0_15,
    n254,
    n253,
    n157,
    n218
  );


  or
  g443
  (
    n609,
    n318,
    n246,
    n178,
    n332
  );


  nand
  g444
  (
    n573,
    n347,
    n194,
    n204,
    n132
  );


  and
  g445
  (
    n450,
    n315,
    n322,
    n296,
    n247
  );


  nor
  g446
  (
    n624,
    n327,
    n240,
    n336,
    n348
  );


  xnor
  g447
  (
    KeyWire_0_12,
    n347,
    n198,
    n242,
    n133
  );


  or
  g448
  (
    n677,
    n303,
    n188,
    n125,
    n340
  );


  and
  g449
  (
    n645,
    n135,
    n342,
    n131,
    n220
  );


  and
  g450
  (
    n656,
    n183,
    n199,
    n252,
    n156
  );


  or
  g451
  (
    n465,
    n330,
    n334,
    n270,
    n253
  );


  nor
  g452
  (
    n554,
    n275,
    n227,
    n342,
    n187
  );


  xnor
  g453
  (
    n579,
    n257,
    n235,
    n181,
    n221
  );


  nand
  g454
  (
    n472,
    n212,
    n222,
    n219,
    n274
  );


  xnor
  g455
  (
    n482,
    n170,
    n211,
    n298,
    n272
  );


  nand
  g456
  (
    n549,
    n159,
    n231,
    n279,
    n206
  );


  nand
  g457
  (
    n592,
    n220,
    n349,
    n187,
    n145
  );


  nand
  g458
  (
    n528,
    n200,
    n204,
    n303,
    n158
  );


  xnor
  g459
  (
    n627,
    n288,
    n170,
    n294,
    n127
  );


  and
  g460
  (
    n564,
    n309,
    n175,
    n155,
    n320
  );


  xnor
  g461
  (
    n565,
    n282,
    n175,
    n225,
    n203
  );


  xor
  g462
  (
    n512,
    n139,
    n326,
    n199,
    n313
  );


  nor
  g463
  (
    n616,
    n278,
    n185,
    n244,
    n146
  );


  nor
  g464
  (
    n605,
    n197,
    n288,
    n239,
    n317
  );


  xnor
  g465
  (
    n496,
    n324,
    n154,
    n220,
    n210
  );


  nand
  g466
  (
    n533,
    n161,
    n343,
    n202,
    n285
  );


  xor
  g467
  (
    KeyWire_0_9,
    n298,
    n261,
    n167,
    n332
  );


  nand
  g468
  (
    n638,
    n204,
    n205,
    n305,
    n196
  );


  xor
  g469
  (
    n668,
    n345,
    n316,
    n218,
    n219
  );


  nor
  g470
  (
    n509,
    n300,
    n343,
    n260,
    n139
  );


  nand
  g471
  (
    n475,
    n266,
    n230,
    n231,
    n167
  );


  or
  g472
  (
    n506,
    n278,
    n182,
    n236,
    n288
  );


  nor
  g473
  (
    n672,
    n289,
    n162,
    n138,
    n333
  );


  nand
  g474
  (
    n484,
    n320,
    n135,
    n308,
    n303
  );


  xor
  g475
  (
    KeyWire_0_2,
    n152,
    n144,
    n331,
    n314
  );


  xnor
  g476
  (
    n562,
    n248,
    n252,
    n189,
    n280
  );


  xor
  g477
  (
    n637,
    n142,
    n209,
    n166,
    n131
  );


  xnor
  g478
  (
    n613,
    n297,
    n200,
    n245,
    n285
  );


  xnor
  g479
  (
    n559,
    n269,
    n283,
    n317,
    n195
  );


  or
  g480
  (
    n649,
    n229,
    n145,
    n173,
    n317
  );


  nand
  g481
  (
    n642,
    n336,
    n267,
    n128,
    n277
  );


  xnor
  g482
  (
    n492,
    n214,
    n198,
    n259,
    n158
  );


  xor
  g483
  (
    n541,
    n339,
    n274,
    n261,
    n301
  );


  xor
  g484
  (
    n658,
    n225,
    n136,
    n333,
    n148
  );


  nor
  g485
  (
    n669,
    n201,
    n219,
    n205
  );


  xnor
  g486
  (
    n454,
    n181,
    n186,
    n241,
    n286
  );


  nor
  g487
  (
    n593,
    n349,
    n171,
    n235,
    n268
  );


  nor
  g488
  (
    n497,
    n234,
    n282,
    n197,
    n241
  );


  or
  g489
  (
    n500,
    n135,
    n334,
    n247,
    n159
  );


  and
  g490
  (
    KeyWire_0_7,
    n226,
    n291,
    n232,
    n306
  );


  nor
  g491
  (
    n557,
    n169,
    n208,
    n353,
    n313
  );


  or
  g492
  (
    n594,
    n207,
    n229,
    n326,
    n213
  );


  nand
  g493
  (
    n458,
    n179,
    n163,
    n281,
    n256
  );


  xor
  g494
  (
    n513,
    n169,
    n217,
    n306,
    n247
  );


  and
  g495
  (
    n653,
    n143,
    n227,
    n133,
    n183
  );


  or
  g496
  (
    n577,
    n147,
    n128,
    n132,
    n174
  );


  nand
  g497
  (
    n670,
    n352,
    n125,
    n207,
    n305
  );


  and
  g498
  (
    n635,
    n292,
    n342,
    n256,
    n216
  );


  xor
  g499
  (
    n617,
    n188,
    n267,
    n339,
    n208
  );


  and
  g500
  (
    n650,
    n226,
    n283,
    n162,
    n285
  );


  and
  g501
  (
    n673,
    n341,
    n341,
    n302,
    n150
  );


  xnor
  g502
  (
    n495,
    n144,
    n327,
    n308,
    n170
  );


  and
  g503
  (
    n568,
    n193,
    n287,
    n320,
    n128
  );


  nor
  g504
  (
    n529,
    n248,
    n273,
    n157,
    n331
  );


  and
  g505
  (
    n536,
    n329,
    n278,
    n238,
    n165
  );


  and
  g506
  (
    n581,
    n216,
    n327,
    n233,
    n315
  );


  nor
  g507
  (
    n504,
    n173,
    n266,
    n318,
    n354
  );


  nand
  g508
  (
    n470,
    n198,
    n217,
    n260,
    n163
  );


  xnor
  g509
  (
    n602,
    n263,
    n147,
    n197,
    n134
  );


  nand
  g510
  (
    n665,
    n174,
    n191,
    n152,
    n238
  );


  and
  g511
  (
    n606,
    n299,
    n250,
    n328,
    n184
  );


  xor
  g512
  (
    n545,
    n336,
    n243,
    n291,
    n186
  );


  nor
  g513
  (
    n567,
    n151,
    n338,
    n165,
    n187
  );


  or
  g514
  (
    n486,
    n225,
    n236,
    n338,
    n286
  );


  and
  g515
  (
    n543,
    n349,
    n192,
    n271,
    n159
  );


  or
  g516
  (
    n571,
    n323,
    n328,
    n143,
    n355
  );


  nand
  g517
  (
    n560,
    n348,
    n330,
    n355,
    n193
  );


  or
  g518
  (
    n548,
    n338,
    n245,
    n189,
    n345
  );


  nor
  g519
  (
    n544,
    n166,
    n293,
    n341,
    n196
  );


  or
  g520
  (
    n518,
    n161,
    n180,
    n296,
    n351
  );


  or
  g521
  (
    n491,
    n139,
    n292,
    n154,
    n251
  );


  nand
  g522
  (
    n574,
    n137,
    n311,
    n291,
    n275
  );


  xor
  g523
  (
    n553,
    n310,
    n271,
    n182,
    n280
  );


  nor
  g524
  (
    n540,
    n151,
    n211,
    n282,
    n294
  );


  or
  g525
  (
    n459,
    n146,
    n315,
    n344,
    n131
  );


  nand
  g526
  (
    n582,
    n276,
    n249,
    n177,
    n189
  );


  and
  g527
  (
    n467,
    n178,
    n336,
    n151,
    n326
  );


  nor
  g528
  (
    n515,
    n261,
    n138,
    n137,
    n142
  );


  xnor
  g529
  (
    n676,
    n223,
    n201,
    n284,
    n130
  );


  xnor
  g530
  (
    n537,
    n327,
    n243,
    n202,
    n350
  );


  nand
  g531
  (
    n471,
    n164,
    n161,
    n329,
    n264
  );


  xnor
  g532
  (
    n631,
    n200,
    n275,
    n150,
    n344
  );


  nor
  g533
  (
    n675,
    n347,
    n352,
    n278,
    n330
  );


  and
  g534
  (
    n614,
    n304,
    n190,
    n153,
    n179
  );


  or
  g535
  (
    n603,
    n140,
    n222,
    n315,
    n249
  );


  xnor
  g536
  (
    n576,
    n245,
    n141,
    n130,
    n357
  );


  nand
  g537
  (
    n476,
    n152,
    n311,
    n321,
    n187
  );


  nand
  g538
  (
    n457,
    n180,
    n211,
    n237,
    n259
  );


  nor
  g539
  (
    n563,
    n276,
    n263,
    n354,
    n246
  );


  nor
  g540
  (
    n644,
    n214,
    n201,
    n266,
    n233
  );


  xor
  g541
  (
    n587,
    n149,
    n189,
    n314,
    n331
  );


  nand
  g542
  (
    n663,
    n256,
    n281,
    n260,
    n199
  );


  nor
  g543
  (
    n654,
    n295,
    n282,
    n168,
    n312
  );


  nor
  g544
  (
    n514,
    n164,
    n270,
    n163,
    n226
  );


  xor
  g545
  (
    n660,
    n340,
    n244,
    n228,
    n269
  );


  or
  g546
  (
    n584,
    n283,
    n288,
    n237,
    n355
  );


  and
  g547
  (
    n626,
    n297,
    n345,
    n262
  );


  xnor
  g548
  (
    n623,
    n222,
    n305,
    n164,
    n346
  );


  xor
  g549
  (
    n583,
    n147,
    n136,
    n219,
    n354
  );


  xnor
  g550
  (
    n566,
    n347,
    n230,
    n133,
    n356
  );


  and
  g551
  (
    n615,
    n323,
    n265,
    n209,
    n337
  );


  xor
  g552
  (
    n640,
    n228,
    n165,
    n353,
    n184
  );


  or
  g553
  (
    n527,
    n265,
    n258,
    n311,
    n263
  );


  and
  g554
  (
    n507,
    n234,
    n346,
    n202,
    n253
  );


  xor
  g555
  (
    n610,
    n248,
    n290,
    n194,
    n236
  );


  xnor
  g556
  (
    n552,
    n150,
    n214,
    n257,
    n190
  );


  xor
  g557
  (
    n633,
    n318,
    n306,
    n274,
    n213
  );


  xnor
  g558
  (
    n569,
    n224,
    n199,
    n194,
    n134
  );


  xnor
  g559
  (
    n511,
    n325,
    n352,
    n249,
    n253
  );


  and
  g560
  (
    n473,
    n246,
    n240,
    n274,
    n335
  );


  xor
  g561
  (
    n517,
    n322,
    n126,
    n334,
    n287
  );


  or
  g562
  (
    n516,
    n140,
    n284,
    n298,
    n233
  );


  and
  g563
  (
    n477,
    n331,
    n264,
    n302,
    n156
  );


  and
  g564
  (
    n505,
    n167,
    n181,
    n129,
    n302
  );


  or
  g565
  (
    n612,
    n166,
    n247,
    n153,
    n246
  );


  xor
  g566
  (
    KeyWire_0_6,
    n176,
    n326,
    n125,
    n175
  );


  nand
  g567
  (
    n588,
    n215,
    n254,
    n228,
    n255
  );


  nand
  g568
  (
    n551,
    n149,
    n129,
    n344,
    n136
  );


  and
  g569
  (
    n461,
    n171,
    n130,
    n240,
    n159
  );


  nand
  g570
  (
    n523,
    n339,
    n157,
    n300,
    n342
  );


  nor
  g571
  (
    n589,
    n337,
    n339,
    n192,
    n303
  );


  xor
  g572
  (
    n498,
    n221,
    n168,
    n138,
    n296
  );


  nand
  g573
  (
    n647,
    n167,
    n272,
    n218,
    n158
  );


  nand
  g574
  (
    n555,
    n232,
    n232,
    n272,
    n290
  );


  xor
  g575
  (
    n530,
    n183,
    n241,
    n212,
    n299
  );


  xor
  g576
  (
    n494,
    n317,
    n190,
    n168,
    n217
  );


  xor
  g577
  (
    n572,
    n188,
    n138,
    n324,
    n280
  );


  and
  g578
  (
    n598,
    n313,
    n248,
    n289,
    n255
  );


  or
  g579
  (
    n595,
    n179,
    n297,
    n174,
    n261
  );


  nor
  g580
  (
    n608,
    n197,
    n193,
    n184,
    n210
  );


  xnor
  g581
  (
    n464,
    n217,
    n169,
    n227,
    n264
  );


  xor
  g582
  (
    n628,
    n188,
    n259,
    n325,
    n295
  );


  nor
  g583
  (
    n558,
    n182,
    n286,
    n283,
    n203
  );


  and
  g584
  (
    n448,
    n224,
    n154,
    n281,
    n126
  );


  nand
  g585
  (
    n570,
    n250,
    n292,
    n352,
    n295
  );


  and
  g586
  (
    n520,
    n324,
    n185,
    n289,
    n242
  );


  and
  g587
  (
    n599,
    n176,
    n223,
    n194,
    n270
  );


  or
  g588
  (
    n630,
    n262,
    n354,
    n250,
    n323
  );


  nand
  g589
  (
    n611,
    n132,
    n277,
    n153
  );


  xnor
  g590
  (
    n590,
    n273,
    n350,
    n353,
    n127
  );


  or
  g591
  (
    n659,
    n218,
    n162,
    n314,
    n185
  );


  nand
  g592
  (
    n478,
    n203,
    n191,
    n142,
    n321
  );


  nor
  g593
  (
    n664,
    n265,
    n172,
    n162,
    n355
  );


  nor
  g594
  (
    n651,
    n299,
    n229,
    n131,
    n258
  );


  nor
  g595
  (
    n535,
    n275,
    n207,
    n312,
    n307
  );


  nand
  g596
  (
    n524,
    n356,
    n216,
    n185,
    n130
  );


  nor
  g597
  (
    n585,
    n134,
    n204,
    n155,
    n136
  );


  nand
  g598
  (
    n678,
    n251,
    n172,
    n307
  );


  or
  g599
  (
    n490,
    n304,
    n216,
    n252,
    n296
  );


  and
  g600
  (
    n632,
    n252,
    n268,
    n329,
    n286
  );


  nor
  g601
  (
    n510,
    n258,
    n277,
    n190,
    n193
  );


  nand
  g602
  (
    n452,
    n178,
    n154,
    n176,
    n287
  );


  xnor
  g603
  (
    n499,
    n196,
    n335,
    n301,
    n353
  );


  nor
  g604
  (
    n521,
    n192,
    n177,
    n147,
    n251
  );


  xor
  g605
  (
    n538,
    n290,
    n279,
    n325,
    n311
  );


  xnor
  g606
  (
    n534,
    n276,
    n156,
    n356,
    n333
  );


  and
  g607
  (
    n586,
    n290,
    n173,
    n329,
    n335
  );


  nand
  g608
  (
    n462,
    n351,
    n267,
    n241,
    n160
  );


  or
  g609
  (
    n655,
    n244,
    n134,
    n165,
    n297
  );


  nand
  g610
  (
    n619,
    n266,
    n206,
    n210,
    n175
  );


  or
  g611
  (
    n666,
    n320,
    n328,
    n206,
    n182
  );


  xnor
  g612
  (
    n493,
    n220,
    n208,
    n295,
    n228
  );


  xor
  g613
  (
    n661,
    n249,
    n254,
    n340,
    n227
  );


  xor
  g614
  (
    n547,
    n239,
    n319,
    n309,
    n203
  );


  or
  g615
  (
    n600,
    n192,
    n186,
    n250,
    n143
  );


  and
  g616
  (
    n546,
    n263,
    n325,
    n314,
    n155
  );


  or
  g617
  (
    n502,
    n133,
    n149,
    n235,
    n160
  );


  or
  g618
  (
    n596,
    n232,
    n350,
    n156,
    n196
  );


  or
  g619
  (
    n578,
    n285,
    n139,
    n143,
    n237
  );


  or
  g620
  (
    n636,
    n276,
    n234,
    n273,
    n260
  );


  and
  g621
  (
    n641,
    n272,
    n356,
    n268,
    n351
  );


  or
  g622
  (
    n539,
    n308,
    n306,
    n191,
    n322
  );


  and
  g623
  (
    n646,
    n294,
    n233,
    n243,
    n135
  );


  and
  g624
  (
    n522,
    n307,
    n301,
    n176,
    n318
  );


  or
  g625
  (
    n451,
    n146,
    n166,
    n144,
    n291
  );


  and
  g626
  (
    n532,
    n284,
    n141,
    n323,
    n148
  );


  and
  g627
  (
    n501,
    n270,
    n198,
    n215,
    n160
  );


  xor
  g628
  (
    n469,
    n181,
    n304,
    n284,
    n330
  );


  nor
  g629
  (
    n468,
    n316,
    n321,
    n257,
    n240
  );


  or
  g630
  (
    n508,
    n126,
    n254,
    n348,
    n281
  );


  or
  g631
  (
    n447,
    n230,
    n236,
    n145,
    n255
  );


  and
  g632
  (
    n556,
    n344,
    n202,
    n225,
    n172
  );


  nand
  g633
  (
    n503,
    n209,
    n226,
    n251,
    n141
  );


  and
  g634
  (
    n526,
    n316,
    n293,
    n255,
    n231
  );


  nand
  g635
  (
    n542,
    n300,
    n335,
    n208,
    n126
  );


  nand
  g636
  (
    n601,
    n142,
    n312,
    n152,
    n259
  );


  nand
  g637
  (
    n639,
    n267,
    n264,
    n258,
    n238
  );


  xnor
  g638
  (
    n618,
    n277,
    n200,
    n316,
    n207
  );


  nand
  g639
  (
    n519,
    n214,
    n337,
    n307,
    n231
  );


  buf
  g640
  (
    n685,
    n458
  );


  not
  g641
  (
    n714,
    n448
  );


  not
  g642
  (
    n738,
    n481
  );


  not
  g643
  (
    n740,
    n464
  );


  buf
  g644
  (
    n696,
    n492
  );


  not
  g645
  (
    n737,
    n502
  );


  buf
  g646
  (
    n718,
    n462
  );


  buf
  g647
  (
    n681,
    n459
  );


  not
  g648
  (
    n728,
    n470
  );


  not
  g649
  (
    n710,
    n499
  );


  buf
  g650
  (
    n734,
    n501
  );


  not
  g651
  (
    n711,
    n456
  );


  not
  g652
  (
    n704,
    n506
  );


  buf
  g653
  (
    n712,
    n488
  );


  buf
  g654
  (
    n707,
    n452
  );


  buf
  g655
  (
    n690,
    n460
  );


  buf
  g656
  (
    n736,
    n447
  );


  buf
  g657
  (
    n684,
    n463
  );


  not
  g658
  (
    n730,
    n467
  );


  buf
  g659
  (
    n689,
    n479
  );


  not
  g660
  (
    n682,
    n454
  );


  buf
  g661
  (
    n698,
    n491
  );


  buf
  g662
  (
    n735,
    n493
  );


  not
  g663
  (
    n683,
    n504
  );


  not
  g664
  (
    n706,
    n466
  );


  not
  g665
  (
    n726,
    n461
  );


  buf
  g666
  (
    n702,
    n472
  );


  not
  g667
  (
    n733,
    n489
  );


  buf
  g668
  (
    n687,
    n476
  );


  buf
  g669
  (
    n703,
    n455
  );


  not
  g670
  (
    n729,
    n453
  );


  buf
  g671
  (
    n731,
    n451
  );


  not
  g672
  (
    n719,
    n505
  );


  buf
  g673
  (
    n709,
    n509
  );


  not
  g674
  (
    n691,
    n465
  );


  buf
  g675
  (
    n686,
    n497
  );


  buf
  g676
  (
    n708,
    n473
  );


  not
  g677
  (
    n695,
    n469
  );


  not
  g678
  (
    n699,
    n468
  );


  not
  g679
  (
    n721,
    n450
  );


  not
  g680
  (
    n701,
    n498
  );


  not
  g681
  (
    n716,
    n508
  );


  buf
  g682
  (
    n679,
    n457
  );


  buf
  g683
  (
    n694,
    n487
  );


  not
  g684
  (
    n725,
    n475
  );


  buf
  g685
  (
    n700,
    n490
  );


  not
  g686
  (
    n717,
    n478
  );


  buf
  g687
  (
    n692,
    n474
  );


  not
  g688
  (
    n713,
    n477
  );


  buf
  g689
  (
    n715,
    n495
  );


  not
  g690
  (
    n688,
    n483
  );


  not
  g691
  (
    n697,
    n484
  );


  not
  g692
  (
    n722,
    n471
  );


  not
  g693
  (
    n724,
    n449
  );


  buf
  g694
  (
    n720,
    n496
  );


  buf
  g695
  (
    n693,
    n480
  );


  not
  g696
  (
    n732,
    n494
  );


  not
  g697
  (
    n741,
    n507
  );


  not
  g698
  (
    n727,
    n510
  );


  not
  g699
  (
    n742,
    n486
  );


  buf
  g700
  (
    n705,
    n503
  );


  buf
  g701
  (
    n680,
    n500
  );


  not
  g702
  (
    n739,
    n482
  );


  not
  g703
  (
    n723,
    n485
  );


  buf
  g704
  (
    n768,
    n387
  );


  buf
  g705
  (
    n796,
    n414
  );


  not
  g706
  (
    n838,
    n409
  );


  buf
  g707
  (
    n851,
    n383
  );


  buf
  g708
  (
    n782,
    n375
  );


  buf
  g709
  (
    n810,
    n32
  );


  not
  g710
  (
    n814,
    n414
  );


  not
  g711
  (
    n816,
    n375
  );


  not
  g712
  (
    n879,
    n711
  );


  buf
  g713
  (
    KeyWire_0_28,
    n719
  );


  buf
  g714
  (
    n813,
    n714
  );


  not
  g715
  (
    n834,
    n27
  );


  not
  g716
  (
    n788,
    n722
  );


  not
  g717
  (
    n797,
    n703
  );


  not
  g718
  (
    n793,
    n382
  );


  not
  g719
  (
    n871,
    n687
  );


  buf
  g720
  (
    n843,
    n724
  );


  buf
  g721
  (
    n846,
    n726
  );


  not
  g722
  (
    n845,
    n369
  );


  not
  g723
  (
    n859,
    n379
  );


  buf
  g724
  (
    n798,
    n364
  );


  nor
  g725
  (
    n850,
    n680,
    n367,
    n695
  );


  xor
  g726
  (
    n882,
    n385,
    n367,
    n709
  );


  or
  g727
  (
    n803,
    n385,
    n428,
    n691
  );


  or
  g728
  (
    n855,
    n424,
    n370,
    n374
  );


  nor
  g729
  (
    n775,
    n390,
    n722,
    n23
  );


  xnor
  g730
  (
    n874,
    n709,
    n31,
    n393
  );


  or
  g731
  (
    n752,
    n404,
    n362,
    n686
  );


  xnor
  g732
  (
    n875,
    n688,
    n721,
    n694
  );


  and
  g733
  (
    n822,
    n679,
    n371,
    n423
  );


  nand
  g734
  (
    n836,
    n358,
    n698,
    n368
  );


  nand
  g735
  (
    n856,
    n692,
    n713,
    n686
  );


  xnor
  g736
  (
    n783,
    n420,
    n385,
    n415
  );


  nor
  g737
  (
    n743,
    n684,
    n714,
    n369
  );


  nor
  g738
  (
    n808,
    n374,
    n695,
    n382
  );


  xnor
  g739
  (
    n864,
    n691,
    n401,
    n385
  );


  xnor
  g740
  (
    n809,
    n31,
    n24,
    n426
  );


  xor
  g741
  (
    n844,
    n368,
    n698,
    n364
  );


  or
  g742
  (
    n772,
    n408,
    n417,
    n412
  );


  xnor
  g743
  (
    n839,
    n379,
    n705,
    n697,
    n706
  );


  or
  g744
  (
    n770,
    n701,
    n421,
    n28,
    n369
  );


  xnor
  g745
  (
    n784,
    n370,
    n380,
    n715,
    n704
  );


  xnor
  g746
  (
    n760,
    n387,
    n720,
    n34,
    n390
  );


  and
  g747
  (
    n755,
    n394,
    n721,
    n393,
    n383
  );


  nor
  g748
  (
    n789,
    n395,
    n34,
    n392,
    n383
  );


  xor
  g749
  (
    n837,
    n416,
    n395,
    n357,
    n360
  );


  and
  g750
  (
    n835,
    n422,
    n426,
    n403,
    n427
  );


  xnor
  g751
  (
    n791,
    n376,
    n377,
    n412,
    n401
  );


  xor
  g752
  (
    n853,
    n397,
    n388,
    n421,
    n684
  );


  or
  g753
  (
    n847,
    n398,
    n373,
    n404,
    n425
  );


  nand
  g754
  (
    n817,
    n378,
    n373,
    n712,
    n407
  );


  xnor
  g755
  (
    n869,
    n30,
    n366,
    n365,
    n361
  );


  xnor
  g756
  (
    n823,
    n364,
    n32,
    n716,
    n33
  );


  and
  g757
  (
    n865,
    n372,
    n379,
    n363
  );


  or
  g758
  (
    n794,
    n28,
    n703,
    n390,
    n692
  );


  or
  g759
  (
    n780,
    n387,
    n716,
    n689
  );


  xnor
  g760
  (
    n781,
    n391,
    n380,
    n34,
    n23
  );


  xor
  g761
  (
    n828,
    n717,
    n371,
    n715,
    n691
  );


  or
  g762
  (
    n756,
    n694,
    n383,
    n715,
    n406
  );


  and
  g763
  (
    KeyWire_0_3,
    n701,
    n26,
    n24,
    n386
  );


  xor
  g764
  (
    n754,
    n419,
    n718,
    n388,
    n395
  );


  xor
  g765
  (
    n763,
    n391,
    n408,
    n693,
    n719
  );


  xnor
  g766
  (
    n748,
    n426,
    n411,
    n381,
    n409
  );


  or
  g767
  (
    n753,
    n685,
    n685,
    n376,
    n33
  );


  or
  g768
  (
    n824,
    n720,
    n406,
    n32,
    n719
  );


  xnor
  g769
  (
    n863,
    n424,
    n367,
    n708,
    n29
  );


  nor
  g770
  (
    n848,
    n386,
    n398,
    n394,
    n370
  );


  nand
  g771
  (
    n866,
    n422,
    n410,
    n361,
    n423
  );


  xnor
  g772
  (
    n769,
    n384,
    n413,
    n372,
    n375
  );


  xnor
  g773
  (
    n870,
    n427,
    n23,
    n406,
    n397
  );


  xor
  g774
  (
    n872,
    n690,
    n31,
    n706,
    n703
  );


  xor
  g775
  (
    n773,
    n359,
    n402,
    n423,
    n26
  );


  xor
  g776
  (
    n873,
    n30,
    n33,
    n710,
    n360
  );


  xnor
  g777
  (
    n881,
    n426,
    n389,
    n702,
    n681
  );


  and
  g778
  (
    n747,
    n406,
    n360,
    n720,
    n707
  );


  xor
  g779
  (
    KeyWire_0_18,
    n709,
    n366,
    n376,
    n373
  );


  nand
  g780
  (
    n861,
    n389,
    n390,
    n379,
    n690
  );


  or
  g781
  (
    n857,
    n425,
    n693,
    n25,
    n712
  );


  xor
  g782
  (
    n867,
    n365,
    n726,
    n417,
    n397
  );


  nor
  g783
  (
    n758,
    n382,
    n371,
    n711,
    n378
  );


  xnor
  g784
  (
    n786,
    n362,
    n419,
    n422,
    n680
  );


  or
  g785
  (
    n815,
    n402,
    n29,
    n369,
    n414
  );


  nand
  g786
  (
    n852,
    n725,
    n377,
    n358
  );


  or
  g787
  (
    n750,
    n415,
    n700,
    n692,
    n359
  );


  xor
  g788
  (
    n764,
    n705,
    n386,
    n416,
    n403
  );


  xnor
  g789
  (
    n830,
    n699,
    n26,
    n380,
    n399
  );


  xor
  g790
  (
    n761,
    n718,
    n380,
    n424,
    n378
  );


  xor
  g791
  (
    n829,
    n381,
    n408,
    n372,
    n714
  );


  and
  g792
  (
    n840,
    n24,
    n27,
    n396,
    n683
  );


  xnor
  g793
  (
    n744,
    n405,
    n27,
    n413,
    n368
  );


  nand
  g794
  (
    n759,
    n717,
    n417,
    n416,
    n398
  );


  xnor
  g795
  (
    n749,
    n403,
    n403,
    n402,
    n409
  );


  xnor
  g796
  (
    n777,
    n367,
    n30,
    n31,
    n710
  );


  xnor
  g797
  (
    n860,
    n366,
    n418,
    n404,
    n396
  );


  or
  g798
  (
    n807,
    n414,
    n25,
    n404,
    n723
  );


  and
  g799
  (
    n787,
    n386,
    n687,
    n419,
    n400
  );


  and
  g800
  (
    n842,
    n407,
    n391,
    n368,
    n377
  );


  nand
  g801
  (
    n785,
    n681,
    n364,
    n712,
    n688
  );


  nand
  g802
  (
    n745,
    n716,
    n686,
    n690,
    n384
  );


  xor
  g803
  (
    n801,
    n710,
    n371,
    n696
  );


  and
  g804
  (
    n868,
    n411,
    n421,
    n698,
    n389
  );


  nor
  g805
  (
    n776,
    n365,
    n411,
    n381,
    n388
  );


  and
  g806
  (
    n766,
    n417,
    n705,
    n27,
    n392
  );


  xor
  g807
  (
    n858,
    n396,
    n384,
    n378,
    n25
  );


  or
  g808
  (
    n806,
    n375,
    n689,
    n422,
    n29
  );


  xor
  g809
  (
    n841,
    n704,
    n708,
    n28,
    n373
  );


  xor
  g810
  (
    n831,
    n685,
    n702,
    n28,
    n413
  );


  nor
  g811
  (
    n854,
    n384,
    n397,
    n424,
    n358
  );


  nor
  g812
  (
    n833,
    n402,
    n411,
    n704,
    n357
  );


  xnor
  g813
  (
    n849,
    n725,
    n22,
    n683,
    n405
  );


  xor
  g814
  (
    n825,
    n372,
    n24,
    n22,
    n400
  );


  nand
  g815
  (
    n826,
    n725,
    n684,
    n423,
    n418
  );


  nand
  g816
  (
    n778,
    n400,
    n724,
    n362,
    n723
  );


  nor
  g817
  (
    n878,
    n34,
    n723,
    n697,
    n410
  );


  nand
  g818
  (
    n877,
    n412,
    n395,
    n683,
    n717
  );


  xor
  g819
  (
    n832,
    n399,
    n362,
    n370,
    n381
  );


  nor
  g820
  (
    n819,
    n412,
    n724,
    n415,
    n700
  );


  xor
  g821
  (
    n799,
    n427,
    n682,
    n699
  );


  xor
  g822
  (
    n800,
    n363,
    n687,
    n708,
    n389
  );


  nand
  g823
  (
    n746,
    n680,
    n702,
    n421,
    n726
  );


  xnor
  g824
  (
    n804,
    n359,
    n718,
    n418,
    n399
  );


  xnor
  g825
  (
    n762,
    n681,
    n713,
    n706,
    n682
  );


  xnor
  g826
  (
    n757,
    n391,
    n427,
    n360,
    n420
  );


  nor
  g827
  (
    n812,
    n30,
    n363,
    n700,
    n407
  );


  xor
  g828
  (
    n876,
    n713,
    n400,
    n394,
    n410
  );


  xnor
  g829
  (
    n767,
    n410,
    n711,
    n361,
    n359
  );


  xnor
  g830
  (
    n751,
    n707,
    n679,
    n420
  );


  xor
  g831
  (
    n792,
    n394,
    n382,
    n396,
    n428
  );


  and
  g832
  (
    n805,
    n405,
    n365,
    n393,
    n413
  );


  nor
  g833
  (
    KeyWire_0_0,
    n694,
    n398,
    n401,
    n696
  );


  nand
  g834
  (
    n811,
    n425,
    n693,
    n682,
    n419
  );


  nor
  g835
  (
    n765,
    n405,
    n688,
    n392,
    n695
  );


  and
  g836
  (
    n820,
    n697,
    n26,
    n29,
    n32
  );


  nor
  g837
  (
    n790,
    n361,
    n409,
    n722,
    n374
  );


  and
  g838
  (
    n821,
    n399,
    n418,
    n721,
    n374
  );


  or
  g839
  (
    n880,
    n707,
    n701,
    n393,
    n407
  );


  xnor
  g840
  (
    n774,
    n358,
    n388,
    n25,
    n401
  );


  nand
  g841
  (
    n862,
    n23,
    n376,
    n425,
    n387
  );


  nand
  g842
  (
    n779,
    n366,
    n416,
    n415,
    n420
  );


  xor
  g843
  (
    n802,
    n357,
    n33,
    n392,
    n408
  );


  and
  g844
  (
    n900,
    n751,
    n525,
    n759,
    n765
  );


  xor
  g845
  (
    n909,
    n559,
    n557,
    n744,
    n764
  );


  nor
  g846
  (
    n908,
    n550,
    n770,
    n511,
    n537
  );


  and
  g847
  (
    n913,
    n755,
    n513,
    n747,
    n746
  );


  nor
  g848
  (
    n886,
    n549,
    n768,
    n766,
    n762
  );


  or
  g849
  (
    n897,
    n564,
    n556,
    n519,
    n758
  );


  and
  g850
  (
    n888,
    n746,
    n757,
    n534,
    n748
  );


  nand
  g851
  (
    KeyWire_0_19,
    n545,
    n560,
    n527,
    n521
  );


  or
  g852
  (
    n918,
    n539,
    n767,
    n768,
    n754
  );


  or
  g853
  (
    n895,
    n773,
    n753,
    n520
  );


  xor
  g854
  (
    n892,
    n750,
    n757,
    n752,
    n761
  );


  xor
  g855
  (
    n904,
    n743,
    n773,
    n771,
    n522
  );


  xor
  g856
  (
    n919,
    n524,
    n749,
    n755,
    n528
  );


  and
  g857
  (
    n891,
    n531,
    n767,
    n555,
    n763
  );


  xnor
  g858
  (
    n914,
    n756,
    n535,
    n530,
    n769
  );


  nand
  g859
  (
    n917,
    n758,
    n551,
    n770,
    n751
  );


  xor
  g860
  (
    KeyWire_0_30,
    n526,
    n749,
    n561,
    n770
  );


  and
  g861
  (
    n885,
    n515,
    n751,
    n744,
    n553
  );


  nor
  g862
  (
    n910,
    n749,
    n544,
    n760,
    n762
  );


  nor
  g863
  (
    n894,
    n761,
    n768,
    n759,
    n750
  );


  nor
  g864
  (
    n893,
    n759,
    n532,
    n754,
    n523
  );


  and
  g865
  (
    n906,
    n516,
    n757,
    n547,
    n546
  );


  nor
  g866
  (
    n915,
    n746,
    n772,
    n536,
    n762
  );


  nor
  g867
  (
    n896,
    n761,
    n767,
    n745,
    n743
  );


  nor
  g868
  (
    n912,
    n552,
    n754,
    n764,
    n771
  );


  nor
  g869
  (
    n887,
    n558,
    n752,
    n533,
    n747
  );


  and
  g870
  (
    n911,
    n769,
    n514,
    n747,
    n766
  );


  or
  g871
  (
    n916,
    n744,
    n764,
    n529,
    n540
  );


  and
  g872
  (
    n883,
    n541,
    n758,
    n548,
    n753
  );


  xnor
  g873
  (
    n902,
    n765,
    n755,
    n774,
    n763
  );


  and
  g874
  (
    n890,
    n543,
    n765,
    n756,
    n563
  );


  xnor
  g875
  (
    n907,
    n512,
    n518,
    n760,
    n748
  );


  nand
  g876
  (
    n889,
    n773,
    n769,
    n772,
    n771
  );


  nand
  g877
  (
    n899,
    n763,
    n562,
    n554,
    n766
  );


  and
  g878
  (
    n905,
    n745,
    n538,
    n750,
    n743
  );


  xor
  g879
  (
    n903,
    n542,
    n756,
    n772,
    n760
  );


  and
  g880
  (
    n901,
    n748,
    n745,
    n517,
    n752
  );


  buf
  g881
  (
    n921,
    n883
  );


  not
  g882
  (
    n920,
    n883
  );


  not
  g883
  (
    n922,
    n921
  );


  not
  g884
  (
    n923,
    n922
  );


  buf
  g885
  (
    n925,
    n922
  );


  not
  g886
  (
    n924,
    n922
  );


  not
  g887
  (
    n927,
    n925
  );


  not
  g888
  (
    n929,
    n923
  );


  buf
  g889
  (
    n930,
    n923
  );


  buf
  g890
  (
    n934,
    n923
  );


  not
  g891
  (
    n931,
    n924
  );


  not
  g892
  (
    n932,
    n924
  );


  buf
  g893
  (
    n926,
    n924
  );


  buf
  g894
  (
    n933,
    n924
  );


  not
  g895
  (
    n928,
    n923
  );


  and
  g896
  (
    n959,
    n626,
    n620,
    n568,
    n602
  );


  or
  g897
  (
    n949,
    n565,
    n929,
    n575,
    n597
  );


  nand
  g898
  (
    n955,
    n615,
    n928,
    n601,
    n609
  );


  nor
  g899
  (
    n946,
    n585,
    n926,
    n574,
    n611
  );


  xor
  g900
  (
    n963,
    n598,
    n618,
    n603,
    n931
  );


  nand
  g901
  (
    n939,
    n887,
    n930,
    n931
  );


  xor
  g902
  (
    n961,
    n595,
    n623,
    n594,
    n629
  );


  nor
  g903
  (
    n953,
    n931,
    n928,
    n569,
    n620
  );


  xor
  g904
  (
    n938,
    n572,
    n929,
    n623,
    n576
  );


  xnor
  g905
  (
    n941,
    n596,
    n584,
    n888,
    n932
  );


  nand
  g906
  (
    n942,
    n933,
    n926,
    n583,
    n929
  );


  or
  g907
  (
    n952,
    n926,
    n573,
    n886,
    n567
  );


  and
  g908
  (
    n940,
    n606,
    n885,
    n600,
    n884
  );


  nand
  g909
  (
    n964,
    n605,
    n885,
    n579,
    n610
  );


  nand
  g910
  (
    n937,
    n586,
    n928,
    n884,
    n593
  );


  or
  g911
  (
    n947,
    n932,
    n625,
    n930,
    n629
  );


  or
  g912
  (
    n944,
    n590,
    n588,
    n591,
    n577
  );


  nor
  g913
  (
    n951,
    n885,
    n604,
    n933,
    n628
  );


  or
  g914
  (
    n958,
    n566,
    n929,
    n630,
    n587
  );


  nand
  g915
  (
    n935,
    n580,
    n932,
    n589,
    n592
  );


  xor
  g916
  (
    n956,
    n926,
    n884,
    n616,
    n621
  );


  or
  g917
  (
    n936,
    n627,
    n883,
    n927,
    n932
  );


  nor
  g918
  (
    n960,
    n624,
    n622,
    n927,
    n626
  );


  nor
  g919
  (
    n943,
    n887,
    n578,
    n599,
    n625
  );


  xnor
  g920
  (
    n962,
    n931,
    n571,
    n627,
    n612
  );


  or
  g921
  (
    n945,
    n608,
    n628,
    n621,
    n607
  );


  xor
  g922
  (
    n957,
    n622,
    n582,
    n886,
    n927
  );


  or
  g923
  (
    n950,
    n928,
    n886,
    n930,
    n570
  );


  xor
  g924
  (
    n948,
    n619,
    n887,
    n617,
    n927
  );


  nand
  g925
  (
    n954,
    n614,
    n624,
    n581,
    n613
  );


  not
  g926
  (
    n966,
    n935
  );


  buf
  g927
  (
    n981,
    n727
  );


  buf
  g928
  (
    n982,
    n938
  );


  buf
  g929
  (
    n979,
    n937
  );


  buf
  g930
  (
    n976,
    n728
  );


  not
  g931
  (
    n975,
    n939
  );


  buf
  g932
  (
    KeyWire_0_20,
    n728
  );


  not
  g933
  (
    n973,
    n936
  );


  buf
  g934
  (
    n965,
    n728
  );


  buf
  g935
  (
    n972,
    n936
  );


  xnor
  g936
  (
    n977,
    n935,
    n937,
    n630
  );


  xnor
  g937
  (
    n969,
    n936,
    n727
  );


  and
  g938
  (
    n968,
    n937,
    n938,
    n935
  );


  and
  g939
  (
    n970,
    n936,
    n729,
    n631
  );


  or
  g940
  (
    n974,
    n727,
    n938,
    n730
  );


  buf
  g941
  (
    n971,
    n729
  );


  nand
  g942
  (
    n978,
    n939,
    n728,
    n938
  );


  xor
  g943
  (
    n980,
    n730,
    n937,
    n935
  );


  not
  g944
  (
    n1001,
    n777
  );


  not
  g945
  (
    n983,
    n777
  );


  buf
  g946
  (
    n1000,
    n776
  );


  not
  g947
  (
    n993,
    n967
  );


  buf
  g948
  (
    n994,
    n966
  );


  buf
  g949
  (
    n986,
    n779
  );


  buf
  g950
  (
    n997,
    n967
  );


  not
  g951
  (
    n987,
    n970
  );


  buf
  g952
  (
    n988,
    n968
  );


  buf
  g953
  (
    n984,
    n971
  );


  nor
  g954
  (
    n991,
    n967,
    n778,
    n968
  );


  and
  g955
  (
    n996,
    n965,
    n776,
    n777
  );


  xor
  g956
  (
    n989,
    n969,
    n970,
    n774
  );


  nand
  g957
  (
    n999,
    n966,
    n778,
    n775
  );


  or
  g958
  (
    n990,
    n969,
    n779,
    n966
  );


  xnor
  g959
  (
    n985,
    n776,
    n775,
    n969
  );


  nand
  g960
  (
    n992,
    n778,
    n968,
    n774
  );


  nor
  g961
  (
    n998,
    n775,
    n965
  );


  and
  g962
  (
    n995,
    n779,
    n780,
    n970
  );


  nand
  g963
  (
    n1007,
    n892,
    n889,
    n891,
    n996
  );


  xor
  g964
  (
    n1003,
    n890,
    n889,
    n893,
    n1000
  );


  and
  g965
  (
    n1002,
    n888,
    n890,
    n894,
    n889
  );


  and
  g966
  (
    n1005,
    n888,
    n891,
    n1001,
    n892
  );


  nor
  g967
  (
    n1006,
    n893,
    n893,
    n999,
    n998
  );


  xor
  g968
  (
    n1004,
    n997,
    n892,
    n890,
    n891
  );


  buf
  g969
  (
    n1008,
    n1002
  );


  not
  g970
  (
    n1011,
    n1002
  );


  buf
  g971
  (
    n1009,
    n1002
  );


  not
  g972
  (
    n1010,
    n1002
  );


  buf
  g973
  (
    n1012,
    n631
  );


  buf
  g974
  (
    n1013,
    n1008
  );


  xnor
  g975
  (
    n1015,
    n785,
    n781,
    n783,
    n784
  );


  and
  g976
  (
    n1016,
    n1013,
    n781,
    n787
  );


  nand
  g977
  (
    n1020,
    n786,
    n786,
    n783,
    n1013
  );


  xor
  g978
  (
    n1018,
    n783,
    n787,
    n788,
    n785
  );


  or
  g979
  (
    n1017,
    n1013,
    n784,
    n788
  );


  nand
  g980
  (
    n1021,
    n1012,
    n787,
    n782
  );


  xor
  g981
  (
    n1019,
    n1012,
    n1013,
    n782,
    n780
  );


  xnor
  g982
  (
    n1014,
    n786,
    n785,
    n1012
  );


  nand
  g983
  (
    n1022,
    n1014,
    n788
  );


  and
  g984
  (
    n1023,
    n895,
    n1022,
    n894
  );


  xnor
  g985
  (
    n1024,
    n894,
    n895,
    n1022
  );


  xnor
  g986
  (
    n1025,
    n976,
    n976,
    n978,
    n1024
  );


  and
  g987
  (
    n1026,
    n975,
    n973,
    n971,
    n1023
  );


  nand
  g988
  (
    n1032,
    n1024,
    n976,
    n1023
  );


  or
  g989
  (
    n1029,
    n974,
    n972,
    n977,
    n975
  );


  or
  g990
  (
    n1031,
    n972,
    n974,
    n977,
    n971
  );


  xnor
  g991
  (
    n1030,
    n979,
    n975,
    n972,
    n978
  );


  and
  g992
  (
    n1027,
    n974,
    n977,
    n1024
  );


  or
  g993
  (
    n1028,
    n978,
    n973,
    n1023
  );


  buf
  g994
  (
    n1037,
    n1030
  );


  buf
  g995
  (
    n1039,
    n1029
  );


  buf
  g996
  (
    n1041,
    n1032
  );


  buf
  g997
  (
    n1038,
    n1028
  );


  and
  g998
  (
    KeyWire_0_11,
    n1025,
    n1026
  );


  and
  g999
  (
    n1033,
    n1028,
    n1028,
    n1029,
    n1031
  );


  and
  g1000
  (
    n1035,
    n1025,
    n1031,
    n1030
  );


  xor
  g1001
  (
    n1040,
    n1029,
    n1030,
    n1027,
    n789
  );


  nand
  g1002
  (
    n1034,
    n1025,
    n1027,
    n1026
  );


  and
  g1003
  (
    n1048,
    n633,
    n638,
    n1036,
    n1034
  );


  or
  g1004
  (
    n1043,
    n634,
    n633,
    n1034,
    n1035
  );


  xnor
  g1005
  (
    n1046,
    n639,
    n638,
    n637,
    n636
  );


  or
  g1006
  (
    n1047,
    n632,
    n429,
    n636,
    n428
  );


  or
  g1007
  (
    n1044,
    n637,
    n632,
    n1033,
    n640
  );


  or
  g1008
  (
    n1045,
    n634,
    n1035,
    n635,
    n1036
  );


  nor
  g1009
  (
    n1042,
    n639,
    n429,
    n635,
    n428
  );


  xnor
  g1010
  (
    n1049,
    n1042,
    n641,
    n640
  );


  not
  g1011
  (
    n1050,
    n1049
  );


  buf
  g1012
  (
    n1051,
    n1049
  );


  not
  g1013
  (
    n1052,
    n1050
  );


  or
  g1014
  (
    n1055,
    n642,
    n1052,
    n896
  );


  xor
  g1015
  (
    n1053,
    n980,
    n980,
    n1052,
    n979
  );


  and
  g1016
  (
    n1054,
    n979,
    n981,
    n980,
    n642
  );


  not
  g1017
  (
    n1058,
    n1054
  );


  xnor
  g1018
  (
    n1057,
    n430,
    n430,
    n429,
    n431
  );


  nor
  g1019
  (
    n1059,
    n430,
    n1053,
    n432
  );


  and
  g1020
  (
    n1056,
    n430,
    n432,
    n431,
    n429
  );


  nand
  g1021
  (
    n1060,
    n1053,
    n432,
    n431
  );


  xnor
  g1022
  (
    n1061,
    n654,
    n652,
    n653,
    n650
  );


  or
  g1023
  (
    n1068,
    n1060,
    n1059,
    n1056,
    n643
  );


  nor
  g1024
  (
    n1064,
    n652,
    n655,
    n646,
    n651
  );


  xor
  g1025
  (
    n1066,
    n1058,
    n651,
    n1057,
    n647
  );


  or
  g1026
  (
    n1067,
    n1059,
    n648,
    n656,
    n649
  );


  nand
  g1027
  (
    n1069,
    n653,
    n1060,
    n654
  );


  nand
  g1028
  (
    KeyWire_0_17,
    n643,
    n649,
    n648,
    n645
  );


  nor
  g1029
  (
    n1062,
    n650,
    n644,
    n647
  );


  nand
  g1030
  (
    n1065,
    n645,
    n646,
    n1060,
    n655
  );


  buf
  g1031
  (
    n1071,
    n1061
  );


  not
  g1032
  (
    n1072,
    n1062
  );


  xnor
  g1033
  (
    n1073,
    n1051,
    n1063
  );


  xor
  g1034
  (
    n1070,
    n1050,
    n1064,
    n1051
  );


  or
  g1035
  (
    n1076,
    n791,
    n789,
    n790
  );


  xnor
  g1036
  (
    KeyWire_0_26,
    n1071,
    n1072,
    n789,
    n792
  );


  nand
  g1037
  (
    n1074,
    n790,
    n1070,
    n791
  );


  and
  g1038
  (
    n1081,
    n1065,
    n902,
    n1075
  );


  nand
  g1039
  (
    n1085,
    n898,
    n901,
    n1074
  );


  xor
  g1040
  (
    n1078,
    n904,
    n1075,
    n900
  );


  xor
  g1041
  (
    n1083,
    n899,
    n904,
    n900
  );


  and
  g1042
  (
    n1080,
    n899,
    n905,
    n896,
    n1076
  );


  nor
  g1043
  (
    n1084,
    n903,
    n905,
    n899,
    n898
  );


  or
  g1044
  (
    n1086,
    n1074,
    n1076,
    n897
  );


  nand
  g1045
  (
    n1082,
    n1076,
    n901,
    n897,
    n1074
  );


  nor
  g1046
  (
    n1079,
    n897,
    n898,
    n896,
    n903
  );


  xnor
  g1047
  (
    n1077,
    n902,
    n905,
    n900,
    n903
  );


  buf
  g1048
  (
    n1088,
    n1086
  );


  not
  g1049
  (
    n1087,
    n1085
  );


  and
  g1050
  (
    n1089,
    n1087,
    n1088,
    n35
  );


  or
  g1051
  (
    n1092,
    n37,
    n38,
    n36,
    n1088
  );


  nor
  g1052
  (
    n1093,
    n38,
    n36,
    n35
  );


  xnor
  g1053
  (
    n1091,
    n35,
    n1088,
    n36,
    n37
  );


  xor
  g1054
  (
    n1090,
    n1087,
    n37,
    n38
  );


  nand
  g1055
  (
    n1110,
    n1055,
    n732,
    n1045
  );


  and
  g1056
  (
    n1105,
    n1047,
    n731,
    n1048,
    n1091
  );


  or
  g1057
  (
    n1108,
    n1046,
    n123,
    n732,
    n1044
  );


  xor
  g1058
  (
    n1095,
    n735,
    n1042,
    n734,
    n123
  );


  nor
  g1059
  (
    n1111,
    n1091,
    n735,
    n733
  );


  xnor
  g1060
  (
    n1102,
    n736,
    n124,
    n1092,
    n731
  );


  nand
  g1061
  (
    n1106,
    n1055,
    n124,
    n733,
    n1090
  );


  nand
  g1062
  (
    n1098,
    n124,
    n1048,
    n736
  );


  or
  g1063
  (
    n1094,
    n1093,
    n731,
    n1090,
    n1043
  );


  and
  g1064
  (
    n1101,
    n1045,
    n1091,
    n730,
    n1089
  );


  xnor
  g1065
  (
    n1097,
    n732,
    n1049,
    n38,
    n735
  );


  and
  g1066
  (
    n1113,
    n734,
    n1091,
    n1093,
    n1046
  );


  xor
  g1067
  (
    n1107,
    n1089,
    n1093,
    n1043
  );


  xor
  g1068
  (
    n1104,
    n1044,
    n1092,
    n736,
    n1042
  );


  xor
  g1069
  (
    n1109,
    n730,
    n1045,
    n736,
    n1089
  );


  xor
  g1070
  (
    n1103,
    n1090,
    n1047,
    n733,
    n1089
  );


  nand
  g1071
  (
    n1099,
    n1092,
    n1073,
    n1044,
    n1048
  );


  nor
  g1072
  (
    n1100,
    n124,
    n735,
    n1054,
    n734
  );


  xor
  g1073
  (
    n1112,
    n1092,
    n1046,
    n731,
    n1090
  );


  nor
  g1074
  (
    n1096,
    n1055,
    n1047,
    n734,
    n1043
  );


  nand
  g1075
  (
    n1127,
    n1095,
    n440
  );


  nor
  g1076
  (
    n1114,
    n439,
    n434,
    n437,
    n433
  );


  and
  g1077
  (
    n1123,
    n1098,
    n437,
    n438,
    n439
  );


  nand
  g1078
  (
    n1117,
    n436,
    n433,
    n435,
    n434
  );


  xnor
  g1079
  (
    KeyWire_0_31,
    n434,
    n437,
    n442,
    n435
  );


  xor
  g1080
  (
    n1120,
    n1095,
    n440,
    n1098,
    n442
  );


  nor
  g1081
  (
    n1128,
    n1094,
    n436,
    n439,
    n1097
  );


  or
  g1082
  (
    n1118,
    n1095,
    n441
  );


  nor
  g1083
  (
    n1125,
    n435,
    n442,
    n1094,
    n433
  );


  nand
  g1084
  (
    n1116,
    n433,
    n1094,
    n438,
    n440
  );


  xor
  g1085
  (
    n1121,
    n1097,
    n441,
    n436,
    n1098
  );


  nor
  g1086
  (
    n1122,
    n438,
    n442,
    n440,
    n437
  );


  and
  g1087
  (
    n1119,
    n1096,
    n1096,
    n435,
    n443
  );


  and
  g1088
  (
    n1115,
    n439,
    n1097,
    n436,
    n434
  );


  and
  g1089
  (
    KeyWire_0_25,
    n432,
    n443,
    n438,
    n1096
  );


  and
  g1090
  (
    n1130,
    n656,
    n657,
    n658
  );


  and
  g1091
  (
    n1129,
    n1114,
    n1114,
    n658,
    n659
  );


  xnor
  g1092
  (
    n1138,
    n737,
    n742,
    n1129,
    n1130
  );


  and
  g1093
  (
    n1132,
    n737,
    n738,
    n739,
    n740
  );


  or
  g1094
  (
    n1134,
    n738,
    n740,
    n1130
  );


  nand
  g1095
  (
    n1137,
    n742,
    n739,
    n1129,
    n741
  );


  or
  g1096
  (
    n1133,
    n737,
    n741,
    n740
  );


  xnor
  g1097
  (
    n1131,
    n740,
    n1129,
    n738,
    n741
  );


  and
  g1098
  (
    n1136,
    n742,
    n1129,
    n739,
    n1130
  );


  xnor
  g1099
  (
    n1135,
    n737,
    n739,
    n742,
    n738
  );


  buf
  g1100
  (
    n1139,
    n1138
  );


  not
  g1101
  (
    n1141,
    n1139
  );


  not
  g1102
  (
    n1140,
    n1139
  );


  or
  g1103
  (
    n1142,
    n1068,
    n1067,
    n1066
  );


  nor
  g1104
  (
    n1145,
    n1068,
    n1140
  );


  xor
  g1105
  (
    n1143,
    n1068,
    n1069,
    n1067
  );


  and
  g1106
  (
    n1144,
    n1067,
    n1066,
    n1140,
    n1069
  );


  not
  g1107
  (
    n1150,
    n1143
  );


  not
  g1108
  (
    n1149,
    n1145
  );


  not
  g1109
  (
    n1148,
    n660
  );


  buf
  g1110
  (
    n1152,
    n661
  );


  and
  g1111
  (
    n1151,
    n662,
    n1143,
    n1144,
    n661
  );


  and
  g1112
  (
    n1146,
    n1145,
    n660,
    n659,
    n1144
  );


  nor
  g1113
  (
    n1147,
    n662,
    n663,
    n1142
  );


  xnor
  g1114
  (
    n1169,
    n982,
    n906,
    n1105,
    n1110
  );


  nor
  g1115
  (
    n1162,
    n1149,
    n913,
    n1103,
    n1105
  );


  xor
  g1116
  (
    n1179,
    n1102,
    n1147,
    n1152,
    n1148
  );


  and
  g1117
  (
    n1178,
    n1152,
    n911,
    n1146,
    n1103
  );


  nor
  g1118
  (
    n1164,
    n1108,
    n1147,
    n907,
    n915
  );


  or
  g1119
  (
    n1168,
    n908,
    n1146,
    n925
  );


  nor
  g1120
  (
    n1173,
    n1112,
    n1151,
    n1149,
    n1150
  );


  and
  g1121
  (
    n1155,
    n909,
    n1109,
    n912,
    n1141
  );


  or
  g1122
  (
    n1160,
    n1099,
    n1104,
    n908,
    n913
  );


  nand
  g1123
  (
    n1157,
    n909,
    n1148,
    n1106,
    n914
  );


  nand
  g1124
  (
    n1161,
    n1148,
    n925,
    n1109,
    n906
  );


  or
  g1125
  (
    n1176,
    n1113,
    n1141,
    n1112,
    n1102
  );


  and
  g1126
  (
    n1180,
    n911,
    n1150,
    n981,
    n1147
  );


  and
  g1127
  (
    n1156,
    n1104,
    n1113,
    n1151,
    n981
  );


  xor
  g1128
  (
    n1177,
    n1105,
    n1113,
    n907,
    n1146
  );


  nor
  g1129
  (
    n1170,
    n1151,
    n1111,
    n1100,
    n1099
  );


  xnor
  g1130
  (
    n1171,
    n913,
    n1102,
    n1150,
    n1107
  );


  or
  g1131
  (
    n1172,
    n1110,
    n914,
    n1106,
    n1111
  );


  or
  g1132
  (
    n1174,
    n911,
    n910,
    n1108,
    n1101
  );


  xor
  g1133
  (
    n1153,
    n1103,
    n1101,
    n909,
    n1141
  );


  xnor
  g1134
  (
    n1154,
    n1141,
    n1149,
    n1106,
    n1109
  );


  nor
  g1135
  (
    n1158,
    n1112,
    n1150,
    n910,
    n1152
  );


  and
  g1136
  (
    n1166,
    n906,
    n1149,
    n1100,
    n1146
  );


  or
  g1137
  (
    n1175,
    n910,
    n912,
    n914,
    n1110
  );


  nor
  g1138
  (
    n1163,
    n1148,
    n1107,
    n912,
    n1104
  );


  or
  g1139
  (
    n1165,
    n1151,
    n908,
    n1147,
    n1100
  );


  xor
  g1140
  (
    n1159,
    n982,
    n1108,
    n1111,
    n907
  );


  nor
  g1141
  (
    n1167,
    n1107,
    n1101,
    n1099,
    n1152
  );


  or
  g1142
  (
    n1187,
    n832,
    n1116,
    n1157,
    n813
  );


  xor
  g1143
  (
    n1286,
    n858,
    n874,
    n668,
    n1119
  );


  or
  g1144
  (
    n1211,
    n1167,
    n1127,
    n850,
    n809
  );


  nand
  g1145
  (
    KeyWire_0_8,
    n834,
    n1128,
    n874,
    n823
  );


  and
  g1146
  (
    n1196,
    n843,
    n1155,
    n1170,
    n1121
  );


  or
  g1147
  (
    n1242,
    n1122,
    n812,
    n829,
    n843
  );


  xor
  g1148
  (
    n1277,
    n1169,
    n829,
    n1126,
    n845
  );


  or
  g1149
  (
    n1214,
    n870,
    n828,
    n1171
  );


  nand
  g1150
  (
    n1195,
    n845,
    n852,
    n849,
    n669
  );


  xor
  g1151
  (
    n1273,
    n878,
    n842,
    n820,
    n831
  );


  xor
  g1152
  (
    n1215,
    n861,
    n835,
    n838,
    n805
  );


  or
  g1153
  (
    n1269,
    n1118,
    n1159,
    n823,
    n836
  );


  and
  g1154
  (
    n1276,
    n837,
    n1160,
    n1179,
    n875
  );


  xnor
  g1155
  (
    n1239,
    n820,
    n879,
    n831,
    n1157
  );


  nor
  g1156
  (
    n1270,
    n827,
    n818,
    n1124,
    n1167
  );


  xor
  g1157
  (
    n1264,
    n856,
    n1121,
    n1176,
    n818
  );


  and
  g1158
  (
    n1223,
    n1166,
    n811,
    n1165,
    n1178
  );


  nand
  g1159
  (
    n1181,
    n1173,
    n877,
    n1158,
    n1127
  );


  xor
  g1160
  (
    n1250,
    n872,
    n668,
    n870,
    n863
  );


  xor
  g1161
  (
    n1197,
    n799,
    n834,
    n839,
    n1155
  );


  xnor
  g1162
  (
    n1237,
    n862,
    n1157,
    n818,
    n872
  );


  xor
  g1163
  (
    n1226,
    n798,
    n837,
    n802,
    n1179
  );


  and
  g1164
  (
    n1288,
    n1165,
    n841,
    n855,
    n847
  );


  xnor
  g1165
  (
    n1228,
    n842,
    n1118,
    n876,
    n857
  );


  nand
  g1166
  (
    n1282,
    n807,
    n669,
    n817,
    n809
  );


  nand
  g1167
  (
    n1240,
    n794,
    n667,
    n811,
    n1163
  );


  and
  g1168
  (
    n1188,
    n803,
    n1180,
    n1178,
    n1156
  );


  xnor
  g1169
  (
    n1259,
    n1166,
    n797,
    n793,
    n870
  );


  and
  g1170
  (
    n1190,
    n858,
    n815,
    n1123,
    n1125
  );


  nand
  g1171
  (
    n1281,
    n1120,
    n1120,
    n815,
    n807
  );


  or
  g1172
  (
    n1201,
    n855,
    n838,
    n826,
    n808
  );


  nor
  g1173
  (
    n1207,
    n812,
    n1158,
    n815,
    n866
  );


  or
  g1174
  (
    n1229,
    n1172,
    n1176,
    n793,
    n840
  );


  xnor
  g1175
  (
    n1262,
    n872,
    n1168,
    n671,
    n1153
  );


  xor
  g1176
  (
    n1283,
    n1115,
    n1173,
    n873,
    n878
  );


  or
  g1177
  (
    n1291,
    n844,
    n810,
    n868,
    n1158
  );


  nand
  g1178
  (
    n1209,
    n848,
    n1171,
    n869,
    n804
  );


  nand
  g1179
  (
    n1184,
    n853,
    n1117,
    n860,
    n1173
  );


  xor
  g1180
  (
    n1183,
    n1162,
    n1174,
    n851,
    n1179
  );


  nand
  g1181
  (
    n1234,
    n831,
    n801,
    n802,
    n851
  );


  xnor
  g1182
  (
    n1292,
    n1178,
    n873,
    n1170,
    n859
  );


  xnor
  g1183
  (
    n1274,
    n667,
    n1171,
    n824,
    n866
  );


  nand
  g1184
  (
    n1265,
    n1124,
    n1114,
    n838,
    n822
  );


  or
  g1185
  (
    n1222,
    n1122,
    n1180,
    n816,
    n846
  );


  and
  g1186
  (
    n1268,
    n803,
    n825,
    n1117,
    n675
  );


  xor
  g1187
  (
    n1224,
    n871,
    n934,
    n868,
    n1177
  );


  xnor
  g1188
  (
    n1266,
    n846,
    n814,
    n867,
    n1174
  );


  and
  g1189
  (
    n1186,
    n852,
    n1154,
    n1156,
    n873
  );


  xnor
  g1190
  (
    n1202,
    n835,
    n878,
    n879,
    n1159
  );


  and
  g1191
  (
    n1235,
    n1161,
    n1162,
    n836,
    n1177
  );


  nand
  g1192
  (
    n1199,
    n861,
    n1166,
    n664,
    n806
  );


  xnor
  g1193
  (
    n1263,
    n1168,
    n1161,
    n862,
    n856
  );


  xnor
  g1194
  (
    n1203,
    n826,
    n1154,
    n839,
    n1173
  );


  nor
  g1195
  (
    n1253,
    n830,
    n674,
    n833,
    n816
  );


  nor
  g1196
  (
    n1252,
    n794,
    n875,
    n877,
    n671
  );


  xnor
  g1197
  (
    n1213,
    n1163,
    n853,
    n796,
    n670
  );


  nand
  g1198
  (
    n1246,
    n1159,
    n821,
    n853,
    n1175
  );


  xor
  g1199
  (
    n1220,
    n1164,
    n825,
    n811,
    n1155
  );


  nor
  g1200
  (
    n1285,
    n1162,
    n828,
    n1163,
    n794
  );


  xnor
  g1201
  (
    n1256,
    n817,
    n856,
    n850,
    n869
  );


  xnor
  g1202
  (
    n1245,
    n1165,
    n1167,
    n673,
    n1123
  );


  or
  g1203
  (
    n1231,
    n1170,
    n1125,
    n805,
    n1172
  );


  nor
  g1204
  (
    n1267,
    n798,
    n1120,
    n855,
    n1157
  );


  or
  g1205
  (
    n1289,
    n810,
    n796,
    n819,
    n857
  );


  nand
  g1206
  (
    n1279,
    n1161,
    n1166,
    n1160,
    n1169
  );


  xnor
  g1207
  (
    n1227,
    n841,
    n1121,
    n1125,
    n837
  );


  nor
  g1208
  (
    n1208,
    n845,
    n1159,
    n808,
    n675
  );


  nor
  g1209
  (
    n1247,
    n847,
    n804,
    n824,
    n830
  );


  and
  g1210
  (
    n1189,
    n1165,
    n800,
    n1160,
    n808
  );


  xor
  g1211
  (
    n1255,
    n1177,
    n859,
    n1164,
    n812
  );


  xor
  g1212
  (
    n1272,
    n672,
    n800,
    n830,
    n871
  );


  or
  g1213
  (
    n1271,
    n1179,
    n1175,
    n799,
    n849
  );


  nor
  g1214
  (
    n1218,
    n665,
    n851,
    n1154,
    n876
  );


  xnor
  g1215
  (
    n1200,
    n840,
    n825,
    n805,
    n814
  );


  nor
  g1216
  (
    n1192,
    n840,
    n817,
    n858,
    n819
  );


  nand
  g1217
  (
    n1210,
    n826,
    n1117,
    n824,
    n1115
  );


  xnor
  g1218
  (
    n1221,
    n792,
    n860,
    n1168,
    n1128
  );


  or
  g1219
  (
    n1284,
    n1126,
    n664,
    n665,
    n933
  );


  xor
  g1220
  (
    n1198,
    n1160,
    n848,
    n1168,
    n800
  );


  nor
  g1221
  (
    n1290,
    n1156,
    n846,
    n1170,
    n864
  );


  or
  g1222
  (
    n1217,
    n803,
    n1162,
    n670,
    n934
  );


  xor
  g1223
  (
    n1248,
    n666,
    n834,
    n797,
    n934
  );


  xor
  g1224
  (
    n1194,
    n1177,
    n833,
    n876,
    n804
  );


  nor
  g1225
  (
    n1243,
    n822,
    n865,
    n857,
    n859
  );


  or
  g1226
  (
    n1233,
    n1176,
    n1127,
    n867,
    n801
  );


  nor
  g1227
  (
    n1206,
    n1115,
    n868,
    n844,
    n934
  );


  nand
  g1228
  (
    n1232,
    n821,
    n1172,
    n832,
    n813
  );


  nor
  g1229
  (
    n1258,
    n666,
    n809,
    n1163,
    n820
  );


  xnor
  g1230
  (
    n1254,
    n814,
    n864,
    n797,
    n1153
  );


  nand
  g1231
  (
    n1287,
    n860,
    n844,
    n1118,
    n827
  );


  or
  g1232
  (
    n1244,
    n1171,
    n854,
    n673,
    n1122
  );


  xnor
  g1233
  (
    n1275,
    n841,
    n795,
    n862,
    n810
  );


  xor
  g1234
  (
    n1219,
    n822,
    n874,
    n1126,
    n1169
  );


  and
  g1235
  (
    n1191,
    n1161,
    n1154,
    n863,
    n1167
  );


  xor
  g1236
  (
    n1212,
    n827,
    n799,
    n848,
    n813
  );


  xnor
  g1237
  (
    n1225,
    n871,
    n1124,
    n806,
    n1172
  );


  and
  g1238
  (
    n1230,
    n842,
    n1164,
    n792,
    n802
  );


  xor
  g1239
  (
    n1216,
    n801,
    n1178,
    n1128,
    n1180
  );


  xor
  g1240
  (
    n1261,
    n1116,
    n816,
    n829,
    n854
  );


  nand
  g1241
  (
    n1238,
    n875,
    n1175,
    n798,
    n821
  );


  nand
  g1242
  (
    n1182,
    n879,
    n865,
    n1175,
    n839
  );


  nor
  g1243
  (
    n1280,
    n793,
    n863,
    n823,
    n877
  );


  xor
  g1244
  (
    n1185,
    n795,
    n869,
    n1174,
    n1116
  );


  or
  g1245
  (
    n1257,
    n843,
    n852,
    n854,
    n861
  );


  or
  g1246
  (
    n1249,
    n865,
    n1119,
    n806,
    n1153
  );


  xnor
  g1247
  (
    n1278,
    n867,
    n836,
    n864,
    n849
  );


  or
  g1248
  (
    n1193,
    n835,
    n1153,
    n674,
    n850
  );


  xor
  g1249
  (
    n1260,
    n819,
    n672,
    n1176,
    n866
  );


  xor
  g1250
  (
    n1236,
    n807,
    n833,
    n1158,
    n1180
  );


  or
  g1251
  (
    n1204,
    n1119,
    n795,
    n1174,
    n847
  );


  nand
  g1252
  (
    n1205,
    n1156,
    n1169,
    n832,
    n796
  );


  nor
  g1253
  (
    n1251,
    n1155,
    n1123,
    n933,
    n1164
  );


  nor
  g1254
  (
    n1317,
    n1269,
    n1196,
    n954,
    n949
  );


  and
  g1255
  (
    n1335,
    n1216,
    n1189,
    n1190,
    n959
  );


  nand
  g1256
  (
    n1366,
    n1258,
    n963,
    n953,
    n1238
  );


  xnor
  g1257
  (
    n1386,
    n1236,
    n1222,
    n958,
    n1231
  );


  xnor
  g1258
  (
    n1323,
    n1199,
    n1203,
    n1192,
    n1254
  );


  xor
  g1259
  (
    n1352,
    n1211,
    n1246,
    n957,
    n1237
  );


  or
  g1260
  (
    n1296,
    n952,
    n1191,
    n1264,
    n1253
  );


  xnor
  g1261
  (
    n1385,
    n1217,
    n1201,
    n1200,
    n1237
  );


  nor
  g1262
  (
    n1380,
    n963,
    n1245,
    n947,
    n945
  );


  nand
  g1263
  (
    n1315,
    n1198,
    n1219,
    n1257,
    n1266
  );


  xnor
  g1264
  (
    n1339,
    n1197,
    n1194,
    n953,
    n1196
  );


  and
  g1265
  (
    n1375,
    n1274,
    n1232,
    n946,
    n1240
  );


  xnor
  g1266
  (
    n1318,
    n1259,
    n1223,
    n1191,
    n1195
  );


  nor
  g1267
  (
    n1320,
    n1267,
    n1249,
    n1226,
    n1197
  );


  and
  g1268
  (
    n1332,
    n947,
    n948,
    n1257,
    n1279
  );


  xnor
  g1269
  (
    n1326,
    n954,
    n1244,
    n1201,
    n1252
  );


  nand
  g1270
  (
    n1354,
    n1236,
    n1193,
    n948,
    n944
  );


  xor
  g1271
  (
    n1294,
    n1274,
    n1189,
    n947,
    n1210
  );


  xnor
  g1272
  (
    n1301,
    n1210,
    n1218,
    n962,
    n1209
  );


  nand
  g1273
  (
    n1378,
    n1255,
    n1253,
    n1266,
    n956
  );


  nand
  g1274
  (
    n1293,
    n1273,
    n960,
    n1227,
    n1212
  );


  nand
  g1275
  (
    n1334,
    n1263,
    n957,
    n1267,
    n948
  );


  xor
  g1276
  (
    n1356,
    n953,
    n964,
    n945,
    n1242
  );


  xor
  g1277
  (
    n1329,
    n1218,
    n1250,
    n956,
    n942
  );


  nor
  g1278
  (
    n1312,
    n1236,
    n1206,
    n1268,
    n963
  );


  nor
  g1279
  (
    n1363,
    n1272,
    n1225,
    n1204,
    n1261
  );


  and
  g1280
  (
    n1316,
    n1231,
    n1232,
    n1196,
    n961
  );


  xor
  g1281
  (
    n1304,
    n1270,
    n1201,
    n1277,
    n1227
  );


  or
  g1282
  (
    n1365,
    n960,
    n1234,
    n1226,
    n949
  );


  xnor
  g1283
  (
    n1377,
    n1202,
    n1229
  );


  nor
  g1284
  (
    n1344,
    n1260,
    n958,
    n957,
    n945
  );


  or
  g1285
  (
    n1343,
    n1213,
    n956,
    n1265,
    n952
  );


  nand
  g1286
  (
    n1349,
    n1184,
    n1248,
    n940,
    n1186
  );


  xor
  g1287
  (
    n1361,
    n1229,
    n950,
    n944,
    n1242
  );


  xnor
  g1288
  (
    n1348,
    n1203,
    n1220,
    n1228,
    n1271
  );


  and
  g1289
  (
    n1303,
    n961,
    n1254,
    n1275,
    n1212
  );


  nor
  g1290
  (
    n1370,
    n1187,
    n942,
    n1228,
    n1233
  );


  and
  g1291
  (
    n1362,
    n1251,
    n1235,
    n954,
    n1209
  );


  xnor
  g1292
  (
    n1298,
    n945,
    n1256,
    n1264,
    n1203
  );


  nor
  g1293
  (
    n1387,
    n1193,
    n1205,
    n939,
    n1255
  );


  or
  g1294
  (
    n1364,
    n1205,
    n1276,
    n1262,
    n946
  );


  xor
  g1295
  (
    n1371,
    n1249,
    n943,
    n1212,
    n956
  );


  and
  g1296
  (
    n1297,
    n955,
    n1263,
    n1199,
    n1183
  );


  and
  g1297
  (
    n1360,
    n960,
    n1268,
    n1262,
    n1225
  );


  xor
  g1298
  (
    n1359,
    n951,
    n1261,
    n1218,
    n1259
  );


  xor
  g1299
  (
    n1383,
    n955,
    n1279,
    n1254,
    n950
  );


  xor
  g1300
  (
    n1372,
    n962,
    n1221,
    n1217,
    n1276
  );


  nor
  g1301
  (
    n1357,
    n1208,
    n964,
    n1270,
    n1279
  );


  nand
  g1302
  (
    n1305,
    n1216,
    n960,
    n1247,
    n1202
  );


  xnor
  g1303
  (
    n1382,
    n1256,
    n1207,
    n1224,
    n951
  );


  xnor
  g1304
  (
    n1358,
    n1246,
    n952,
    n1258,
    n1233
  );


  or
  g1305
  (
    n1327,
    n1206,
    n944,
    n962,
    n1198
  );


  xor
  g1306
  (
    n1353,
    n1269,
    n1239,
    n1273
  );


  xnor
  g1307
  (
    n1330,
    n1241,
    n943,
    n1259,
    n946
  );


  or
  g1308
  (
    n1342,
    n1192,
    n1239,
    n946,
    n961
  );


  and
  g1309
  (
    n1345,
    n1219,
    n1195,
    n1265,
    n1227
  );


  xnor
  g1310
  (
    n1347,
    n1266,
    n955,
    n943,
    n1239
  );


  xnor
  g1311
  (
    n1299,
    n941,
    n1240,
    n1222,
    n953
  );


  or
  g1312
  (
    n1341,
    n1257,
    n1213,
    n1270,
    n942
  );


  xor
  g1313
  (
    n1311,
    n1246,
    n1219,
    n1278,
    n1205
  );


  xor
  g1314
  (
    n1346,
    n1217,
    n1197,
    n1243,
    n1238
  );


  or
  g1315
  (
    n1328,
    n1275,
    n1247,
    n1265,
    n1200
  );


  nand
  g1316
  (
    n1369,
    n1260,
    n1249,
    n1272,
    n1220
  );


  or
  g1317
  (
    n1355,
    n1261,
    n1263,
    n951,
    n1244
  );


  xor
  g1318
  (
    n1314,
    n1280,
    n942,
    n951,
    n961
  );


  or
  g1319
  (
    n1307,
    n1211,
    n1188,
    n1274,
    n1216
  );


  or
  g1320
  (
    n1374,
    n1235,
    n949,
    n1243
  );


  nor
  g1321
  (
    n1302,
    n1234,
    n959,
    n1269,
    n1235
  );


  nor
  g1322
  (
    n1350,
    n948,
    n1238,
    n941,
    n1210
  );


  or
  g1323
  (
    n1308,
    n950,
    n1278,
    n963,
    n1230
  );


  and
  g1324
  (
    n1313,
    n1213,
    n964,
    n1225,
    n1240
  );


  xnor
  g1325
  (
    n1309,
    n1233,
    n1231,
    n1208,
    n1262
  );


  nor
  g1326
  (
    n1340,
    n1258,
    n1275,
    n944,
    n1230
  );


  xor
  g1327
  (
    n1373,
    n1272,
    n1267,
    n1250,
    n1230
  );


  and
  g1328
  (
    n1381,
    n1215,
    n1215,
    n1214,
    n1271
  );


  or
  g1329
  (
    n1319,
    n962,
    n1208,
    n1181,
    n1255
  );


  xnor
  g1330
  (
    n1331,
    n952,
    n940,
    n1251
  );


  nand
  g1331
  (
    n1376,
    n947,
    n1185,
    n1253,
    n1204
  );


  nand
  g1332
  (
    n1336,
    n955,
    n1199,
    n1245
  );


  nand
  g1333
  (
    n1310,
    n1237,
    n1209,
    n1226,
    n941
  );


  xor
  g1334
  (
    n1325,
    n1232,
    n1182,
    n1276,
    n1242
  );


  nand
  g1335
  (
    n1379,
    n1280,
    n1211,
    n1247,
    n959
  );


  xor
  g1336
  (
    n1384,
    n1221,
    n957,
    n1277,
    n940
  );


  xor
  g1337
  (
    n1351,
    n1223,
    n1224,
    n1207,
    n1220
  );


  xor
  g1338
  (
    n1333,
    n1198,
    n1251,
    n1271,
    n1215
  );


  xor
  g1339
  (
    n1324,
    n1206,
    n1264,
    n1195,
    n1200
  );


  xnor
  g1340
  (
    n1367,
    n943,
    n954,
    n1241,
    n950
  );


  xor
  g1341
  (
    n1368,
    n958,
    n1188,
    n1243,
    n1252
  );


  or
  g1342
  (
    n1300,
    n1244,
    n959,
    n1250,
    n958
  );


  nor
  g1343
  (
    n1306,
    n1204,
    n1252,
    n1214,
    n1221
  );


  nand
  g1344
  (
    n1322,
    n1234,
    n1207,
    n1241,
    n1214
  );


  xor
  g1345
  (
    n1295,
    n964,
    n1256,
    n1277,
    n1194
  );


  xor
  g1346
  (
    n1338,
    n1228,
    n1222,
    n1278,
    n1190
  );


  xor
  g1347
  (
    n1321,
    n1260,
    n941,
    n1223,
    n1224
  );


  nor
  g1348
  (
    n1337,
    n1268,
    n1248,
    n939
  );


  nand
  g1349
  (
    n1388,
    n982,
    n1293
  );


  nor
  g1350
  (
    n1390,
    n676,
    n1388
  );


  nor
  g1351
  (
    n1389,
    n1388,
    n676
  );


  nor
  g1352
  (
    n1396,
    n1003,
    n1003,
    n1004,
    n1390
  );


  nand
  g1353
  (
    n1391,
    n1006,
    n1005,
    n1004
  );


  and
  g1354
  (
    n1397,
    n1389,
    n1004,
    n1390,
    n1005
  );


  nor
  g1355
  (
    n1398,
    n1007,
    n1296,
    n1390,
    n1005
  );


  nor
  g1356
  (
    n1395,
    n1294,
    n1006,
    n1003,
    n1389
  );


  nand
  g1357
  (
    n1394,
    n1389,
    n1007,
    n1390
  );


  nor
  g1358
  (
    n1393,
    n1389,
    n1003,
    n1006
  );


  xnor
  g1359
  (
    n1392,
    n1007,
    n1005,
    n1297,
    n1295
  );


  xor
  g1360
  (
    n1414,
    n1283,
    n1284,
    n1303,
    n1011
  );


  nand
  g1361
  (
    n1421,
    n1313,
    n677,
    n1311,
    n1010
  );


  nor
  g1362
  (
    n1409,
    n1010,
    n1009,
    n1395,
    n1290
  );


  xnor
  g1363
  (
    KeyWire_0_16,
    n1011,
    n1291,
    n1396,
    n1392
  );


  or
  g1364
  (
    n1419,
    n1283,
    n1302,
    n1009,
    n1395
  );


  xor
  g1365
  (
    n1416,
    n1304,
    n1392,
    n1397,
    n1286
  );


  nand
  g1366
  (
    n1399,
    n1282,
    n1393,
    n1287
  );


  nand
  g1367
  (
    n1422,
    n1299,
    n1305,
    n1309,
    n1281
  );


  nor
  g1368
  (
    n1405,
    n1282,
    n677,
    n1310,
    n1285
  );


  nand
  g1369
  (
    n1403,
    n1397,
    n1008,
    n1391,
    n1394
  );


  nor
  g1370
  (
    n1418,
    n1292,
    n1280,
    n1394,
    n1009
  );


  nor
  g1371
  (
    n1408,
    n1308,
    n1391,
    n1301
  );


  nand
  g1372
  (
    n1412,
    n1287,
    n1282,
    n1396
  );


  and
  g1373
  (
    n1415,
    n1397,
    n1288,
    n1300,
    n1292
  );


  nand
  g1374
  (
    n1401,
    n1290,
    n1011,
    n1288
  );


  nor
  g1375
  (
    n1402,
    n1394,
    n1281,
    n1010,
    n1009
  );


  xor
  g1376
  (
    n1407,
    n1314,
    n1286,
    n1008,
    n1398
  );


  xnor
  g1377
  (
    n1413,
    n1289,
    n1306,
    n1315,
    n1312
  );


  nor
  g1378
  (
    n1417,
    n1287,
    n1283,
    n1289,
    n1307
  );


  or
  g1379
  (
    n1410,
    n678,
    n1285,
    n1291,
    n1398
  );


  xnor
  g1380
  (
    n1404,
    n1010,
    n1395,
    n1298,
    n1281
  );


  nand
  g1381
  (
    n1411,
    n1286,
    n1284,
    n1398
  );


  xnor
  g1382
  (
    n1420,
    n1392,
    n1288,
    n1291,
    n678
  );


  nor
  g1383
  (
    n1400,
    n1393,
    n1290,
    n1289,
    n1285
  );


  not
  g1384
  (
    n1430,
    n1345
  );


  and
  g1385
  (
    n1435,
    n1407,
    n1341,
    n1404,
    n1356
  );


  xor
  g1386
  (
    n1423,
    n1355,
    n1403,
    n1326,
    n1323
  );


  nand
  g1387
  (
    n1424,
    n1327,
    n1410,
    n1332,
    n1357
  );


  xnor
  g1388
  (
    n1437,
    n1412,
    n1411,
    n1330,
    n1317
  );


  or
  g1389
  (
    n1432,
    n1316,
    n1324,
    n1401,
    n1320
  );


  and
  g1390
  (
    KeyWire_0_23,
    n1335,
    n1318,
    n1344,
    n1346
  );


  and
  g1391
  (
    n1434,
    n1405,
    n1410,
    n1408,
    n1351
  );


  nand
  g1392
  (
    n1429,
    n1410,
    n1412,
    n1338,
    n1340
  );


  xnor
  g1393
  (
    n1426,
    n1333,
    n1321,
    n1411,
    n1349
  );


  nand
  g1394
  (
    n1431,
    n1348,
    n1337,
    n1319,
    n1328
  );


  nor
  g1395
  (
    n1436,
    n1352,
    n1411,
    n1334,
    n1350
  );


  xnor
  g1396
  (
    n1427,
    n1409,
    n1336,
    n1331,
    n1343
  );


  xor
  g1397
  (
    n1425,
    n1339,
    n1329,
    n1342,
    n1402
  );


  nor
  g1398
  (
    n1433,
    n1322,
    n1353,
    n1325,
    n1412
  );


  and
  g1399
  (
    n1428,
    n1354,
    n1413,
    n1347,
    n1406
  );


  xnor
  g1400
  (
    n1446,
    n917,
    n1425,
    n1429,
    n1415
  );


  xor
  g1401
  (
    KeyWire_0_14,
    n1016,
    n916,
    n1427,
    n1015
  );


  nor
  g1402
  (
    n1450,
    n1021,
    n1020,
    n444,
    n880
  );


  nor
  g1403
  (
    n1445,
    n1017,
    n1014,
    n1416,
    n919
  );


  xnor
  g1404
  (
    n1439,
    n1437,
    n444,
    n1413,
    n1436
  );


  xor
  g1405
  (
    n1443,
    n443,
    n1363,
    n882,
    n1014
  );


  or
  g1406
  (
    n1444,
    n1434,
    n1413,
    n1438,
    n1437
  );


  nand
  g1407
  (
    n1463,
    n443,
    n1015,
    n1414,
    n444
  );


  or
  g1408
  (
    n1466,
    n1018,
    n915,
    n1425,
    n1417
  );


  nor
  g1409
  (
    n1451,
    n1016,
    n1427,
    n1424,
    n1432
  );


  or
  g1410
  (
    n1452,
    n1414,
    n445,
    n1361,
    n446
  );


  xor
  g1411
  (
    n1465,
    n1019,
    n1414,
    n880,
    n1434
  );


  xnor
  g1412
  (
    n1453,
    n1360,
    n1020,
    n915,
    n446
  );


  nor
  g1413
  (
    n1464,
    n881,
    n1020,
    n1428,
    n1021
  );


  nand
  g1414
  (
    n1447,
    n918,
    n1430,
    n1433,
    n1415
  );


  xor
  g1415
  (
    n1457,
    n1426,
    n1430,
    n1416,
    n882
  );


  nand
  g1416
  (
    n1449,
    n918,
    n1016,
    n1019,
    n1431
  );


  xnor
  g1417
  (
    n1441,
    n444,
    n445,
    n1015,
    n881
  );


  and
  g1418
  (
    n1458,
    n1019,
    n1438,
    n1021,
    n1292
  );


  nand
  g1419
  (
    n1448,
    n446,
    n1416,
    n1417,
    n1359
  );


  and
  g1420
  (
    KeyWire_0_22,
    n1018,
    n918,
    n1429,
    n445
  );


  and
  g1421
  (
    n1462,
    n916,
    n881,
    n1018,
    n1014
  );


  nand
  g1422
  (
    n1468,
    n919,
    n919,
    n1016,
    n1432
  );


  xnor
  g1423
  (
    n1456,
    n1435,
    n917
  );


  and
  g1424
  (
    n1440,
    n1017,
    n880,
    n1362,
    n916
  );


  nor
  g1425
  (
    n1461,
    n445,
    n1015,
    n1417,
    n1423
  );


  and
  g1426
  (
    n1460,
    n1428,
    n1431,
    n1358,
    n1436
  );


  xnor
  g1427
  (
    n1455,
    n446,
    n1426,
    n1020,
    n1017
  );


  xnor
  g1428
  (
    n1467,
    n1433,
    n1021,
    n882,
    n1019
  );


  nor
  g1429
  (
    n1454,
    n1418,
    n1017,
    n1415,
    n1018
  );


  buf
  g1430
  (
    n1470,
    n1440
  );


  not
  g1431
  (
    n1469,
    n1439
  );


  xor
  g1432
  (
    n1471,
    n1373,
    n1367,
    n1377,
    n1469
  );


  xnor
  g1433
  (
    n1474,
    n1365,
    n1380,
    n1470,
    n1378
  );


  nand
  g1434
  (
    n1476,
    n1470,
    n1385,
    n1469,
    n1384
  );


  or
  g1435
  (
    n1477,
    n1387,
    n1370,
    n1470,
    n1374
  );


  xor
  g1436
  (
    n1475,
    n1375,
    n1369,
    n1364,
    n1383
  );


  or
  g1437
  (
    n1472,
    n1469,
    n1368,
    n1366,
    n1470
  );


  and
  g1438
  (
    n1473,
    n1469,
    n1371,
    n1381,
    n1372
  );


  nand
  g1439
  (
    n1478,
    n1376,
    n1382,
    n1386,
    n1379
  );


  xnor
  g1440
  (
    n1484,
    n1452,
    n1419,
    n1418,
    n1420
  );


  nor
  g1441
  (
    n1489,
    n1450,
    n1419,
    n1441,
    n1455
  );


  xor
  g1442
  (
    n1486,
    n1421,
    n1472,
    n1471,
    n1419
  );


  xor
  g1443
  (
    n1485,
    n1420,
    n1421,
    n1446
  );


  xnor
  g1444
  (
    n1481,
    n1476,
    n1444,
    n1475,
    n1448
  );


  and
  g1445
  (
    n1487,
    n1445,
    n1442,
    n1477,
    n1473
  );


  or
  g1446
  (
    n1480,
    n1422,
    n1476,
    n1454,
    n1032
  );


  xor
  g1447
  (
    n1488,
    n1422,
    n1443,
    n1420,
    n1418
  );


  nor
  g1448
  (
    n1479,
    n1449,
    n1453,
    n1422,
    n1478
  );


  xor
  g1449
  (
    n1482,
    n1451,
    n1447,
    n1457,
    n1477
  );


  and
  g1450
  (
    n1483,
    n1456,
    n1478,
    n1474,
    n1032
  );


  and
  g1451
  (
    n1491,
    n1480,
    n1489,
    n1038,
    n1485
  );


  or
  g1452
  (
    n1493,
    n1458,
    n1484,
    n1483,
    n1481
  );


  xor
  g1453
  (
    n1492,
    n1461,
    n1464,
    n1038,
    n1039
  );


  nor
  g1454
  (
    n1497,
    n1039,
    n1459,
    n1037,
    n1487
  );


  and
  g1455
  (
    n1490,
    n1040,
    n1040,
    n1467,
    n1037
  );


  nor
  g1456
  (
    n1496,
    n1466,
    n1468,
    n1460,
    n1462
  );


  and
  g1457
  (
    KeyWire_0_27,
    n1463,
    n1482,
    n1479,
    n1465
  );


  nor
  g1458
  (
    n1494,
    n1486,
    n1488,
    n1041
  );


  xor
  KeyGate_0_0
  (
    n795,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n252,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n456,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n818,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n216,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n120,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n629,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n671,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1241,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n621,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n343,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1036,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n625,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n51,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1459,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n622,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1406,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1063,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n771,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n898,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n967,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n443,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1442,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1438,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n118,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1126,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1075,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1495,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n827,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n244,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n884,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1124,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


