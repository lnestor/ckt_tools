

module Stat_1215_51_5
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n780,
  n773,
  n839,
  n840,
  n835,
  n838,
  n859,
  n856,
  n858,
  n868,
  n857,
  n972,
  n978,
  n981,
  n974,
  n1052,
  n1065,
  n1249,
  n1248,
  n1247,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input n33;
  input n34;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n780;
  output n773;
  output n839;
  output n840;
  output n835;
  output n838;
  output n859;
  output n856;
  output n858;
  output n868;
  output n857;
  output n972;
  output n978;
  output n981;
  output n974;
  output n1052;
  output n1065;
  output n1249;
  output n1248;
  output n1247;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n836;
  wire n837;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n973;
  wire n975;
  wire n976;
  wire n977;
  wire n979;
  wire n980;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n166,
    n24
  );


  buf
  g1
  (
    n86,
    n9
  );


  not
  g2
  (
    n80,
    n3
  );


  not
  g3
  (
    n137,
    n19
  );


  buf
  g4
  (
    n38,
    n31
  );


  buf
  g5
  (
    n78,
    n28
  );


  buf
  g6
  (
    n129,
    n21
  );


  not
  g7
  (
    n114,
    n27
  );


  not
  g8
  (
    n74,
    n25
  );


  buf
  g9
  (
    n64,
    n18
  );


  not
  g10
  (
    n119,
    n33
  );


  buf
  g11
  (
    n68,
    n2
  );


  not
  g12
  (
    n106,
    n15
  );


  not
  g13
  (
    n93,
    n29
  );


  buf
  g14
  (
    n104,
    n27
  );


  buf
  g15
  (
    n92,
    n34
  );


  buf
  g16
  (
    n134,
    n28
  );


  not
  g17
  (
    n118,
    n29
  );


  not
  g18
  (
    n72,
    n12
  );


  buf
  g19
  (
    n51,
    n14
  );


  not
  g20
  (
    n130,
    n13
  );


  buf
  g21
  (
    n67,
    n5
  );


  buf
  g22
  (
    n105,
    n18
  );


  not
  g23
  (
    n35,
    n1
  );


  not
  g24
  (
    n108,
    n14
  );


  buf
  g25
  (
    n124,
    n11
  );


  buf
  g26
  (
    n40,
    n33
  );


  buf
  g27
  (
    n76,
    n10
  );


  not
  g28
  (
    n155,
    n24
  );


  buf
  g29
  (
    n98,
    n3
  );


  buf
  g30
  (
    n44,
    n22
  );


  buf
  g31
  (
    n123,
    n1
  );


  buf
  g32
  (
    n82,
    n26
  );


  not
  g33
  (
    n60,
    n8
  );


  buf
  g34
  (
    n157,
    n8
  );


  buf
  g35
  (
    n90,
    n19
  );


  not
  g36
  (
    n136,
    n23
  );


  not
  g37
  (
    n53,
    n28
  );


  not
  g38
  (
    n79,
    n23
  );


  not
  g39
  (
    n135,
    n13
  );


  not
  g40
  (
    n160,
    n15
  );


  not
  g41
  (
    n65,
    n32
  );


  buf
  g42
  (
    n63,
    n22
  );


  buf
  g43
  (
    n138,
    n16
  );


  buf
  g44
  (
    n47,
    n33
  );


  not
  g45
  (
    n91,
    n7
  );


  not
  g46
  (
    n109,
    n25
  );


  not
  g47
  (
    n112,
    n23
  );


  buf
  g48
  (
    n120,
    n21
  );


  not
  g49
  (
    n77,
    n16
  );


  buf
  g50
  (
    n59,
    n19
  );


  not
  g51
  (
    n69,
    n5
  );


  buf
  g52
  (
    n122,
    n9
  );


  buf
  g53
  (
    n107,
    n18
  );


  buf
  g54
  (
    n139,
    n9
  );


  buf
  g55
  (
    n132,
    n30
  );


  not
  g56
  (
    n146,
    n9
  );


  not
  g57
  (
    n52,
    n11
  );


  buf
  g58
  (
    n161,
    n20
  );


  buf
  g59
  (
    n87,
    n32
  );


  buf
  g60
  (
    n127,
    n15
  );


  buf
  g61
  (
    n152,
    n32
  );


  not
  g62
  (
    n71,
    n21
  );


  buf
  g63
  (
    KeyWire_0_27,
    n20
  );


  buf
  g64
  (
    n164,
    n21
  );


  buf
  g65
  (
    n97,
    n1
  );


  not
  g66
  (
    n151,
    n16
  );


  buf
  g67
  (
    n54,
    n31
  );


  not
  g68
  (
    n143,
    n22
  );


  buf
  g69
  (
    n154,
    n32
  );


  buf
  g70
  (
    n125,
    n30
  );


  not
  g71
  (
    n66,
    n25
  );


  not
  g72
  (
    n95,
    n2
  );


  not
  g73
  (
    n149,
    n14
  );


  buf
  g74
  (
    n156,
    n2
  );


  not
  g75
  (
    n46,
    n25
  );


  buf
  g76
  (
    KeyWire_0_1,
    n15
  );


  buf
  g77
  (
    n45,
    n5
  );


  buf
  g78
  (
    n126,
    n31
  );


  not
  g79
  (
    n163,
    n2
  );


  buf
  g80
  (
    n170,
    n22
  );


  not
  g81
  (
    n103,
    n26
  );


  buf
  g82
  (
    n148,
    n10
  );


  buf
  g83
  (
    n111,
    n24
  );


  not
  g84
  (
    n70,
    n17
  );


  not
  g85
  (
    n147,
    n7
  );


  not
  g86
  (
    n85,
    n31
  );


  buf
  g87
  (
    n158,
    n11
  );


  not
  g88
  (
    n96,
    n18
  );


  not
  g89
  (
    n159,
    n8
  );


  buf
  g90
  (
    n84,
    n6
  );


  not
  g91
  (
    n101,
    n24
  );


  not
  g92
  (
    n58,
    n13
  );


  buf
  g93
  (
    n117,
    n10
  );


  not
  g94
  (
    n141,
    n1
  );


  buf
  g95
  (
    n133,
    n17
  );


  buf
  g96
  (
    n142,
    n3
  );


  buf
  g97
  (
    n145,
    n5
  );


  not
  g98
  (
    n41,
    n6
  );


  buf
  g99
  (
    n115,
    n4
  );


  buf
  g100
  (
    n73,
    n16
  );


  not
  g101
  (
    KeyWire_0_14,
    n17
  );


  not
  g102
  (
    n121,
    n10
  );


  not
  g103
  (
    n37,
    n34
  );


  not
  g104
  (
    n83,
    n34
  );


  not
  g105
  (
    n50,
    n7
  );


  not
  g106
  (
    n165,
    n34
  );


  not
  g107
  (
    n94,
    n6
  );


  buf
  g108
  (
    n55,
    n27
  );


  buf
  g109
  (
    n167,
    n29
  );


  buf
  g110
  (
    n153,
    n4
  );


  buf
  g111
  (
    n43,
    n8
  );


  buf
  g112
  (
    n61,
    n12
  );


  not
  g113
  (
    n62,
    n3
  );


  not
  g114
  (
    n169,
    n20
  );


  not
  g115
  (
    n48,
    n27
  );


  buf
  g116
  (
    n36,
    n7
  );


  not
  g117
  (
    n81,
    n26
  );


  buf
  g118
  (
    n168,
    n23
  );


  not
  g119
  (
    n128,
    n11
  );


  buf
  g120
  (
    n75,
    n13
  );


  buf
  g121
  (
    n110,
    n14
  );


  buf
  g122
  (
    n140,
    n26
  );


  buf
  g123
  (
    n99,
    n33
  );


  not
  g124
  (
    n162,
    n19
  );


  buf
  g125
  (
    n89,
    n28
  );


  not
  g126
  (
    n100,
    n12
  );


  buf
  g127
  (
    n57,
    n6
  );


  not
  g128
  (
    n144,
    n30
  );


  not
  g129
  (
    n113,
    n17
  );


  buf
  g130
  (
    n116,
    n4
  );


  buf
  g131
  (
    n56,
    n20
  );


  buf
  g132
  (
    n42,
    n12
  );


  buf
  g133
  (
    n131,
    n29
  );


  not
  g134
  (
    n49,
    n30
  );


  buf
  g135
  (
    n88,
    n4
  );


  buf
  g136
  (
    n371,
    n99
  );


  not
  g137
  (
    n194,
    n96
  );


  buf
  g138
  (
    n605,
    n133
  );


  buf
  g139
  (
    n290,
    n38
  );


  buf
  g140
  (
    n382,
    n130
  );


  not
  g141
  (
    n603,
    n116
  );


  buf
  g142
  (
    n196,
    n159
  );


  not
  g143
  (
    n575,
    n95
  );


  buf
  g144
  (
    n553,
    n142
  );


  not
  g145
  (
    n499,
    n98
  );


  not
  g146
  (
    n611,
    n160
  );


  buf
  g147
  (
    KeyWire_0_23,
    n106
  );


  buf
  g148
  (
    n483,
    n64
  );


  buf
  g149
  (
    n375,
    n149
  );


  not
  g150
  (
    n265,
    n119
  );


  not
  g151
  (
    n458,
    n161
  );


  buf
  g152
  (
    KeyWire_0_31,
    n62
  );


  not
  g153
  (
    n470,
    n129
  );


  not
  g154
  (
    n231,
    n61
  );


  buf
  g155
  (
    n192,
    n78
  );


  buf
  g156
  (
    n369,
    n45
  );


  buf
  g157
  (
    n443,
    n152
  );


  not
  g158
  (
    n552,
    n167
  );


  not
  g159
  (
    n267,
    n79
  );


  buf
  g160
  (
    n448,
    n115
  );


  not
  g161
  (
    n631,
    n42
  );


  buf
  g162
  (
    n434,
    n119
  );


  not
  g163
  (
    n590,
    n129
  );


  not
  g164
  (
    n461,
    n149
  );


  not
  g165
  (
    n280,
    n108
  );


  buf
  g166
  (
    n294,
    n155
  );


  not
  g167
  (
    n396,
    n69
  );


  buf
  g168
  (
    n404,
    n40
  );


  not
  g169
  (
    n179,
    n138
  );


  not
  g170
  (
    n416,
    n71
  );


  not
  g171
  (
    n279,
    n114
  );


  buf
  g172
  (
    n329,
    n152
  );


  buf
  g173
  (
    n627,
    n40
  );


  buf
  g174
  (
    n365,
    n107
  );


  buf
  g175
  (
    n452,
    n80
  );


  not
  g176
  (
    n506,
    n44
  );


  buf
  g177
  (
    n255,
    n167
  );


  not
  g178
  (
    n409,
    n88
  );


  not
  g179
  (
    n507,
    n157
  );


  buf
  g180
  (
    n312,
    n126
  );


  buf
  g181
  (
    n395,
    n102
  );


  buf
  g182
  (
    n521,
    n109
  );


  not
  g183
  (
    n264,
    n59
  );


  buf
  g184
  (
    n426,
    n44
  );


  buf
  g185
  (
    n393,
    n98
  );


  buf
  g186
  (
    n348,
    n105
  );


  not
  g187
  (
    n191,
    n140
  );


  not
  g188
  (
    n573,
    n102
  );


  not
  g189
  (
    n341,
    n77
  );


  not
  g190
  (
    n175,
    n73
  );


  buf
  g191
  (
    n218,
    n124
  );


  not
  g192
  (
    n459,
    n43
  );


  not
  g193
  (
    n569,
    n101
  );


  buf
  g194
  (
    n204,
    n144
  );


  buf
  g195
  (
    n322,
    n98
  );


  not
  g196
  (
    n556,
    n68
  );


  not
  g197
  (
    n334,
    n97
  );


  buf
  g198
  (
    n311,
    n115
  );


  buf
  g199
  (
    n230,
    n90
  );


  buf
  g200
  (
    n594,
    n87
  );


  not
  g201
  (
    n328,
    n56
  );


  buf
  g202
  (
    n563,
    n63
  );


  buf
  g203
  (
    n445,
    n67
  );


  buf
  g204
  (
    n424,
    n46
  );


  buf
  g205
  (
    n560,
    n113
  );


  buf
  g206
  (
    n597,
    n104
  );


  buf
  g207
  (
    n622,
    n155
  );


  not
  g208
  (
    n368,
    n66
  );


  not
  g209
  (
    n363,
    n135
  );


  buf
  g210
  (
    n487,
    n153
  );


  buf
  g211
  (
    KeyWire_0_18,
    n58
  );


  buf
  g212
  (
    n270,
    n88
  );


  buf
  g213
  (
    n567,
    n123
  );


  buf
  g214
  (
    n219,
    n126
  );


  buf
  g215
  (
    n326,
    n55
  );


  buf
  g216
  (
    n378,
    n101
  );


  buf
  g217
  (
    n374,
    n55
  );


  not
  g218
  (
    n324,
    n92
  );


  buf
  g219
  (
    n298,
    n117
  );


  buf
  g220
  (
    n319,
    n132
  );


  not
  g221
  (
    n640,
    n121
  );


  buf
  g222
  (
    n353,
    n91
  );


  not
  g223
  (
    n178,
    n94
  );


  buf
  g224
  (
    n357,
    n164
  );


  buf
  g225
  (
    n377,
    n165
  );


  not
  g226
  (
    n480,
    n36
  );


  not
  g227
  (
    n269,
    n134
  );


  not
  g228
  (
    n596,
    n143
  );


  not
  g229
  (
    n238,
    n42
  );


  not
  g230
  (
    n593,
    n161
  );


  not
  g231
  (
    n481,
    n81
  );


  not
  g232
  (
    n519,
    n60
  );


  buf
  g233
  (
    n228,
    n131
  );


  buf
  g234
  (
    n388,
    n159
  );


  not
  g235
  (
    n384,
    n83
  );


  buf
  g236
  (
    n526,
    n132
  );


  buf
  g237
  (
    n190,
    n133
  );


  buf
  g238
  (
    n187,
    n139
  );


  buf
  g239
  (
    n632,
    n137
  );


  not
  g240
  (
    n288,
    n131
  );


  not
  g241
  (
    n577,
    n35
  );


  buf
  g242
  (
    n243,
    n144
  );


  buf
  g243
  (
    n239,
    n80
  );


  buf
  g244
  (
    n435,
    n62
  );


  not
  g245
  (
    n197,
    n137
  );


  not
  g246
  (
    n300,
    n135
  );


  not
  g247
  (
    n297,
    n39
  );


  buf
  g248
  (
    n213,
    n57
  );


  not
  g249
  (
    KeyWire_0_0,
    n65
  );


  buf
  g250
  (
    n216,
    n51
  );


  not
  g251
  (
    n614,
    n138
  );


  not
  g252
  (
    n466,
    n111
  );


  buf
  g253
  (
    n250,
    n61
  );


  buf
  g254
  (
    n413,
    n48
  );


  buf
  g255
  (
    n580,
    n45
  );


  buf
  g256
  (
    n366,
    n158
  );


  not
  g257
  (
    n380,
    n70
  );


  buf
  g258
  (
    n513,
    n39
  );


  not
  g259
  (
    n209,
    n107
  );


  buf
  g260
  (
    n578,
    n136
  );


  buf
  g261
  (
    n538,
    n49
  );


  not
  g262
  (
    n340,
    n124
  );


  not
  g263
  (
    n635,
    n165
  );


  not
  g264
  (
    n402,
    n163
  );


  not
  g265
  (
    n257,
    n152
  );


  not
  g266
  (
    n345,
    n165
  );


  not
  g267
  (
    n464,
    n150
  );


  not
  g268
  (
    n282,
    n82
  );


  not
  g269
  (
    n359,
    n164
  );


  not
  g270
  (
    n325,
    n136
  );


  buf
  g271
  (
    n376,
    n129
  );


  buf
  g272
  (
    n339,
    n85
  );


  not
  g273
  (
    n619,
    n148
  );


  buf
  g274
  (
    n455,
    n115
  );


  not
  g275
  (
    n431,
    n125
  );


  not
  g276
  (
    n346,
    n167
  );


  not
  g277
  (
    n226,
    n42
  );


  not
  g278
  (
    n212,
    n137
  );


  not
  g279
  (
    n227,
    n132
  );


  not
  g280
  (
    n246,
    n120
  );


  buf
  g281
  (
    n283,
    n108
  );


  buf
  g282
  (
    n529,
    n144
  );


  buf
  g283
  (
    n547,
    n106
  );


  not
  g284
  (
    n182,
    n140
  );


  buf
  g285
  (
    n561,
    n161
  );


  buf
  g286
  (
    n587,
    n157
  );


  buf
  g287
  (
    n472,
    n92
  );


  not
  g288
  (
    n309,
    n77
  );


  not
  g289
  (
    n200,
    n148
  );


  buf
  g290
  (
    n386,
    n162
  );


  not
  g291
  (
    n181,
    n59
  );


  buf
  g292
  (
    KeyWire_0_11,
    n49
  );


  buf
  g293
  (
    n258,
    n95
  );


  buf
  g294
  (
    n555,
    n168
  );


  buf
  g295
  (
    n412,
    n76
  );


  buf
  g296
  (
    n358,
    n64
  );


  not
  g297
  (
    n420,
    n136
  );


  buf
  g298
  (
    n638,
    n127
  );


  not
  g299
  (
    n543,
    n132
  );


  buf
  g300
  (
    n360,
    n83
  );


  buf
  g301
  (
    n222,
    n135
  );


  buf
  g302
  (
    n469,
    n67
  );


  not
  g303
  (
    n186,
    n145
  );


  buf
  g304
  (
    KeyWire_0_20,
    n122
  );


  buf
  g305
  (
    n321,
    n157
  );


  buf
  g306
  (
    n281,
    n75
  );


  buf
  g307
  (
    n524,
    n97
  );


  buf
  g308
  (
    n432,
    n95
  );


  buf
  g309
  (
    n475,
    n117
  );


  not
  g310
  (
    n188,
    n103
  );


  not
  g311
  (
    n407,
    n143
  );


  buf
  g312
  (
    n602,
    n114
  );


  not
  g313
  (
    n439,
    n43
  );


  buf
  g314
  (
    n438,
    n76
  );


  buf
  g315
  (
    n399,
    n118
  );


  buf
  g316
  (
    KeyWire_0_4,
    n156
  );


  not
  g317
  (
    n276,
    n119
  );


  not
  g318
  (
    n236,
    n66
  );


  not
  g319
  (
    n589,
    n36
  );


  not
  g320
  (
    n306,
    n43
  );


  buf
  g321
  (
    n198,
    n149
  );


  not
  g322
  (
    n541,
    n158
  );


  not
  g323
  (
    n624,
    n156
  );


  not
  g324
  (
    n639,
    n55
  );


  buf
  g325
  (
    n446,
    n53
  );


  buf
  g326
  (
    n351,
    n37
  );


  buf
  g327
  (
    n485,
    n78
  );


  buf
  g328
  (
    n266,
    n69
  );


  not
  g329
  (
    n471,
    n154
  );


  buf
  g330
  (
    n444,
    n109
  );


  buf
  g331
  (
    n462,
    n44
  );


  buf
  g332
  (
    n565,
    n101
  );


  buf
  g333
  (
    n308,
    n54
  );


  buf
  g334
  (
    n566,
    n112
  );


  not
  g335
  (
    n608,
    n147
  );


  not
  g336
  (
    n356,
    n72
  );


  buf
  g337
  (
    n383,
    n63
  );


  not
  g338
  (
    n549,
    n118
  );


  not
  g339
  (
    n583,
    n134
  );


  buf
  g340
  (
    n241,
    n122
  );


  buf
  g341
  (
    n582,
    n134
  );


  buf
  g342
  (
    n338,
    n139
  );


  not
  g343
  (
    n189,
    n50
  );


  not
  g344
  (
    n623,
    n63
  );


  not
  g345
  (
    n545,
    n168
  );


  not
  g346
  (
    n584,
    n38
  );


  buf
  g347
  (
    n535,
    n86
  );


  not
  g348
  (
    n299,
    n61
  );


  buf
  g349
  (
    n394,
    n168
  );


  buf
  g350
  (
    n331,
    n146
  );


  not
  g351
  (
    n527,
    n105
  );


  not
  g352
  (
    n457,
    n150
  );


  not
  g353
  (
    n307,
    n52
  );


  not
  g354
  (
    n482,
    n78
  );


  buf
  g355
  (
    n429,
    n107
  );


  not
  g356
  (
    n491,
    n85
  );


  not
  g357
  (
    n441,
    n74
  );


  buf
  g358
  (
    n595,
    n109
  );


  not
  g359
  (
    n440,
    n113
  );


  not
  g360
  (
    n343,
    n41
  );


  not
  g361
  (
    n320,
    n86
  );


  not
  g362
  (
    n367,
    n131
  );


  not
  g363
  (
    KeyWire_0_9,
    n43
  );


  not
  g364
  (
    n261,
    n36
  );


  not
  g365
  (
    n533,
    n165
  );


  buf
  g366
  (
    n296,
    n52
  );


  buf
  g367
  (
    n564,
    n102
  );


  buf
  g368
  (
    n303,
    n110
  );


  buf
  g369
  (
    n389,
    n65
  );


  buf
  g370
  (
    n579,
    n51
  );


  buf
  g371
  (
    n317,
    n162
  );


  buf
  g372
  (
    n613,
    n106
  );


  not
  g373
  (
    n373,
    n68
  );


  buf
  g374
  (
    n460,
    n65
  );


  not
  g375
  (
    n505,
    n63
  );


  buf
  g376
  (
    n530,
    n125
  );


  not
  g377
  (
    n173,
    n139
  );


  not
  g378
  (
    n528,
    n158
  );


  not
  g379
  (
    n370,
    n56
  );


  buf
  g380
  (
    n456,
    n150
  );


  buf
  g381
  (
    n601,
    n114
  );


  not
  g382
  (
    n304,
    n55
  );


  not
  g383
  (
    n474,
    n99
  );


  buf
  g384
  (
    n410,
    n141
  );


  buf
  g385
  (
    n233,
    n79
  );


  buf
  g386
  (
    n315,
    n128
  );


  not
  g387
  (
    n406,
    n145
  );


  not
  g388
  (
    n558,
    n151
  );


  not
  g389
  (
    n174,
    n155
  );


  not
  g390
  (
    n478,
    n72
  );


  buf
  g391
  (
    n606,
    n135
  );


  not
  g392
  (
    n592,
    n81
  );


  not
  g393
  (
    n636,
    n113
  );


  buf
  g394
  (
    n571,
    n103
  );


  not
  g395
  (
    n260,
    n105
  );


  not
  g396
  (
    n272,
    n87
  );


  buf
  g397
  (
    n405,
    n142
  );


  buf
  g398
  (
    n522,
    n51
  );


  not
  g399
  (
    n408,
    n147
  );


  not
  g400
  (
    n537,
    n140
  );


  buf
  g401
  (
    n295,
    n133
  );


  buf
  g402
  (
    n422,
    n116
  );


  not
  g403
  (
    n428,
    n166
  );


  buf
  g404
  (
    n292,
    n71
  );


  not
  g405
  (
    n512,
    n88
  );


  not
  g406
  (
    n557,
    n99
  );


  not
  g407
  (
    n335,
    n141
  );


  not
  g408
  (
    n559,
    n87
  );


  not
  g409
  (
    n286,
    n41
  );


  buf
  g410
  (
    n391,
    n112
  );


  buf
  g411
  (
    n489,
    n148
  );


  not
  g412
  (
    n332,
    n92
  );


  buf
  g413
  (
    n415,
    n116
  );


  not
  g414
  (
    n277,
    n59
  );


  buf
  g415
  (
    n305,
    n94
  );


  buf
  g416
  (
    n607,
    n133
  );


  buf
  g417
  (
    n253,
    n157
  );


  buf
  g418
  (
    n473,
    n145
  );


  buf
  g419
  (
    n516,
    n99
  );


  buf
  g420
  (
    n201,
    n164
  );


  not
  g421
  (
    n411,
    n97
  );


  buf
  g422
  (
    n554,
    n100
  );


  buf
  g423
  (
    n504,
    n39
  );


  buf
  g424
  (
    n525,
    n128
  );


  not
  g425
  (
    n349,
    n66
  );


  buf
  g426
  (
    n629,
    n93
  );


  buf
  g427
  (
    n425,
    n134
  );


  buf
  g428
  (
    n254,
    n83
  );


  buf
  g429
  (
    n436,
    n153
  );


  not
  g430
  (
    n450,
    n162
  );


  not
  g431
  (
    n498,
    n73
  );


  buf
  g432
  (
    n621,
    n127
  );


  not
  g433
  (
    n493,
    n111
  );


  not
  g434
  (
    n249,
    n48
  );


  not
  g435
  (
    n625,
    n66
  );


  buf
  g436
  (
    n634,
    n72
  );


  buf
  g437
  (
    n454,
    n53
  );


  buf
  g438
  (
    n514,
    n117
  );


  buf
  g439
  (
    n548,
    n85
  );


  buf
  g440
  (
    n278,
    n86
  );


  buf
  g441
  (
    n207,
    n147
  );


  buf
  g442
  (
    n501,
    n96
  );


  not
  g443
  (
    n199,
    n48
  );


  buf
  g444
  (
    n235,
    n89
  );


  not
  g445
  (
    n523,
    n108
  );


  buf
  g446
  (
    KeyWire_0_21,
    n81
  );


  not
  g447
  (
    n215,
    n117
  );


  buf
  g448
  (
    n479,
    n57
  );


  not
  g449
  (
    n172,
    n46
  );


  buf
  g450
  (
    n248,
    n131
  );


  not
  g451
  (
    n562,
    n123
  );


  not
  g452
  (
    n615,
    n152
  );


  buf
  g453
  (
    n252,
    n110
  );


  buf
  g454
  (
    n568,
    n112
  );


  not
  g455
  (
    n546,
    n116
  );


  not
  g456
  (
    n609,
    n82
  );


  not
  g457
  (
    n495,
    n84
  );


  not
  g458
  (
    n220,
    n121
  );


  not
  g459
  (
    n620,
    n47
  );


  buf
  g460
  (
    n510,
    n121
  );


  not
  g461
  (
    n502,
    n123
  );


  not
  g462
  (
    n210,
    n54
  );


  not
  g463
  (
    n217,
    n130
  );


  buf
  g464
  (
    n289,
    n110
  );


  buf
  g465
  (
    KeyWire_0_26,
    n94
  );


  not
  g466
  (
    n275,
    n160
  );


  buf
  g467
  (
    n397,
    n167
  );


  not
  g468
  (
    n496,
    n130
  );


  not
  g469
  (
    n400,
    n50
  );


  buf
  g470
  (
    n293,
    n100
  );


  not
  g471
  (
    n232,
    n166
  );


  buf
  g472
  (
    n262,
    n108
  );


  buf
  g473
  (
    n520,
    n91
  );


  not
  g474
  (
    n500,
    n37
  );


  not
  g475
  (
    n310,
    n71
  );


  not
  g476
  (
    n347,
    n49
  );


  not
  g477
  (
    n453,
    n158
  );


  buf
  g478
  (
    n185,
    n98
  );


  not
  g479
  (
    n362,
    n163
  );


  not
  g480
  (
    n302,
    n143
  );


  not
  g481
  (
    n390,
    n47
  );


  not
  g482
  (
    n193,
    n153
  );


  buf
  g483
  (
    n628,
    n126
  );


  not
  g484
  (
    n534,
    n83
  );


  buf
  g485
  (
    n271,
    n90
  );


  not
  g486
  (
    n223,
    n156
  );


  buf
  g487
  (
    n221,
    n84
  );


  not
  g488
  (
    n626,
    n153
  );


  buf
  g489
  (
    n171,
    n97
  );


  buf
  g490
  (
    n214,
    n89
  );


  buf
  g491
  (
    n225,
    n79
  );


  not
  g492
  (
    n342,
    n84
  );


  buf
  g493
  (
    n544,
    n50
  );


  buf
  g494
  (
    KeyWire_0_28,
    n57
  );


  buf
  g495
  (
    n385,
    n53
  );


  buf
  g496
  (
    n419,
    n93
  );


  not
  g497
  (
    n447,
    n129
  );


  not
  g498
  (
    n503,
    n46
  );


  not
  g499
  (
    n313,
    n119
  );


  buf
  g500
  (
    n612,
    n100
  );


  buf
  g501
  (
    n344,
    n156
  );


  not
  g502
  (
    n392,
    n107
  );


  buf
  g503
  (
    n323,
    n75
  );


  buf
  g504
  (
    n437,
    n124
  );


  not
  g505
  (
    n540,
    n139
  );


  not
  g506
  (
    n387,
    n70
  );


  not
  g507
  (
    n418,
    n56
  );


  buf
  g508
  (
    n518,
    n113
  );


  not
  g509
  (
    n234,
    n122
  );


  not
  g510
  (
    n355,
    n146
  );


  buf
  g511
  (
    n586,
    n75
  );


  buf
  g512
  (
    n245,
    n40
  );


  not
  g513
  (
    n291,
    n159
  );


  not
  g514
  (
    n274,
    n154
  );


  not
  g515
  (
    n333,
    n69
  );


  not
  g516
  (
    n531,
    n58
  );


  buf
  g517
  (
    n183,
    n151
  );


  not
  g518
  (
    n268,
    n96
  );


  not
  g519
  (
    n379,
    n162
  );


  not
  g520
  (
    n517,
    n124
  );


  buf
  g521
  (
    n361,
    n143
  );


  buf
  g522
  (
    n421,
    n76
  );


  not
  g523
  (
    n449,
    n154
  );


  not
  g524
  (
    n488,
    n54
  );


  buf
  g525
  (
    n494,
    n103
  );


  buf
  g526
  (
    n633,
    n91
  );


  buf
  g527
  (
    n539,
    n65
  );


  buf
  g528
  (
    n515,
    n123
  );


  buf
  g529
  (
    n442,
    n74
  );


  buf
  g530
  (
    n484,
    n140
  );


  not
  g531
  (
    n414,
    n68
  );


  not
  g532
  (
    n352,
    n79
  );


  not
  g533
  (
    n600,
    n74
  );


  not
  g534
  (
    n463,
    n58
  );


  buf
  g535
  (
    n430,
    n50
  );


  not
  g536
  (
    n263,
    n144
  );


  not
  g537
  (
    n401,
    n89
  );


  buf
  g538
  (
    n314,
    n56
  );


  not
  g539
  (
    n465,
    n100
  );


  nand
  g540
  (
    n381,
    n159,
    n91
  );


  and
  g541
  (
    n195,
    n70,
    n87
  );


  xor
  g542
  (
    n251,
    n80,
    n67
  );


  xor
  g543
  (
    n427,
    n52,
    n109
  );


  nand
  g544
  (
    n202,
    n138,
    n60
  );


  xnor
  g545
  (
    n604,
    n40,
    n64
  );


  xnor
  g546
  (
    n316,
    n93,
    n51
  );


  xor
  g547
  (
    n327,
    n37,
    n125
  );


  nor
  g548
  (
    n208,
    n61,
    n160
  );


  xor
  g549
  (
    n336,
    n154,
    n121
  );


  xnor
  g550
  (
    n287,
    n57,
    n89
  );


  nand
  g551
  (
    n364,
    n130,
    n141
  );


  nand
  g552
  (
    n177,
    n114,
    n127
  );


  nor
  g553
  (
    KeyWire_0_24,
    n128,
    n102
  );


  nand
  g554
  (
    n301,
    n101,
    n59
  );


  and
  g555
  (
    n330,
    n82,
    n62
  );


  xor
  g556
  (
    n598,
    n120,
    n95
  );


  nor
  g557
  (
    n617,
    n39,
    n110
  );


  and
  g558
  (
    n184,
    n60,
    n73
  );


  nand
  g559
  (
    n203,
    n126,
    n118
  );


  xor
  g560
  (
    n490,
    n46,
    n52
  );


  or
  g561
  (
    n417,
    n151,
    n96
  );


  nand
  g562
  (
    n242,
    n136,
    n77
  );


  xnor
  g563
  (
    n468,
    n81,
    n41
  );


  or
  g564
  (
    n244,
    n49,
    n90
  );


  xnor
  g565
  (
    KeyWire_0_12,
    n111,
    n146
  );


  xor
  g566
  (
    n467,
    n163,
    n160
  );


  xor
  g567
  (
    n477,
    n148,
    n88
  );


  nor
  g568
  (
    n247,
    n103,
    n111
  );


  buf
  g569
  (
    KeyWire_0_16,
    n35
  );


  or
  g570
  (
    n511,
    n76,
    n73
  );


  xor
  g571
  (
    n536,
    n105,
    n118
  );


  and
  g572
  (
    KeyWire_0_19,
    n164,
    n147
  );


  nor
  g573
  (
    n451,
    n60,
    n70
  );


  xor
  g574
  (
    n237,
    n120,
    n122
  );


  or
  g575
  (
    n256,
    n104,
    n54
  );


  xor
  g576
  (
    n570,
    n168,
    n45
  );


  and
  g577
  (
    n486,
    n47,
    n150
  );


  nor
  g578
  (
    n176,
    n86,
    n82
  );


  nor
  g579
  (
    n476,
    n151,
    n69
  );


  xor
  g580
  (
    n318,
    n38,
    n74
  );


  nor
  g581
  (
    n229,
    n35,
    n163
  );


  xor
  g582
  (
    n637,
    n145,
    n80
  );


  or
  g583
  (
    n372,
    n155,
    n72
  );


  xor
  g584
  (
    n581,
    n161,
    n42
  );


  nor
  g585
  (
    n354,
    n45,
    n104
  );


  nand
  g586
  (
    n532,
    n41,
    n71
  );


  xnor
  g587
  (
    n588,
    n47,
    n146
  );


  nor
  g588
  (
    n273,
    n92,
    n84
  );


  or
  g589
  (
    n542,
    n85,
    n166
  );


  nor
  g590
  (
    n259,
    n128,
    n68
  );


  nand
  g591
  (
    n551,
    n78,
    n112
  );


  xor
  g592
  (
    n497,
    n142,
    n125
  );


  xnor
  g593
  (
    n211,
    n138,
    n137
  );


  xor
  g594
  (
    n224,
    n77,
    n67
  );


  xor
  g595
  (
    n508,
    n106,
    n62
  );


  and
  g596
  (
    n240,
    n53,
    n149
  );


  xor
  g597
  (
    n350,
    n94,
    n166
  );


  nand
  g598
  (
    n610,
    n75,
    n44
  );


  nand
  g599
  (
    n585,
    n36,
    n90
  );


  and
  g600
  (
    n206,
    n127,
    n93
  );


  xor
  g601
  (
    n630,
    n64,
    n38
  );


  nand
  g602
  (
    n616,
    n104,
    n58
  );


  nand
  g603
  (
    n509,
    n142,
    n48
  );


  xor
  g604
  (
    KeyWire_0_25,
    n115,
    n120
  );


  nand
  g605
  (
    n572,
    n37,
    n141
  );


  buf
  g606
  (
    n647,
    n173
  );


  not
  g607
  (
    n646,
    n178
  );


  not
  g608
  (
    n651,
    n182
  );


  buf
  g609
  (
    n653,
    n179
  );


  not
  g610
  (
    KeyWire_0_10,
    n171
  );


  not
  g611
  (
    n642,
    n181
  );


  buf
  g612
  (
    n643,
    n172
  );


  not
  g613
  (
    n644,
    n175
  );


  not
  g614
  (
    n641,
    n174
  );


  buf
  g615
  (
    n648,
    n176
  );


  buf
  g616
  (
    n650,
    n180
  );


  buf
  g617
  (
    n649,
    n183
  );


  buf
  g618
  (
    n645,
    n177
  );


  not
  g619
  (
    n658,
    n649
  );


  buf
  g620
  (
    n691,
    n650
  );


  not
  g621
  (
    n665,
    n645
  );


  not
  g622
  (
    n674,
    n191
  );


  not
  g623
  (
    KeyWire_0_13,
    n641
  );


  not
  g624
  (
    n671,
    n194
  );


  not
  g625
  (
    n685,
    n200
  );


  not
  g626
  (
    n684,
    n646
  );


  not
  g627
  (
    n693,
    n651
  );


  not
  g628
  (
    n673,
    n648
  );


  not
  g629
  (
    n675,
    n642
  );


  buf
  g630
  (
    n661,
    n651
  );


  buf
  g631
  (
    n659,
    n185
  );


  buf
  g632
  (
    n694,
    n202
  );


  buf
  g633
  (
    n682,
    n196
  );


  not
  g634
  (
    n660,
    n645
  );


  buf
  g635
  (
    n668,
    n649
  );


  buf
  g636
  (
    n677,
    n197
  );


  not
  g637
  (
    n656,
    n189
  );


  buf
  g638
  (
    n690,
    n641
  );


  not
  g639
  (
    n696,
    n186
  );


  buf
  g640
  (
    n667,
    n649
  );


  buf
  g641
  (
    n672,
    n647
  );


  buf
  g642
  (
    n695,
    n645
  );


  buf
  g643
  (
    n681,
    n644
  );


  not
  g644
  (
    n669,
    n642
  );


  not
  g645
  (
    n678,
    n646
  );


  buf
  g646
  (
    n663,
    n643
  );


  buf
  g647
  (
    n679,
    n199
  );


  not
  g648
  (
    n664,
    n643
  );


  not
  g649
  (
    n686,
    n193
  );


  not
  g650
  (
    n654,
    n188
  );


  buf
  g651
  (
    n687,
    n646
  );


  buf
  g652
  (
    KeyWire_0_8,
    n644
  );


  buf
  g653
  (
    n670,
    n641
  );


  buf
  g654
  (
    n680,
    n641
  );


  or
  g655
  (
    n688,
    n643,
    n201,
    n642,
    n644
  );


  nand
  g656
  (
    n692,
    n650,
    n650,
    n647,
    n648
  );


  xnor
  g657
  (
    n666,
    n648,
    n644,
    n204,
    n647
  );


  nand
  g658
  (
    n655,
    n190,
    n642,
    n650,
    n184
  );


  xnor
  g659
  (
    n662,
    n647,
    n651,
    n649,
    n646
  );


  nand
  g660
  (
    n689,
    n648,
    n195,
    n192,
    n645
  );


  xor
  g661
  (
    n683,
    n203,
    n198,
    n187,
    n643
  );


  and
  g662
  (
    n708,
    n253,
    n222,
    n241,
    n251
  );


  nand
  g663
  (
    n705,
    n658,
    n228,
    n231,
    n657
  );


  and
  g664
  (
    n698,
    n225,
    n256,
    n218,
    n239
  );


  or
  g665
  (
    n701,
    n244,
    n224,
    n654
  );


  or
  g666
  (
    n710,
    n658,
    n240,
    n233,
    n654
  );


  xor
  g667
  (
    n706,
    n657,
    n208,
    n211,
    n258
  );


  xor
  g668
  (
    n714,
    n657,
    n216,
    n238,
    n656
  );


  or
  g669
  (
    n699,
    n230,
    n219,
    n221,
    n235
  );


  nor
  g670
  (
    n713,
    n214,
    n207,
    n655,
    n237
  );


  xor
  g671
  (
    n712,
    n217,
    n226,
    n210,
    n227
  );


  nor
  g672
  (
    n697,
    n249,
    n220,
    n656,
    n655
  );


  and
  g673
  (
    n702,
    n236,
    n257,
    n252,
    n657
  );


  xor
  g674
  (
    n711,
    n656,
    n243,
    n248,
    n247
  );


  or
  g675
  (
    n707,
    n206,
    n212,
    n209,
    n656
  );


  and
  g676
  (
    n703,
    n245,
    n215,
    n234,
    n654
  );


  xnor
  g677
  (
    n700,
    n250,
    n246,
    n232,
    n205
  );


  xor
  g678
  (
    n709,
    n223,
    n254,
    n242,
    n655
  );


  and
  g679
  (
    n704,
    n255,
    n229,
    n655,
    n213
  );


  and
  g680
  (
    n728,
    n279,
    n703,
    n260,
    n262
  );


  xnor
  g681
  (
    n723,
    n711,
    n284,
    n298,
    n307
  );


  or
  g682
  (
    n725,
    n708,
    n297,
    n706,
    n288
  );


  xnor
  g683
  (
    n724,
    n308,
    n302,
    n713,
    n304
  );


  or
  g684
  (
    n717,
    n281,
    n712,
    n309,
    n264
  );


  or
  g685
  (
    n731,
    n266,
    n709,
    n280,
    n710
  );


  nor
  g686
  (
    n721,
    n292,
    n275,
    n259,
    n296
  );


  nand
  g687
  (
    n716,
    n293,
    n295,
    n289,
    n268
  );


  xnor
  g688
  (
    n729,
    n300,
    n702,
    n704,
    n272
  );


  and
  g689
  (
    n719,
    n303,
    n700,
    n701,
    n698
  );


  nor
  g690
  (
    n722,
    n261,
    n286,
    n285,
    n291
  );


  xnor
  g691
  (
    n718,
    n276,
    n270,
    n267,
    n283
  );


  nand
  g692
  (
    n726,
    n271,
    n265,
    n274,
    n299
  );


  nor
  g693
  (
    n720,
    n301,
    n699,
    n697,
    n282
  );


  nor
  g694
  (
    n727,
    n290,
    n269,
    n294,
    n273
  );


  xor
  g695
  (
    n730,
    n306,
    n278,
    n305,
    n705
  );


  xnor
  g696
  (
    n715,
    n263,
    n707,
    n277,
    n287
  );


  xnor
  g697
  (
    n736,
    n381,
    n718,
    n369,
    n336
  );


  nand
  g698
  (
    n734,
    n344,
    n366,
    n728,
    n323
  );


  nor
  g699
  (
    n749,
    n353,
    n383,
    n722,
    n346
  );


  xor
  g700
  (
    n747,
    n339,
    n322,
    n367,
    n725
  );


  xor
  g701
  (
    n754,
    n311,
    n347,
    n331,
    n335
  );


  nand
  g702
  (
    n755,
    n320,
    n330,
    n316,
    n325
  );


  nand
  g703
  (
    n745,
    n314,
    n368,
    n723,
    n360
  );


  nand
  g704
  (
    n742,
    n376,
    n378,
    n319,
    n310
  );


  and
  g705
  (
    n746,
    n334,
    n387,
    n730,
    n727
  );


  nor
  g706
  (
    n740,
    n727,
    n384,
    n377,
    n328
  );


  and
  g707
  (
    n748,
    n716,
    n327,
    n349,
    n312
  );


  or
  g708
  (
    n752,
    n371,
    n340,
    n313,
    n374
  );


  or
  g709
  (
    n735,
    n726,
    n720,
    n722,
    n321
  );


  or
  g710
  (
    n738,
    n364,
    n342,
    n317,
    n373
  );


  xor
  g711
  (
    n744,
    n375,
    n361,
    n356,
    n370
  );


  nand
  g712
  (
    n751,
    n724,
    n318,
    n365,
    n729
  );


  xor
  g713
  (
    n757,
    n338,
    n329,
    n354,
    n385
  );


  nor
  g714
  (
    n750,
    n351,
    n332,
    n352,
    n386
  );


  xnor
  g715
  (
    n733,
    n348,
    n359,
    n717,
    n719
  );


  xor
  g716
  (
    n739,
    n357,
    n343,
    n382,
    n731
  );


  nand
  g717
  (
    n743,
    n324,
    n729,
    n341,
    n337
  );


  nand
  g718
  (
    n753,
    n715,
    n362,
    n326,
    n315
  );


  and
  g719
  (
    n741,
    n372,
    n379,
    n730,
    n726
  );


  xnor
  g720
  (
    n756,
    n380,
    n333,
    n724,
    n721
  );


  nand
  g721
  (
    n737,
    n350,
    n355,
    n728,
    n345
  );


  and
  g722
  (
    n732,
    n358,
    n725,
    n723,
    n363
  );


  and
  g723
  (
    n759,
    n732,
    n659
  );


  xor
  g724
  (
    KeyWire_0_15,
    n659,
    n658,
    n733
  );


  xnor
  g725
  (
    n765,
    n661,
    n734
  );


  and
  g726
  (
    n760,
    n661,
    n660,
    n759
  );


  nor
  g727
  (
    n761,
    n759,
    n661,
    n662,
    n758
  );


  xnor
  g728
  (
    n764,
    n389,
    n663,
    n758,
    n759
  );


  nand
  g729
  (
    n766,
    n660,
    n662,
    n659
  );


  nor
  g730
  (
    n763,
    n663,
    n662,
    n758,
    n388
  );


  xor
  g731
  (
    n762,
    n662,
    n661,
    n660,
    n759
  );


  buf
  g732
  (
    n768,
    n760
  );


  buf
  g733
  (
    n767,
    n760
  );


  buf
  g734
  (
    n769,
    n760
  );


  not
  g735
  (
    n770,
    n767
  );


  not
  g736
  (
    n772,
    n770
  );


  buf
  g737
  (
    n771,
    n770
  );


  nor
  g738
  (
    n778,
    n763,
    n764,
    n772
  );


  nor
  g739
  (
    n773,
    n766,
    n771,
    n772,
    n762
  );


  xor
  g740
  (
    n779,
    n771,
    n761,
    n765,
    n763
  );


  nand
  g741
  (
    n777,
    n763,
    n760,
    n761,
    n764
  );


  or
  g742
  (
    n776,
    n772,
    n764,
    n765,
    n762
  );


  nor
  g743
  (
    n780,
    n169,
    n766,
    n765,
    n771
  );


  or
  g744
  (
    n775,
    n762,
    n771,
    n772,
    n761
  );


  xor
  g745
  (
    n774,
    n762,
    n761,
    n765,
    n763
  );


  nor
  g746
  (
    n783,
    n394,
    n398,
    n775,
    n400
  );


  xor
  g747
  (
    n782,
    n403,
    n778,
    n399,
    n777
  );


  xor
  g748
  (
    n786,
    n405,
    n780,
    n779,
    n393
  );


  and
  g749
  (
    n784,
    n395,
    n401,
    n397,
    n402
  );


  xnor
  g750
  (
    n785,
    n406,
    n391,
    n396,
    n390
  );


  and
  g751
  (
    n781,
    n407,
    n404,
    n776,
    n392
  );


  not
  g752
  (
    n788,
    n781
  );


  not
  g753
  (
    n789,
    n781
  );


  buf
  g754
  (
    n790,
    n781
  );


  not
  g755
  (
    n787,
    n781
  );


  and
  g756
  (
    n792,
    n412,
    n410,
    n424,
    n428
  );


  nor
  g757
  (
    n794,
    n782,
    n789,
    n418,
    n663
  );


  nor
  g758
  (
    n797,
    n665,
    n787,
    n415,
    n788
  );


  and
  g759
  (
    n791,
    n664,
    n416,
    n413,
    n788
  );


  xor
  g760
  (
    n800,
    n417,
    n408,
    n411,
    n421
  );


  xnor
  g761
  (
    n793,
    n789,
    n409,
    n787,
    n664
  );


  nor
  g762
  (
    n796,
    n664,
    n788,
    n414,
    n420
  );


  nand
  g763
  (
    n798,
    n426,
    n663,
    n422,
    n788
  );


  nand
  g764
  (
    n799,
    n427,
    n782,
    n664,
    n425
  );


  xnor
  g765
  (
    n795,
    n423,
    n787,
    n419
  );


  buf
  g766
  (
    n813,
    n796
  );


  not
  g767
  (
    n807,
    n798
  );


  buf
  g768
  (
    n804,
    n800
  );


  buf
  g769
  (
    n815,
    n795
  );


  not
  g770
  (
    n809,
    n795
  );


  not
  g771
  (
    n806,
    n794
  );


  not
  g772
  (
    n808,
    n791
  );


  not
  g773
  (
    n802,
    n797
  );


  not
  g774
  (
    n818,
    n797
  );


  buf
  g775
  (
    n801,
    n796
  );


  not
  g776
  (
    n811,
    n799
  );


  buf
  g777
  (
    n817,
    n794
  );


  not
  g778
  (
    n803,
    n793
  );


  buf
  g779
  (
    n805,
    n800
  );


  not
  g780
  (
    n816,
    n798
  );


  not
  g781
  (
    n814,
    n792
  );


  buf
  g782
  (
    n810,
    n799
  );


  not
  g783
  (
    n812,
    n793
  );


  buf
  g784
  (
    n820,
    n809
  );


  buf
  g785
  (
    n824,
    n806
  );


  buf
  g786
  (
    n819,
    n802
  );


  not
  g787
  (
    n826,
    n805
  );


  not
  g788
  (
    n827,
    n805
  );


  not
  g789
  (
    n832,
    n804
  );


  not
  g790
  (
    n821,
    n782
  );


  not
  g791
  (
    n823,
    n809
  );


  not
  g792
  (
    n828,
    n807
  );


  buf
  g793
  (
    n833,
    n803
  );


  not
  g794
  (
    n834,
    n784
  );


  buf
  g795
  (
    n831,
    n783
  );


  not
  g796
  (
    n825,
    n783
  );


  xor
  g797
  (
    n822,
    n806,
    n801,
    n784
  );


  nor
  g798
  (
    n829,
    n804,
    n807,
    n803,
    n808
  );


  xor
  g799
  (
    n830,
    n783,
    n808,
    n784,
    n782
  );


  or
  g800
  (
    n839,
    n821,
    n439,
    n438,
    n819
  );


  xnor
  g801
  (
    n835,
    n435,
    n436,
    n430,
    n445
  );


  xnor
  g802
  (
    n837,
    n431,
    n442,
    n444,
    n443
  );


  xnor
  g803
  (
    n836,
    n819,
    n810,
    n441,
    n440
  );


  nor
  g804
  (
    n840,
    n434,
    n432,
    n820
  );


  or
  g805
  (
    n838,
    n437,
    n433,
    n821,
    n429
  );


  nand
  g806
  (
    n841,
    n169,
    n170
  );


  nor
  g807
  (
    n842,
    n840,
    n839,
    n169
  );


  xor
  g808
  (
    n843,
    n841,
    n446
  );


  not
  g809
  (
    n845,
    n843
  );


  and
  g810
  (
    n844,
    n652,
    n843,
    n651
  );


  not
  g811
  (
    n852,
    n844
  );


  not
  g812
  (
    n848,
    n845
  );


  not
  g813
  (
    n846,
    n844
  );


  buf
  g814
  (
    n849,
    n845
  );


  not
  g815
  (
    n851,
    n845
  );


  not
  g816
  (
    n853,
    n845
  );


  not
  g817
  (
    n847,
    n844
  );


  buf
  g818
  (
    n850,
    n844
  );


  nor
  g819
  (
    n859,
    n822,
    n745,
    n754,
    n738
  );


  xnor
  g820
  (
    n869,
    n846,
    n824,
    n814,
    n811
  );


  or
  g821
  (
    n855,
    n848,
    n848,
    n847,
    n849
  );


  or
  g822
  (
    n860,
    n812,
    n815,
    n749,
    n742
  );


  nor
  g823
  (
    n868,
    n652,
    n846,
    n750,
    n811
  );


  nand
  g824
  (
    n854,
    n847,
    n755,
    n752,
    n746
  );


  and
  g825
  (
    n867,
    n823,
    n736,
    n748,
    n848
  );


  or
  g826
  (
    n857,
    n824,
    n813,
    n822,
    n812
  );


  and
  g827
  (
    n866,
    n756,
    n744,
    n849,
    n741
  );


  nand
  g828
  (
    KeyWire_0_29,
    n848,
    n816,
    n846
  );


  and
  g829
  (
    n863,
    n842,
    n818,
    n739,
    n751
  );


  and
  g830
  (
    n858,
    n846,
    n737,
    n813,
    n847
  );


  nand
  g831
  (
    n864,
    n743,
    n753,
    n849,
    n815
  );


  nor
  g832
  (
    n862,
    n817,
    n714,
    n735,
    n849
  );


  nand
  g833
  (
    n861,
    n747,
    n847,
    n740,
    n817
  );


  nand
  g834
  (
    n856,
    n757,
    n823,
    n810,
    n814
  );


  and
  g835
  (
    n875,
    n867,
    n851
  );


  and
  g836
  (
    n879,
    n850,
    n852
  );


  nand
  g837
  (
    n873,
    n865,
    n850
  );


  nand
  g838
  (
    n874,
    n852,
    n851
  );


  or
  g839
  (
    n877,
    n851,
    n731
  );


  nand
  g840
  (
    n871,
    n853,
    n868
  );


  and
  g841
  (
    n880,
    n863,
    n850,
    n853
  );


  nor
  g842
  (
    n872,
    n850,
    n852,
    n859
  );


  nor
  g843
  (
    n870,
    n170,
    n860,
    n869,
    n861
  );


  xor
  g844
  (
    n876,
    n864,
    n851,
    n853,
    n862
  );


  xor
  g845
  (
    n878,
    n866,
    n852,
    n853,
    n818
  );


  not
  g846
  (
    n882,
    n870
  );


  not
  g847
  (
    n881,
    n871
  );


  nor
  g848
  (
    n883,
    n881,
    n873,
    n872
  );


  nand
  g849
  (
    n885,
    n766,
    n883
  );


  or
  g850
  (
    n884,
    n766,
    n883
  );


  buf
  g851
  (
    n887,
    n767
  );


  nor
  g852
  (
    n886,
    n875,
    n884,
    n874,
    n885
  );


  xor
  g853
  (
    n891,
    n881,
    n887,
    n882
  );


  and
  g854
  (
    n888,
    n881,
    n881,
    n886,
    n448
  );


  xnor
  g855
  (
    n890,
    n887,
    n882,
    n447
  );


  and
  g856
  (
    n889,
    n451,
    n450,
    n886,
    n449
  );


  nand
  g857
  (
    n895,
    n466,
    n456,
    n495,
    n485
  );


  xnor
  g858
  (
    n903,
    n482,
    n470,
    n473,
    n475
  );


  and
  g859
  (
    n894,
    n483,
    n890,
    n476,
    n498
  );


  xor
  g860
  (
    n901,
    n888,
    n477,
    n454,
    n890
  );


  nand
  g861
  (
    n898,
    n888,
    n490,
    n460,
    n499
  );


  nand
  g862
  (
    n899,
    n890,
    n468,
    n462,
    n486
  );


  nand
  g863
  (
    n900,
    n453,
    n452,
    n491,
    n890
  );


  xor
  g864
  (
    n905,
    n889,
    n464,
    n484,
    n472
  );


  or
  g865
  (
    n902,
    n891,
    n458,
    n487,
    n888
  );


  xnor
  g866
  (
    n896,
    n471,
    n891,
    n457,
    n481
  );


  xnor
  g867
  (
    KeyWire_0_5,
    n489,
    n479,
    n889,
    n494
  );


  xor
  g868
  (
    n893,
    n474,
    n465,
    n497,
    n492
  );


  xnor
  g869
  (
    n904,
    n889,
    n488,
    n463,
    n891
  );


  nand
  g870
  (
    n897,
    n459,
    n480,
    n493,
    n478
  );


  nand
  g871
  (
    n892,
    n889,
    n888,
    n891,
    n467
  );


  nor
  g872
  (
    n907,
    n496,
    n461,
    n455,
    n469
  );


  and
  g873
  (
    n927,
    n507,
    n544,
    n524,
    n512
  );


  xnor
  g874
  (
    n937,
    n548,
    n901,
    n899,
    n530
  );


  and
  g875
  (
    n924,
    n896,
    n577,
    n893,
    n574
  );


  nand
  g876
  (
    n931,
    n561,
    n897,
    n515,
    n568
  );


  nand
  g877
  (
    n935,
    n893,
    n900,
    n571,
    n525
  );


  xnor
  g878
  (
    n921,
    n579,
    n902,
    n904,
    n571
  );


  nor
  g879
  (
    n918,
    n520,
    n562,
    n573,
    n904
  );


  or
  g880
  (
    n915,
    n900,
    n567,
    n550,
    n899
  );


  nand
  g881
  (
    n914,
    n564,
    n536,
    n905,
    n521
  );


  or
  g882
  (
    n913,
    n907,
    n531,
    n905,
    n501
  );


  nor
  g883
  (
    n908,
    n566,
    n527,
    n506,
    n532
  );


  xnor
  g884
  (
    n912,
    n553,
    n529,
    n517,
    n535
  );


  nor
  g885
  (
    n936,
    n897,
    n513,
    n551,
    n565
  );


  xnor
  g886
  (
    n934,
    n577,
    n511,
    n540,
    n522
  );


  and
  g887
  (
    n917,
    n895,
    n528,
    n533,
    n574
  );


  or
  g888
  (
    n920,
    n552,
    n541,
    n503,
    n526
  );


  xor
  g889
  (
    n916,
    n538,
    n896,
    n543,
    n894
  );


  xor
  g890
  (
    n910,
    n901,
    n570,
    n903,
    n898
  );


  xor
  g891
  (
    n938,
    n523,
    n572,
    n568,
    n510
  );


  nor
  g892
  (
    n933,
    n559,
    n578,
    n563,
    n519
  );


  nor
  g893
  (
    n932,
    n555,
    n566,
    n547,
    n902
  );


  or
  g894
  (
    n939,
    n502,
    n518,
    n567,
    n514
  );


  nand
  g895
  (
    n930,
    n539,
    n565,
    n895,
    n569
  );


  xor
  g896
  (
    n925,
    n569,
    n505,
    n575,
    n573
  );


  nand
  g897
  (
    n928,
    n542,
    n907,
    n576
  );


  and
  g898
  (
    n911,
    n556,
    n575,
    n892,
    n537
  );


  xor
  g899
  (
    n923,
    n516,
    n580,
    n508,
    n560
  );


  or
  g900
  (
    n926,
    n906,
    n545,
    n894,
    n898
  );


  xnor
  g901
  (
    n929,
    n549,
    n500,
    n554,
    n546
  );


  nor
  g902
  (
    n909,
    n558,
    n572,
    n903,
    n509
  );


  xor
  g903
  (
    n919,
    n579,
    n570,
    n504,
    n578
  );


  and
  g904
  (
    n922,
    n534,
    n906,
    n557,
    n892
  );


  buf
  g905
  (
    n940,
    n916
  );


  buf
  g906
  (
    n960,
    n919
  );


  not
  g907
  (
    n950,
    n920
  );


  buf
  g908
  (
    n959,
    n915
  );


  not
  g909
  (
    n949,
    n786
  );


  not
  g910
  (
    n946,
    n914
  );


  not
  g911
  (
    n956,
    n917
  );


  not
  g912
  (
    n942,
    n786
  );


  buf
  g913
  (
    n948,
    n913
  );


  buf
  g914
  (
    n944,
    n918
  );


  buf
  g915
  (
    n951,
    n913
  );


  not
  g916
  (
    n945,
    n909
  );


  not
  g917
  (
    n955,
    n785
  );


  buf
  g918
  (
    n962,
    n918
  );


  not
  g919
  (
    n961,
    n911
  );


  not
  g920
  (
    n957,
    n910
  );


  xnor
  g921
  (
    n953,
    n910,
    n917
  );


  and
  g922
  (
    n943,
    n914,
    n786
  );


  xnor
  g923
  (
    n941,
    n785,
    n911
  );


  or
  g924
  (
    n963,
    n915,
    n785
  );


  xor
  g925
  (
    n952,
    n919,
    n786
  );


  and
  g926
  (
    n958,
    n785,
    n912
  );


  xor
  g927
  (
    n947,
    n916,
    n912
  );


  nor
  g928
  (
    n954,
    n908,
    n920
  );


  and
  g929
  (
    n965,
    n926,
    n940,
    n945,
    n946
  );


  xor
  g930
  (
    n981,
    n941,
    n924,
    n942,
    n921
  );


  nand
  g931
  (
    n978,
    n932,
    n943,
    n937,
    n941
  );


  or
  g932
  (
    n964,
    n939,
    n926,
    n936,
    n934
  );


  nor
  g933
  (
    n975,
    n586,
    n948,
    n928,
    n921
  );


  xor
  g934
  (
    n969,
    n931,
    n587,
    n584,
    n947
  );


  or
  g935
  (
    n967,
    n925,
    n933,
    n582,
    n929
  );


  and
  g936
  (
    n971,
    n927,
    n934,
    n930,
    n581
  );


  xnor
  g937
  (
    n979,
    n938,
    n587,
    n584,
    n922
  );


  and
  g938
  (
    n972,
    n925,
    n933,
    n586,
    n944
  );


  and
  g939
  (
    n980,
    n949,
    n585,
    n935
  );


  and
  g940
  (
    n970,
    n927,
    n938,
    n946,
    n945
  );


  nand
  g941
  (
    n974,
    n942,
    n936,
    n939,
    n940
  );


  nor
  g942
  (
    n976,
    n947,
    n931,
    n582,
    n924
  );


  nor
  g943
  (
    KeyWire_0_17,
    n930,
    n932,
    n928,
    n923
  );


  or
  g944
  (
    n973,
    n943,
    n923,
    n583,
    n922
  );


  or
  g945
  (
    n977,
    n580,
    n583,
    n929,
    n935
  );


  or
  g946
  (
    n966,
    n937,
    n581,
    n948,
    n944
  );


  nand
  g947
  (
    n994,
    n592,
    n595,
    n951,
    n979
  );


  and
  g948
  (
    n983,
    n952,
    n975,
    n971,
    n593
  );


  nor
  g949
  (
    n984,
    n952,
    n980,
    n589,
    n597
  );


  xor
  g950
  (
    n990,
    n968,
    n593,
    n592,
    n599
  );


  or
  g951
  (
    n987,
    n949,
    n598,
    n601,
    n594
  );


  nand
  g952
  (
    n989,
    n590,
    n588,
    n597,
    n969
  );


  or
  g953
  (
    n991,
    n953,
    n596,
    n603,
    n970
  );


  and
  g954
  (
    n982,
    n972,
    n603,
    n973,
    n974
  );


  nand
  g955
  (
    n986,
    n589,
    n600,
    n981,
    n602
  );


  and
  g956
  (
    n988,
    n599,
    n590,
    n595,
    n976
  );


  or
  g957
  (
    n985,
    n978,
    n953,
    n596,
    n598
  );


  or
  g958
  (
    n995,
    n600,
    n602,
    n591,
    n950
  );


  and
  g959
  (
    n993,
    n591,
    n977,
    n950,
    n588
  );


  nand
  g960
  (
    n992,
    n601,
    n951,
    n954,
    n594
  );


  buf
  g961
  (
    n1006,
    n982
  );


  not
  g962
  (
    n999,
    n987
  );


  buf
  g963
  (
    KeyWire_0_30,
    n986
  );


  buf
  g964
  (
    n1000,
    n987
  );


  buf
  g965
  (
    n998,
    n986
  );


  buf
  g966
  (
    n1001,
    n985
  );


  not
  g967
  (
    n997,
    n983
  );


  not
  g968
  (
    n1004,
    n985
  );


  not
  g969
  (
    n1003,
    n984
  );


  buf
  g970
  (
    n996,
    n983
  );


  not
  g971
  (
    n1005,
    n984
  );


  buf
  g972
  (
    n1007,
    n982
  );


  buf
  g973
  (
    n1040,
    n999
  );


  not
  g974
  (
    n1008,
    n997
  );


  buf
  g975
  (
    n1018,
    n998
  );


  not
  g976
  (
    n1037,
    n1002
  );


  buf
  g977
  (
    n1043,
    n997
  );


  not
  g978
  (
    n1013,
    n997
  );


  buf
  g979
  (
    n1036,
    n998
  );


  not
  g980
  (
    n1032,
    n996
  );


  buf
  g981
  (
    n1026,
    n1003
  );


  buf
  g982
  (
    n1024,
    n1003
  );


  not
  g983
  (
    KeyWire_0_7,
    n997
  );


  not
  g984
  (
    n1034,
    n998
  );


  buf
  g985
  (
    n1027,
    n996
  );


  buf
  g986
  (
    n1021,
    n998
  );


  buf
  g987
  (
    n1019,
    n1000
  );


  buf
  g988
  (
    KeyWire_0_22,
    n996
  );


  not
  g989
  (
    n1015,
    n1003
  );


  not
  g990
  (
    n1039,
    n1003
  );


  not
  g991
  (
    n1030,
    n1002
  );


  buf
  g992
  (
    n1035,
    n1000
  );


  buf
  g993
  (
    n1009,
    n1004
  );


  buf
  g994
  (
    n1025,
    n1004
  );


  buf
  g995
  (
    n1012,
    n999
  );


  buf
  g996
  (
    n1014,
    n1001
  );


  buf
  g997
  (
    n1023,
    n955
  );


  buf
  g998
  (
    n1022,
    n999
  );


  buf
  g999
  (
    n1011,
    n1001
  );


  buf
  g1000
  (
    n1016,
    n1002
  );


  buf
  g1001
  (
    n1041,
    n1004
  );


  buf
  g1002
  (
    n1028,
    n1004
  );


  buf
  g1003
  (
    n1020,
    n999
  );


  buf
  g1004
  (
    n1033,
    n996
  );


  buf
  g1005
  (
    n1038,
    n1001
  );


  not
  g1006
  (
    n1031,
    n1002
  );


  xor
  g1007
  (
    n1017,
    n1001,
    n954
  );


  buf
  g1008
  (
    n1010,
    n1000
  );


  xor
  g1009
  (
    n1045,
    n959,
    n958
  );


  not
  g1010
  (
    n1047,
    n960
  );


  and
  g1011
  (
    n1048,
    n956,
    n1008,
    n958,
    n959
  );


  or
  g1012
  (
    n1046,
    n1008,
    n957,
    n956
  );


  nor
  g1013
  (
    n1044,
    n955,
    n1008,
    n1009
  );


  buf
  g1014
  (
    n1049,
    n1044
  );


  nand
  g1015
  (
    n1050,
    n1009,
    n1046,
    n1045
  );


  xnor
  g1016
  (
    n1052,
    n1009,
    n1049
  );


  nor
  g1017
  (
    n1051,
    n1044,
    n1009,
    n1010,
    n1046
  );


  nand
  g1018
  (
    n1054,
    n1051,
    n1010,
    n1011
  );


  xnor
  g1019
  (
    n1053,
    n1052,
    n1010,
    n1011
  );


  or
  g1020
  (
    n1058,
    n1013,
    n1053,
    n1014,
    n1015
  );


  not
  g1021
  (
    n1061,
    n1012
  );


  and
  g1022
  (
    n1060,
    n1015,
    n1048,
    n1053
  );


  and
  g1023
  (
    n1057,
    n1048,
    n1015,
    n1013
  );


  nand
  g1024
  (
    n1056,
    n1014,
    n1047,
    n1016
  );


  xor
  g1025
  (
    n1055,
    n1014,
    n1053,
    n1015,
    n1011
  );


  and
  g1026
  (
    n1062,
    n1014,
    n1054,
    n1053
  );


  and
  g1027
  (
    n1059,
    n1013,
    n1054,
    n1047
  );


  not
  g1028
  (
    n1063,
    n1055
  );


  nand
  g1029
  (
    n1066,
    n877,
    n879,
    n1063
  );


  xor
  g1030
  (
    n1065,
    n880,
    n878,
    n1063,
    n879
  );


  xor
  g1031
  (
    n1064,
    n876,
    n880,
    n877,
    n878
  );


  xor
  g1032
  (
    n1068,
    n1065,
    n963,
    n962
  );


  nor
  g1033
  (
    n1067,
    n1066,
    n961,
    n962
  );


  nand
  g1034
  (
    n1071,
    n1067,
    n1058,
    n1059
  );


  or
  g1035
  (
    n1075,
    n1068,
    n1056,
    n1057,
    n1060
  );


  nor
  g1036
  (
    n1076,
    n1057,
    n1067,
    n1058
  );


  and
  g1037
  (
    n1072,
    n1059,
    n1068,
    n1056,
    n604
  );


  or
  g1038
  (
    n1070,
    n1068,
    n1059,
    n1067,
    n1057
  );


  or
  g1039
  (
    n1069,
    n605,
    n1055,
    n1059
  );


  nand
  g1040
  (
    n1074,
    n1056,
    n1058,
    n883,
    n1068
  );


  xor
  g1041
  (
    n1073,
    n605,
    n1057,
    n604,
    n1060
  );


  or
  g1042
  (
    n1089,
    n608,
    n614,
    n990,
    n634
  );


  nand
  g1043
  (
    n1078,
    n1074,
    n610,
    n638,
    n1073
  );


  or
  g1044
  (
    n1091,
    n633,
    n990,
    n1070,
    n611
  );


  nand
  g1045
  (
    n1094,
    n619,
    n611,
    n992,
    n618
  );


  and
  g1046
  (
    n1105,
    n613,
    n626,
    n1071,
    n1070
  );


  xnor
  g1047
  (
    n1095,
    n637,
    n991,
    n608,
    n1073
  );


  or
  g1048
  (
    n1093,
    n988,
    n626,
    n609,
    n1073
  );


  nor
  g1049
  (
    n1084,
    n991,
    n606,
    n621,
    n990
  );


  xnor
  g1050
  (
    n1102,
    n1074,
    n617,
    n630,
    n624
  );


  xor
  g1051
  (
    n1082,
    n1069,
    n616,
    n635
  );


  nand
  g1052
  (
    n1100,
    n638,
    n616,
    n606,
    n628
  );


  nor
  g1053
  (
    n1077,
    n624,
    n993,
    n636,
    n630
  );


  or
  g1054
  (
    n1103,
    n612,
    n637,
    n1071,
    n1075
  );


  xnor
  g1055
  (
    n1096,
    n625,
    n622,
    n1069,
    n623
  );


  xor
  g1056
  (
    n1097,
    n1072,
    n988,
    n1075,
    n614
  );


  nor
  g1057
  (
    n1101,
    n1070,
    n622,
    n1071,
    n988
  );


  or
  g1058
  (
    n1099,
    n636,
    n1072,
    n621,
    n1075
  );


  nand
  g1059
  (
    n1083,
    n615,
    n1071,
    n633,
    n620
  );


  and
  g1060
  (
    n1098,
    n632,
    n612,
    n989,
    n617
  );


  nand
  g1061
  (
    n1085,
    n639,
    n1074,
    n1072,
    n628
  );


  or
  g1062
  (
    n1092,
    n991,
    n1073,
    n639,
    n629
  );


  and
  g1063
  (
    n1086,
    n989,
    n1076,
    n1072,
    n615
  );


  nand
  g1064
  (
    n1081,
    n625,
    n1070,
    n1069,
    n609
  );


  nor
  g1065
  (
    n1080,
    n634,
    n627,
    n993,
    n1075
  );


  xnor
  g1066
  (
    n1087,
    n613,
    n607,
    n620,
    n1069
  );


  and
  g1067
  (
    n1088,
    n1074,
    n631,
    n610,
    n629
  );


  or
  g1068
  (
    n1104,
    n619,
    n627,
    n992
  );


  or
  g1069
  (
    n1079,
    n989,
    n640,
    n623
  );


  nand
  g1070
  (
    KeyWire_0_6,
    n632,
    n631,
    n618,
    n607
  );


  or
  g1071
  (
    n1137,
    n670,
    n653,
    n689,
    n1103
  );


  xor
  g1072
  (
    n1117,
    n1077,
    n683,
    n1084
  );


  xor
  g1073
  (
    n1155,
    n653,
    n676,
    n1076,
    n1094
  );


  xor
  g1074
  (
    n1173,
    n789,
    n691,
    n652,
    n694
  );


  nor
  g1075
  (
    n1141,
    n1007,
    n768,
    n1103,
    n671
  );


  xor
  g1076
  (
    n1180,
    n1096,
    n1089,
    n790,
    n692
  );


  nand
  g1077
  (
    n1157,
    n790,
    n1082,
    n689,
    n676
  );


  and
  g1078
  (
    n1166,
    n692,
    n688,
    n678,
    n666
  );


  and
  g1079
  (
    n1140,
    n1101,
    n1105,
    n1079,
    n1097
  );


  and
  g1080
  (
    n1130,
    n1080,
    n681,
    n1101,
    n1082
  );


  xor
  g1081
  (
    n1182,
    n1005,
    n1077,
    n995,
    n680
  );


  or
  g1082
  (
    n1176,
    n1088,
    n695,
    n1060,
    n693
  );


  nand
  g1083
  (
    n1167,
    n790,
    n832,
    n1093,
    n695
  );


  nand
  g1084
  (
    n1148,
    n670,
    n690,
    n1061,
    n677
  );


  xnor
  g1085
  (
    n1147,
    n690,
    n690,
    n1083,
    n830
  );


  or
  g1086
  (
    n1106,
    n673,
    n691,
    n1097,
    n832
  );


  nor
  g1087
  (
    n1135,
    n1086,
    n1083,
    n769,
    n672
  );


  nand
  g1088
  (
    n1112,
    n993,
    n669,
    n1100,
    n833
  );


  or
  g1089
  (
    n1132,
    n689,
    n687,
    n1084,
    n995
  );


  nor
  g1090
  (
    n1126,
    n963,
    n1088,
    n1094,
    n675
  );


  xor
  g1091
  (
    n1174,
    n1093,
    n685,
    n1060
  );


  nand
  g1092
  (
    n1110,
    n831,
    n666,
    n1099,
    n681
  );


  or
  g1093
  (
    n1160,
    n1089,
    n682,
    n677,
    n1081
  );


  xnor
  g1094
  (
    n1114,
    n680,
    n678,
    n826,
    n1098
  );


  or
  g1095
  (
    n1165,
    n1088,
    n834,
    n668,
    n696
  );


  xor
  g1096
  (
    n1158,
    n1090,
    n1091,
    n1006,
    n768
  );


  xnor
  g1097
  (
    n1113,
    n680,
    n693,
    n1089,
    n1092
  );


  xor
  g1098
  (
    n1125,
    n676,
    n1061,
    n1086,
    n829
  );


  xnor
  g1099
  (
    n1116,
    n670,
    n686,
    n834,
    n667
  );


  or
  g1100
  (
    n1149,
    n694,
    n1092,
    n769,
    n828
  );


  xor
  g1101
  (
    n1153,
    n1086,
    n825,
    n1105,
    n1089
  );


  xnor
  g1102
  (
    n1139,
    n1061,
    n677,
    n682,
    n670
  );


  nand
  g1103
  (
    n1181,
    n1091,
    n830,
    n1087,
    n825
  );


  xor
  g1104
  (
    n1136,
    n1102,
    n687,
    n675,
    n1098
  );


  or
  g1105
  (
    n1115,
    n833,
    n829,
    n1105,
    n674
  );


  nand
  g1106
  (
    n1169,
    n1080,
    n691,
    n685,
    n834
  );


  nand
  g1107
  (
    n1119,
    n1098,
    n1095,
    n684,
    n1085
  );


  xnor
  g1108
  (
    n1152,
    n1093,
    n684,
    n769,
    n669
  );


  nand
  g1109
  (
    n1163,
    n1087,
    n684,
    n668,
    n665
  );


  nand
  g1110
  (
    n1127,
    n790,
    n1101,
    n688,
    n1097
  );


  and
  g1111
  (
    n1120,
    n1078,
    n676,
    n831,
    n667
  );


  or
  g1112
  (
    n1134,
    n1104,
    n692,
    n768,
    n827
  );


  xor
  g1113
  (
    n1164,
    n682,
    n686,
    n1082,
    n1061
  );


  xnor
  g1114
  (
    n1138,
    n829,
    n652,
    n681,
    n830
  );


  xor
  g1115
  (
    n1144,
    n831,
    n692,
    n1088,
    n1090
  );


  xor
  g1116
  (
    n1133,
    n693,
    n672,
    n1092,
    n688
  );


  nor
  g1117
  (
    n1122,
    n679,
    n1101,
    n1076,
    n668
  );


  or
  g1118
  (
    n1109,
    n828,
    n1095,
    n690,
    n695
  );


  nand
  g1119
  (
    n1121,
    n1099,
    n675,
    n678,
    n1086
  );


  xor
  g1120
  (
    n1184,
    n665,
    n1006,
    n1099,
    n687
  );


  or
  g1121
  (
    n1143,
    n674,
    n685,
    n1104,
    n653
  );


  and
  g1122
  (
    n1156,
    n675,
    n666,
    n1005,
    n1078
  );


  and
  g1123
  (
    n1128,
    n1099,
    n1094,
    n1079,
    n683
  );


  nand
  g1124
  (
    n1170,
    n667,
    n1096,
    n665,
    n1105
  );


  xnor
  g1125
  (
    n1131,
    n1087,
    n1062,
    n669,
    n1095
  );


  nor
  g1126
  (
    n1154,
    n1091,
    n1085,
    n1096,
    n684
  );


  nor
  g1127
  (
    n1177,
    n995,
    n1077,
    n1083,
    n691
  );


  nor
  g1128
  (
    n1161,
    n696,
    n1103,
    n681,
    n672
  );


  and
  g1129
  (
    n1129,
    n1079,
    n1095,
    n994,
    n1080
  );


  nor
  g1130
  (
    n1107,
    n1096,
    n680,
    n767,
    n827
  );


  or
  g1131
  (
    n1168,
    n1077,
    n832,
    n994,
    n1007
  );


  or
  g1132
  (
    n1108,
    n674,
    n673,
    n1104,
    n679
  );


  or
  g1133
  (
    n1124,
    n1097,
    n679,
    n689,
    n1104
  );


  nor
  g1134
  (
    n1111,
    n767,
    n683,
    n1006,
    n696
  );


  xnor
  g1135
  (
    n1162,
    n1082,
    n1007,
    n677,
    n1087
  );


  nor
  g1136
  (
    n1172,
    n1091,
    n1102,
    n1100,
    n833
  );


  or
  g1137
  (
    n1123,
    n694,
    n666,
    n1100,
    n768
  );


  and
  g1138
  (
    n1118,
    n1080,
    n683,
    n994,
    n1090
  );


  and
  g1139
  (
    n1185,
    n695,
    n1062,
    n671,
    n1085
  );


  or
  g1140
  (
    n1142,
    n1079,
    n826,
    n682,
    n1081
  );


  and
  g1141
  (
    n1175,
    n1081,
    n678,
    n668,
    n673
  );


  xnor
  g1142
  (
    n1159,
    n1007,
    n789,
    n686,
    n1084
  );


  xor
  g1143
  (
    n1171,
    n1085,
    n693,
    n679,
    n769
  );


  nand
  g1144
  (
    n1150,
    n1078,
    n1081,
    n1100,
    n1094
  );


  xor
  g1145
  (
    n1179,
    n1098,
    n1078,
    n1076,
    n669
  );


  xnor
  g1146
  (
    KeyWire_0_3,
    n1103,
    n696,
    n674,
    n1062
  );


  or
  g1147
  (
    n1183,
    n1005,
    n671,
    n687,
    n1083
  );


  nand
  g1148
  (
    n1151,
    n1102,
    n673,
    n672,
    n1062
  );


  nand
  g1149
  (
    n1146,
    n1005,
    n686,
    n671,
    n1102
  );


  xor
  g1150
  (
    n1178,
    n1006,
    n694,
    n688,
    n1092
  );


  nor
  g1151
  (
    n1145,
    n653,
    n667,
    n1093,
    n1090
  );


  xnor
  g1152
  (
    n1192,
    n1037,
    n1020,
    n1024,
    n1131
  );


  nand
  g1153
  (
    n1230,
    n1038,
    n1034,
    n1031,
    n1170
  );


  nor
  g1154
  (
    n1216,
    n1153,
    n1030,
    n1032,
    n1171
  );


  nand
  g1155
  (
    n1229,
    n1016,
    n1157,
    n1127,
    n1160
  );


  nor
  g1156
  (
    n1227,
    n1020,
    n1040,
    n1114,
    n1030
  );


  or
  g1157
  (
    n1219,
    n1147,
    n1023,
    n1151,
    n1025
  );


  or
  g1158
  (
    n1211,
    n1038,
    n1163,
    n1020,
    n1155
  );


  nand
  g1159
  (
    n1200,
    n1132,
    n1154,
    n1036,
    n1119
  );


  xor
  g1160
  (
    n1197,
    n1134,
    n1035,
    n1039
  );


  xnor
  g1161
  (
    n1222,
    n1025,
    n1040,
    n1024,
    n1112
  );


  or
  g1162
  (
    n1205,
    n1027,
    n1123,
    n1106,
    n1016
  );


  nor
  g1163
  (
    n1215,
    n1041,
    n1031,
    n1025,
    n1034
  );


  nand
  g1164
  (
    n1206,
    n1121,
    n1166,
    n1019,
    n1028
  );


  xnor
  g1165
  (
    n1187,
    n1032,
    n1038,
    n1035,
    n1041
  );


  nand
  g1166
  (
    n1218,
    n1181,
    n1034,
    n1023,
    n1136
  );


  nand
  g1167
  (
    n1203,
    n1019,
    n1018,
    n1037,
    n1032
  );


  and
  g1168
  (
    n1234,
    n1149,
    n1036,
    n1043
  );


  xnor
  g1169
  (
    n1225,
    n1029,
    n1145,
    n1152,
    n1018
  );


  and
  g1170
  (
    n1214,
    n1159,
    n1107,
    n1043,
    n1041
  );


  nand
  g1171
  (
    n1208,
    n1180,
    n1028,
    n1019,
    n1026
  );


  nand
  g1172
  (
    n1228,
    n1037,
    n1021,
    n1169,
    n1024
  );


  nor
  g1173
  (
    n1191,
    n1022,
    n1033,
    n1030,
    n1115
  );


  or
  g1174
  (
    n1231,
    n1175,
    n1109,
    n1018,
    n1017
  );


  or
  g1175
  (
    n1202,
    n1024,
    n1122,
    n1138,
    n1164
  );


  or
  g1176
  (
    n1212,
    n1028,
    n1150,
    n1033,
    n1022
  );


  nor
  g1177
  (
    n1220,
    n1117,
    n1186,
    n1034,
    n1146
  );


  and
  g1178
  (
    n1198,
    n1130,
    n1177,
    n1184,
    n1026
  );


  nor
  g1179
  (
    n1213,
    n1144,
    n1037,
    n1035,
    n1137
  );


  or
  g1180
  (
    KeyWire_0_2,
    n1029,
    n1040,
    n1042,
    n1026
  );


  nor
  g1181
  (
    n1224,
    n1043,
    n1029,
    n1124
  );


  nor
  g1182
  (
    n1190,
    n1125,
    n1156,
    n1025,
    n1141
  );


  or
  g1183
  (
    n1233,
    n1135,
    n1167,
    n1022,
    n1030
  );


  and
  g1184
  (
    n1195,
    n1027,
    n1128,
    n1113,
    n1039
  );


  and
  g1185
  (
    n1188,
    n1023,
    n1027,
    n1021
  );


  xnor
  g1186
  (
    n1194,
    n1168,
    n1133,
    n1040,
    n1039
  );


  and
  g1187
  (
    n1217,
    n1142,
    n1031,
    n1139,
    n1038
  );


  xnor
  g1188
  (
    n1207,
    n1162,
    n1173,
    n1126,
    n1174
  );


  xor
  g1189
  (
    n1210,
    n1111,
    n1023,
    n1021,
    n1016
  );


  nand
  g1190
  (
    n1199,
    n1027,
    n1179,
    n1143,
    n1018
  );


  nor
  g1191
  (
    n1223,
    n1116,
    n1118,
    n1017,
    n1120
  );


  nor
  g1192
  (
    n1204,
    n1036,
    n1158,
    n1161,
    n1028
  );


  xor
  g1193
  (
    n1201,
    n1031,
    n1042,
    n1185,
    n1178
  );


  or
  g1194
  (
    n1226,
    n1041,
    n1033,
    n1176
  );


  xnor
  g1195
  (
    n1189,
    n1140,
    n1110,
    n1019,
    n1039
  );


  nor
  g1196
  (
    n1232,
    n1043,
    n1017,
    n1042
  );


  nand
  g1197
  (
    n1196,
    n1172,
    n1032,
    n1182,
    n1017
  );


  nor
  g1198
  (
    n1209,
    n1026,
    n1020,
    n1183,
    n1165
  );


  nor
  g1199
  (
    n1193,
    n1108,
    n1022,
    n1129,
    n1148
  );


  or
  g1200
  (
    n1244,
    n1224,
    n1211,
    n1193,
    n1208
  );


  nand
  g1201
  (
    n1236,
    n1226,
    n1201,
    n1221,
    n1217
  );


  xnor
  g1202
  (
    n1237,
    n1190,
    n1204,
    n1189,
    n1228
  );


  and
  g1203
  (
    n1240,
    n1218,
    n1216,
    n1234,
    n1200
  );


  nor
  g1204
  (
    n1241,
    n1225,
    n1212,
    n1209,
    n1207
  );


  and
  g1205
  (
    n1246,
    n1222,
    n1220,
    n1202,
    n1232
  );


  xnor
  g1206
  (
    n1245,
    n1187,
    n1213,
    n1194,
    n1205
  );


  xnor
  g1207
  (
    n1243,
    n1230,
    n1215,
    n1198,
    n1214
  );


  nand
  g1208
  (
    n1242,
    n1197,
    n1196,
    n1219,
    n1231
  );


  and
  g1209
  (
    n1239,
    n1223,
    n1188,
    n1206,
    n1203
  );


  nand
  g1210
  (
    n1238,
    n1227,
    n1210,
    n1233,
    n1199
  );


  or
  g1211
  (
    n1235,
    n1229,
    n1191,
    n1192,
    n1195
  );


  or
  g1212
  (
    n1249,
    n1241,
    n1235,
    n1237,
    n1240
  );


  or
  g1213
  (
    n1247,
    n1238,
    n1239,
    n1246,
    n1244
  );


  or
  g1214
  (
    n1248,
    n1242,
    n1243,
    n1236,
    n1245
  );


  xnor
  KeyGate_0_0
  (
    n180,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n39,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1221,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1186,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n618,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n906,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1090,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1042,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n676,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n403,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n652,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n433,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n550,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n657,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n150,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n758,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n591,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n968,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n574,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n284,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n337,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n398,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n1029,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n423,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n285,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n492,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n599,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n102,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n205,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n865,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1002,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n576,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

