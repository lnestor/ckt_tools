

module Stat_996_1734
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n847,
  n853,
  n859,
  n861,
  n823,
  n829,
  n822,
  n854,
  n825,
  n851,
  n839,
  n858,
  n846,
  n855,
  n833,
  n824,
  n845,
  n996,
  n1003,
  n1002,
  n1006,
  n1001,
  n1010,
  n1008,
  n1011,
  n1012,
  n1014,
  n1013,
  n1015,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n847;
  output n853;
  output n859;
  output n861;
  output n823;
  output n829;
  output n822;
  output n854;
  output n825;
  output n851;
  output n839;
  output n858;
  output n846;
  output n855;
  output n833;
  output n824;
  output n845;
  output n996;
  output n1003;
  output n1002;
  output n1006;
  output n1001;
  output n1010;
  output n1008;
  output n1011;
  output n1012;
  output n1014;
  output n1013;
  output n1015;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n826;
  wire n827;
  wire n828;
  wire n830;
  wire n831;
  wire n832;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n848;
  wire n849;
  wire n850;
  wire n852;
  wire n856;
  wire n857;
  wire n860;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1004;
  wire n1005;
  wire n1007;
  wire n1009;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    n90,
    n14
  );


  buf
  g1
  (
    n65,
    n2
  );


  buf
  g2
  (
    n54,
    n18
  );


  buf
  g3
  (
    n21,
    n4
  );


  not
  g4
  (
    n20,
    n12
  );


  not
  g5
  (
    n69,
    n12
  );


  not
  g6
  (
    n82,
    n3
  );


  buf
  g7
  (
    n52,
    n3
  );


  not
  g8
  (
    n92,
    n16
  );


  buf
  g9
  (
    KeyWire_0_18,
    n6
  );


  not
  g10
  (
    n76,
    n2
  );


  buf
  g11
  (
    n67,
    n17
  );


  not
  g12
  (
    n41,
    n6
  );


  not
  g13
  (
    n38,
    n11
  );


  not
  g14
  (
    n79,
    n6
  );


  buf
  g15
  (
    n93,
    n3
  );


  buf
  g16
  (
    n36,
    n3
  );


  buf
  g17
  (
    n40,
    n18
  );


  buf
  g18
  (
    n68,
    n1
  );


  not
  g19
  (
    n45,
    n12
  );


  buf
  g20
  (
    n29,
    n5
  );


  not
  g21
  (
    n72,
    n7
  );


  not
  g22
  (
    n56,
    n9
  );


  not
  g23
  (
    n87,
    n11
  );


  buf
  g24
  (
    n74,
    n2
  );


  buf
  g25
  (
    KeyWire_0_6,
    n10
  );


  buf
  g26
  (
    n31,
    n16
  );


  buf
  g27
  (
    n35,
    n19
  );


  not
  g28
  (
    n64,
    n17
  );


  not
  g29
  (
    n62,
    n5
  );


  not
  g30
  (
    n60,
    n8
  );


  buf
  g31
  (
    n51,
    n15
  );


  not
  g32
  (
    n77,
    n15
  );


  not
  g33
  (
    n37,
    n10
  );


  buf
  g34
  (
    n33,
    n14
  );


  not
  g35
  (
    n94,
    n16
  );


  buf
  g36
  (
    n50,
    n9
  );


  buf
  g37
  (
    n26,
    n13
  );


  buf
  g38
  (
    n73,
    n10
  );


  not
  g39
  (
    n63,
    n16
  );


  buf
  g40
  (
    n42,
    n13
  );


  buf
  g41
  (
    n66,
    n7
  );


  buf
  g42
  (
    n22,
    n13
  );


  not
  g43
  (
    n75,
    n19
  );


  buf
  g44
  (
    n95,
    n5
  );


  buf
  g45
  (
    n47,
    n8
  );


  not
  g46
  (
    n25,
    n4
  );


  not
  g47
  (
    n58,
    n7
  );


  not
  g48
  (
    n32,
    n4
  );


  not
  g49
  (
    n30,
    n12
  );


  not
  g50
  (
    n89,
    n5
  );


  not
  g51
  (
    n24,
    n1
  );


  not
  g52
  (
    n61,
    n13
  );


  buf
  g53
  (
    n49,
    n15
  );


  not
  g54
  (
    n43,
    n17
  );


  not
  g55
  (
    n53,
    n7
  );


  buf
  g56
  (
    n78,
    n2
  );


  not
  g57
  (
    n23,
    n17
  );


  buf
  g58
  (
    n84,
    n19
  );


  buf
  g59
  (
    n57,
    n14
  );


  not
  g60
  (
    n59,
    n9
  );


  buf
  g61
  (
    n71,
    n1
  );


  buf
  g62
  (
    n70,
    n18
  );


  buf
  g63
  (
    n83,
    n1
  );


  buf
  g64
  (
    n34,
    n11
  );


  buf
  g65
  (
    n80,
    n4
  );


  not
  g66
  (
    n48,
    n15
  );


  not
  g67
  (
    n91,
    n9
  );


  not
  g68
  (
    n44,
    n10
  );


  not
  g69
  (
    n55,
    n18
  );


  buf
  g70
  (
    n88,
    n8
  );


  buf
  g71
  (
    n27,
    n19
  );


  not
  g72
  (
    n39,
    n6
  );


  not
  g73
  (
    n46,
    n11
  );


  buf
  g74
  (
    KeyWire_0_12,
    n8
  );


  buf
  g75
  (
    n86,
    n14
  );


  buf
  g76
  (
    n170,
    n54
  );


  not
  g77
  (
    n128,
    n28
  );


  not
  g78
  (
    n138,
    n32
  );


  not
  g79
  (
    n123,
    n66
  );


  buf
  g80
  (
    n219,
    n90
  );


  buf
  g81
  (
    n236,
    n68
  );


  buf
  g82
  (
    n206,
    n24
  );


  not
  g83
  (
    n186,
    n42
  );


  buf
  g84
  (
    n241,
    n39
  );


  not
  g85
  (
    n243,
    n80
  );


  buf
  g86
  (
    n133,
    n85
  );


  not
  g87
  (
    n254,
    n61
  );


  buf
  g88
  (
    n146,
    n73
  );


  not
  g89
  (
    n118,
    n89
  );


  not
  g90
  (
    n106,
    n79
  );


  buf
  g91
  (
    n177,
    n86
  );


  buf
  g92
  (
    n176,
    n95
  );


  not
  g93
  (
    n226,
    n51
  );


  buf
  g94
  (
    n126,
    n31
  );


  buf
  g95
  (
    n141,
    n72
  );


  not
  g96
  (
    n114,
    n94
  );


  not
  g97
  (
    n131,
    n88
  );


  buf
  g98
  (
    n101,
    n77
  );


  buf
  g99
  (
    n215,
    n29
  );


  not
  g100
  (
    n143,
    n86
  );


  buf
  g101
  (
    n213,
    n83
  );


  buf
  g102
  (
    n129,
    n49
  );


  not
  g103
  (
    n160,
    n35
  );


  buf
  g104
  (
    n223,
    n85
  );


  not
  g105
  (
    n127,
    n92
  );


  not
  g106
  (
    n192,
    n20
  );


  buf
  g107
  (
    n159,
    n91
  );


  buf
  g108
  (
    n258,
    n74
  );


  not
  g109
  (
    n207,
    n53
  );


  buf
  g110
  (
    n154,
    n50
  );


  not
  g111
  (
    n224,
    n36
  );


  buf
  g112
  (
    n252,
    n74
  );


  not
  g113
  (
    n181,
    n83
  );


  buf
  g114
  (
    n193,
    n84
  );


  not
  g115
  (
    n105,
    n85
  );


  buf
  g116
  (
    n257,
    n85
  );


  not
  g117
  (
    n102,
    n22
  );


  buf
  g118
  (
    n250,
    n79
  );


  buf
  g119
  (
    n124,
    n26
  );


  not
  g120
  (
    n247,
    n42
  );


  not
  g121
  (
    n104,
    n71
  );


  not
  g122
  (
    n256,
    n42
  );


  not
  g123
  (
    n168,
    n73
  );


  buf
  g124
  (
    n240,
    n62
  );


  not
  g125
  (
    n117,
    n48
  );


  not
  g126
  (
    n98,
    n94
  );


  buf
  g127
  (
    n245,
    n56
  );


  not
  g128
  (
    n188,
    n95
  );


  not
  g129
  (
    n122,
    n43
  );


  buf
  g130
  (
    n116,
    n56
  );


  not
  g131
  (
    KeyWire_0_1,
    n29
  );


  not
  g132
  (
    n136,
    n23
  );


  buf
  g133
  (
    n169,
    n88
  );


  not
  g134
  (
    n121,
    n80
  );


  not
  g135
  (
    n230,
    n29
  );


  not
  g136
  (
    n195,
    n39
  );


  not
  g137
  (
    n175,
    n90
  );


  not
  g138
  (
    n189,
    n42
  );


  buf
  g139
  (
    n130,
    n36
  );


  not
  g140
  (
    n179,
    n67
  );


  buf
  g141
  (
    n199,
    n65
  );


  not
  g142
  (
    n210,
    n54
  );


  not
  g143
  (
    n182,
    n59
  );


  buf
  g144
  (
    n161,
    n89
  );


  buf
  g145
  (
    n261,
    n71
  );


  buf
  g146
  (
    n209,
    n23
  );


  not
  g147
  (
    n204,
    n47
  );


  buf
  g148
  (
    n184,
    n32
  );


  not
  g149
  (
    n144,
    n27
  );


  not
  g150
  (
    KeyWire_0_20,
    n76
  );


  not
  g151
  (
    n246,
    n89
  );


  buf
  g152
  (
    n191,
    n78
  );


  buf
  g153
  (
    n142,
    n20
  );


  not
  g154
  (
    n125,
    n48
  );


  not
  g155
  (
    n231,
    n46
  );


  not
  g156
  (
    n132,
    n81
  );


  not
  g157
  (
    n180,
    n52
  );


  not
  g158
  (
    n155,
    n36
  );


  buf
  g159
  (
    n242,
    n67
  );


  buf
  g160
  (
    n200,
    n95
  );


  not
  g161
  (
    n233,
    n67
  );


  not
  g162
  (
    n218,
    n81
  );


  not
  g163
  (
    n238,
    n39
  );


  buf
  g164
  (
    n194,
    n87
  );


  buf
  g165
  (
    n96,
    n75
  );


  buf
  g166
  (
    n119,
    n21
  );


  not
  g167
  (
    n147,
    n62
  );


  not
  g168
  (
    n244,
    n45
  );


  buf
  g169
  (
    n251,
    n63
  );


  not
  g170
  (
    n97,
    n94
  );


  not
  g171
  (
    n100,
    n76
  );


  not
  g172
  (
    n197,
    n34
  );


  not
  g173
  (
    n260,
    n69
  );


  not
  g174
  (
    n151,
    n66
  );


  buf
  g175
  (
    n112,
    n64
  );


  buf
  g176
  (
    n221,
    n57
  );


  not
  g177
  (
    KeyWire_0_25,
    n86
  );


  not
  g178
  (
    n157,
    n61
  );


  not
  g179
  (
    n145,
    n75
  );


  buf
  g180
  (
    n173,
    n60
  );


  buf
  g181
  (
    n263,
    n90
  );


  buf
  g182
  (
    n178,
    n48
  );


  not
  g183
  (
    n205,
    n93
  );


  not
  g184
  (
    n220,
    n74
  );


  not
  g185
  (
    n115,
    n37
  );


  not
  g186
  (
    n139,
    n64
  );


  not
  g187
  (
    n212,
    n57
  );


  not
  g188
  (
    n248,
    n94
  );


  buf
  g189
  (
    n167,
    n80
  );


  buf
  g190
  (
    n137,
    n59
  );


  not
  g191
  (
    n201,
    n74
  );


  not
  g192
  (
    n267,
    n34
  );


  buf
  g193
  (
    n196,
    n59
  );


  buf
  g194
  (
    n152,
    n80
  );


  buf
  g195
  (
    n158,
    n40
  );


  not
  g196
  (
    n214,
    n55
  );


  buf
  g197
  (
    n149,
    n75
  );


  buf
  g198
  (
    n107,
    n68
  );


  buf
  g199
  (
    n172,
    n53
  );


  not
  g200
  (
    n111,
    n31
  );


  buf
  g201
  (
    n163,
    n62
  );


  not
  g202
  (
    n264,
    n92
  );


  not
  g203
  (
    n183,
    n26
  );


  nor
  g204
  (
    n140,
    n37,
    n72,
    n40,
    n45
  );


  and
  g205
  (
    n185,
    n92,
    n31,
    n69,
    n70
  );


  or
  g206
  (
    n265,
    n83,
    n76,
    n23,
    n32
  );


  or
  g207
  (
    n208,
    n86,
    n28,
    n46,
    n21
  );


  xor
  g208
  (
    n110,
    n88,
    n22,
    n64,
    n50
  );


  nand
  g209
  (
    n255,
    n44,
    n55,
    n45,
    n53
  );


  xnor
  g210
  (
    n203,
    n28,
    n37,
    n81,
    n51
  );


  and
  g211
  (
    n135,
    n79,
    n25,
    n20,
    n78
  );


  xnor
  g212
  (
    n156,
    n39,
    n63,
    n26,
    n65
  );


  nor
  g213
  (
    n259,
    n65,
    n89,
    n82,
    n41
  );


  or
  g214
  (
    n217,
    n47,
    n63,
    n55,
    n52
  );


  xor
  g215
  (
    n109,
    n62,
    n34,
    n56,
    n55
  );


  xnor
  g216
  (
    n150,
    n40,
    n81,
    n72,
    n38
  );


  xor
  g217
  (
    n162,
    n30,
    n51,
    n46,
    n24
  );


  nand
  g218
  (
    n229,
    n67,
    n84,
    n25,
    n50
  );


  nor
  g219
  (
    n235,
    n58,
    n75,
    n43,
    n69
  );


  xor
  g220
  (
    n171,
    n38,
    n88,
    n47,
    n34
  );


  nor
  g221
  (
    n198,
    n71,
    n31,
    n49,
    n52
  );


  nand
  g222
  (
    KeyWire_0_0,
    n60,
    n35,
    n30
  );


  or
  g223
  (
    n239,
    n33,
    n87,
    n23
  );


  xor
  g224
  (
    n222,
    n91,
    n30,
    n63,
    n20
  );


  nor
  g225
  (
    KeyWire_0_10,
    n93,
    n51,
    n37,
    n49
  );


  nand
  g226
  (
    n266,
    n48,
    n57,
    n95,
    n32
  );


  and
  g227
  (
    n237,
    n79,
    n92,
    n70,
    n49
  );


  xor
  g228
  (
    n190,
    n68,
    n72,
    n60,
    n84
  );


  and
  g229
  (
    n216,
    n70,
    n22,
    n93,
    n43
  );


  xor
  g230
  (
    n249,
    n47,
    n27,
    n35,
    n21
  );


  or
  g231
  (
    n120,
    n46,
    n93,
    n50,
    n84
  );


  nor
  g232
  (
    n228,
    n41,
    n44,
    n54,
    n33
  );


  nor
  g233
  (
    n113,
    n25,
    n54,
    n22,
    n52
  );


  nand
  g234
  (
    n153,
    n78,
    n24,
    n69,
    n73
  );


  or
  g235
  (
    n234,
    n27,
    n36,
    n82,
    n45
  );


  nand
  g236
  (
    n202,
    n66,
    n44,
    n24,
    n77
  );


  xor
  g237
  (
    n166,
    n91,
    n91,
    n64,
    n38
  );


  xnor
  g238
  (
    n148,
    n35,
    n66,
    n38,
    n25
  );


  xnor
  g239
  (
    n134,
    n56,
    n83,
    n78,
    n76
  );


  and
  g240
  (
    n227,
    n58,
    n58,
    n28,
    n73
  );


  xnor
  g241
  (
    n262,
    n71,
    n87,
    n82,
    n33
  );


  nor
  g242
  (
    n165,
    n41,
    n58,
    n57,
    n65
  );


  xnor
  g243
  (
    n211,
    n61,
    n77,
    n43,
    n59
  );


  and
  g244
  (
    n253,
    n70,
    n82,
    n60,
    n41
  );


  or
  g245
  (
    n232,
    n33,
    n53,
    n26,
    n90
  );


  xor
  g246
  (
    n99,
    n68,
    n21,
    n77,
    n27
  );


  nand
  g247
  (
    n108,
    n29,
    n40,
    n44,
    n61
  );


  buf
  g248
  (
    n320,
    n113
  );


  buf
  g249
  (
    n402,
    n228
  );


  buf
  g250
  (
    n341,
    n163
  );


  buf
  g251
  (
    n376,
    n171
  );


  buf
  g252
  (
    n325,
    n178
  );


  buf
  g253
  (
    n358,
    n97
  );


  not
  g254
  (
    n279,
    n167
  );


  not
  g255
  (
    n385,
    n168
  );


  buf
  g256
  (
    n407,
    n188
  );


  not
  g257
  (
    n367,
    n225
  );


  not
  g258
  (
    n274,
    n239
  );


  buf
  g259
  (
    n433,
    n174
  );


  buf
  g260
  (
    n340,
    n237
  );


  buf
  g261
  (
    n375,
    n99
  );


  buf
  g262
  (
    n398,
    n184
  );


  and
  g263
  (
    n276,
    n236,
    n96
  );


  and
  g264
  (
    n396,
    n172,
    n119,
    n97,
    n187
  );


  xnor
  g265
  (
    n374,
    n122,
    n247,
    n175,
    n134
  );


  nand
  g266
  (
    n302,
    n192,
    n151,
    n169,
    n229
  );


  or
  g267
  (
    n424,
    n216,
    n236,
    n229,
    n153
  );


  xnor
  g268
  (
    n361,
    n194,
    n217,
    n111,
    n181
  );


  nand
  g269
  (
    n287,
    n175,
    n241,
    n205,
    n135
  );


  nand
  g270
  (
    n411,
    n206,
    n137,
    n99,
    n249
  );


  and
  g271
  (
    n270,
    n183,
    n148,
    n109,
    n116
  );


  xor
  g272
  (
    n326,
    n199,
    n143,
    n215,
    n123
  );


  nor
  g273
  (
    n432,
    n185,
    n190,
    n114,
    n215
  );


  xor
  g274
  (
    n271,
    n236,
    n230,
    n181,
    n136
  );


  nand
  g275
  (
    n405,
    n162,
    n249,
    n195,
    n173
  );


  xor
  g276
  (
    n351,
    n138,
    n96,
    n165,
    n222
  );


  or
  g277
  (
    n364,
    n112,
    n153,
    n128,
    n133
  );


  xnor
  g278
  (
    n386,
    n174,
    n222,
    n111,
    n235
  );


  or
  g279
  (
    n378,
    n240,
    n245,
    n209,
    n230
  );


  or
  g280
  (
    n395,
    n202,
    n158,
    n107
  );


  nor
  g281
  (
    n331,
    n243,
    n167,
    n116,
    n113
  );


  nand
  g282
  (
    n418,
    n98,
    n140,
    n244,
    n189
  );


  nand
  g283
  (
    n359,
    n241,
    n121,
    n128,
    n103
  );


  or
  g284
  (
    n306,
    n120,
    n185,
    n176,
    n195
  );


  nor
  g285
  (
    n350,
    n168,
    n145,
    n108,
    n191
  );


  and
  g286
  (
    n362,
    n147,
    n197,
    n110,
    n192
  );


  xnor
  g287
  (
    n322,
    n211,
    n231,
    n208,
    n108
  );


  nand
  g288
  (
    n428,
    n230,
    n196,
    n99,
    n156
  );


  nand
  g289
  (
    n346,
    n234,
    n240,
    n249,
    n159
  );


  nand
  g290
  (
    n363,
    n109,
    n227,
    n200,
    n151
  );


  nand
  g291
  (
    n409,
    n121,
    n103,
    n193,
    n170
  );


  xor
  g292
  (
    n408,
    n240,
    n219,
    n118
  );


  or
  g293
  (
    n347,
    n242,
    n235,
    n111,
    n155
  );


  nor
  g294
  (
    n368,
    n177,
    n115,
    n119,
    n158
  );


  or
  g295
  (
    n397,
    n198,
    n98,
    n213,
    n138
  );


  nand
  g296
  (
    n399,
    n197,
    n229,
    n231,
    n221
  );


  or
  g297
  (
    n284,
    n221,
    n247,
    n212,
    n220
  );


  xnor
  g298
  (
    n419,
    n150,
    n151,
    n189
  );


  and
  g299
  (
    n312,
    n137,
    n225,
    n199,
    n119
  );


  xor
  g300
  (
    n327,
    n130,
    n240,
    n113,
    n194
  );


  nand
  g301
  (
    n308,
    n223,
    n96,
    n221,
    n210
  );


  and
  g302
  (
    n328,
    n135,
    n142,
    n213,
    n150
  );


  or
  g303
  (
    n373,
    n165,
    n202,
    n195,
    n196
  );


  nand
  g304
  (
    n281,
    n134,
    n106,
    n180,
    n205
  );


  or
  g305
  (
    n336,
    n132,
    n237,
    n172,
    n158
  );


  and
  g306
  (
    n289,
    n188,
    n217,
    n155,
    n128
  );


  xnor
  g307
  (
    n348,
    n232,
    n171,
    n234,
    n250
  );


  or
  g308
  (
    n272,
    n126,
    n124,
    n242,
    n233
  );


  and
  g309
  (
    n382,
    n126,
    n181,
    n215,
    n216
  );


  and
  g310
  (
    n410,
    n231,
    n179,
    n131,
    n187
  );


  nand
  g311
  (
    n329,
    n149,
    n248,
    n244,
    n126
  );


  or
  g312
  (
    n377,
    n206,
    n113,
    n176,
    n104
  );


  xnor
  g313
  (
    n427,
    n161,
    n100,
    n132,
    n196
  );


  xor
  g314
  (
    n422,
    n221,
    n174,
    n130,
    n208
  );


  nand
  g315
  (
    n273,
    n227,
    n209,
    n120,
    n219
  );


  and
  g316
  (
    n269,
    n140,
    n106,
    n129,
    n114
  );


  and
  g317
  (
    n290,
    n211,
    n145,
    n232,
    n212
  );


  nand
  g318
  (
    n318,
    n201,
    n124,
    n169,
    n212
  );


  xor
  g319
  (
    n416,
    n228,
    n164,
    n222,
    n200
  );


  and
  g320
  (
    n390,
    n237,
    n157,
    n108,
    n97
  );


  xnor
  g321
  (
    n349,
    n142,
    n248,
    n239,
    n227
  );


  nor
  g322
  (
    n356,
    n143,
    n225,
    n144,
    n114
  );


  nand
  g323
  (
    n389,
    n238,
    n127,
    n122,
    n149
  );


  nor
  g324
  (
    n426,
    n201,
    n244,
    n156,
    n188
  );


  nor
  g325
  (
    n342,
    n117,
    n131,
    n190,
    n139
  );


  and
  g326
  (
    n299,
    n243,
    n248,
    n152,
    n239
  );


  nand
  g327
  (
    n414,
    n204,
    n152,
    n186,
    n238
  );


  or
  g328
  (
    n310,
    n105,
    n123,
    n144,
    n203
  );


  nand
  g329
  (
    n429,
    n233,
    n206,
    n183,
    n179
  );


  nand
  g330
  (
    n425,
    n160,
    n136,
    n138,
    n139
  );


  or
  g331
  (
    n335,
    n235,
    n249,
    n125,
    n115
  );


  xnor
  g332
  (
    n415,
    n200,
    n224,
    n198,
    n176
  );


  xnor
  g333
  (
    n420,
    n218,
    n131,
    n127,
    n183
  );


  nand
  g334
  (
    n365,
    n107,
    n142,
    n190,
    n116
  );


  nor
  g335
  (
    KeyWire_0_28,
    n223,
    n134,
    n122,
    n129
  );


  xor
  g336
  (
    n288,
    n167,
    n178,
    n155,
    n106
  );


  nand
  g337
  (
    n295,
    n193,
    n118,
    n112,
    n245
  );


  or
  g338
  (
    n304,
    n130,
    n191,
    n134,
    n166
  );


  or
  g339
  (
    n417,
    n212,
    n170,
    n104,
    n100
  );


  nand
  g340
  (
    n309,
    n124,
    n157,
    n173,
    n120
  );


  nand
  g341
  (
    n394,
    n125,
    n195,
    n144,
    n185
  );


  or
  g342
  (
    n391,
    n206,
    n207,
    n238,
    n104
  );


  and
  g343
  (
    n285,
    n204,
    n151,
    n178,
    n172
  );


  or
  g344
  (
    n303,
    n99,
    n148,
    n140,
    n107
  );


  nand
  g345
  (
    n400,
    n216,
    n147,
    n235,
    n196
  );


  nor
  g346
  (
    n380,
    n220,
    n182,
    n203,
    n210
  );


  xor
  g347
  (
    n423,
    n105,
    n141,
    n107,
    n121
  );


  xnor
  g348
  (
    n401,
    n191,
    n149,
    n245,
    n180
  );


  nand
  g349
  (
    n317,
    n236,
    n193,
    n157,
    n216
  );


  or
  g350
  (
    n421,
    n173,
    n186,
    n140,
    n241
  );


  or
  g351
  (
    n297,
    n142,
    n184,
    n226,
    n137
  );


  nand
  g352
  (
    n323,
    n244,
    n157,
    n116,
    n115
  );


  or
  g353
  (
    n360,
    n210,
    n123,
    n171,
    n177
  );


  and
  g354
  (
    n333,
    n174,
    n207,
    n169,
    n233
  );


  nor
  g355
  (
    n313,
    n159,
    n154,
    n160,
    n138
  );


  nor
  g356
  (
    n379,
    n180,
    n209,
    n127,
    n125
  );


  xnor
  g357
  (
    n275,
    n145,
    n143,
    n246,
    n126
  );


  xor
  g358
  (
    n352,
    n163,
    n154,
    n207,
    n143
  );


  and
  g359
  (
    n283,
    n121,
    n178,
    n227,
    n193
  );


  or
  g360
  (
    n381,
    n135,
    n247,
    n191,
    n110
  );


  xor
  g361
  (
    n301,
    n208,
    n161,
    n164,
    n246
  );


  nor
  g362
  (
    n372,
    n199,
    n186,
    n213,
    n228
  );


  and
  g363
  (
    n314,
    n203,
    n229,
    n243,
    n175
  );


  and
  g364
  (
    n332,
    n132,
    n234,
    n130,
    n164
  );


  xor
  g365
  (
    n343,
    n213,
    n214,
    n101,
    n118
  );


  and
  g366
  (
    n315,
    n205,
    n117,
    n232,
    n187
  );


  nand
  g367
  (
    n334,
    n183,
    n96,
    n167,
    n112
  );


  xor
  g368
  (
    n307,
    n160,
    n146,
    n141,
    n132
  );


  xor
  g369
  (
    n393,
    n131,
    n112,
    n128,
    n148
  );


  and
  g370
  (
    n311,
    n246,
    n208,
    n220,
    n172
  );


  nand
  g371
  (
    n406,
    n241,
    n146,
    n101,
    n98
  );


  nor
  g372
  (
    n371,
    n207,
    n170,
    n139,
    n190
  );


  xor
  g373
  (
    n292,
    n225,
    n100,
    n127,
    n173
  );


  and
  g374
  (
    n366,
    n110,
    n156,
    n129,
    n217
  );


  nor
  g375
  (
    n280,
    n189,
    n226,
    n243,
    n168
  );


  or
  g376
  (
    n337,
    n204,
    n161,
    n109,
    n197
  );


  nand
  g377
  (
    n268,
    n146,
    n232,
    n182,
    n169
  );


  or
  g378
  (
    n321,
    n171,
    n218,
    n161,
    n175
  );


  and
  g379
  (
    n330,
    n163,
    n106,
    n210,
    n164
  );


  or
  g380
  (
    n413,
    n205,
    n188,
    n129,
    n153
  );


  or
  g381
  (
    n404,
    n214,
    n123,
    n102,
    n226
  );


  xnor
  g382
  (
    n344,
    n181,
    n150,
    n147,
    n204
  );


  xor
  g383
  (
    n384,
    n159,
    n199,
    n153,
    n160
  );


  xnor
  g384
  (
    n277,
    n197,
    n226,
    n176,
    n103
  );


  and
  g385
  (
    n282,
    n223,
    n246,
    n149,
    n168
  );


  xor
  g386
  (
    n392,
    n192,
    n109,
    n177,
    n101
  );


  or
  g387
  (
    n319,
    n186,
    n159,
    n133,
    n102
  );


  or
  g388
  (
    n357,
    n180,
    n201,
    n148,
    n152
  );


  or
  g389
  (
    n388,
    n105,
    n145,
    n192,
    n104
  );


  xnor
  g390
  (
    n345,
    n166,
    n202,
    n141
  );


  and
  g391
  (
    KeyWire_0_19,
    n214,
    n117,
    n165,
    n162
  );


  and
  g392
  (
    n300,
    n211,
    n184,
    n119,
    n182
  );


  nor
  g393
  (
    n369,
    n154,
    n214,
    n217,
    n179
  );


  xor
  g394
  (
    n298,
    n224,
    n242,
    n245,
    n248
  );


  xnor
  g395
  (
    n286,
    n200,
    n233,
    n154,
    n194
  );


  or
  g396
  (
    n412,
    n102,
    n110,
    n111,
    n156
  );


  or
  g397
  (
    n296,
    n215,
    n97,
    n218,
    n166
  );


  and
  g398
  (
    n278,
    n211,
    n194,
    n184,
    n150
  );


  and
  g399
  (
    n324,
    n115,
    n155,
    n165,
    n146
  );


  nor
  g400
  (
    n305,
    n179,
    n247,
    n242,
    n124
  );


  xnor
  g401
  (
    n387,
    n101,
    n222,
    n218,
    n135
  );


  xnor
  g402
  (
    n353,
    n170,
    n182,
    n98,
    n220
  );


  nor
  g403
  (
    n370,
    n201,
    n163,
    n108,
    n238
  );


  xnor
  g404
  (
    n294,
    n139,
    n147,
    n137,
    n144
  );


  xor
  g405
  (
    n293,
    n162,
    n224,
    n231,
    n102
  );


  xnor
  g406
  (
    n339,
    n122,
    n185,
    n228,
    n219
  );


  nand
  g407
  (
    n338,
    n105,
    n187,
    n136,
    n162
  );


  or
  g408
  (
    n383,
    n209,
    n223,
    n203,
    n198
  );


  or
  g409
  (
    n431,
    n103,
    n133,
    n224,
    n230
  );


  and
  g410
  (
    n403,
    n166,
    n136,
    n125,
    n120
  );


  or
  g411
  (
    n316,
    n100,
    n152,
    n239,
    n117
  );


  and
  g412
  (
    n355,
    n234,
    n237,
    n202,
    n219
  );


  and
  g413
  (
    n430,
    n114,
    n133,
    n198,
    n177
  );


  nor
  g414
  (
    n576,
    n422,
    n277,
    n362,
    n358
  );


  nor
  g415
  (
    n465,
    n303,
    n414,
    n318,
    n270
  );


  nor
  g416
  (
    n533,
    n424,
    n425,
    n415,
    n364
  );


  or
  g417
  (
    n595,
    n336,
    n420,
    n361,
    n365
  );


  nor
  g418
  (
    n475,
    n366,
    n425,
    n303,
    n417
  );


  xnor
  g419
  (
    n457,
    n410,
    n270,
    n407,
    n318
  );


  nor
  g420
  (
    n538,
    n345,
    n301,
    n408
  );


  xnor
  g421
  (
    n524,
    n276,
    n334,
    n320,
    n286
  );


  xnor
  g422
  (
    n478,
    n301,
    n355,
    n348,
    n376
  );


  xnor
  g423
  (
    n547,
    n329,
    n380,
    n333,
    n353
  );


  xnor
  g424
  (
    n572,
    n420,
    n407,
    n311,
    n275
  );


  xor
  g425
  (
    n593,
    n388,
    n284,
    n339,
    n316
  );


  or
  g426
  (
    n550,
    n386,
    n294,
    n344,
    n379
  );


  nor
  g427
  (
    n471,
    n281,
    n300,
    n292,
    n311
  );


  xor
  g428
  (
    n558,
    n287,
    n403,
    n409,
    n380
  );


  xor
  g429
  (
    n539,
    n373,
    n268,
    n311,
    n306
  );


  nor
  g430
  (
    n561,
    n413,
    n344,
    n281,
    n384
  );


  nand
  g431
  (
    KeyWire_0_13,
    n321,
    n375,
    n406,
    n427
  );


  and
  g432
  (
    n563,
    n345,
    n293,
    n404,
    n353
  );


  and
  g433
  (
    n520,
    n271,
    n281,
    n385,
    n374
  );


  xor
  g434
  (
    n540,
    n365,
    n352,
    n393,
    n346
  );


  and
  g435
  (
    n575,
    n413,
    n399,
    n283,
    n341
  );


  xor
  g436
  (
    n489,
    n409,
    n298,
    n421,
    n299
  );


  nand
  g437
  (
    n522,
    n398,
    n402,
    n416,
    n341
  );


  xnor
  g438
  (
    n440,
    n360,
    n290,
    n400,
    n394
  );


  nor
  g439
  (
    n488,
    n282,
    n382,
    n284,
    n394
  );


  and
  g440
  (
    n565,
    n291,
    n347,
    n379,
    n367
  );


  xor
  g441
  (
    n509,
    n418,
    n338,
    n345,
    n323
  );


  xnor
  g442
  (
    n467,
    n358,
    n285,
    n269,
    n385
  );


  xnor
  g443
  (
    n458,
    n298,
    n346,
    n309,
    n423
  );


  nor
  g444
  (
    n573,
    n368,
    n365,
    n327,
    n424
  );


  xor
  g445
  (
    n439,
    n293,
    n343,
    n362,
    n397
  );


  xnor
  g446
  (
    n577,
    n309,
    n337,
    n310,
    n389
  );


  xnor
  g447
  (
    n508,
    n296,
    n285,
    n393,
    n395
  );


  and
  g448
  (
    n555,
    n375,
    n392,
    n272,
    n282
  );


  and
  g449
  (
    n463,
    n392,
    n315,
    n279,
    n383
  );


  xnor
  g450
  (
    KeyWire_0_24,
    n308,
    n361,
    n284,
    n375
  );


  or
  g451
  (
    n579,
    n427,
    n277,
    n426,
    n394
  );


  or
  g452
  (
    n443,
    n297,
    n293,
    n316,
    n429
  );


  xnor
  g453
  (
    n557,
    n294,
    n382,
    n373,
    n333
  );


  nand
  g454
  (
    n446,
    n383,
    n417,
    n324,
    n271
  );


  nor
  g455
  (
    n525,
    n411,
    n348,
    n363,
    n390
  );


  xor
  g456
  (
    n462,
    n399,
    n347,
    n415,
    n328
  );


  nor
  g457
  (
    n476,
    n307,
    n272,
    n395,
    n278
  );


  xnor
  g458
  (
    n474,
    n352,
    n339,
    n283,
    n369
  );


  xor
  g459
  (
    n542,
    n380,
    n392,
    n402,
    n397
  );


  or
  g460
  (
    n571,
    n422,
    n355,
    n325,
    n419
  );


  xnor
  g461
  (
    n590,
    n318,
    n377,
    n287,
    n289
  );


  xnor
  g462
  (
    n583,
    n381,
    n426,
    n291,
    n377
  );


  xnor
  g463
  (
    n527,
    n335,
    n378,
    n391,
    n390
  );


  xor
  g464
  (
    n456,
    n305,
    n416,
    n357,
    n332
  );


  or
  g465
  (
    n518,
    n321,
    n317,
    n272,
    n428
  );


  xnor
  g466
  (
    n480,
    n370,
    n355,
    n308,
    n388
  );


  nor
  g467
  (
    n578,
    n412,
    n404,
    n385,
    n429
  );


  nand
  g468
  (
    n535,
    n328,
    n367,
    n318,
    n301
  );


  nor
  g469
  (
    KeyWire_0_4,
    n268,
    n290,
    n312,
    n428
  );


  or
  g470
  (
    n551,
    n275,
    n331,
    n414,
    n366
  );


  and
  g471
  (
    n447,
    n311,
    n402,
    n338,
    n280
  );


  nand
  g472
  (
    n452,
    n299,
    n426,
    n353,
    n370
  );


  nor
  g473
  (
    n486,
    n368,
    n349,
    n343,
    n361
  );


  and
  g474
  (
    n500,
    n342,
    n330,
    n427,
    n376
  );


  and
  g475
  (
    n506,
    n303,
    n299,
    n379,
    n315
  );


  and
  g476
  (
    n549,
    n405,
    n427,
    n390,
    n314
  );


  or
  g477
  (
    n581,
    n273,
    n332,
    n280,
    n363
  );


  or
  g478
  (
    n530,
    n386,
    n339,
    n324,
    n389
  );


  nand
  g479
  (
    n441,
    n396,
    n319,
    n351,
    n275
  );


  nand
  g480
  (
    n580,
    n340,
    n411,
    n269,
    n335
  );


  or
  g481
  (
    n544,
    n401,
    n373,
    n366,
    n326
  );


  or
  g482
  (
    n587,
    n273,
    n412,
    n337,
    n350
  );


  nor
  g483
  (
    n564,
    n420,
    n360,
    n313,
    n368
  );


  or
  g484
  (
    n507,
    n313,
    n361,
    n345,
    n350
  );


  xor
  g485
  (
    n556,
    n321,
    n425,
    n421,
    n300
  );


  xnor
  g486
  (
    n513,
    n335,
    n383,
    n419,
    n269
  );


  nor
  g487
  (
    n460,
    n327,
    n341,
    n338,
    n404
  );


  xnor
  g488
  (
    n455,
    n428,
    n384,
    n308,
    n406
  );


  xor
  g489
  (
    n503,
    n331,
    n306,
    n363,
    n408
  );


  nand
  g490
  (
    n562,
    n340,
    n346,
    n369,
    n357
  );


  and
  g491
  (
    n588,
    n331,
    n335,
    n408,
    n422
  );


  xnor
  g492
  (
    n519,
    n307,
    n295,
    n390,
    n328
  );


  or
  g493
  (
    n434,
    n377,
    n421,
    n297,
    n417
  );


  xor
  g494
  (
    KeyWire_0_21,
    n288,
    n391,
    n339,
    n409
  );


  nor
  g495
  (
    n537,
    n384,
    n349,
    n269,
    n274
  );


  nand
  g496
  (
    n566,
    n410,
    n278,
    n358,
    n394
  );


  xor
  g497
  (
    n492,
    n397,
    n312,
    n285,
    n314
  );


  xor
  g498
  (
    n499,
    n415,
    n279,
    n291,
    n275
  );


  and
  g499
  (
    n502,
    n403,
    n371,
    n327,
    n360
  );


  xnor
  g500
  (
    n490,
    n349,
    n406,
    n389,
    n398
  );


  xnor
  g501
  (
    n444,
    n316,
    n387,
    n277,
    n337
  );


  or
  g502
  (
    n505,
    n290,
    n322,
    n372,
    n326
  );


  nor
  g503
  (
    n451,
    n306,
    n276,
    n330,
    n305
  );


  nor
  g504
  (
    n495,
    n272,
    n322,
    n355,
    n372
  );


  nand
  g505
  (
    n472,
    n278,
    n369,
    n326,
    n286
  );


  nor
  g506
  (
    n477,
    n386,
    n319,
    n332,
    n424
  );


  and
  g507
  (
    n449,
    n312,
    n297,
    n388,
    n268
  );


  and
  g508
  (
    n560,
    n289,
    n419,
    n399,
    n411
  );


  and
  g509
  (
    n515,
    n270,
    n364,
    n282,
    n276
  );


  xor
  g510
  (
    n438,
    n296,
    n405,
    n313,
    n416
  );


  xor
  g511
  (
    n512,
    n323,
    n294,
    n333,
    n380
  );


  nand
  g512
  (
    n559,
    n391,
    n279,
    n317,
    n413
  );


  and
  g513
  (
    n483,
    n304,
    n348,
    n396,
    n417
  );


  nor
  g514
  (
    n589,
    n292,
    n403,
    n413,
    n388
  );


  nor
  g515
  (
    n568,
    n333,
    n283,
    n342,
    n423
  );


  nor
  g516
  (
    n491,
    n416,
    n396,
    n295,
    n327
  );


  xor
  g517
  (
    n496,
    n378,
    n344,
    n285,
    n325
  );


  nand
  g518
  (
    n459,
    n400,
    n294,
    n348,
    n293
  );


  nand
  g519
  (
    n554,
    n337,
    n295,
    n330,
    n290
  );


  and
  g520
  (
    n482,
    n407,
    n347,
    n381,
    n324
  );


  xnor
  g521
  (
    n454,
    n325,
    n356,
    n378,
    n332
  );


  xor
  g522
  (
    n511,
    n302,
    n429,
    n374,
    n401
  );


  xnor
  g523
  (
    n531,
    n320,
    n287,
    n407,
    n397
  );


  nand
  g524
  (
    n484,
    n279,
    n396,
    n422,
    n315
  );


  xor
  g525
  (
    n567,
    n300,
    n386,
    n304,
    n336
  );


  nor
  g526
  (
    n493,
    n334,
    n313,
    n280,
    n370
  );


  nand
  g527
  (
    KeyWire_0_16,
    n286,
    n382,
    n357,
    n352
  );


  and
  g528
  (
    n570,
    n296,
    n382,
    n360,
    n398
  );


  or
  g529
  (
    n528,
    n377,
    n391,
    n400,
    n302
  );


  and
  g530
  (
    n497,
    n372,
    n326,
    n280,
    n354
  );


  or
  g531
  (
    n469,
    n354,
    n317,
    n289,
    n329
  );


  nor
  g532
  (
    n501,
    n387,
    n393,
    n298,
    n303
  );


  xor
  g533
  (
    n470,
    n395,
    n274,
    n383,
    n304
  );


  or
  g534
  (
    n529,
    n317,
    n297,
    n309,
    n336
  );


  and
  g535
  (
    n494,
    n343,
    n359,
    n367,
    n306
  );


  xnor
  g536
  (
    n514,
    n310,
    n387,
    n357,
    n274
  );


  xor
  g537
  (
    n584,
    n322,
    n369,
    n329,
    n410
  );


  xnor
  g538
  (
    n523,
    n403,
    n420,
    n364,
    n334
  );


  or
  g539
  (
    n453,
    n322,
    n412,
    n271,
    n286
  );


  and
  g540
  (
    n592,
    n319,
    n418,
    n421
  );


  xor
  g541
  (
    n543,
    n271,
    n315,
    n347,
    n373
  );


  xnor
  g542
  (
    n516,
    n412,
    n328,
    n268,
    n342
  );


  and
  g543
  (
    n510,
    n314,
    n395,
    n295,
    n371
  );


  and
  g544
  (
    n481,
    n273,
    n302,
    n405,
    n291
  );


  xor
  g545
  (
    n586,
    n324,
    n385,
    n277,
    n288
  );


  nand
  g546
  (
    n473,
    n281,
    n278,
    n401,
    n352
  );


  xnor
  g547
  (
    n545,
    n350,
    n425,
    n288,
    n375
  );


  and
  g548
  (
    n485,
    n410,
    n371,
    n378,
    n296
  );


  xnor
  g549
  (
    n552,
    n310,
    n288,
    n374,
    n398
  );


  xnor
  g550
  (
    n591,
    n366,
    n359,
    n309,
    n392
  );


  xor
  g551
  (
    n487,
    n340,
    n423,
    n305,
    n304
  );


  nor
  g552
  (
    n532,
    n344,
    n346,
    n405,
    n406
  );


  or
  g553
  (
    n468,
    n325,
    n389,
    n323,
    n273
  );


  and
  g554
  (
    n517,
    n356,
    n354,
    n351,
    n310
  );


  nor
  g555
  (
    n504,
    n323,
    n282,
    n354,
    n356
  );


  nand
  g556
  (
    n445,
    n367,
    n418,
    n287,
    n319
  );


  nand
  g557
  (
    n498,
    n270,
    n409,
    n342,
    n384
  );


  nand
  g558
  (
    n569,
    n340,
    n381,
    n312,
    n374
  );


  or
  g559
  (
    n436,
    n370,
    n320,
    n419,
    n316
  );


  or
  g560
  (
    n582,
    n362,
    n301,
    n302,
    n365
  );


  or
  g561
  (
    n450,
    n298,
    n411,
    n426,
    n364
  );


  nor
  g562
  (
    n526,
    n321,
    n343,
    n401,
    n353
  );


  and
  g563
  (
    n548,
    n307,
    n371,
    n314,
    n349
  );


  xnor
  g564
  (
    n585,
    n379,
    n320,
    n423,
    n387
  );


  and
  g565
  (
    n521,
    n341,
    n331,
    n338,
    n329
  );


  nor
  g566
  (
    n536,
    n283,
    n351,
    n414,
    n358
  );


  or
  g567
  (
    n541,
    n276,
    n402,
    n292
  );


  or
  g568
  (
    n546,
    n376,
    n429,
    n404,
    n305
  );


  xnor
  g569
  (
    n437,
    n274,
    n381,
    n399,
    n300
  );


  xnor
  g570
  (
    n574,
    n362,
    n372,
    n400,
    n284
  );


  xor
  g571
  (
    n448,
    n289,
    n415,
    n330,
    n414
  );


  or
  g572
  (
    n442,
    n307,
    n359,
    n308,
    n368
  );


  xor
  g573
  (
    n594,
    n376,
    n356,
    n299,
    n424
  );


  and
  g574
  (
    n464,
    n393,
    n363,
    n428,
    n350
  );


  or
  g575
  (
    n466,
    n351,
    n334,
    n359,
    n336
  );


  and
  g576
  (
    n601,
    n494,
    n463,
    n516,
    n448
  );


  nor
  g577
  (
    n679,
    n523,
    n492,
    n466,
    n536
  );


  nor
  g578
  (
    n685,
    n251,
    n552,
    n524
  );


  and
  g579
  (
    n618,
    n250,
    n253,
    n470,
    n554
  );


  xor
  g580
  (
    n716,
    n555,
    n538,
    n519,
    n497
  );


  xor
  g581
  (
    n612,
    n454,
    n512,
    n497,
    n467
  );


  xnor
  g582
  (
    n604,
    n476,
    n444,
    n543,
    n549
  );


  and
  g583
  (
    n674,
    n447,
    n534,
    n482,
    n469
  );


  or
  g584
  (
    n724,
    n452,
    n485,
    n498,
    n513
  );


  and
  g585
  (
    n714,
    n499,
    n467,
    n448,
    n436
  );


  xor
  g586
  (
    n683,
    n463,
    n490,
    n545,
    n496
  );


  or
  g587
  (
    n627,
    n550,
    n542,
    n440,
    n494
  );


  nand
  g588
  (
    n639,
    n506,
    n521,
    n450,
    n500
  );


  xor
  g589
  (
    n655,
    n533,
    n531,
    n447,
    n451
  );


  nor
  g590
  (
    n725,
    n457,
    n538,
    n491,
    n509
  );


  and
  g591
  (
    n731,
    n547,
    n477,
    n472,
    n448
  );


  and
  g592
  (
    n718,
    n483,
    n517,
    n455,
    n536
  );


  xor
  g593
  (
    n622,
    n511,
    n526,
    n501,
    n494
  );


  xor
  g594
  (
    n675,
    n253,
    n446,
    n434
  );


  and
  g595
  (
    n607,
    n454,
    n258,
    n435,
    n492
  );


  nor
  g596
  (
    n626,
    n444,
    n517,
    n546,
    n474
  );


  nor
  g597
  (
    n654,
    n503,
    n542,
    n547,
    n513
  );


  and
  g598
  (
    n713,
    n479,
    n449,
    n516,
    n523
  );


  nor
  g599
  (
    n688,
    n441,
    n483,
    n512,
    n487
  );


  xnor
  g600
  (
    n641,
    n260,
    n496,
    n478,
    n537
  );


  or
  g601
  (
    n723,
    n545,
    n550,
    n453,
    n512
  );


  xnor
  g602
  (
    n602,
    n502,
    n257,
    n533,
    n252
  );


  or
  g603
  (
    n599,
    n492,
    n488,
    n472,
    n470
  );


  xnor
  g604
  (
    n705,
    n554,
    n261,
    n478,
    n489
  );


  nand
  g605
  (
    KeyWire_0_7,
    n514,
    n462,
    n471,
    n490
  );


  or
  g606
  (
    n659,
    n552,
    n526,
    n456,
    n458
  );


  nor
  g607
  (
    n667,
    n510,
    n507,
    n474,
    n263
  );


  nor
  g608
  (
    n682,
    n516,
    n440,
    n450,
    n250
  );


  nor
  g609
  (
    n665,
    n544,
    n539,
    n507,
    n452
  );


  or
  g610
  (
    n636,
    n518,
    n445,
    n552,
    n528
  );


  and
  g611
  (
    n696,
    n461,
    n527,
    n530,
    n518
  );


  or
  g612
  (
    n681,
    n257,
    n449,
    n451,
    n551
  );


  or
  g613
  (
    n709,
    n445,
    n455,
    n489,
    n530
  );


  xnor
  g614
  (
    n598,
    n438,
    n477,
    n519,
    n262
  );


  xnor
  g615
  (
    n608,
    n253,
    n473,
    n517,
    n264
  );


  nand
  g616
  (
    n614,
    n499,
    n525,
    n445,
    n444
  );


  nand
  g617
  (
    n643,
    n477,
    n466,
    n459,
    n460
  );


  xor
  g618
  (
    n623,
    n439,
    n265,
    n493,
    n465
  );


  xnor
  g619
  (
    n666,
    n510,
    n522,
    n555,
    n475
  );


  xor
  g620
  (
    n633,
    n511,
    n460,
    n478,
    n456
  );


  nand
  g621
  (
    n669,
    n464,
    n544,
    n546,
    n541
  );


  and
  g622
  (
    n662,
    n457,
    n527,
    n538,
    n543
  );


  or
  g623
  (
    n640,
    n541,
    n484,
    n259,
    n452
  );


  xnor
  g624
  (
    n689,
    n258,
    n520,
    n555,
    n535
  );


  nand
  g625
  (
    n596,
    n525,
    n508,
    n255,
    n465
  );


  nor
  g626
  (
    n663,
    n464,
    n535,
    n531,
    n440
  );


  or
  g627
  (
    n671,
    n480,
    n554,
    n260,
    n502
  );


  xnor
  g628
  (
    KeyWire_0_15,
    n485,
    n488,
    n515,
    n256
  );


  nand
  g629
  (
    n649,
    n515,
    n518,
    n553,
    n264
  );


  or
  g630
  (
    KeyWire_0_26,
    n514,
    n453,
    n450,
    n440
  );


  xnor
  g631
  (
    n605,
    n442,
    n539,
    n259,
    n541
  );


  xnor
  g632
  (
    n656,
    n548,
    n251,
    n464,
    n537
  );


  nand
  g633
  (
    n597,
    n534,
    n434,
    n553,
    n257
  );


  xnor
  g634
  (
    n680,
    n467,
    n513,
    n495,
    n497
  );


  nand
  g635
  (
    n632,
    n439,
    n498,
    n509,
    n260
  );


  xor
  g636
  (
    n697,
    n438,
    n521,
    n499,
    n490
  );


  xor
  g637
  (
    n648,
    n480,
    n546,
    n481,
    n522
  );


  nand
  g638
  (
    n706,
    n436,
    n543,
    n473,
    n437
  );


  nand
  g639
  (
    KeyWire_0_30,
    n509,
    n550,
    n442,
    n265
  );


  nor
  g640
  (
    n646,
    n468,
    n500,
    n540,
    n522
  );


  xor
  g641
  (
    n609,
    n536,
    n526,
    n485,
    n505
  );


  and
  g642
  (
    n645,
    n532,
    n484,
    n489,
    n512
  );


  nor
  g643
  (
    n732,
    n537,
    n448,
    n264,
    n500
  );


  or
  g644
  (
    n712,
    n462,
    n435,
    n548,
    n530
  );


  nand
  g645
  (
    n722,
    n466,
    n262,
    n253,
    n506
  );


  nand
  g646
  (
    n733,
    n265,
    n502,
    n479,
    n547
  );


  nand
  g647
  (
    n701,
    n526,
    n265,
    n550,
    n474
  );


  and
  g648
  (
    n625,
    n459,
    n503,
    n534,
    n264
  );


  nand
  g649
  (
    n700,
    n539,
    n515,
    n554,
    n520
  );


  and
  g650
  (
    n691,
    n484,
    n546,
    n533,
    n528
  );


  nor
  g651
  (
    n631,
    n464,
    n540,
    n491,
    n446
  );


  nand
  g652
  (
    n613,
    n254,
    n436,
    n471,
    n466
  );


  nand
  g653
  (
    n699,
    n443,
    n549,
    n452,
    n538
  );


  nor
  g654
  (
    n684,
    n436,
    n539,
    n474,
    n486
  );


  xor
  g655
  (
    n687,
    n525,
    n483,
    n495,
    n458
  );


  nor
  g656
  (
    n710,
    n505,
    n252,
    n257,
    n519
  );


  and
  g657
  (
    n628,
    n531,
    n261,
    n520,
    n553
  );


  or
  g658
  (
    n698,
    n443,
    n458,
    n486,
    n439
  );


  nor
  g659
  (
    n637,
    n498,
    n496,
    n449,
    n437
  );


  nand
  g660
  (
    n711,
    n258,
    n545,
    n445,
    n514
  );


  or
  g661
  (
    n630,
    n529,
    n497,
    n531,
    n517
  );


  and
  g662
  (
    n606,
    n455,
    n470,
    n439
  );


  xor
  g663
  (
    n670,
    n256,
    n450,
    n460,
    n441
  );


  or
  g664
  (
    n615,
    n548,
    n457,
    n504,
    n500
  );


  and
  g665
  (
    n635,
    n551,
    n459,
    n489,
    n509
  );


  or
  g666
  (
    n728,
    n525,
    n529,
    n472,
    n501
  );


  xnor
  g667
  (
    n603,
    n513,
    n541,
    n442,
    n460
  );


  and
  g668
  (
    n726,
    n481,
    n259,
    n444,
    n488
  );


  and
  g669
  (
    n730,
    n522,
    n480,
    n437,
    n493
  );


  xor
  g670
  (
    n673,
    n508,
    n461,
    n495,
    n469
  );


  nand
  g671
  (
    n727,
    n442,
    n478,
    n521,
    n549
  );


  nand
  g672
  (
    n692,
    n487,
    n529,
    n485,
    n251
  );


  and
  g673
  (
    n600,
    n503,
    n456,
    n468,
    n477
  );


  xor
  g674
  (
    n660,
    n453,
    n551,
    n481,
    n482
  );


  and
  g675
  (
    n638,
    n447,
    n508,
    n530,
    n487
  );


  nor
  g676
  (
    n694,
    n486,
    n462,
    n254,
    n434
  );


  xnor
  g677
  (
    n704,
    n475,
    n535,
    n508,
    n457
  );


  xnor
  g678
  (
    n664,
    n532,
    n528,
    n524,
    n501
  );


  xor
  g679
  (
    n677,
    n449,
    n528,
    n434,
    n441
  );


  nand
  g680
  (
    n657,
    n475,
    n537,
    n551,
    n463
  );


  and
  g681
  (
    n647,
    n454,
    n256,
    n555
  );


  nand
  g682
  (
    n653,
    n499,
    n456,
    n482,
    n263
  );


  and
  g683
  (
    n678,
    n533,
    n543,
    n549,
    n540
  );


  nand
  g684
  (
    n621,
    n471,
    n523,
    n506,
    n475
  );


  xor
  g685
  (
    n715,
    n505,
    n438,
    n521,
    n462
  );


  xnor
  g686
  (
    n644,
    n536,
    n469,
    n473,
    n507
  );


  or
  g687
  (
    n695,
    n435,
    n518,
    n454,
    n535
  );


  xnor
  g688
  (
    n617,
    n453,
    n519,
    n510,
    n259
  );


  nand
  g689
  (
    n661,
    n446,
    n524,
    n502,
    n480
  );


  xnor
  g690
  (
    n721,
    n435,
    n250,
    n491,
    n451
  );


  nor
  g691
  (
    n707,
    n520,
    n472,
    n498,
    n262
  );


  xor
  g692
  (
    n620,
    n534,
    n492,
    n527,
    n547
  );


  nand
  g693
  (
    n717,
    n540,
    n510,
    n254,
    n504
  );


  xnor
  g694
  (
    n619,
    n488,
    n251,
    n458,
    n254
  );


  nand
  g695
  (
    n693,
    n468,
    n255,
    n501,
    n451
  );


  nor
  g696
  (
    n672,
    n465,
    n461,
    n495,
    n514
  );


  xor
  g697
  (
    n720,
    n476,
    n511,
    n490,
    n261
  );


  and
  g698
  (
    n729,
    n491,
    n544,
    n493,
    n479
  );


  xnor
  g699
  (
    n610,
    n441,
    n511,
    n532,
    n266
  );


  or
  g700
  (
    n702,
    n262,
    n252,
    n481,
    n482
  );


  xor
  g701
  (
    n708,
    n542,
    n471,
    n504,
    n486
  );


  and
  g702
  (
    n624,
    n487,
    n553,
    n255,
    n483
  );


  xor
  g703
  (
    n719,
    n494,
    n496,
    n516,
    n515
  );


  and
  g704
  (
    n686,
    n506,
    n548,
    n258,
    n467
  );


  nand
  g705
  (
    KeyWire_0_11,
    n529,
    n255,
    n544,
    n484
  );


  or
  g706
  (
    n651,
    n532,
    n473,
    n505,
    n443
  );


  or
  g707
  (
    KeyWire_0_17,
    n504,
    n260,
    n261,
    n476
  );


  or
  g708
  (
    n658,
    n545,
    n437,
    n542,
    n468
  );


  xor
  g709
  (
    KeyWire_0_3,
    n524,
    n443,
    n438,
    n463
  );


  nor
  g710
  (
    n611,
    n469,
    n461,
    n455,
    n252
  );


  xnor
  g711
  (
    n676,
    n459,
    n493,
    n479,
    n447
  );


  and
  g712
  (
    n652,
    n503,
    n523,
    n465,
    n476
  );


  and
  g713
  (
    n634,
    n527,
    n507,
    n263
  );


  xnor
  g714
  (
    n798,
    n662,
    n672,
    n700,
    n686
  );


  and
  g715
  (
    n792,
    n678,
    n629,
    n728,
    n691
  );


  and
  g716
  (
    n794,
    n721,
    n646,
    n682,
    n601
  );


  nand
  g717
  (
    n748,
    n725,
    n661,
    n675,
    n668
  );


  and
  g718
  (
    n804,
    n668,
    n691,
    n673,
    n704
  );


  or
  g719
  (
    n754,
    n596,
    n714,
    n651,
    n660
  );


  nand
  g720
  (
    n783,
    n699,
    n718,
    n692,
    n717
  );


  nand
  g721
  (
    n764,
    n610,
    n684,
    n677,
    n685
  );


  xor
  g722
  (
    n785,
    n687,
    n702,
    n611,
    n665
  );


  or
  g723
  (
    n745,
    n625,
    n710,
    n679,
    n648
  );


  xnor
  g724
  (
    n807,
    n674,
    n641,
    n722,
    n654
  );


  nand
  g725
  (
    n737,
    n615,
    n665,
    n720,
    n680
  );


  xnor
  g726
  (
    n808,
    n679,
    n707,
    n618
  );


  and
  g727
  (
    n779,
    n609,
    n728,
    n711,
    n689
  );


  nand
  g728
  (
    n744,
    n702,
    n656,
    n627,
    n680
  );


  and
  g729
  (
    n775,
    n667,
    n694,
    n712,
    n662
  );


  nor
  g730
  (
    n801,
    n683,
    n727,
    n695,
    n718
  );


  xor
  g731
  (
    n781,
    n673,
    n698,
    n696,
    n727
  );


  xor
  g732
  (
    n773,
    n675,
    n692,
    n669,
    n724
  );


  xor
  g733
  (
    n816,
    n717,
    n721,
    n709
  );


  and
  g734
  (
    n740,
    n701,
    n706,
    n693,
    n717
  );


  nor
  g735
  (
    n802,
    n597,
    n681,
    n686,
    n703
  );


  nor
  g736
  (
    n819,
    n704,
    n660,
    n666
  );


  xor
  g737
  (
    n810,
    n681,
    n679,
    n690,
    n613
  );


  or
  g738
  (
    n789,
    n673,
    n685,
    n672,
    n689
  );


  nand
  g739
  (
    n780,
    n695,
    n713,
    n644,
    n701
  );


  or
  g740
  (
    n753,
    n669,
    n685,
    n642,
    n632
  );


  or
  g741
  (
    n734,
    n688,
    n686,
    n718,
    n638
  );


  nand
  g742
  (
    n788,
    n712,
    n680,
    n726,
    n619
  );


  and
  g743
  (
    n760,
    n702,
    n669,
    n728,
    n633
  );


  xor
  g744
  (
    n736,
    n672,
    n682,
    n649,
    n657
  );


  and
  g745
  (
    n813,
    n713,
    n647,
    n703,
    n696
  );


  nor
  g746
  (
    n741,
    n681,
    n698,
    n715
  );


  xnor
  g747
  (
    n782,
    n715,
    n688,
    n700,
    n723
  );


  nor
  g748
  (
    n809,
    n674,
    n684,
    n640,
    n706
  );


  nand
  g749
  (
    n750,
    n668,
    n684,
    n626,
    n710
  );


  nand
  g750
  (
    n784,
    n722,
    n661,
    n721,
    n694
  );


  xor
  g751
  (
    n817,
    n673,
    n714,
    n667,
    n704
  );


  xor
  g752
  (
    n815,
    n691,
    n678,
    n705,
    n695
  );


  and
  g753
  (
    n790,
    n708,
    n703,
    n678,
    n612
  );


  nand
  g754
  (
    n738,
    n635,
    n724,
    n723,
    n670
  );


  nor
  g755
  (
    n756,
    n700,
    n614,
    n726,
    n716
  );


  xnor
  g756
  (
    n755,
    n693,
    n726,
    n668,
    n712
  );


  xnor
  g757
  (
    KeyWire_0_9,
    n664,
    n643,
    n674,
    n620
  );


  xor
  g758
  (
    n742,
    n616,
    n621,
    n671,
    n692
  );


  and
  g759
  (
    n803,
    n624,
    n698,
    n697,
    n713
  );


  and
  g760
  (
    n757,
    n645,
    n608,
    n684,
    n697
  );


  xor
  g761
  (
    n766,
    n725,
    n711,
    n672,
    n659
  );


  xor
  g762
  (
    n747,
    n652,
    n690,
    n699,
    n727
  );


  nand
  g763
  (
    n818,
    n690,
    n693,
    n698,
    n605
  );


  nor
  g764
  (
    n746,
    n665,
    n688,
    n660,
    n679
  );


  nor
  g765
  (
    n735,
    n676,
    n722,
    n670,
    n660
  );


  xor
  g766
  (
    n771,
    n705,
    n696,
    n694,
    n691
  );


  nand
  g767
  (
    n805,
    n726,
    n695,
    n617,
    n653
  );


  or
  g768
  (
    n772,
    n699,
    n715,
    n659,
    n687
  );


  xnor
  g769
  (
    n791,
    n696,
    n655,
    n603,
    n606
  );


  nor
  g770
  (
    n765,
    n703,
    n664,
    n689,
    n708
  );


  or
  g771
  (
    n770,
    n663,
    n711,
    n688,
    n713
  );


  nand
  g772
  (
    n774,
    n682,
    n710,
    n675,
    n725
  );


  xnor
  g773
  (
    n806,
    n711,
    n663,
    n639,
    n705
  );


  nor
  g774
  (
    n811,
    n663,
    n669,
    n607,
    n727
  );


  nand
  g775
  (
    n797,
    n720,
    n721,
    n709,
    n604
  );


  xor
  g776
  (
    n749,
    n630,
    n694,
    n677,
    n701
  );


  and
  g777
  (
    n767,
    n600,
    n671,
    n661,
    n722
  );


  xor
  g778
  (
    n768,
    n723,
    n701,
    n712,
    n702
  );


  or
  g779
  (
    n752,
    n677,
    n700,
    n634,
    n716
  );


  nor
  g780
  (
    n795,
    n705,
    n675,
    n658,
    n719
  );


  or
  g781
  (
    n787,
    n678,
    n683,
    n724,
    n697
  );


  and
  g782
  (
    n800,
    n670,
    n687,
    n637,
    n693
  );


  and
  g783
  (
    n761,
    n631,
    n706,
    n671,
    n659
  );


  or
  g784
  (
    n758,
    n685,
    n725,
    n724,
    n699
  );


  xor
  g785
  (
    n763,
    n663,
    n662,
    n686,
    n665
  );


  xnor
  g786
  (
    n762,
    n661,
    n666,
    n720,
    n708
  );


  or
  g787
  (
    n793,
    n683,
    n674,
    n666,
    n704
  );


  xnor
  g788
  (
    n786,
    n670,
    n659,
    n719,
    n729
  );


  nor
  g789
  (
    n777,
    n690,
    n598,
    n716,
    n602
  );


  and
  g790
  (
    n776,
    n623,
    n680,
    n714,
    n697
  );


  xnor
  g791
  (
    n759,
    n664,
    n599,
    n667,
    n719
  );


  nand
  g792
  (
    n778,
    n728,
    n662,
    n714,
    n671
  );


  nor
  g793
  (
    n769,
    n664,
    n717,
    n636,
    n692
  );


  nor
  g794
  (
    KeyWire_0_22,
    n650,
    n719,
    n622,
    n682
  );


  xor
  g795
  (
    n814,
    n628,
    n667,
    n676
  );


  and
  g796
  (
    n739,
    n681,
    n709,
    n706,
    n683
  );


  nor
  g797
  (
    KeyWire_0_31,
    n687,
    n718,
    n716,
    n707
  );


  or
  g798
  (
    n751,
    n707,
    n720,
    n689,
    n723
  );


  xor
  g799
  (
    n812,
    n676,
    n677,
    n708,
    n710
  );


  xnor
  g800
  (
    n833,
    n576,
    n565,
    n587,
    n585
  );


  or
  g801
  (
    n862,
    n769,
    n764,
    n577,
    n578
  );


  or
  g802
  (
    n837,
    n765,
    n581,
    n558
  );


  and
  g803
  (
    n839,
    n577,
    n766,
    n566,
    n561
  );


  nand
  g804
  (
    n831,
    n574,
    n739,
    n563,
    n583
  );


  nand
  g805
  (
    n843,
    n570,
    n557,
    n585
  );


  or
  g806
  (
    n847,
    n569,
    n775,
    n571,
    n586
  );


  or
  g807
  (
    n822,
    n574,
    n737,
    n563,
    n745
  );


  xor
  g808
  (
    n851,
    n585,
    n560,
    n580
  );


  and
  g809
  (
    n844,
    n565,
    n577,
    n560,
    n744
  );


  or
  g810
  (
    n854,
    n582,
    n581,
    n572,
    n557
  );


  nand
  g811
  (
    n857,
    n758,
    n558,
    n559,
    n586
  );


  nand
  g812
  (
    n859,
    n743,
    n556,
    n563,
    n742
  );


  and
  g813
  (
    n836,
    n556,
    n741,
    n562,
    n559
  );


  and
  g814
  (
    n855,
    n576,
    n572,
    n568,
    n573
  );


  and
  g815
  (
    n841,
    n564,
    n750,
    n558,
    n580
  );


  or
  g816
  (
    n845,
    n586,
    n578,
    n559,
    n579
  );


  or
  g817
  (
    KeyWire_0_8,
    n574,
    n760,
    n576,
    n756
  );


  xnor
  g818
  (
    n827,
    n583,
    n568,
    n746,
    n574
  );


  nand
  g819
  (
    n856,
    n754,
    n573,
    n562,
    n749
  );


  or
  g820
  (
    n840,
    n573,
    n587,
    n562,
    n565
  );


  and
  g821
  (
    n821,
    n556,
    n582,
    n560,
    n575
  );


  nor
  g822
  (
    n858,
    n736,
    n571,
    n759,
    n569
  );


  or
  g823
  (
    n846,
    n584,
    n578,
    n580
  );


  and
  g824
  (
    n832,
    n757,
    n738,
    n579,
    n564
  );


  nor
  g825
  (
    n825,
    n569,
    n740,
    n572,
    n570
  );


  or
  g826
  (
    n826,
    n570,
    n768,
    n564,
    n561
  );


  and
  g827
  (
    n834,
    n556,
    n587,
    n565,
    n751
  );


  xnor
  g828
  (
    n860,
    n761,
    n563,
    n579,
    n567
  );


  nand
  g829
  (
    n829,
    n776,
    n747,
    n575,
    n564
  );


  nor
  g830
  (
    n842,
    n559,
    n562,
    n770,
    n558
  );


  or
  g831
  (
    n835,
    n753,
    n584,
    n582,
    n570
  );


  xor
  g832
  (
    n849,
    n583,
    n571,
    n734,
    n584
  );


  xnor
  g833
  (
    n828,
    n572,
    n581,
    n585,
    n767
  );


  or
  g834
  (
    KeyWire_0_5,
    n566,
    n748,
    n774,
    n569
  );


  and
  g835
  (
    n861,
    n763,
    n762,
    n561,
    n582
  );


  or
  g836
  (
    n830,
    n566,
    n561,
    n573,
    n576
  );


  nand
  g837
  (
    n820,
    n567,
    n571,
    n584,
    n735
  );


  xnor
  g838
  (
    n823,
    n579,
    n575,
    n752,
    n560
  );


  nand
  g839
  (
    n838,
    n772,
    n567,
    n587,
    n588
  );


  nor
  g840
  (
    n850,
    n566,
    n586,
    n568,
    n557
  );


  nor
  g841
  (
    n824,
    n577,
    n755,
    n773,
    n568
  );


  nand
  g842
  (
    n848,
    n771,
    n575,
    n567,
    n583
  );


  buf
  g843
  (
    n863,
    n730
  );


  buf
  g844
  (
    n867,
    n839
  );


  xnor
  g845
  (
    n866,
    n838,
    n730
  );


  nand
  g846
  (
    n865,
    n840,
    n837,
    n729
  );


  and
  g847
  (
    n864,
    n729,
    n841,
    n731
  );


  buf
  g848
  (
    n871,
    n867
  );


  buf
  g849
  (
    n876,
    n781
  );


  buf
  g850
  (
    n882,
    n864
  );


  buf
  g851
  (
    n875,
    n866
  );


  not
  g852
  (
    n877,
    n865
  );


  buf
  g853
  (
    n870,
    n863
  );


  not
  g854
  (
    n868,
    n779
  );


  not
  g855
  (
    n869,
    n777
  );


  not
  g856
  (
    n883,
    n865
  );


  not
  g857
  (
    n878,
    n866
  );


  buf
  g858
  (
    n880,
    n782
  );


  xnor
  g859
  (
    n879,
    n866,
    n867
  );


  or
  g860
  (
    n873,
    n782,
    n781,
    n778
  );


  nor
  g861
  (
    n872,
    n866,
    n865,
    n780
  );


  or
  g862
  (
    n881,
    n865,
    n781,
    n864
  );


  xnor
  g863
  (
    n874,
    n867,
    n781,
    n863
  );


  nor
  g864
  (
    n887,
    n807,
    n808,
    n874,
    n879
  );


  or
  g865
  (
    n906,
    n815,
    n813,
    n872,
    n818
  );


  xor
  g866
  (
    n897,
    n807,
    n868,
    n794
  );


  and
  g867
  (
    n931,
    n802,
    n805,
    n879,
    n784
  );


  xor
  g868
  (
    n938,
    n872,
    n788,
    n876,
    n871
  );


  nor
  g869
  (
    n902,
    n870,
    n804,
    n791
  );


  xor
  g870
  (
    n940,
    n875,
    n790,
    n796,
    n793
  );


  or
  g871
  (
    n933,
    n880,
    n810,
    n882,
    n878
  );


  xnor
  g872
  (
    n904,
    n430,
    n875,
    n801,
    n812
  );


  or
  g873
  (
    n919,
    n819,
    n798,
    n870,
    n809
  );


  and
  g874
  (
    n942,
    n795,
    n783,
    n800,
    n818
  );


  or
  g875
  (
    n939,
    n791,
    n799,
    n812,
    n804
  );


  and
  g876
  (
    n895,
    n854,
    n813,
    n882,
    n850
  );


  nand
  g877
  (
    n899,
    n877,
    n800,
    n801,
    n818
  );


  nor
  g878
  (
    KeyWire_0_23,
    n784,
    n805,
    n806,
    n816
  );


  xor
  g879
  (
    n889,
    n787,
    n844,
    n883,
    n873
  );


  xnor
  g880
  (
    n893,
    n813,
    n859,
    n785,
    n811
  );


  xnor
  g881
  (
    n921,
    n797,
    n788,
    n816,
    n807
  );


  nand
  g882
  (
    n929,
    n792,
    n879,
    n872,
    n789
  );


  xnor
  g883
  (
    n913,
    n869,
    n783,
    n862,
    n786
  );


  xnor
  g884
  (
    n937,
    n795,
    n785,
    n798,
    n816
  );


  nand
  g885
  (
    n886,
    n791,
    n843,
    n812,
    n814
  );


  or
  g886
  (
    n898,
    n811,
    n787,
    n799,
    n870
  );


  xor
  g887
  (
    n935,
    n817,
    n797,
    n782,
    n798
  );


  nand
  g888
  (
    n918,
    n874,
    n788,
    n845,
    n784
  );


  xnor
  g889
  (
    n920,
    n803,
    n852,
    n876,
    n883
  );


  nand
  g890
  (
    n892,
    n794,
    n873,
    n795,
    n868
  );


  xor
  g891
  (
    n888,
    n787,
    n797,
    n871,
    n796
  );


  and
  g892
  (
    n924,
    n815,
    n875,
    n810,
    n883
  );


  xnor
  g893
  (
    n884,
    n811,
    n797,
    n851,
    n860
  );


  nor
  g894
  (
    n903,
    n806,
    n794,
    n883,
    n881
  );


  xnor
  g895
  (
    n915,
    n789,
    n877,
    n812,
    n809
  );


  nand
  g896
  (
    n896,
    n873,
    n804,
    n792,
    n786
  );


  xor
  g897
  (
    n928,
    n800,
    n861,
    n791,
    n785
  );


  or
  g898
  (
    n936,
    n882,
    n782,
    n847,
    n880
  );


  and
  g899
  (
    n930,
    n813,
    n799,
    n809,
    n869
  );


  xnor
  g900
  (
    n900,
    n787,
    n878,
    n881,
    n815
  );


  xnor
  g901
  (
    n901,
    n876,
    n800,
    n877,
    n814
  );


  xnor
  g902
  (
    n941,
    n783,
    n789,
    n806,
    n871
  );


  and
  g903
  (
    n914,
    n855,
    n817,
    n868,
    n858
  );


  nand
  g904
  (
    n917,
    n793,
    n842,
    n816,
    n790
  );


  or
  g905
  (
    n908,
    n806,
    n793,
    n879,
    n784
  );


  xnor
  g906
  (
    n922,
    n882,
    n805,
    n876,
    n874
  );


  and
  g907
  (
    n912,
    n803,
    n788,
    n807,
    n805
  );


  nor
  g908
  (
    n885,
    n880,
    n814,
    n802
  );


  xor
  g909
  (
    n909,
    n869,
    n808,
    n870,
    n798
  );


  xnor
  g910
  (
    n894,
    n817,
    n881,
    n878,
    n811
  );


  and
  g911
  (
    n907,
    n786,
    n801,
    n796,
    n789
  );


  xnor
  g912
  (
    n927,
    n849,
    n795,
    n793,
    n869
  );


  or
  g913
  (
    n891,
    n792,
    n803,
    n848,
    n808
  );


  or
  g914
  (
    n934,
    n796,
    n819,
    n873,
    n874
  );


  nor
  g915
  (
    n905,
    n803,
    n799,
    n786,
    n846
  );


  nor
  g916
  (
    n925,
    n878,
    n810,
    n815,
    n875
  );


  nor
  g917
  (
    n932,
    n794,
    n802,
    n783,
    n817
  );


  xor
  g918
  (
    n910,
    n809,
    n856,
    n801,
    n880
  );


  or
  g919
  (
    n911,
    n790,
    n792,
    n785,
    n818
  );


  xnor
  g920
  (
    n926,
    n810,
    n819,
    n857
  );


  nand
  g921
  (
    n916,
    n881,
    n853,
    n790,
    n808
  );


  nand
  g922
  (
    n923,
    n802,
    n877,
    n872,
    n871
  );


  and
  g923
  (
    n943,
    n905,
    n903,
    n267,
    n900
  );


  nand
  g924
  (
    n959,
    n895,
    n933,
    n898,
    n588
  );


  and
  g925
  (
    n962,
    n929,
    n915,
    n936,
    n920
  );


  xor
  g926
  (
    n958,
    n913,
    n890,
    n930,
    n906
  );


  nand
  g927
  (
    n973,
    n918,
    n931,
    n934,
    n940
  );


  and
  g928
  (
    n968,
    n913,
    n910,
    n591,
    n888
  );


  nand
  g929
  (
    n947,
    n892,
    n939,
    n902
  );


  nor
  g930
  (
    n974,
    n884,
    n589,
    n942,
    n901
  );


  xor
  g931
  (
    n965,
    n916,
    n906,
    n589,
    n918
  );


  nand
  g932
  (
    n948,
    n939,
    n893,
    n908,
    n923
  );


  xnor
  g933
  (
    n944,
    n926,
    n900,
    n940,
    n898
  );


  nor
  g934
  (
    n954,
    n911,
    n266,
    n932,
    n904
  );


  xor
  g935
  (
    n976,
    n927,
    n938,
    n590,
    n935
  );


  nor
  g936
  (
    n964,
    n922,
    n927,
    n940,
    n939
  );


  or
  g937
  (
    n953,
    n589,
    n917,
    n590,
    n588
  );


  or
  g938
  (
    n952,
    n931,
    n910,
    n923,
    n921
  );


  xor
  g939
  (
    n951,
    n936,
    n589,
    n592,
    n938
  );


  or
  g940
  (
    n961,
    n909,
    n267,
    n935,
    n926
  );


  and
  g941
  (
    n975,
    n267,
    n887,
    n907,
    n912
  );


  xnor
  g942
  (
    n967,
    n920,
    n908,
    n889,
    n924
  );


  xnor
  g943
  (
    n950,
    n937,
    n588,
    n904,
    n915
  );


  nor
  g944
  (
    n955,
    n886,
    n590,
    n896,
    n924
  );


  nand
  g945
  (
    n966,
    n903,
    n899,
    n941,
    n266
  );


  xor
  g946
  (
    n969,
    n592,
    n896,
    n919,
    n591
  );


  or
  g947
  (
    n970,
    n921,
    n897,
    n912,
    n942
  );


  and
  g948
  (
    n956,
    n899,
    n909,
    n914,
    n941
  );


  nand
  g949
  (
    n946,
    n266,
    n940,
    n917,
    n934
  );


  or
  g950
  (
    n949,
    n919,
    n905,
    n928,
    n938
  );


  xor
  g951
  (
    n977,
    n941,
    n894,
    n901,
    n938
  );


  nand
  g952
  (
    n963,
    n897,
    n591,
    n925,
    n907
  );


  xor
  g953
  (
    n972,
    n922,
    n885,
    n925,
    n916
  );


  xor
  g954
  (
    n945,
    n930,
    n902,
    n929,
    n942
  );


  nand
  g955
  (
    n960,
    n267,
    n891,
    n911,
    n941
  );


  xor
  g956
  (
    n971,
    n590,
    n933,
    n932,
    n591
  );


  and
  g957
  (
    n957,
    n937,
    n928,
    n942,
    n914
  );


  not
  g958
  (
    n988,
    n971
  );


  not
  g959
  (
    n982,
    n957
  );


  not
  g960
  (
    n987,
    n964
  );


  xnor
  g961
  (
    KeyWire_0_2,
    n974,
    n959,
    n960
  );


  xor
  g962
  (
    n985,
    n947,
    n953,
    n955,
    n975
  );


  and
  g963
  (
    n981,
    n968,
    n430,
    n944,
    n946
  );


  and
  g964
  (
    n980,
    n969,
    n954,
    n952,
    n966
  );


  nand
  g965
  (
    n979,
    n956,
    n961,
    n972,
    n948
  );


  nand
  g966
  (
    n984,
    n943,
    n951,
    n963,
    n958
  );


  xor
  g967
  (
    n983,
    n965,
    n973,
    n950,
    n967
  );


  and
  g968
  (
    n986,
    n949,
    n945,
    n970,
    n962
  );


  nor
  g969
  (
    n990,
    n980,
    n980,
    n979,
    n982
  );


  xnor
  g970
  (
    n993,
    n981,
    n979,
    n980,
    n592
  );


  xnor
  g971
  (
    KeyWire_0_29,
    n978,
    n979,
    n982
  );


  or
  g972
  (
    n992,
    n982,
    n978,
    n981
  );


  nand
  g973
  (
    n989,
    n592,
    n979,
    n980,
    n981
  );


  xor
  g974
  (
    n995,
    n732,
    n976,
    n733
  );


  and
  g975
  (
    n997,
    n989,
    n731,
    n732
  );


  or
  g976
  (
    KeyWire_0_27,
    n732,
    n733,
    n992
  );


  and
  g977
  (
    n994,
    n977,
    n732,
    n991,
    n990
  );


  xor
  g978
  (
    n999,
    n997,
    n996,
    n984
  );


  nor
  g979
  (
    n1000,
    n984,
    n983,
    n985
  );


  xor
  g980
  (
    n998,
    n983,
    n983,
    n995,
    n984
  );


  and
  g981
  (
    n1006,
    n431,
    n986
  );


  and
  g982
  (
    n1009,
    n988,
    n985,
    n1000,
    n432
  );


  nor
  g983
  (
    n1011,
    n993,
    n988,
    n985,
    n986
  );


  nor
  g984
  (
    KeyWire_0_14,
    n986,
    n999,
    n432,
    n430
  );


  nand
  g985
  (
    n1004,
    n433,
    n1000,
    n431,
    n998
  );


  nand
  g986
  (
    n1001,
    n433,
    n1000,
    n999,
    n987
  );


  nor
  g987
  (
    n1005,
    n1000,
    n987,
    n431,
    n432
  );


  nor
  g988
  (
    n1008,
    n999,
    n985,
    n987,
    n432
  );


  xor
  g989
  (
    n1003,
    n988,
    n431,
    n993,
    n433
  );


  xnor
  g990
  (
    n1007,
    n430,
    n998,
    n999,
    n433
  );


  xnor
  g991
  (
    n1010,
    n988,
    n998,
    n987
  );


  xnor
  g992
  (
    n1015,
    n594,
    n1010,
    n593
  );


  nand
  g993
  (
    n1014,
    n593,
    n594,
    n595
  );


  nor
  g994
  (
    n1013,
    n594,
    n1011,
    n595,
    n593
  );


  or
  g995
  (
    n1012,
    n1009,
    n1008,
    n595
  );


  xnor
  KeyGate_0_0
  (
    n174,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n187,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n978,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n616,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n553,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n853,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n85,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n690,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n852,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n743,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n164,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n703,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n28,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n435,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1002,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n629,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n479,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n668,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n81,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n354,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n225,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n461,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n799,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n890,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n534,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n103,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n650,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n996,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n291,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n991,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n642,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n796,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

