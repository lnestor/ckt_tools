// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_305 written by SynthGen on 2021/04/05 11:24:14
module Stat_3000_305( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1538, n2983, n2981, n2989, n2980, n2986, n2985, n2988,
 n2982, n2984, n3019, n3026, n3013, n3032, n3020, n3018,
 n3022, n3015, n3027, n3017, n3012, n3024, n3021, n3016,
 n3029, n3011, n3025, n3014, n3028, n3023, n3031, n3030);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1538, n2983, n2981, n2989, n2980, n2986, n2985, n2988,
 n2982, n2984, n3019, n3026, n3013, n3032, n3020, n3018,
 n3022, n3015, n3027, n3017, n3012, n3024, n3021, n3016,
 n3029, n3011, n3025, n3014, n3028, n3023, n3031, n3030;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
 n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
 n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
 n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
 n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
 n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
 n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
 n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
 n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
 n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
 n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
 n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
 n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
 n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
 n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
 n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
 n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
 n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
 n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
 n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
 n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
 n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
 n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
 n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
 n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
 n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
 n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
 n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
 n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
 n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
 n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
 n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
 n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
 n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
 n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
 n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
 n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
 n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
 n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
 n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
 n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
 n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
 n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
 n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
 n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
 n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
 n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
 n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
 n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
 n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
 n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
 n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
 n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
 n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
 n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
 n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
 n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
 n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
 n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
 n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
 n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
 n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
 n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
 n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
 n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
 n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
 n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
 n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
 n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
 n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
 n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
 n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
 n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
 n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
 n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
 n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
 n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
 n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
 n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
 n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
 n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
 n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
 n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
 n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
 n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
 n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
 n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
 n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
 n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
 n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
 n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
 n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
 n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
 n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
 n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
 n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
 n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
 n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
 n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
 n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
 n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
 n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
 n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
 n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
 n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
 n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
 n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
 n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
 n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
 n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
 n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
 n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
 n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
 n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
 n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
 n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
 n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
 n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
 n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
 n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
 n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
 n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
 n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
 n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
 n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
 n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
 n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
 n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
 n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
 n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
 n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
 n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
 n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
 n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
 n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
 n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
 n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
 n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
 n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
 n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
 n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
 n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
 n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
 n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
 n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
 n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
 n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
 n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
 n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
 n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
 n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
 n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
 n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
 n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
 n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
 n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
 n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
 n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
 n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
 n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
 n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
 n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
 n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
 n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
 n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
 n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
 n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
 n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
 n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
 n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
 n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
 n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
 n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
 n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
 n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
 n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
 n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
 n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
 n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
 n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
 n2978, n2979, n2987, n2990, n2991, n2992, n2993, n2994,
 n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
 n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010;

buf  g0 (n74, n13);
not  g1 (n56, n8);
not  g2 (n52, n1);
not  g3 (n55, n2);
not  g4 (n79, n1);
buf  g5 (n92, n7);
buf  g6 (n82, n17);
buf  g7 (n36, n3);
buf  g8 (n85, n2);
buf  g9 (n95, n13);
not  g10 (n46, n10);
not  g11 (n66, n3);
buf  g12 (n65, n16);
not  g13 (n96, n15);
not  g14 (n60, n16);
not  g15 (n70, n10);
not  g16 (n86, n7);
buf  g17 (n48, n17);
buf  g18 (n83, n12);
buf  g19 (n64, n13);
not  g20 (n37, n1);
buf  g21 (n59, n10);
not  g22 (n87, n2);
not  g23 (n51, n3);
buf  g24 (n54, n4);
buf  g25 (n98, n13);
not  g26 (n97, n6);
buf  g27 (n80, n14);
buf  g28 (n40, n2);
not  g29 (n71, n11);
buf  g30 (n76, n5);
buf  g31 (n49, n3);
buf  g32 (n63, n7);
buf  g33 (n43, n6);
buf  g34 (n90, n12);
not  g35 (n39, n5);
buf  g36 (n45, n14);
buf  g37 (n69, n8);
not  g38 (n75, n6);
not  g39 (n73, n9);
not  g40 (n34, n4);
not  g41 (n38, n12);
not  g42 (n77, n16);
buf  g43 (n47, n16);
buf  g44 (n57, n9);
buf  g45 (n41, n9);
not  g46 (n33, n4);
not  g47 (n78, n14);
buf  g48 (n67, n4);
buf  g49 (n62, n14);
not  g50 (n91, n5);
buf  g51 (n58, n8);
not  g52 (n35, n12);
buf  g53 (n61, n10);
buf  g54 (n42, n11);
buf  g55 (n84, n15);
not  g56 (n72, n7);
buf  g57 (n94, n5);
buf  g58 (n81, n15);
buf  g59 (n89, n8);
not  g60 (n68, n11);
not  g61 (n50, n6);
buf  g62 (n44, n15);
not  g63 (n53, n1);
not  g64 (n88, n9);
not  g65 (n93, n11);
not  g66 (n172, n44);
not  g67 (n275, n48);
buf  g68 (n244, n60);
buf  g69 (n139, n33);
not  g70 (n138, n75);
not  g71 (n196, n64);
buf  g72 (n214, n67);
buf  g73 (n204, n49);
not  g74 (n140, n34);
not  g75 (n248, n77);
not  g76 (n199, n47);
not  g77 (n239, n45);
not  g78 (n185, n74);
buf  g79 (n187, n71);
buf  g80 (n141, n55);
not  g81 (n205, n74);
not  g82 (n175, n53);
buf  g83 (n206, n72);
buf  g84 (n266, n76);
buf  g85 (n112, n46);
buf  g86 (n170, n61);
buf  g87 (n146, n47);
buf  g88 (n237, n55);
buf  g89 (n260, n63);
not  g90 (n166, n36);
buf  g91 (n182, n37);
not  g92 (n270, n50);
not  g93 (n156, n36);
buf  g94 (n122, n39);
buf  g95 (n202, n41);
not  g96 (n251, n63);
buf  g97 (n176, n69);
buf  g98 (n255, n38);
buf  g99 (n119, n65);
buf  g100 (n236, n52);
not  g101 (n179, n63);
not  g102 (n133, n78);
buf  g103 (n144, n60);
not  g104 (n128, n45);
buf  g105 (n274, n47);
buf  g106 (n190, n73);
buf  g107 (n269, n34);
buf  g108 (n117, n77);
not  g109 (n136, n73);
not  g110 (n225, n70);
not  g111 (n167, n43);
not  g112 (n178, n61);
not  g113 (n118, n38);
buf  g114 (n265, n71);
buf  g115 (n183, n68);
buf  g116 (n177, n42);
not  g117 (n189, n76);
buf  g118 (n252, n65);
buf  g119 (n249, n33);
not  g120 (n180, n66);
buf  g121 (n173, n51);
not  g122 (n123, n75);
not  g123 (n147, n37);
buf  g124 (n273, n54);
not  g125 (n134, n43);
buf  g126 (n235, n58);
buf  g127 (n191, n36);
not  g128 (n253, n69);
not  g129 (n192, n45);
buf  g130 (n105, n77);
not  g131 (n127, n65);
not  g132 (n151, n39);
not  g133 (n233, n50);
not  g134 (n109, n42);
buf  g135 (n110, n48);
buf  g136 (n230, n51);
buf  g137 (n115, n78);
buf  g138 (n247, n70);
buf  g139 (n242, n46);
not  g140 (n164, n52);
buf  g141 (n238, n33);
not  g142 (n174, n36);
not  g143 (n203, n38);
not  g144 (n113, n52);
buf  g145 (n246, n58);
not  g146 (n223, n38);
not  g147 (n227, n63);
not  g148 (n121, n70);
not  g149 (n142, n74);
not  g150 (n220, n62);
buf  g151 (n217, n56);
not  g152 (n152, n76);
not  g153 (n163, n37);
buf  g154 (n207, n68);
not  g155 (n259, n46);
buf  g156 (n268, n71);
not  g157 (n278, n35);
not  g158 (n150, n53);
not  g159 (n194, n45);
buf  g160 (n120, n76);
not  g161 (n267, n66);
buf  g162 (n261, n75);
not  g163 (n102, n41);
not  g164 (n100, n35);
not  g165 (n201, n46);
buf  g166 (n271, n72);
not  g167 (n245, n71);
not  g168 (n221, n48);
buf  g169 (n155, n54);
buf  g170 (n148, n68);
not  g171 (n211, n62);
buf  g172 (n103, n39);
buf  g173 (n243, n42);
buf  g174 (n209, n67);
buf  g175 (n130, n73);
not  g176 (n162, n54);
buf  g177 (n272, n35);
not  g178 (n250, n47);
not  g179 (n226, n66);
not  g180 (n215, n58);
not  g181 (n108, n41);
buf  g182 (n143, n59);
not  g183 (n281, n64);
buf  g184 (n213, n69);
buf  g185 (n137, n34);
buf  g186 (n101, n57);
buf  g187 (n193, n64);
not  g188 (n234, n34);
not  g189 (n208, n59);
buf  g190 (n228, n57);
buf  g191 (n241, n78);
not  g192 (n184, n42);
not  g193 (n212, n43);
not  g194 (n124, n74);
not  g195 (n181, n62);
buf  g196 (n104, n64);
not  g197 (n231, n48);
not  g198 (n129, n59);
buf  g199 (n279, n37);
not  g200 (n111, n54);
not  g201 (n264, n51);
not  g202 (n145, n50);
not  g203 (n126, n73);
buf  g204 (n276, n70);
buf  g205 (n216, n57);
not  g206 (n280, n69);
buf  g207 (n149, n41);
buf  g208 (n263, n52);
not  g209 (n218, n44);
not  g210 (n200, n58);
buf  g211 (n107, n60);
buf  g212 (n169, n56);
buf  g213 (n198, n43);
buf  g214 (n116, n77);
not  g215 (n186, n33);
not  g216 (n258, n57);
not  g217 (n114, n44);
buf  g218 (n229, n68);
not  g219 (n240, n40);
not  g220 (n224, n39);
not  g221 (n135, n50);
buf  g222 (n153, n40);
not  g223 (n106, n72);
not  g224 (n262, n40);
not  g225 (n171, n56);
buf  g226 (n232, n53);
buf  g227 (n159, n59);
buf  g228 (n277, n35);
buf  g229 (n188, n72);
buf  g230 (n254, n44);
buf  g231 (n158, n75);
not  g232 (n131, n66);
not  g233 (n195, n65);
buf  g234 (n168, n60);
buf  g235 (n125, n40);
not  g236 (n99, n51);
buf  g237 (n210, n55);
not  g238 (n165, n49);
buf  g239 (n197, n62);
not  g240 (n222, n55);
not  g241 (n256, n49);
buf  g242 (n161, n53);
not  g243 (n160, n56);
not  g244 (n157, n61);
buf  g245 (n154, n67);
not  g246 (n219, n61);
not  g247 (n132, n67);
not  g248 (n257, n49);
not  g249 (n851, n164);
not  g250 (n798, n107);
not  g251 (n536, n204);
not  g252 (n677, n142);
buf  g253 (n881, n137);
buf  g254 (n746, n101);
buf  g255 (n491, n184);
not  g256 (n443, n200);
buf  g257 (n825, n223);
not  g258 (n291, n126);
buf  g259 (n815, n207);
not  g260 (n880, n208);
not  g261 (n644, n178);
buf  g262 (n841, n173);
buf  g263 (n460, n237);
not  g264 (n831, n119);
not  g265 (n296, n162);
buf  g266 (n767, n238);
not  g267 (n415, n207);
buf  g268 (n540, n170);
buf  g269 (n305, n203);
not  g270 (n956, n255);
not  g271 (n959, n120);
buf  g272 (n449, n148);
buf  g273 (n522, n138);
buf  g274 (n393, n174);
not  g275 (n555, n179);
buf  g276 (n696, n145);
not  g277 (n930, n214);
not  g278 (n572, n105);
not  g279 (n423, n130);
buf  g280 (n576, n248);
not  g281 (n725, n187);
not  g282 (n863, n175);
buf  g283 (n949, n240);
not  g284 (n721, n239);
buf  g285 (n727, n216);
buf  g286 (n285, n138);
not  g287 (n699, n100);
not  g288 (n665, n176);
not  g289 (n331, n218);
buf  g290 (n704, n131);
not  g291 (n861, n227);
not  g292 (n361, n181);
not  g293 (n712, n255);
buf  g294 (n913, n231);
buf  g295 (n312, n177);
buf  g296 (n821, n249);
buf  g297 (n806, n106);
not  g298 (n934, n197);
buf  g299 (n364, n232);
buf  g300 (n655, n263);
not  g301 (n669, n110);
buf  g302 (n664, n102);
buf  g303 (n474, n250);
buf  g304 (n805, n123);
not  g305 (n390, n135);
buf  g306 (n611, n165);
not  g307 (n420, n260);
not  g308 (n589, n163);
not  g309 (n952, n135);
buf  g310 (n330, n163);
buf  g311 (n634, n253);
buf  g312 (n919, n158);
buf  g313 (n747, n216);
not  g314 (n594, n243);
not  g315 (n631, n154);
buf  g316 (n528, n106);
not  g317 (n609, n137);
not  g318 (n450, n186);
not  g319 (n297, n219);
not  g320 (n355, n250);
buf  g321 (n288, n225);
buf  g322 (n958, n165);
buf  g323 (n516, n175);
buf  g324 (n541, n102);
buf  g325 (n463, n185);
buf  g326 (n652, n118);
not  g327 (n781, n264);
buf  g328 (n858, n178);
buf  g329 (n695, n166);
buf  g330 (n636, n160);
not  g331 (n846, n256);
buf  g332 (n398, n242);
buf  g333 (n283, n238);
buf  g334 (n549, n235);
buf  g335 (n809, n252);
not  g336 (n627, n151);
buf  g337 (n584, n263);
buf  g338 (n345, n152);
not  g339 (n910, n203);
buf  g340 (n748, n133);
not  g341 (n726, n196);
not  g342 (n843, n124);
not  g343 (n466, n167);
not  g344 (n356, n150);
not  g345 (n803, n148);
not  g346 (n388, n121);
buf  g347 (n744, n260);
not  g348 (n922, n142);
not  g349 (n828, n233);
buf  g350 (n383, n221);
buf  g351 (n945, n150);
buf  g352 (n392, n173);
buf  g353 (n898, n144);
not  g354 (n893, n142);
not  g355 (n412, n144);
not  g356 (n947, n250);
not  g357 (n710, n210);
not  g358 (n943, n253);
not  g359 (n944, n207);
not  g360 (n292, n209);
not  g361 (n562, n99);
not  g362 (n658, n146);
not  g363 (n765, n262);
buf  g364 (n926, n145);
not  g365 (n857, n132);
buf  g366 (n351, n199);
not  g367 (n845, n254);
not  g368 (n328, n241);
not  g369 (n534, n147);
not  g370 (n564, n146);
buf  g371 (n946, n194);
buf  g372 (n810, n101);
not  g373 (n539, n130);
not  g374 (n569, n120);
buf  g375 (n357, n179);
not  g376 (n754, n175);
buf  g377 (n801, n253);
not  g378 (n384, n251);
buf  g379 (n618, n140);
not  g380 (n724, n208);
not  g381 (n509, n164);
buf  g382 (n406, n243);
buf  g383 (n366, n247);
buf  g384 (n577, n161);
not  g385 (n855, n259);
buf  g386 (n619, n166);
buf  g387 (n788, n190);
not  g388 (n447, n139);
not  g389 (n394, n187);
not  g390 (n313, n157);
buf  g391 (n344, n128);
buf  g392 (n306, n115);
not  g393 (n827, n99);
not  g394 (n349, n170);
not  g395 (n775, n100);
buf  g396 (n853, n202);
buf  g397 (n340, n135);
buf  g398 (n322, n125);
not  g399 (n593, n152);
not  g400 (n896, n213);
not  g401 (n751, n161);
not  g402 (n914, n231);
buf  g403 (n650, n174);
buf  g404 (n335, n182);
buf  g405 (n923, n113);
not  g406 (n703, n265);
buf  g407 (n583, n226);
buf  g408 (n647, n232);
not  g409 (n396, n177);
not  g410 (n755, n226);
not  g411 (n282, n217);
not  g412 (n284, n116);
not  g413 (n342, n259);
buf  g414 (n370, n190);
not  g415 (n502, n176);
not  g416 (n659, n201);
buf  g417 (n505, n248);
buf  g418 (n918, n214);
not  g419 (n615, n200);
buf  g420 (n854, n252);
buf  g421 (n741, n262);
buf  g422 (n503, n199);
not  g423 (n738, n121);
not  g424 (n362, n105);
buf  g425 (n425, n256);
not  g426 (n911, n212);
buf  g427 (n929, n227);
not  g428 (n433, n223);
not  g429 (n544, n228);
buf  g430 (n360, n217);
not  g431 (n909, n163);
not  g432 (n777, n102);
buf  g433 (n641, n149);
not  g434 (n599, n157);
not  g435 (n849, n137);
not  g436 (n739, n248);
buf  g437 (n906, n242);
not  g438 (n728, n188);
buf  g439 (n617, n103);
not  g440 (n596, n205);
buf  g441 (n445, n107);
buf  g442 (n733, n194);
buf  g443 (n882, n118);
not  g444 (n640, n249);
not  g445 (n796, n246);
buf  g446 (n490, n249);
buf  g447 (n471, n123);
not  g448 (n878, n216);
not  g449 (n797, n157);
not  g450 (n686, n108);
not  g451 (n737, n149);
buf  g452 (n614, n197);
not  g453 (n424, n214);
not  g454 (n916, n225);
not  g455 (n713, n126);
not  g456 (n921, n206);
not  g457 (n558, n104);
buf  g458 (n729, n265);
not  g459 (n604, n127);
buf  g460 (n864, n244);
not  g461 (n711, n168);
buf  g462 (n592, n206);
buf  g463 (n512, n178);
buf  g464 (n761, n105);
not  g465 (n568, n111);
not  g466 (n338, n169);
buf  g467 (n648, n200);
not  g468 (n465, n147);
buf  g469 (n308, n126);
not  g470 (n417, n264);
buf  g471 (n680, n136);
not  g472 (n481, n248);
not  g473 (n295, n144);
buf  g474 (n377, n172);
not  g475 (n674, n140);
buf  g476 (n920, n268);
not  g477 (n372, n211);
buf  g478 (n877, n158);
not  g479 (n553, n178);
buf  g480 (n839, n244);
not  g481 (n936, n132);
not  g482 (n753, n205);
not  g483 (n286, n117);
not  g484 (n673, n158);
buf  g485 (n879, n167);
not  g486 (n298, n268);
buf  g487 (n687, n241);
not  g488 (n832, n115);
buf  g489 (n942, n128);
not  g490 (n698, n159);
buf  g491 (n875, n144);
not  g492 (n459, n226);
buf  g493 (n679, n108);
buf  g494 (n381, n268);
not  g495 (n787, n245);
buf  g496 (n758, n217);
buf  g497 (n626, n215);
not  g498 (n535, n259);
not  g499 (n409, n242);
buf  g500 (n657, n258);
buf  g501 (n666, n233);
buf  g502 (n578, n191);
buf  g503 (n817, n133);
buf  g504 (n427, n142);
buf  g505 (n354, n154);
buf  g506 (n760, n103);
buf  g507 (n551, n235);
buf  g508 (n435, n247);
not  g509 (n925, n136);
buf  g510 (n519, n174);
not  g511 (n421, n146);
buf  g512 (n337, n180);
not  g513 (n570, n172);
not  g514 (n763, n205);
buf  g515 (n780, n173);
not  g516 (n649, n130);
not  g517 (n363, n215);
not  g518 (n499, n154);
buf  g519 (n823, n184);
not  g520 (n902, n217);
not  g521 (n319, n112);
not  g522 (n542, n202);
not  g523 (n772, n160);
buf  g524 (n957, n129);
buf  g525 (n579, n229);
buf  g526 (n822, n168);
buf  g527 (n932, n247);
not  g528 (n660, n193);
buf  g529 (n489, n106);
not  g530 (n903, n102);
buf  g531 (n715, n236);
buf  g532 (n327, n254);
not  g533 (n667, n181);
buf  g534 (n613, n183);
buf  g535 (n847, n103);
not  g536 (n299, n147);
buf  g537 (n938, n261);
buf  g538 (n560, n235);
not  g539 (n386, n183);
buf  g540 (n812, n169);
buf  g541 (n718, n186);
not  g542 (n336, n182);
buf  g543 (n480, n114);
buf  g544 (n301, n175);
not  g545 (n819, n212);
buf  g546 (n820, n195);
buf  g547 (n454, n198);
buf  g548 (n643, n241);
buf  g549 (n402, n107);
buf  g550 (n961, n215);
buf  g551 (n411, n156);
not  g552 (n483, n187);
buf  g553 (n353, n141);
not  g554 (n482, n143);
buf  g555 (n374, n189);
buf  g556 (n321, n187);
not  g557 (n689, n148);
not  g558 (n743, n171);
buf  g559 (n380, n199);
not  g560 (n639, n199);
buf  g561 (n397, n149);
not  g562 (n468, n239);
buf  g563 (n529, n192);
not  g564 (n448, n197);
buf  g565 (n808, n208);
not  g566 (n456, n229);
buf  g567 (n838, n134);
not  g568 (n317, n254);
not  g569 (n559, n143);
buf  g570 (n789, n218);
not  g571 (n430, n161);
not  g572 (n418, n246);
not  g573 (n874, n214);
not  g574 (n759, n132);
buf  g575 (n314, n140);
buf  g576 (n813, n128);
buf  g577 (n811, n127);
not  g578 (n757, n237);
buf  g579 (n690, n234);
buf  g580 (n414, n211);
buf  g581 (n464, n166);
not  g582 (n734, n250);
buf  g583 (n642, n151);
buf  g584 (n469, n227);
not  g585 (n325, n222);
buf  g586 (n706, n236);
buf  g587 (n586, n252);
buf  g588 (n300, n111);
not  g589 (n403, n182);
buf  g590 (n735, n246);
not  g591 (n511, n186);
not  g592 (n622, n244);
not  g593 (n740, n202);
not  g594 (n520, n136);
buf  g595 (n745, n258);
buf  g596 (n441, n129);
not  g597 (n561, n239);
not  g598 (n782, n123);
not  g599 (n645, n117);
not  g600 (n473, n172);
buf  g601 (n897, n267);
buf  g602 (n694, n205);
buf  g603 (n341, n222);
buf  g604 (n701, n218);
buf  g605 (n506, n161);
not  g606 (n510, n213);
buf  g607 (n707, n193);
not  g608 (n543, n186);
buf  g609 (n307, n195);
buf  g610 (n426, n172);
not  g611 (n367, n154);
not  g612 (n554, n204);
not  g613 (n462, n231);
buf  g614 (n868, n156);
not  g615 (n401, n109);
not  g616 (n799, n174);
buf  g617 (n479, n198);
buf  g618 (n610, n245);
buf  g619 (n895, n254);
buf  g620 (n369, n155);
not  g621 (n742, n147);
not  g622 (n530, n165);
not  g623 (n478, n156);
buf  g624 (n873, n107);
buf  g625 (n883, n150);
buf  g626 (n311, n251);
buf  g627 (n507, n188);
buf  g628 (n616, n169);
not  g629 (n612, n234);
not  g630 (n867, n141);
buf  g631 (n457, n213);
not  g632 (n783, n134);
buf  g633 (n395, n256);
not  g634 (n623, n166);
not  g635 (n842, n219);
buf  g636 (n684, n188);
buf  g637 (n598, n244);
buf  g638 (n807, n110);
buf  g639 (n571, n264);
not  g640 (n485, n140);
buf  g641 (n630, n245);
not  g642 (n440, n201);
not  g643 (n635, n221);
buf  g644 (n702, n104);
not  g645 (n859, n208);
not  g646 (n316, n153);
not  g647 (n872, n218);
buf  g648 (n527, n141);
not  g649 (n494, n101);
not  g650 (n590, n139);
buf  g651 (n442, n111);
buf  g652 (n359, n192);
not  g653 (n347, n230);
not  g654 (n829, n157);
not  g655 (n912, n249);
not  g656 (n683, n266);
buf  g657 (n682, n176);
buf  g658 (n416, n143);
not  g659 (n840, n151);
not  g660 (n455, n130);
not  g661 (n472, n225);
not  g662 (n470, n189);
not  g663 (n632, n203);
not  g664 (n352, n257);
buf  g665 (n885, n204);
not  g666 (n939, n238);
buf  g667 (n672, n266);
not  g668 (n904, n189);
not  g669 (n884, n104);
not  g670 (n488, n209);
buf  g671 (n582, n128);
buf  g672 (n324, n201);
buf  g673 (n575, n264);
not  g674 (n818, n183);
buf  g675 (n770, n112);
buf  g676 (n326, n159);
not  g677 (n792, n265);
not  g678 (n567, n262);
not  g679 (n786, n223);
buf  g680 (n638, n184);
not  g681 (n907, n100);
buf  g682 (n670, n190);
not  g683 (n302, n192);
not  g684 (n439, n230);
buf  g685 (n931, n118);
buf  g686 (n685, n253);
not  g687 (n368, n153);
not  g688 (n581, n194);
buf  g689 (n793, n197);
buf  g690 (n869, n262);
not  g691 (n515, n220);
buf  g692 (n557, n221);
not  g693 (n804, n160);
buf  g694 (n941, n139);
buf  g695 (n764, n260);
not  g696 (n940, n222);
buf  g697 (n310, n133);
not  g698 (n496, n256);
buf  g699 (n816, n258);
not  g700 (n476, n233);
buf  g701 (n732, n185);
buf  g702 (n436, n206);
buf  g703 (n661, n149);
not  g704 (n376, n124);
buf  g705 (n607, n236);
buf  g706 (n837, n101);
not  g707 (n891, n226);
buf  g708 (n834, n242);
buf  g709 (n960, n203);
buf  g710 (n814, n234);
not  g711 (n538, n160);
buf  g712 (n752, n171);
not  g713 (n563, n237);
buf  g714 (n924, n243);
not  g715 (n784, n230);
not  g716 (n526, n131);
not  g717 (n651, n195);
buf  g718 (n730, n169);
buf  g719 (n768, n117);
not  g720 (n603, n252);
not  g721 (n444, n105);
buf  g722 (n332, n191);
buf  g723 (n315, n127);
buf  g724 (n866, n119);
not  g725 (n320, n236);
buf  g726 (n550, n180);
buf  g727 (n573, n261);
buf  g728 (n547, n162);
buf  g729 (n856, n228);
not  g730 (n766, n193);
not  g731 (n446, n230);
not  g732 (n387, n200);
not  g733 (n654, n131);
not  g734 (n408, n145);
buf  g735 (n844, n198);
not  g736 (n717, n167);
buf  g737 (n373, n126);
buf  g738 (n574, n221);
buf  g739 (n750, n224);
not  g740 (n776, n152);
not  g741 (n705, n122);
not  g742 (n605, n210);
buf  g743 (n375, n116);
buf  g744 (n871, n246);
not  g745 (n899, n158);
buf  g746 (n693, n257);
buf  g747 (n517, n251);
buf  g748 (n365, n191);
buf  g749 (n431, n258);
buf  g750 (n467, n193);
not  g751 (n865, n133);
buf  g752 (n722, n117);
not  g753 (n429, n150);
buf  g754 (n399, n159);
buf  g755 (n692, n148);
not  g756 (n495, n211);
not  g757 (n438, n247);
buf  g758 (n954, n109);
buf  g759 (n587, n112);
buf  g760 (n769, n119);
buf  g761 (n346, n240);
buf  g762 (n836, n177);
buf  g763 (n452, n224);
buf  g764 (n537, n121);
buf  g765 (n802, n104);
buf  g766 (n791, n103);
buf  g767 (n477, n257);
not  g768 (n566, n155);
buf  g769 (n458, n196);
buf  g770 (n546, n198);
not  g771 (n716, n227);
buf  g772 (n329, n204);
buf  g773 (n422, n216);
not  g774 (n620, n220);
buf  g775 (n790, n261);
not  g776 (n628, n116);
not  g777 (n862, n196);
buf  g778 (n714, n191);
buf  g779 (n876, n113);
not  g780 (n900, n263);
not  g781 (n432, n241);
buf  g782 (n545, n164);
not  g783 (n889, n145);
not  g784 (n595, n125);
buf  g785 (n531, n225);
not  g786 (n892, n163);
buf  g787 (n826, n109);
not  g788 (n294, n219);
buf  g789 (n585, n210);
buf  g790 (n629, n106);
not  g791 (n933, n189);
not  g792 (n548, n115);
not  g793 (n498, n156);
not  g794 (n400, n112);
buf  g795 (n835, n220);
not  g796 (n608, n170);
not  g797 (n289, n215);
buf  g798 (n407, n267);
not  g799 (n688, n232);
not  g800 (n475, n229);
not  g801 (n624, n125);
not  g802 (n580, n129);
not  g803 (n334, n164);
not  g804 (n637, n232);
buf  g805 (n795, n108);
buf  g806 (n908, n211);
buf  g807 (n556, n136);
buf  g808 (n833, n195);
buf  g809 (n600, n132);
not  g810 (n830, n155);
buf  g811 (n656, n113);
not  g812 (n762, n179);
buf  g813 (n385, n182);
not  g814 (n453, n100);
buf  g815 (n410, n229);
not  g816 (n736, n176);
not  g817 (n333, n114);
not  g818 (n662, n228);
not  g819 (n779, n259);
not  g820 (n513, n124);
buf  g821 (n287, n235);
buf  g822 (n532, n180);
not  g823 (n708, n238);
not  g824 (n824, n194);
not  g825 (n887, n138);
not  g826 (n497, n231);
not  g827 (n437, n240);
not  g828 (n675, n113);
buf  g829 (n773, n121);
not  g830 (n565, n224);
not  g831 (n723, n129);
buf  g832 (n493, n152);
not  g833 (n697, n228);
not  g834 (n886, n170);
not  g835 (n653, n131);
not  g836 (n428, n181);
buf  g837 (n621, n179);
not  g838 (n800, n138);
not  g839 (n434, n224);
not  g840 (n348, n108);
buf  g841 (n293, n266);
not  g842 (n749, n141);
buf  g843 (n518, n135);
not  g844 (n358, n168);
buf  g845 (n785, n257);
not  g846 (n860, n122);
buf  g847 (n552, n114);
not  g848 (n484, n122);
buf  g849 (n591, n151);
buf  g850 (n486, n209);
not  g851 (n413, n155);
not  g852 (n720, n109);
not  g853 (n508, n124);
buf  g854 (n523, n118);
not  g855 (n848, n99);
buf  g856 (n774, n219);
buf  g857 (n597, n223);
buf  g858 (n378, n139);
buf  g859 (n382, n237);
buf  g860 (n905, n99);
buf  g861 (n935, n266);
not  g862 (n888, n213);
not  g863 (n678, n180);
not  g864 (n951, n212);
buf  g865 (n700, n267);
buf  g866 (n343, n120);
buf  g867 (n461, n122);
buf  g868 (n756, n255);
not  g869 (n487, n159);
buf  g870 (n709, n162);
not  g871 (n524, n134);
buf  g872 (n691, n206);
not  g873 (n318, n123);
not  g874 (n719, n167);
buf  g875 (n339, n201);
buf  g876 (n602, n125);
not  g877 (n500, n261);
buf  g878 (n501, n267);
buf  g879 (n633, n268);
buf  g880 (n955, n165);
not  g881 (n304, n234);
buf  g882 (n405, n134);
buf  g883 (n950, n220);
buf  g884 (n915, n177);
buf  g885 (n371, n190);
buf  g886 (n379, n185);
not  g887 (n668, n260);
not  g888 (n525, n114);
buf  g889 (n601, n240);
buf  g890 (n533, n153);
not  g891 (n350, n110);
buf  g892 (n937, n239);
buf  g893 (n917, n162);
buf  g894 (n389, n181);
not  g895 (n521, n127);
not  g896 (n492, n184);
not  g897 (n778, n222);
not  g898 (n681, n110);
not  g899 (n504, n183);
buf  g900 (n391, n196);
not  g901 (n309, n146);
not  g902 (n928, n116);
buf  g903 (n303, n171);
not  g904 (n870, n137);
not  g905 (n514, n120);
buf  g906 (n290, n251);
not  g907 (n588, n115);
not  g908 (n890, n255);
buf  g909 (n850, n168);
not  g910 (n323, n111);
not  g911 (n771, n265);
buf  g912 (n663, n207);
buf  g913 (n927, n119);
buf  g914 (n451, n210);
not  g915 (n953, n192);
not  g916 (n901, n263);
not  g917 (n404, n245);
buf  g918 (n794, n212);
not  g919 (n852, n153);
buf  g920 (n894, n143);
buf  g921 (n625, n185);
buf  g922 (n948, n171);
buf  g923 (n671, n243);
not  g924 (n606, n233);
not  g925 (n676, n188);
not  g926 (n646, n202);
not  g927 (n419, n209);
not  g928 (n731, n173);
xnor g929 (n1052, n791, n793, n792, n432);
xnor g930 (n1241, n331, n828, n461, n579);
xor  g931 (n975, n901, n397, n825, n730);
nand g932 (n1267, n746, n327, n924, n323);
or   g933 (n993, n758, n894, n936, n875);
nor  g934 (n1323, n695, n342, n626, n913);
and  g935 (n990, n472, n895, n707, n911);
and  g936 (n1132, n479, n317, n846, n935);
xnor g937 (n1125, n672, n724, n919, n584);
nor  g938 (n1047, n916, n463, n471, n943);
and  g939 (n1246, n802, n741, n695, n591);
nor  g940 (n1135, n897, n763, n853, n911);
or   g941 (n1143, n877, n818, n382, n808);
xnor g942 (n983, n865, n577, n784, n765);
nor  g943 (n1328, n357, n734, n779, n856);
and  g944 (n1302, n941, n343, n711, n908);
or   g945 (n1096, n467, n878, n812, n893);
or   g946 (n1128, n745, n598, n942, n685);
nand g947 (n1129, n326, n418, n557, n908);
or   g948 (n1330, n858, n283, n771, n820);
xnor g949 (n1153, n482, n572, n541, n699);
and  g950 (n1083, n516, n606, n402, n387);
and  g951 (n1119, n440, n766, n459, n840);
nand g952 (n1259, n467, n813, n389, n344);
and  g953 (n1090, n688, n892, n633, n391);
xnor g954 (n1173, n582, n405, n855, n625);
xor  g955 (n1053, n934, n929, n719, n485);
xnor g956 (n985, n513, n901, n407, n898);
and  g957 (n1284, n514, n806, n887, n392);
xnor g958 (n1195, n656, n603, n943, n925);
xnor g959 (n1237, n892, n933, n514, n828);
nor  g960 (n1326, n503, n589, n418, n308);
nor  g961 (n1170, n372, n833, n653, n603);
nand g962 (n1198, n740, n400, n838, n886);
xnor g963 (n1130, n317, n721, n383, n345);
xnor g964 (n1319, n596, n369, n673, n493);
xnor g965 (n1234, n350, n687, n359, n473);
xnor g966 (n963, n913, n748, n507, n298);
or   g967 (n966, n848, n301, n484, n727);
or   g968 (n968, n878, n947, n509, n302);
xnor g969 (n1276, n940, n666, n368, n702);
xor  g970 (n1278, n346, n656, n515, n904);
xor  g971 (n1308, n503, n399, n365, n919);
and  g972 (n1050, n755, n639, n526, n558);
and  g973 (n1268, n940, n768, n915, n735);
and  g974 (n1254, n930, n677, n652, n636);
xnor g975 (n1188, n783, n611, n825, n502);
xnor g976 (n1157, n699, n832, n751, n932);
and  g977 (n1131, n856, n419, n642, n664);
nand g978 (n1318, n294, n906, n829, n632);
and  g979 (n1035, n445, n443, n413, n714);
xor  g980 (n1257, n573, n920, n415, n702);
xor  g981 (n1235, n316, n333, n399, n332);
xor  g982 (n1048, n737, n456, n653, n460);
nand g983 (n1098, n874, n466, n551, n906);
or   g984 (n1008, n640, n852, n923, n760);
xor  g985 (n1043, n615, n704, n804, n926);
xor  g986 (n1317, n380, n629, n532, n396);
nor  g987 (n1097, n906, n686, n403, n290);
and  g988 (n1179, n482, n608, n321, n668);
xnor g989 (n987, n663, n618, n512, n710);
and  g990 (n1189, n383, n464, n705, n886);
xor  g991 (n1113, n761, n554, n469, n487);
xor  g992 (n1309, n388, n291, n858, n701);
nor  g993 (n1068, n847, n738, n506, n854);
nand g994 (n1277, n942, n841, n934, n463);
nor  g995 (n1306, n620, n434, n876, n379);
and  g996 (n1218, n569, n867, n406, n470);
and  g997 (n1071, n422, n904, n564, n842);
nand g998 (n1212, n893, n849, n426, n674);
and  g999 (n1169, n824, n877, n841, n917);
nor  g1000 (n1226, n813, n769, n511, n632);
or   g1001 (n1031, n911, n922, n935, n421);
and  g1002 (n1185, n946, n629, n574, n690);
and  g1003 (n1066, n822, n914, n519, n559);
nor  g1004 (n1209, n348, n700, n854, n926);
xnor g1005 (n1229, n901, n910, n410, n387);
and  g1006 (n1332, n707, n788, n661, n453);
nand g1007 (n1089, n769, n293, n394, n592);
nor  g1008 (n1099, n742, n344, n759, n377);
xnor g1009 (n1194, n433, n912, n924, n933);
and  g1010 (n965, n698, n891, n823, n648);
xnor g1011 (n1263, n771, n351, n663, n808);
or   g1012 (n1206, n430, n926, n568, n680);
nor  g1013 (n1281, n893, n805, n307, n874);
or   g1014 (n1296, n749, n594, n869, n907);
or   g1015 (n1011, n447, n930, n845, n875);
xor  g1016 (n1165, n554, n921, n339, n403);
or   g1017 (n1149, n581, n341, n907, n883);
xor  g1018 (n1145, n733, n936, n730, n433);
or   g1019 (n972, n728, n376, n325, n303);
xor  g1020 (n1019, n920, n648, n543, n923);
xor  g1021 (n973, n853, n367, n406, n366);
xor  g1022 (n1168, n349, n907, n558, n539);
xor  g1023 (n1134, n944, n782, n835, n912);
nand g1024 (n1193, n660, n807, n889, n703);
and  g1025 (n1091, n819, n505, n453, n634);
nand g1026 (n1018, n347, n932, n490, n676);
or   g1027 (n1010, n884, n805, n659, n547);
xnor g1028 (n967, n583, n551, n913, n521);
xor  g1029 (n1270, n887, n465, n798, n462);
and  g1030 (n1126, n502, n476, n946, n927);
xor  g1031 (n1067, n376, n786, n824, n292);
xnor g1032 (n1311, n939, n290, n927, n649);
xor  g1033 (n1219, n549, n938, n322, n839);
and  g1034 (n1022, n915, n510, n809, n429);
xnor g1035 (n1070, n869, n362, n896, n488);
nor  g1036 (n1014, n799, n356, n526, n887);
nor  g1037 (n1073, n651, n299, n597, n712);
xor  g1038 (n1217, n720, n422, n739, n889);
and  g1039 (n1211, n303, n844, n607, n309);
and  g1040 (n1002, n899, n829, n888, n325);
and  g1041 (n1294, n716, n935, n790, n696);
and  g1042 (n1264, n581, n507, n834, n555);
xnor g1043 (n964, n661, n739, n896, n615);
or   g1044 (n1285, n937, n938, n452, n857);
xnor g1045 (n1140, n548, n747, n600, n449);
and  g1046 (n1141, n416, n870, n884, n887);
and  g1047 (n1147, n381, n620, n334, n420);
nand g1048 (n1148, n647, n322, n448, n614);
xor  g1049 (n1144, n340, n677, n878, n882);
and  g1050 (n986, n518, n566, n890, n571);
or   g1051 (n1292, n836, n381, n886, n590);
nor  g1052 (n978, n300, n535, n922, n773);
or   g1053 (n1085, n587, n691, n608, n349);
and  g1054 (n1321, n872, n338, n457, n818);
xnor g1055 (n1046, n757, n832, n791, n684);
or   g1056 (n1075, n304, n394, n880, n756);
nor  g1057 (n1327, n427, n560, n764, n901);
nand g1058 (n1081, n888, n793, n670, n881);
and  g1059 (n1286, n446, n770, n500, n426);
or   g1060 (n1084, n857, n546, n943, n754);
nand g1061 (n1183, n937, n566, n800, n814);
nor  g1062 (n1177, n944, n908, n869, n922);
or   g1063 (n1271, n401, n836, n811, n543);
nand g1064 (n1005, n594, n391, n649, n537);
and  g1065 (n1182, n936, n643, n909, n517);
xor  g1066 (n1248, n882, n302, n741, n917);
nor  g1067 (n1155, n652, n900, n843, n395);
xnor g1068 (n1110, n714, n816, n918, n930);
or   g1069 (n1095, n569, n419, n497, n540);
and  g1070 (n1315, n870, n922, n413, n794);
and  g1071 (n1262, n619, n464, n868, n664);
or   g1072 (n1100, n390, n844, n693, n885);
nand g1073 (n1162, n942, n535, n438, n301);
nor  g1074 (n1175, n339, n328, n885, n903);
xnor g1075 (n1205, n866, n720, n564, n616);
xor  g1076 (n1251, n428, n533, n732, n436);
nand g1077 (n1334, n506, n444, n921, n319);
nor  g1078 (n1051, n855, n318, n667, n492);
xor  g1079 (n1108, n536, n811, n884, n890);
or   g1080 (n1054, n420, n903, n585, n284);
xor  g1081 (n1304, n495, n446, n777, n670);
nor  g1082 (n1045, n423, n635, n774, n488);
and  g1083 (n1214, n560, n571, n417, n723);
nor  g1084 (n1142, n897, n368, n561, n874);
or   g1085 (n1191, n886, n683, n402, n788);
and  g1086 (n1106, n941, n912, n938, n404);
or   g1087 (n998, n545, n852, n925, n645);
nor  g1088 (n1015, n414, n424, n873, n489);
nand g1089 (n1065, n498, n477, n550, n519);
or   g1090 (n1289, n431, n712, n528, n792);
xor  g1091 (n1228, n545, n644, n817, n487);
xnor g1092 (n1138, n665, n523, n425, n331);
nor  g1093 (n1210, n647, n917, n916, n679);
or   g1094 (n979, n579, n530, n354, n480);
nand g1095 (n1017, n946, n787, n342, n561);
xnor g1096 (n962, n917, n745, n537, n782);
nand g1097 (n1024, n444, n588, n622, n496);
xnor g1098 (n1056, n891, n622, n845, n689);
nor  g1099 (n1030, n304, n449, n364, n341);
and  g1100 (n1290, n731, n565, n905, n732);
or   g1101 (n1034, n481, n333, n868, n915);
and  g1102 (n1023, n610, n327, n797, n762);
nor  g1103 (n988, n599, n531, n296, n686);
nor  g1104 (n1280, n758, n640, n870, n826);
nand g1105 (n1049, n688, n931, n678, n725);
and  g1106 (n1080, n491, n578, n708, n434);
xor  g1107 (n991, n362, n534, n754, n542);
nor  g1108 (n1061, n763, n822, n837, n892);
xnor g1109 (n971, n582, n697, n624, n494);
xnor g1110 (n1305, n334, n515, n628, n494);
and  g1111 (n1094, n382, n455, n466, n616);
and  g1112 (n996, n925, n862, n430, n803);
and  g1113 (n1310, n945, n477, n892, n736);
nand g1114 (n1301, n873, n484, n459, n722);
nand g1115 (n1320, n617, n796, n881, n934);
nand g1116 (n994, n796, n363, n777, n923);
or   g1117 (n1322, n842, n861, n612, n838);
xnor g1118 (n1295, n693, n929, n447, n520);
xnor g1119 (n1006, n914, n921, n289, n475);
nor  g1120 (n1167, n440, n312, n690, n789);
nand g1121 (n1037, n809, n562, n940, n883);
xor  g1122 (n1112, n784, n912, n438, n872);
and  g1123 (n995, n933, n723, n814, n356);
or   g1124 (n1032, n641, n867, n348, n744);
nor  g1125 (n1044, n860, n637, n575, n884);
xnor g1126 (n1057, n384, n709, n743, n539);
xor  g1127 (n1062, n337, n945, n498, n553);
nor  g1128 (n1275, n928, n896, n345, n889);
nor  g1129 (n1216, n340, n445, n871, n898);
nand g1130 (n1256, n850, n454, n657, n928);
nand g1131 (n1039, n613, n933, n353, n305);
or   g1132 (n1076, n363, n920, n885, n937);
and  g1133 (n977, n454, n735, n683, n655);
xnor g1134 (n1184, n897, n409, n696, n417);
nand g1135 (n1133, n563, n567, n767, n821);
and  g1136 (n1250, n353, n311, n801, n902);
and  g1137 (n1324, n481, n778, n352, n429);
nor  g1138 (n1004, n877, n604, n587, n531);
xor  g1139 (n1215, n727, n329, n654, n918);
and  g1140 (n1137, n914, n728, n586, n337);
or   g1141 (n1114, n726, n442, n874, n937);
nor  g1142 (n1000, n715, n504, n918, n324);
xor  g1143 (n1291, n635, n837, n516, n634);
and  g1144 (n1158, n680, n380, n588, n352);
xor  g1145 (n974, n785, n803, n609, n525);
nor  g1146 (n1058, n493, n909, n592, n295);
and  g1147 (n1253, n815, n896, n485, n807);
nor  g1148 (n1120, n606, n398, n734, n604);
xnor g1149 (n1020, n324, n500, n935, n736);
nand g1150 (n1252, n889, n880, n673, n795);
and  g1151 (n1087, n760, n330, n717, n575);
xnor g1152 (n992, n655, n768, n873, n666);
xor  g1153 (n1163, n522, n725, n369, n450);
nor  g1154 (n1104, n492, n715, n878, n286);
xnor g1155 (n1124, n806, n286, n416, n318);
nand g1156 (n1118, n607, n724, n678, n552);
or   g1157 (n1203, n659, n567, n495, n326);
nor  g1158 (n1026, n871, n310, n396, n752);
nand g1159 (n1016, n512, n532, n877, n800);
xor  g1160 (n976, n827, n895, n389, n457);
nand g1161 (n1260, n627, n718, n578, n573);
or   g1162 (n1176, n753, n287, n315, n713);
nand g1163 (n1266, n522, n795, n883, n411);
and  g1164 (n1060, n848, n704, n370, n291);
xnor g1165 (n1078, n431, n859, n562, n586);
and  g1166 (n1288, n755, n443, n613, n521);
and  g1167 (n1220, n472, n833, n802, n684);
nand g1168 (n1086, n870, n625, n305, n407);
and  g1169 (n999, n650, n930, n751, n733);
nand g1170 (n1072, n785, n395, n513, n703);
nand g1171 (n1159, n478, n415, n750, n942);
and  g1172 (n1204, n692, n293, n595, n458);
nand g1173 (n1160, n524, n929, n523, n408);
xnor g1174 (n1283, n633, n491, n421, n423);
xnor g1175 (n1223, n336, n682, n830, n306);
or   g1176 (n1021, n899, n576, n905, n546);
or   g1177 (n1154, n602, n474, n820, n898);
nor  g1178 (n1139, n501, n789, n931, n910);
xnor g1179 (n1093, n919, n536, n772, n471);
xnor g1180 (n1064, n913, n907, n939, n614);
xnor g1181 (n1303, n372, n469, n580, n583);
or   g1182 (n1101, n883, n740, n359, n367);
nor  g1183 (n1146, n297, n497, n478, n888);
or   g1184 (n1238, n748, n486, n691, n294);
xnor g1185 (n1115, n462, n780, n749, n315);
nor  g1186 (n1233, n511, n903, n412, n335);
and  g1187 (n1243, n787, n375, n669, n746);
xnor g1188 (n1186, n282, n400, n328, n672);
and  g1189 (n1261, n876, n631, n894, n350);
xnor g1190 (n1029, n398, n557, n320, n931);
xnor g1191 (n1293, n427, n726, n899, n593);
xnor g1192 (n1152, n773, n761, n776, n743);
nor  g1193 (n1279, n530, n504, n489, n774);
xnor g1194 (n1282, n881, n775, n864, n890);
nand g1195 (n1009, n770, n297, n520, n534);
and  g1196 (n1249, n364, n849, n347, n882);
xnor g1197 (n1213, n641, n627, n517, n801);
nand g1198 (n1069, n668, n601, n645, n939);
xnor g1199 (n1123, n451, n458, n924, n414);
or   g1200 (n1240, n941, n388, n541, n810);
nand g1201 (n1150, n871, n742, n288, n374);
xor  g1202 (n1105, n750, n900, n729, n411);
xnor g1203 (n1221, n863, n909, n626, n437);
or   g1204 (n1325, n378, n623, n639, n624);
xnor g1205 (n1127, n658, n692, n804, n556);
nand g1206 (n1224, n306, n775, n361, n570);
xor  g1207 (n1231, n358, n835, n599, n916);
xnor g1208 (n1027, n662, n617, n335, n605);
nand g1209 (n1273, n872, n373, n483, n563);
or   g1210 (n1181, n662, n450, n799, n932);
nand g1211 (n1225, n529, n729, n611, n598);
and  g1212 (n1007, n898, n860, n851, n397);
xnor g1213 (n969, n766, n840, n357, n947);
or   g1214 (n1025, n374, n393, n320, n580);
or   g1215 (n1088, n638, n867, n709, n671);
nand g1216 (n1180, n285, n867, n694, n918);
or   g1217 (n1190, n527, n631, n900, n931);
nor  g1218 (n1274, n378, n473, n881, n612);
nand g1219 (n1297, n605, n559, n810, n321);
nand g1220 (n982, n392, n865, n819, n895);
or   g1221 (n1079, n584, n409, n821, n719);
xor  g1222 (n1255, n371, n448, n437, n283);
or   g1223 (n1116, n425, n570, n548, n910);
nor  g1224 (n1202, n675, n474, n650, n556);
or   g1225 (n1196, n676, n547, n934, n718);
or   g1226 (n1156, n946, n816, n851, n897);
xor  g1227 (n1111, n879, n314, n875, n385);
xor  g1228 (n1329, n783, n284, n373, n839);
nor  g1229 (n1207, n486, n895, n823, n916);
xor  g1230 (n984, n772, n619, n894, n921);
xor  g1231 (n1287, n314, n442, n928, n738);
nand g1232 (n1316, n651, n282, n831, n424);
and  g1233 (n1121, n843, n377, n550, n596);
or   g1234 (n1299, n929, n576, n759, n681);
and  g1235 (n1313, n891, n875, n379, n872);
nor  g1236 (n1122, n358, n927, n386, n371);
xor  g1237 (n1222, n906, n628, n757, n831);
xnor g1238 (n1172, n295, n595, n289, n879);
nor  g1239 (n1300, n885, n710, n568, n764);
xor  g1240 (n997, n939, n574, n441, n744);
nor  g1241 (n1033, n540, n846, n553, n296);
xnor g1242 (n1117, n452, n470, n786, n682);
nand g1243 (n1164, n351, n610, n700, n869);
xnor g1244 (n1187, n412, n890, n637, n309);
nor  g1245 (n1208, n355, n505, n509, n313);
nor  g1246 (n1001, n826, n847, n319, n904);
nand g1247 (n1244, n941, n667, n508, n589);
xor  g1248 (n1236, n671, n902, n882, n393);
xnor g1249 (n1171, n924, n893, n657, n873);
xnor g1250 (n1227, n490, n479, n797, n602);
or   g1251 (n989, n375, n465, n527, n518);
and  g1252 (n1109, n863, n868, n287, n879);
nor  g1253 (n1103, n945, n944, n790, n850);
xor  g1254 (n1200, n765, n756, n601, n830);
nor  g1255 (n1232, n525, n630, n310, n336);
nand g1256 (n981, n798, n646, n880, n544);
xnor g1257 (n1063, n642, n476, n905, n552);
nand g1258 (n1242, n538, n544, n524, n355);
xor  g1259 (n1272, n292, n674, n323, n542);
nand g1260 (n1245, n915, n685, n410, n779);
or   g1261 (n1042, n468, n722, n711, n689);
xnor g1262 (n1013, n827, n914, n386, n834);
nand g1263 (n1036, n299, n909, n899, n721);
nand g1264 (n1201, n572, n555, n902, n565);
and  g1265 (n1178, n920, n288, n585, n330);
xnor g1266 (n1077, n577, n591, n510, n903);
nand g1267 (n1230, n908, n940, n864, n496);
and  g1268 (n1247, n475, n499, n675, n483);
xnor g1269 (n1074, n436, n747, n285, n638);
nor  g1270 (n1239, n752, n919, n621, n900);
xor  g1271 (n1174, n461, n776, n538, n354);
nand g1272 (n1055, n932, n817, n346, n928);
xnor g1273 (n1258, n902, n360, n658, n366);
xor  g1274 (n1028, n300, n508, n911, n861);
or   g1275 (n1333, n435, n528, n643, n868);
xnor g1276 (n1298, n938, n307, n439, n600);
xnor g1277 (n1161, n338, n706, n549, n456);
and  g1278 (n1041, n439, n298, n862, n501);
nor  g1279 (n980, n390, n737, n408, n316);
or   g1280 (n1082, n687, n361, n708, n329);
and  g1281 (n970, n694, n894, n891, n468);
nand g1282 (n1059, n480, n405, n313, n879);
xor  g1283 (n1038, n597, n451, n701, n384);
xor  g1284 (n1312, n880, n762, n753, n593);
nand g1285 (n1102, n665, n630, n590, n697);
xnor g1286 (n1107, n660, n654, n778, n428);
xor  g1287 (n1003, n716, n781, n888, n529);
or   g1288 (n1265, n717, n432, n876, n360);
or   g1289 (n1166, n623, n401, n370, n926);
xnor g1290 (n1012, n646, n332, n441, n943);
and  g1291 (n1040, n343, n644, n910, n871);
or   g1292 (n1269, n308, n927, n669, n713);
nand g1293 (n1197, n618, n767, n904, n812);
xnor g1294 (n1199, n533, n945, n780, n876);
or   g1295 (n1307, n731, n636, n621, n460);
nor  g1296 (n1092, n925, n706, n385, n866);
nor  g1297 (n1331, n923, n311, n365, n499);
xor  g1298 (n1151, n435, n781, n794, n815);
nor  g1299 (n1314, n698, n905, n609, n681);
and  g1300 (n1136, n936, n404, n705, n455);
and  g1301 (n1192, n859, n944, n679, n312);
nand g1302 (n1340, n982, n1023, n974, n1005);
xor  g1303 (n1336, n969, n986, n1031, n981);
or   g1304 (n1345, n1010, n991, n1014, n966);
or   g1305 (n1335, n979, n1026, n985, n1000);
xnor g1306 (n1350, n1018, n1020, n983, n1006);
xor  g1307 (n1348, n964, n1007, n977, n1016);
xnor g1308 (n1343, n992, n1012, n1025, n976);
and  g1309 (n1344, n989, n1009, n980, n995);
or   g1310 (n1352, n1029, n1001, n963, n1022);
xnor g1311 (n1339, n997, n1003, n971, n962);
or   g1312 (n1337, n987, n993, n1024, n968);
nor  g1313 (n1342, n1019, n1015, n984, n996);
xor  g1314 (n1341, n978, n1011, n988, n994);
xor  g1315 (n1338, n967, n1032, n972, n1027);
or   g1316 (n1347, n973, n998, n1030, n975);
nor  g1317 (n1346, n990, n999, n1017, n1002);
nor  g1318 (n1351, n1033, n1004, n970, n1028);
nor  g1319 (n1349, n1021, n1008, n1013, n965);
buf  g1320 (n1358, n1342);
buf  g1321 (n1356, n1341);
not  g1322 (n1354, n1339);
not  g1323 (n1353, n1348);
buf  g1324 (n1363, n1343);
not  g1325 (n1355, n1336);
not  g1326 (n1366, n269);
not  g1327 (n1362, n1346);
buf  g1328 (n1359, n1338);
not  g1329 (n1357, n269);
buf  g1330 (n1365, n1344);
buf  g1331 (n1364, n1347);
or   g1332 (n1361, n1340, n1335);
nand g1333 (n1360, n1345, n1337, n269);
buf  g1334 (n1377, n1354);
not  g1335 (n1371, n1358);
buf  g1336 (n1379, n1359);
buf  g1337 (n1372, n1353);
buf  g1338 (n1380, n1357);
buf  g1339 (n1368, n1356);
buf  g1340 (n1382, n1355);
not  g1341 (n1383, n1355);
not  g1342 (n1381, n1359);
not  g1343 (n1386, n1357);
buf  g1344 (n1374, n1358);
buf  g1345 (n1373, n1358);
buf  g1346 (n1367, n1357);
buf  g1347 (n1369, n1359);
buf  g1348 (n1370, n1359);
not  g1349 (n1375, n1357);
not  g1350 (n1384, n1354);
buf  g1351 (n1385, n1353);
buf  g1352 (n1376, n1358);
buf  g1353 (n1378, n1356);
or   g1354 (n1456, n1173, n1369, n1241, n1270);
xnor g1355 (n1462, n1368, n1236, n1232, n1071);
and  g1356 (n1443, n1145, n1378, n1374, n1182);
nor  g1357 (n1450, n1062, n1257, n1226, n1197);
nor  g1358 (n1455, n1181, n1227, n1177, n1120);
nand g1359 (n1444, n1101, n1104, n1114, n1382);
xnor g1360 (n1440, n1386, n1235, n1196, n1269);
xnor g1361 (n1417, n1133, n1155, n1371, n1213);
nand g1362 (n1405, n1260, n1147, n1249, n1386);
or   g1363 (n1449, n1372, n1384, n1050, n1191);
xor  g1364 (n1411, n1125, n1262, n1385, n1228);
xnor g1365 (n1453, n1080, n1201, n1045, n1156);
nor  g1366 (n1421, n1242, n1383, n1251, n1246);
xnor g1367 (n1427, n1074, n1183, n1381, n1141);
xor  g1368 (n1437, n1167, n1069, n1384, n1377);
and  g1369 (n1429, n1038, n1068, n1093, n1157);
xnor g1370 (n1424, n1385, n1189, n1130, n1134);
nor  g1371 (n1412, n1372, n1371, n1165, n1253);
nor  g1372 (n1413, n1161, n1057, n1188, n1386);
and  g1373 (n1396, n1267, n1090, n1209, n1218);
nand g1374 (n1409, n1273, n1124, n1210, n1233);
nor  g1375 (n1401, n1138, n1372, n1265, n1162);
xnor g1376 (n1419, n1149, n1375, n1166, n1059);
xnor g1377 (n1416, n1041, n1373, n1383, n1217);
or   g1378 (n1394, n1216, n1136, n1379, n1077);
nor  g1379 (n1432, n1386, n1179, n1103, n1379);
xor  g1380 (n1447, n1252, n1144, n1040, n1194);
or   g1381 (n1466, n1370, n1374, n1375, n1271);
nor  g1382 (n1457, n1369, n1231, n1368, n1079);
xnor g1383 (n1403, n1121, n1107, n1379, n1072);
nor  g1384 (n1465, n1087, n1139, n1172, n1272);
xor  g1385 (n1398, n1369, n1203, n1099, n1094);
nand g1386 (n1441, n1381, n1110, n1206, n1065);
and  g1387 (n1423, n1067, n1381, n1176, n1380);
or   g1388 (n1387, n1132, n1192, n1234, n1160);
xor  g1389 (n1436, n1108, n1106, n1143, n1053);
nand g1390 (n1404, n1111, n1381, n1046, n1034);
nand g1391 (n1393, n1150, n1043, n1223, n1054);
xor  g1392 (n1418, n1086, n1377, n1075, n1088);
nand g1393 (n1428, n1118, n1367, n1247, n1230);
xor  g1394 (n1452, n1174, n1140, n1225, n1255);
nand g1395 (n1431, n1379, n1168, n1212, n1367);
xnor g1396 (n1407, n1055, n1219, n1187, n1229);
or   g1397 (n1420, n1371, n1078, n1119, n1044);
or   g1398 (n1392, n1100, n1142, n1238, n1244);
nand g1399 (n1425, n1169, n1377, n1215, n1385);
xnor g1400 (n1395, n1383, n1035, n1378);
xor  g1401 (n1446, n1070, n1186, n1175, n1375);
or   g1402 (n1430, n1367, n1049, n1259, n1116);
and  g1403 (n1410, n1250, n1066, n1131, n1063);
xnor g1404 (n1458, n1370, n1254, n1221, n1185);
xor  g1405 (n1426, n1380, n1170, n1383, n1064);
nand g1406 (n1454, n1382, n1266, n1037, n1243);
xnor g1407 (n1445, n1105, n1039, n1091, n1369);
nor  g1408 (n1415, n1089, n1085, n1384);
xor  g1409 (n1463, n1372, n1382, n1220, n1098);
nand g1410 (n1389, n1152, n1268, n1258, n1052);
and  g1411 (n1399, n1109, n1199, n1204, n1153);
xnor g1412 (n1397, n1135, n1376, n1081, n1158);
or   g1413 (n1461, n1373, n1073, n1375, n1083);
xor  g1414 (n1435, n1163, n1123, n1376, n1082);
xnor g1415 (n1434, n1382, n1126, n1048, n1127);
xor  g1416 (n1422, n1190, n1376, n1198, n1151);
xor  g1417 (n1459, n1148, n1261, n1237, n1373);
or   g1418 (n1460, n1096, n1211, n1154, n1263);
nor  g1419 (n1406, n1092, n1380, n1368, n1222);
nor  g1420 (n1433, n1245, n1129, n1380, n1180);
or   g1421 (n1390, n1264, n1117, n1239, n1195);
xnor g1422 (n1402, n1047, n1256, n1368, n1128);
nor  g1423 (n1451, n1208, n1376, n1373, n1171);
xnor g1424 (n1391, n1371, n1112, n1370, n1248);
or   g1425 (n1408, n1200, n1060, n1178, n1122);
xnor g1426 (n1448, n1370, n1137, n1056, n1385);
and  g1427 (n1439, n1042, n1207, n1193, n1084);
and  g1428 (n1388, n1240, n1377, n1214, n1097);
xor  g1429 (n1414, n1374, n1367, n1115, n1146);
nor  g1430 (n1438, n1374, n1378, n1061, n1224);
or   g1431 (n1400, n1051, n1159, n1184, n1058);
nor  g1432 (n1464, n1113, n1202, n1076, n1095);
xor  g1433 (n1442, n1036, n1164, n1205, n1102);
not  g1434 (n1467, n1387);
not  g1435 (n1468, n1387);
not  g1436 (n1470, n1387);
buf  g1437 (n1469, n1387);
buf  g1438 (n1477, n1362);
not  g1439 (n1472, n1467);
nor  g1440 (n1478, n1467, n1280, n1363, n1468);
xnor g1441 (n1476, n1363, n1276, n1360);
and  g1442 (n1473, n1361, n1360, n1275, n1362);
or   g1443 (n1475, n1362, n1467, n1468);
or   g1444 (n1471, n1468, n1277, n1469, n1360);
xnor g1445 (n1474, n1362, n1274, n1361, n1279);
xnor g1446 (n1479, n1278, n1361, n1468);
buf  g1447 (n1484, n1473);
buf  g1448 (n1493, n1471);
not  g1449 (n1487, n1474);
buf  g1450 (n1489, n1472);
not  g1451 (n1480, n1471);
not  g1452 (n1485, n1473);
buf  g1453 (n1495, n1471);
buf  g1454 (n1481, n1472);
not  g1455 (n1494, n1474);
buf  g1456 (n1491, n1473);
not  g1457 (n1482, n1474);
not  g1458 (n1492, n1474);
not  g1459 (n1483, n1472);
buf  g1460 (n1488, n1472);
buf  g1461 (n1486, n1471);
not  g1462 (n1490, n1473);
xor  g1463 (n1543, n1390, n1401);
nor  g1464 (n1522, n1394, n1483);
xnor g1465 (n1540, n1487, n1397, n1396, n1489);
nor  g1466 (n1536, n1487, n1389, n1416, n1415);
xor  g1467 (n1496, n1480, n1416, n1402, n1418);
or   g1468 (n1535, n1481, n1424, n1389, n1409);
nor  g1469 (n1519, n1486, n1402, n1415, n1406);
xnor g1470 (n1542, n1420, n1409, n1413, n1423);
nand g1471 (n1499, n1424, n1488, n1413, n1421);
or   g1472 (n1548, n1400, n1426, n1412, n1401);
xor  g1473 (n1529, n1484, n1401, n1392, n1490);
nand g1474 (n1504, n1407, n1490, n1417, n1418);
nand g1475 (n1538, n1400, n1397, n1414, n1491);
xnor g1476 (n1526, n1420, n1408, n1391);
nand g1477 (n1505, n1486, n1487, n1392, n1388);
nand g1478 (n1516, n1413, n1420, n1492, n1402);
or   g1479 (n1518, n1411, n1481, n1491, n1393);
nor  g1480 (n1501, n1482, n1485);
xor  g1481 (n1531, n1416, n1488, n1412, n1398);
xnor g1482 (n1506, n1489, n1423, n1491, n1481);
xnor g1483 (n1527, n1417, n1421, n1422, n1426);
or   g1484 (n1503, n1395, n1417, n1413, n1406);
nand g1485 (n1515, n1425, n1419, n1426, n1395);
xor  g1486 (n1517, n1410, n1402, n1419, n1398);
or   g1487 (n1544, n1483, n1421, n1492, n1404);
xnor g1488 (n1547, n1405, n1412, n1411, n1418);
and  g1489 (n1546, n1483, n1425, n1396, n1410);
xnor g1490 (n1500, n1403, n1399, n1480, n1391);
xnor g1491 (n1502, n1486, n1392, n1412, n1485);
or   g1492 (n1534, n1398, n1422, n1405, n1484);
xor  g1493 (n1514, n1425, n1489, n1391, n1388);
nor  g1494 (n1507, n1408, n1482, n1394, n1400);
xor  g1495 (n1508, n1492, n1480, n1484, n1406);
xnor g1496 (n1523, n1396, n1425, n1400, n1390);
xnor g1497 (n1509, n1422, n1489, n1420, n1394);
xnor g1498 (n1545, n1417, n1492, n1423, n1406);
nor  g1499 (n1537, n1486, n1396, n1415, n1407);
or   g1500 (n1497, n1424, n1403, n1405, n1388);
nand g1501 (n1530, n1482, n1399, n1401, n1421);
nand g1502 (n1511, n1408, n1393, n1488, n1480);
or   g1503 (n1521, n1410, n1393, n1414, n1394);
nand g1504 (n1512, n1397, n1483, n1399, n1391);
nor  g1505 (n1524, n1393, n1414, n1399, n1423);
xnor g1506 (n1541, n1424, n1411, n1487, n1490);
xor  g1507 (n1539, n1397, n1407, n1404, n1410);
xnor g1508 (n1533, n1403, n1398, n1411, n1390);
xor  g1509 (n1510, n1419, n1409, n1392, n1488);
nor  g1510 (n1520, n1390, n1404, n1389, n1409);
nor  g1511 (n1513, n1490, n1407, n1395, n1493);
and  g1512 (n1498, n1419, n1416, n1405, n1491);
and  g1513 (n1525, n1422, n1484, n1485, n1418);
and  g1514 (n1532, n1389, n1404, n1403, n1414);
nor  g1515 (n1528, n1481, n1415, n1388, n1395);
and  g1516 (n1582, n1432, n950, n1469, n1296);
nor  g1517 (n1560, n1438, n948, n1493, n1508);
nor  g1518 (n1585, n274, n1517, n1526, n949);
xnor g1519 (n1565, n1527, n271, n1497, n1520);
nand g1520 (n1562, n1441, n1435, n1439, n270);
or   g1521 (n1594, n1288, n1547, n272, n1427);
and  g1522 (n1584, n1430, n1364, n1516, n1284);
nor  g1523 (n1579, n271, n1429, n273, n270);
xor  g1524 (n1592, n1428, n1365, n1293, n1431);
nand g1525 (n1598, n950, n270, n1433, n1427);
nand g1526 (n1570, n1470, n1535, n1503, n1439);
or   g1527 (n1596, n274, n1430, n1439, n1499);
nor  g1528 (n1549, n1429, n1437, n271, n1442);
xor  g1529 (n1587, n270, n1532, n949, n1443);
or   g1530 (n1571, n1438, n1364, n79, n1510);
or   g1531 (n1595, n1435, n952, n950, n1436);
nand g1532 (n1589, n1506, n1282, n1544, n1364);
xnor g1533 (n1553, n1285, n1430, n1438, n950);
nor  g1534 (n1593, n1530, n1437, n1513, n1469);
or   g1535 (n1550, n951, n1435, n949, n1363);
or   g1536 (n1563, n1540, n1433, n1294, n1502);
nand g1537 (n1578, n1507, n1439, n275);
nand g1538 (n1559, n1546, n1519, n272, n1529);
and  g1539 (n1590, n79, n1289, n1543, n951);
nor  g1540 (n1574, n1469, n1434, n1426, n274);
nand g1541 (n1557, n1537, n1363, n1524, n1431);
xnor g1542 (n1575, n1435, n1433, n947, n1440);
xnor g1543 (n1558, n1545, n1470, n79);
nor  g1544 (n1581, n1440, n1505, n273, n1427);
xnor g1545 (n1586, n1523, n1290, n1428, n1538);
xnor g1546 (n1597, n1522, n1500, n1365, n1350);
and  g1547 (n1568, n1432, n1364, n1531, n1440);
nand g1548 (n1577, n1352, n272, n1436, n1509);
or   g1549 (n1573, n1501, n1431, n949, n273);
nor  g1550 (n1564, n1287, n1470, n1431, n1514);
xor  g1551 (n1566, n1281, n1541, n1512, n1365);
and  g1552 (n1555, n1441, n1428, n951);
xor  g1553 (n1599, n1351, n1434, n1436, n1536);
xor  g1554 (n1583, n276, n273, n1432, n1442);
xnor g1555 (n1556, n1441, n1493, n1427, n1498);
xnor g1556 (n1561, n1292, n1525, n1434, n1438);
xnor g1557 (n1569, n1286, n1440, n271, n1542);
xor  g1558 (n1591, n948, n1295, n1548, n1518);
or   g1559 (n1572, n1429, n1437, n948, n1494);
nand g1560 (n1551, n947, n1442, n274, n1430);
xor  g1561 (n1552, n1349, n1442, n1429, n1493);
nand g1562 (n1580, n1534, n1515, n275, n78);
or   g1563 (n1600, n272, n1432, n1437, n1521);
and  g1564 (n1576, n1433, n948, n951, n1434);
xnor g1565 (n1554, n275, n1365, n1511, n1436);
nor  g1566 (n1567, n1283, n79, n1504, n1528);
or   g1567 (n1588, n1533, n1291, n1441, n1539);
buf  g1568 (n1626, n1570);
not  g1569 (n1672, n1575);
buf  g1570 (n1794, n1593);
buf  g1571 (n1690, n1551);
buf  g1572 (n1748, n1586);
buf  g1573 (n1782, n1559);
buf  g1574 (n1606, n1553);
not  g1575 (n1753, n1597);
buf  g1576 (n1714, n1587);
buf  g1577 (n1670, n1557);
not  g1578 (n1668, n1571);
not  g1579 (n1736, n1565);
not  g1580 (n1603, n1579);
buf  g1581 (n1750, n1560);
not  g1582 (n1702, n1596);
buf  g1583 (n1747, n1572);
buf  g1584 (n1665, n1568);
buf  g1585 (n1757, n1569);
not  g1586 (n1646, n1575);
buf  g1587 (n1725, n1597);
not  g1588 (n1790, n1588);
not  g1589 (n1696, n1579);
not  g1590 (n1742, n1575);
buf  g1591 (n1614, n1584);
not  g1592 (n1629, n1554);
not  g1593 (n1662, n1585);
not  g1594 (n1632, n1558);
not  g1595 (n1608, n1551);
not  g1596 (n1723, n1479);
not  g1597 (n1621, n1554);
buf  g1598 (n1617, n1600);
not  g1599 (n1688, n1567);
buf  g1600 (n1805, n1476);
buf  g1601 (n1631, n1479);
buf  g1602 (n1795, n1566);
buf  g1603 (n1746, n1592);
buf  g1604 (n1800, n1562);
not  g1605 (n1735, n1476);
not  g1606 (n1673, n1600);
buf  g1607 (n1604, n1560);
buf  g1608 (n1793, n1561);
buf  g1609 (n1726, n1577);
buf  g1610 (n1781, n1598);
not  g1611 (n1756, n1599);
buf  g1612 (n1709, n1576);
not  g1613 (n1738, n1580);
buf  g1614 (n1787, n1571);
buf  g1615 (n1745, n1583);
buf  g1616 (n1763, n1590);
buf  g1617 (n1715, n1584);
buf  g1618 (n1737, n1552);
not  g1619 (n1788, n1574);
buf  g1620 (n1661, n1580);
not  g1621 (n1642, n1478);
buf  g1622 (n1773, n1557);
not  g1623 (n1767, n1598);
not  g1624 (n1752, n1569);
not  g1625 (n1691, n1567);
buf  g1626 (n1612, n1562);
not  g1627 (n1644, n1552);
not  g1628 (n1601, n1591);
buf  g1629 (n1666, n1592);
not  g1630 (n1679, n1550);
buf  g1631 (n1743, n1589);
not  g1632 (n1692, n1563);
not  g1633 (n1807, n1549);
not  g1634 (n1769, n1598);
buf  g1635 (n1766, n1590);
buf  g1636 (n1719, n1566);
buf  g1637 (n1609, n1561);
not  g1638 (n1799, n1561);
not  g1639 (n1657, n1585);
not  g1640 (n1768, n1597);
not  g1641 (n1624, n1588);
not  g1642 (n1703, n1574);
not  g1643 (n1710, n1567);
not  g1644 (n1754, n1572);
buf  g1645 (n1681, n1564);
buf  g1646 (n1802, n1596);
buf  g1647 (n1722, n1589);
buf  g1648 (n1732, n1569);
not  g1649 (n1650, n1581);
not  g1650 (n1651, n1558);
buf  g1651 (n1783, n1564);
buf  g1652 (n1697, n1551);
buf  g1653 (n1700, n1576);
buf  g1654 (n1640, n1557);
not  g1655 (n1694, n1475);
not  g1656 (n1716, n1573);
buf  g1657 (n1731, n1568);
buf  g1658 (n1762, n1577);
buf  g1659 (n1619, n1567);
not  g1660 (n1605, n1577);
not  g1661 (n1647, n1556);
not  g1662 (n1622, n1565);
buf  g1663 (n1695, n1560);
not  g1664 (n1680, n1478);
not  g1665 (n1740, n1478);
buf  g1666 (n1765, n1556);
buf  g1667 (n1789, n1593);
not  g1668 (n1777, n1582);
buf  g1669 (n1685, n1560);
not  g1670 (n1636, n1568);
not  g1671 (n1620, n1599);
not  g1672 (n1751, n1477);
buf  g1673 (n1669, n1594);
buf  g1674 (n1711, n1591);
buf  g1675 (n1728, n1581);
not  g1676 (n1659, n1600);
not  g1677 (n1638, n1563);
buf  g1678 (n1775, n1591);
buf  g1679 (n1618, n1565);
buf  g1680 (n1734, n1578);
not  g1681 (n1804, n1593);
not  g1682 (n1806, n1570);
not  g1683 (n1607, n1558);
buf  g1684 (n1671, n1551);
buf  g1685 (n1796, n1595);
not  g1686 (n1760, n1578);
buf  g1687 (n1724, n1577);
not  g1688 (n1705, n1591);
not  g1689 (n1641, n1549);
not  g1690 (n1625, n1479);
buf  g1691 (n1759, n1574);
not  g1692 (n1771, n1555);
not  g1693 (n1602, n1571);
not  g1694 (n1718, n1552);
not  g1695 (n1613, n1477);
not  g1696 (n1678, n1596);
not  g1697 (n1634, n1593);
not  g1698 (n1628, n1565);
not  g1699 (n1676, n1581);
not  g1700 (n1664, n1595);
buf  g1701 (n1761, n1554);
buf  g1702 (n1713, n1588);
buf  g1703 (n1675, n1581);
not  g1704 (n1656, n1582);
buf  g1705 (n1798, n1562);
buf  g1706 (n1610, n1475);
buf  g1707 (n1635, n1573);
buf  g1708 (n1730, n1552);
buf  g1709 (n1706, n1590);
not  g1710 (n1776, n1583);
buf  g1711 (n1755, n1550);
not  g1712 (n1654, n1600);
not  g1713 (n1689, n1555);
not  g1714 (n1683, n1597);
not  g1715 (n1637, n1590);
buf  g1716 (n1686, n1578);
buf  g1717 (n1648, n1476);
not  g1718 (n1627, n1575);
buf  g1719 (n1733, n1587);
buf  g1720 (n1785, n1477);
buf  g1721 (n1797, n1599);
buf  g1722 (n1630, n1550);
buf  g1723 (n1687, n1475);
buf  g1724 (n1720, n1569);
buf  g1725 (n1643, n1563);
not  g1726 (n1653, n1598);
not  g1727 (n1698, n1579);
not  g1728 (n1774, n1555);
buf  g1729 (n1803, n1572);
buf  g1730 (n1633, n1587);
buf  g1731 (n1699, n1596);
buf  g1732 (n1704, n1595);
buf  g1733 (n1749, n1559);
not  g1734 (n1727, n1586);
buf  g1735 (n1663, n1566);
buf  g1736 (n1615, n1561);
buf  g1737 (n1729, n1583);
not  g1738 (n1721, n1573);
buf  g1739 (n1791, n1564);
not  g1740 (n1712, n1579);
not  g1741 (n1707, n1571);
not  g1742 (n1677, n1586);
not  g1743 (n1652, n1554);
buf  g1744 (n1764, n1568);
not  g1745 (n1779, n1559);
not  g1746 (n1684, n1594);
not  g1747 (n1801, n1595);
not  g1748 (n1772, n1576);
buf  g1749 (n1744, n1564);
buf  g1750 (n1616, n1553);
not  g1751 (n1649, n1563);
buf  g1752 (n1784, n1588);
buf  g1753 (n1778, n1592);
not  g1754 (n1758, n1553);
buf  g1755 (n1739, n1592);
buf  g1756 (n1658, n1599);
buf  g1757 (n1682, n1562);
buf  g1758 (n1741, n1570);
not  g1759 (n1693, n1594);
not  g1760 (n1717, n1550);
not  g1761 (n1780, n1585);
buf  g1762 (n1611, n1589);
not  g1763 (n1667, n1478);
not  g1764 (n1808, n1584);
buf  g1765 (n1792, n1589);
not  g1766 (n1701, n1576);
not  g1767 (n1623, n1574);
not  g1768 (n1786, n1479);
or   g1769 (n1645, n1582, n1573, n1557);
xor  g1770 (n1674, n1558, n1475, n1559, n1549);
and  g1771 (n1639, n1549, n1584, n1594, n1578);
nor  g1772 (n1708, n1476, n1587, n1585, n1580);
and  g1773 (n1660, n1582, n1583, n1566, n1570);
xor  g1774 (n1655, n1553, n1555, n1580, n1572);
nand g1775 (n1770, n1477, n1556, n1586);
buf  g1776 (n1853, n1650);
not  g1777 (n2134, n1646);
buf  g1778 (n2092, n1715);
not  g1779 (n2375, n1695);
not  g1780 (n2244, n1668);
not  g1781 (n2069, n1693);
not  g1782 (n2296, n1726);
buf  g1783 (n1887, n1792);
buf  g1784 (n2107, n1763);
buf  g1785 (n1996, n1730);
buf  g1786 (n2185, n1778);
not  g1787 (n2288, n1729);
not  g1788 (n1925, n1495);
buf  g1789 (n2114, n1728);
not  g1790 (n1992, n1723);
not  g1791 (n2062, n1684);
not  g1792 (n2262, n1714);
not  g1793 (n1895, n1673);
buf  g1794 (n1972, n1763);
not  g1795 (n2111, n1632);
not  g1796 (n1981, n1671);
not  g1797 (n2106, n1603);
buf  g1798 (n1826, n1776);
buf  g1799 (n2089, n1696);
buf  g1800 (n1913, n1678);
not  g1801 (n1933, n1737);
not  g1802 (n2316, n1794);
buf  g1803 (n2327, n1637);
not  g1804 (n2266, n1658);
not  g1805 (n2036, n1715);
not  g1806 (n2238, n1629);
not  g1807 (n2030, n1724);
buf  g1808 (n2359, n1807);
buf  g1809 (n2142, n1724);
not  g1810 (n2085, n1749);
not  g1811 (n2053, n1750);
not  g1812 (n2306, n1638);
not  g1813 (n2381, n1665);
buf  g1814 (n1898, n1682);
buf  g1815 (n2127, n1746);
buf  g1816 (n2215, n1735);
not  g1817 (n1849, n1644);
buf  g1818 (n1980, n1705);
not  g1819 (n2105, n1746);
buf  g1820 (n2044, n1792);
not  g1821 (n2257, n1655);
not  g1822 (n2251, n1608);
buf  g1823 (n1984, n1724);
buf  g1824 (n2309, n1748);
buf  g1825 (n2050, n1623);
buf  g1826 (n2035, n1748);
buf  g1827 (n2122, n1767);
buf  g1828 (n2297, n1694);
not  g1829 (n1985, n1603);
buf  g1830 (n2131, n1608);
not  g1831 (n2322, n1667);
not  g1832 (n1882, n1661);
not  g1833 (n1840, n1798);
buf  g1834 (n2038, n1806);
buf  g1835 (n2292, n1629);
buf  g1836 (n2370, n1785);
buf  g1837 (n2263, n1716);
not  g1838 (n2135, n1627);
not  g1839 (n2249, n1745);
not  g1840 (n2016, n1634);
not  g1841 (n2311, n1640);
not  g1842 (n2214, n1764);
buf  g1843 (n2285, n1690);
not  g1844 (n2002, n1791);
not  g1845 (n1909, n1746);
not  g1846 (n1944, n1770);
buf  g1847 (n1920, n1736);
buf  g1848 (n2197, n1783);
not  g1849 (n2243, n1646);
buf  g1850 (n2178, n1754);
buf  g1851 (n2155, n1770);
buf  g1852 (n2293, n1753);
buf  g1853 (n1934, n1677);
buf  g1854 (n1941, n1778);
not  g1855 (n2174, n1715);
buf  g1856 (n1998, n1620);
not  g1857 (n2103, n1719);
not  g1858 (n1891, n1647);
buf  g1859 (n1879, n1666);
not  g1860 (n2290, n1756);
buf  g1861 (n2113, n1625);
buf  g1862 (n2312, n1621);
buf  g1863 (n2136, n1695);
not  g1864 (n2310, n1685);
buf  g1865 (n1931, n1777);
not  g1866 (n1819, n1611);
buf  g1867 (n1923, n1621);
buf  g1868 (n1885, n1793);
buf  g1869 (n2137, n1772);
buf  g1870 (n1912, n1755);
not  g1871 (n1864, n1673);
not  g1872 (n2330, n1709);
not  g1873 (n2274, n1640);
buf  g1874 (n2203, n1643);
not  g1875 (n2331, n1757);
buf  g1876 (n1815, n1804);
not  g1877 (n2216, n1638);
buf  g1878 (n1971, n1725);
buf  g1879 (n2004, n1663);
not  g1880 (n2321, n1787);
not  g1881 (n2011, n1751);
not  g1882 (n2065, n1681);
buf  g1883 (n1940, n1607);
buf  g1884 (n2273, n1667);
not  g1885 (n2230, n1765);
not  g1886 (n2098, n1495);
buf  g1887 (n2080, n1776);
not  g1888 (n1862, n1606);
buf  g1889 (n1818, n1649);
buf  g1890 (n1926, n1631);
not  g1891 (n2032, n1774);
buf  g1892 (n1850, n1765);
not  g1893 (n2110, n1622);
not  g1894 (n1869, n1784);
not  g1895 (n1811, n1603);
buf  g1896 (n1835, n1684);
buf  g1897 (n1861, n1768);
buf  g1898 (n2099, n1779);
not  g1899 (n2350, n1712);
not  g1900 (n2094, n1618);
not  g1901 (n2188, n1619);
not  g1902 (n1969, n1750);
buf  g1903 (n1859, n1792);
not  g1904 (n2121, n1679);
buf  g1905 (n2328, n1665);
not  g1906 (n2169, n1699);
buf  g1907 (n2353, n1793);
buf  g1908 (n1899, n1658);
buf  g1909 (n1883, n1762);
not  g1910 (n1950, n1639);
buf  g1911 (n1884, n1617);
buf  g1912 (n2366, n1760);
buf  g1913 (n2100, n1660);
buf  g1914 (n2138, n1619);
buf  g1915 (n2021, n1639);
not  g1916 (n2252, n1709);
not  g1917 (n2338, n1655);
not  g1918 (n2160, n1625);
buf  g1919 (n2031, n1603);
not  g1920 (n1994, n1732);
not  g1921 (n2242, n1723);
not  g1922 (n2182, n1737);
buf  g1923 (n2084, n1721);
not  g1924 (n2347, n1610);
not  g1925 (n1823, n1762);
buf  g1926 (n2161, n1674);
not  g1927 (n1977, n1722);
buf  g1928 (n2170, n1790);
not  g1929 (n2333, n1636);
not  g1930 (n1962, n1628);
buf  g1931 (n1852, n1787);
buf  g1932 (n1890, n1768);
not  g1933 (n2248, n1686);
not  g1934 (n2298, n1673);
not  g1935 (n2097, n1648);
buf  g1936 (n1902, n1651);
buf  g1937 (n2163, n1795);
buf  g1938 (n2219, n1777);
not  g1939 (n2074, n1741);
not  g1940 (n1824, n1792);
not  g1941 (n2237, n1615);
not  g1942 (n2229, n1781);
buf  g1943 (n2010, n1715);
not  g1944 (n2042, n1782);
not  g1945 (n2017, n1732);
buf  g1946 (n2264, n1707);
not  g1947 (n2102, n1683);
not  g1948 (n2341, n1741);
not  g1949 (n1841, n1666);
not  g1950 (n1905, n1689);
buf  g1951 (n2019, n1602);
buf  g1952 (n1914, n1743);
buf  g1953 (n2172, n1730);
not  g1954 (n2192, n1711);
not  g1955 (n1903, n1727);
not  g1956 (n2008, n1720);
not  g1957 (n2077, n1663);
not  g1958 (n1873, n1602);
not  g1959 (n2014, n1636);
buf  g1960 (n2147, n1801);
buf  g1961 (n1911, n1776);
buf  g1962 (n1904, n1684);
buf  g1963 (n2057, n1655);
not  g1964 (n1893, n1739);
not  g1965 (n2278, n1734);
not  g1966 (n2360, n1614);
buf  g1967 (n2261, n1801);
not  g1968 (n2159, n1601);
buf  g1969 (n2104, n1806);
not  g1970 (n1888, n1699);
buf  g1971 (n2209, n1652);
buf  g1972 (n2168, n1670);
buf  g1973 (n2270, n1678);
not  g1974 (n2046, n1648);
not  g1975 (n2294, n1765);
buf  g1976 (n2060, n1702);
buf  g1977 (n1810, n1691);
not  g1978 (n1922, n1620);
buf  g1979 (n2139, n1622);
not  g1980 (n2018, n1788);
not  g1981 (n1851, n1766);
not  g1982 (n1907, n1664);
buf  g1983 (n2207, n1780);
not  g1984 (n1865, n1738);
buf  g1985 (n2167, n1760);
buf  g1986 (n1866, n1775);
buf  g1987 (n2211, n1805);
not  g1988 (n2049, n1644);
not  g1989 (n2090, n1687);
not  g1990 (n1896, n1721);
not  g1991 (n2007, n1642);
buf  g1992 (n2256, n1781);
not  g1993 (n1827, n1706);
buf  g1994 (n2279, n1743);
buf  g1995 (n2189, n1797);
not  g1996 (n2344, n1771);
buf  g1997 (n1820, n1655);
buf  g1998 (n2096, n1677);
not  g1999 (n2054, n1646);
not  g2000 (n2156, n1656);
buf  g2001 (n2283, n1675);
buf  g2002 (n2368, n1613);
buf  g2003 (n2003, n1728);
not  g2004 (n1863, n1768);
buf  g2005 (n2371, n1617);
buf  g2006 (n2220, n1747);
not  g2007 (n2227, n1748);
not  g2008 (n2233, n1656);
not  g2009 (n2115, n1728);
not  g2010 (n1976, n1630);
not  g2011 (n2040, n1748);
buf  g2012 (n2091, n1662);
buf  g2013 (n2141, n1691);
buf  g2014 (n1844, n1745);
not  g2015 (n2145, n1807);
not  g2016 (n2171, n1740);
buf  g2017 (n2028, n1758);
buf  g2018 (n2340, n1785);
not  g2019 (n1966, n1767);
not  g2020 (n2128, n1799);
buf  g2021 (n2276, n1649);
not  g2022 (n1817, n1494);
not  g2023 (n2346, n1646);
not  g2024 (n1886, n1724);
not  g2025 (n2314, n1644);
not  g2026 (n1952, n1704);
buf  g2027 (n2177, n1806);
not  g2028 (n2058, n1612);
buf  g2029 (n1943, n1604);
not  g2030 (n2152, n1774);
buf  g2031 (n1982, n1638);
buf  g2032 (n2223, n1788);
buf  g2033 (n1834, n1691);
buf  g2034 (n2006, n1756);
buf  g2035 (n1878, n1690);
buf  g2036 (n2318, n1668);
buf  g2037 (n1937, n1690);
buf  g2038 (n2076, n1669);
not  g2039 (n2175, n1674);
buf  g2040 (n2225, n1672);
not  g2041 (n1857, n1776);
not  g2042 (n1874, n1681);
buf  g2043 (n2180, n1630);
not  g2044 (n1845, n1751);
buf  g2045 (n2260, n1701);
buf  g2046 (n1870, n1624);
not  g2047 (n1846, n1628);
buf  g2048 (n1921, n1742);
buf  g2049 (n2315, n1789);
buf  g2050 (n2123, n1636);
not  g2051 (n2253, n1761);
not  g2052 (n2001, n1752);
buf  g2053 (n2281, n1773);
not  g2054 (n2027, n1781);
buf  g2055 (n1954, n1630);
not  g2056 (n2358, n1758);
buf  g2057 (n1945, n1794);
not  g2058 (n2117, n1711);
buf  g2059 (n1928, n1772);
buf  g2060 (n1961, n1676);
buf  g2061 (n2034, n1804);
buf  g2062 (n2070, n1714);
not  g2063 (n2047, n1685);
buf  g2064 (n2342, n1659);
buf  g2065 (n2277, n1606);
buf  g2066 (n2250, n1641);
buf  g2067 (n1831, n1606);
not  g2068 (n1892, n1788);
not  g2069 (n2148, n1805);
not  g2070 (n2164, n1726);
not  g2071 (n1848, n1667);
not  g2072 (n2267, n1619);
not  g2073 (n2140, n1766);
buf  g2074 (n2205, n1673);
not  g2075 (n2324, n1752);
buf  g2076 (n2093, n1624);
buf  g2077 (n1986, n1743);
not  g2078 (n2120, n1694);
buf  g2079 (n1953, n1689);
buf  g2080 (n1894, n1747);
buf  g2081 (n1935, n1632);
buf  g2082 (n2023, n1664);
buf  g2083 (n2087, n1769);
not  g2084 (n1919, n1754);
buf  g2085 (n2239, n1649);
not  g2086 (n2146, n1635);
not  g2087 (n2291, n1702);
not  g2088 (n2334, n1637);
buf  g2089 (n2116, n1651);
buf  g2090 (n2025, n1612);
not  g2091 (n2201, n1733);
not  g2092 (n2247, n1651);
buf  g2093 (n2235, n1744);
buf  g2094 (n1938, n1756);
not  g2095 (n2063, n1706);
not  g2096 (n2218, n1722);
buf  g2097 (n2165, n1610);
not  g2098 (n1814, n1763);
buf  g2099 (n1897, n1688);
buf  g2100 (n2191, n1761);
not  g2101 (n1880, n1602);
buf  g2102 (n1837, n1800);
not  g2103 (n1833, n1767);
buf  g2104 (n2039, n1620);
not  g2105 (n2304, n1601);
buf  g2106 (n2383, n1739);
not  g2107 (n2108, n1648);
buf  g2108 (n1990, n1800);
buf  g2109 (n2020, n1708);
not  g2110 (n1989, n1678);
not  g2111 (n2269, n1757);
buf  g2112 (n2012, n1803);
not  g2113 (n1936, n1666);
not  g2114 (n2367, n1802);
buf  g2115 (n1918, n1641);
not  g2116 (n2061, n1749);
not  g2117 (n2086, n1745);
buf  g2118 (n2119, n1678);
buf  g2119 (n1963, n1626);
not  g2120 (n1917, n1618);
not  g2121 (n2326, n1624);
buf  g2122 (n1856, n1744);
not  g2123 (n1939, n1789);
not  g2124 (n2271, n1706);
buf  g2125 (n1958, n1746);
buf  g2126 (n1974, n1793);
buf  g2127 (n2037, n1659);
buf  g2128 (n2213, n1738);
not  g2129 (n2287, n1623);
not  g2130 (n2190, n1736);
not  g2131 (n2289, n1616);
not  g2132 (n2362, n1719);
buf  g2133 (n2354, n1791);
buf  g2134 (n1900, n1606);
buf  g2135 (n1983, n1692);
buf  g2136 (n1999, n1679);
not  g2137 (n1838, n1687);
buf  g2138 (n2335, n1726);
not  g2139 (n1942, n1692);
not  g2140 (n2282, n1689);
not  g2141 (n2343, n1702);
buf  g2142 (n1965, n1727);
not  g2143 (n2373, n1779);
not  g2144 (n1924, n1714);
not  g2145 (n1951, n1645);
buf  g2146 (n2319, n1791);
buf  g2147 (n2272, n1798);
buf  g2148 (n2206, n1798);
not  g2149 (n2355, n1607);
buf  g2150 (n2245, n1763);
not  g2151 (n2382, n1676);
not  g2152 (n1988, n1668);
buf  g2153 (n1855, n1716);
buf  g2154 (n2313, n1661);
buf  g2155 (n2064, n1731);
not  g2156 (n2345, n1650);
not  g2157 (n2051, n1657);
not  g2158 (n1967, n1654);
not  g2159 (n1872, n1682);
buf  g2160 (n2194, n1680);
buf  g2161 (n2236, n1663);
not  g2162 (n2079, n1657);
not  g2163 (n1847, n1701);
not  g2164 (n2153, n1708);
not  g2165 (n2255, n1712);
not  g2166 (n2348, n1642);
buf  g2167 (n2339, n1796);
not  g2168 (n2082, n1604);
not  g2169 (n1816, n1679);
not  g2170 (n2379, n1605);
buf  g2171 (n2055, n1653);
buf  g2172 (n1927, n1667);
buf  g2173 (n2176, n1635);
not  g2174 (n2222, n1695);
not  g2175 (n2349, n1697);
not  g2176 (n2217, n1618);
not  g2177 (n2068, n1685);
not  g2178 (n2181, n1764);
not  g2179 (n2284, n1773);
not  g2180 (n1829, n1607);
buf  g2181 (n2200, n1634);
buf  g2182 (n1975, n1656);
buf  g2183 (n2369, n1752);
buf  g2184 (n2000, n1710);
not  g2185 (n2024, n1664);
not  g2186 (n2081, n1654);
buf  g2187 (n2118, n1783);
not  g2188 (n1906, n1633);
buf  g2189 (n1868, n1643);
buf  g2190 (n1915, n1669);
not  g2191 (n1860, n1725);
buf  g2192 (n1991, n1604);
not  g2193 (n2124, n1653);
not  g2194 (n1959, n1660);
buf  g2195 (n1960, n1784);
not  g2196 (n2212, n1801);
buf  g2197 (n2356, n1802);
buf  g2198 (n1987, n1750);
not  g2199 (n1875, n1707);
buf  g2200 (n1854, n1622);
buf  g2201 (n1955, n1613);
not  g2202 (n2022, n1637);
buf  g2203 (n2363, n1742);
not  g2204 (n2158, n1607);
not  g2205 (n1948, n1722);
not  g2206 (n1947, n1615);
buf  g2207 (n1932, n1743);
buf  g2208 (n1809, n1711);
not  g2209 (n1901, n1622);
not  g2210 (n2029, n1784);
not  g2211 (n1949, n1777);
not  g2212 (n2378, n1774);
buf  g2213 (n2320, n1718);
not  g2214 (n2280, n1796);
buf  g2215 (n2196, n1632);
not  g2216 (n1889, n1771);
buf  g2217 (n2073, n1740);
not  g2218 (n2183, n1609);
buf  g2219 (n1970, n1787);
buf  g2220 (n1842, n1757);
not  g2221 (n1836, n1681);
buf  g2222 (n2202, n1762);
not  g2223 (n1916, n1658);
buf  g2224 (n2009, n1627);
buf  g2225 (n1964, n1705);
not  g2226 (n2208, n1601);
buf  g2227 (n2224, n1616);
not  g2228 (n1973, n1778);
not  g2229 (n2275, n1697);
not  g2230 (n1979, n1680);
not  g2231 (n2286, n1728);
not  g2232 (n2240, n1674);
not  g2233 (n2336, n1675);
not  g2234 (n1812, n1719);
not  g2235 (n2154, n1713);
buf  g2236 (n1968, n1739);
not  g2237 (n2365, n1796);
buf  g2238 (n2337, n1789);
not  g2239 (n2048, n1717);
buf  g2240 (n2162, n1608);
buf  g2241 (n2083, n1770);
not  g2242 (n1858, n1804);
buf  g2243 (n2072, n1692);
buf  g2244 (n2013, n1744);
not  g2245 (n1821, n1720);
buf  g2246 (n2317, n1805);
not  g2247 (n2043, n1790);
not  g2248 (n2268, n1775);
not  g2249 (n2130, n1786);
buf  g2250 (n1813, n1704);
not  g2251 (n2352, n1621);
not  g2252 (n2198, n1664);
not  g2253 (n1871, n1653);
not  g2254 (n2125, n1722);
buf  g2255 (n2143, n1653);
not  g2256 (n2033, n1617);
not  g2257 (n2151, n1702);
buf  g2258 (n2150, n1761);
not  g2259 (n2231, n1623);
not  g2260 (n2026, n1712);
buf  g2261 (n2308, n1703);
buf  g2262 (n2210, n1785);
xnor g2263 (n2259, n1609, n1613, n1684, n1805);
nand g2264 (n2015, n1700, n1707, n1494, n1657);
and  g2265 (n2364, n1780, n1495, n1726, n1803);
or   g2266 (n2246, n1661, n1688, n1654);
and  g2267 (n2075, n1753, n1786, n1740, n1700);
xor  g2268 (n2195, n1734, n1671, n1619, n1700);
nand g2269 (n2301, n1708, n1808, n1755, n1769);
nor  g2270 (n2193, n1808, n1662, n1645, n1677);
and  g2271 (n2041, n1716, n1672, n1723, n1804);
or   g2272 (n2173, n1638, n1808, n1701, n1794);
xnor g2273 (n2095, n1698, n1627, n1799, n1682);
nand g2274 (n2234, n1797, n1758, n1775, n1676);
xor  g2275 (n2226, n1759, n1745, n1741, n1610);
nand g2276 (n2052, n1661, n1760, n1685, n1624);
xor  g2277 (n2241, n1742, n1634, n1635, n1800);
xnor g2278 (n2179, n1688, n1733, n1693, n1658);
and  g2279 (n2299, n1633, n1790, n1800, n1629);
xor  g2280 (n2129, n1696, n1697, n1744, n1615);
and  g2281 (n1978, n1761, n1747, n1771, n1694);
xor  g2282 (n1828, n1793, n1611, n1635, n1705);
xnor g2283 (n2204, n1647, n1704, n1730, n1618);
nor  g2284 (n2071, n1682, n1713, n1650, n1773);
and  g2285 (n2067, n1628, n1758, n1614, n1799);
xnor g2286 (n1956, n1768, n1778, n1640, n1698);
and  g2287 (n2066, n1672, n1747, n1753, n1795);
nor  g2288 (n1881, n1791, n1721, n1626, n1713);
nand g2289 (n2109, n1704, n1641, n1495, n1628);
or   g2290 (n2059, n1601, n1656, n1643, n1755);
or   g2291 (n2133, n1639, n1672, n1634, n1679);
xnor g2292 (n2254, n1762, n1786, n1612, n1771);
or   g2293 (n2005, n1799, n1604, n1764, n1788);
nand g2294 (n2332, n1759, n1693, n1610, n1803);
xor  g2295 (n2258, n1654, n1641, n1719, n1696);
xnor g2296 (n2157, n1782, n1705, n1769, n1707);
nand g2297 (n2228, n1738, n1730, n1689, n1754);
xnor g2298 (n1930, n1650, n1720, n1725, n1659);
or   g2299 (n1822, n1670, n1727, n1644, n1657);
xnor g2300 (n2325, n1637, n1605, n1642, n1611);
nand g2301 (n2144, n1766, n1611, n1765, n1782);
nor  g2302 (n2361, n1671, n1602, n1736, n1700);
nand g2303 (n2303, n1716, n1732, n1779, n1665);
and  g2304 (n2166, n1701, n1647, n1731, n1677);
nor  g2305 (n1946, n1723, n1621, n1683, n1735);
or   g2306 (n2088, n1750, n1609, n1642, n1652);
xor  g2307 (n2186, n1749, n1784, n1627, n1797);
nand g2308 (n2149, n1692, n1729, n1698, n1735);
xnor g2309 (n1867, n1652, n1615, n1608, n1710);
xor  g2310 (n2045, n1660, n1721, n1733, n1645);
and  g2311 (n2132, n1731, n1751, n1753, n1680);
or   g2312 (n1877, n1687, n1703, n1787, n1669);
xnor g2313 (n1830, n1737, n1742, n1752, n1494);
and  g2314 (n2372, n1648, n1749, n1633, n1803);
xor  g2315 (n1997, n1782, n1785, n1786, n1760);
or   g2316 (n1832, n1740, n1614, n1790, n1717);
xor  g2317 (n2329, n1739, n1732, n1625, n1623);
or   g2318 (n2302, n1796, n1645, n1683, n1718);
xor  g2319 (n1995, n1706, n1717, n1783, n1686);
xnor g2320 (n1839, n1759, n1777, n1639, n1681);
nand g2321 (n1825, n1731, n1769, n1620, n1725);
xnor g2322 (n2126, n1659, n1662, n1729, n1691);
or   g2323 (n1876, n1718, n1798, n1647, n1770);
xnor g2324 (n2199, n1712, n1708, n1767, n1697);
xor  g2325 (n2112, n1773, n1616, n1808, n1714);
and  g2326 (n1843, n1737, n1698, n1780, n1806);
xnor g2327 (n2265, n1690, n1687, n1713, n1631);
nand g2328 (n2232, n1674, n1801, n1751, n1670);
nor  g2329 (n1908, n1640, n1669, n1802, n1703);
and  g2330 (n2295, n1631, n1613, n1626);
xnor g2331 (n2307, n1676, n1660, n1652, n1757);
nand g2332 (n2056, n1675, n1605, n1754, n1699);
xnor g2333 (n2357, n1703, n1631, n1633, n1614);
and  g2334 (n2300, n1780, n1774, n1709, n1741);
xor  g2335 (n1957, n1797, n1665, n1779, n1617);
and  g2336 (n2351, n1663, n1710, n1795, n1772);
or   g2337 (n2184, n1695, n1729, n1783, n1781);
xor  g2338 (n2380, n1605, n1759, n1693, n1775);
nor  g2339 (n1929, n1794, n1756, n1720, n1643);
or   g2340 (n2187, n1651, n1807, n1764, n1680);
nor  g2341 (n2323, n1670, n1694, n1649, n1807);
xnor g2342 (n2221, n1636, n1662, n1735, n1625);
xnor g2343 (n2377, n1696, n1734, n1717, n1699);
and  g2344 (n2101, n1686, n1711, n1789, n1612);
and  g2345 (n1910, n1772, n1727, n1630, n1738);
xnor g2346 (n2376, n1755, n1616, n1718, n1686);
xnor g2347 (n2374, n1736, n1802, n1733, n1666);
xor  g2348 (n1993, n1675, n1632, n1683, n1734);
nor  g2349 (n2305, n1766, n1629, n1710, n1609);
nand g2350 (n2078, n1671, n1709, n1795, n1668);
and  g2351 (n2495, n2210, n1838, n1945, n2181);
nand g2352 (n2443, n1987, n2342, n2308, n2171);
nand g2353 (n2388, n2080, n2045, n1990, n2085);
xor  g2354 (n2561, n2170, n1995, n2275, n2050);
or   g2355 (n2488, n2321, n2262, n2309, n1973);
and  g2356 (n2420, n2278, n2355, n2037, n2146);
or   g2357 (n2585, n1823, n1912, n2254, n2202);
and  g2358 (n2427, n2359, n2169, n2086, n2082);
xor  g2359 (n2541, n2326, n2336, n2292, n1937);
xnor g2360 (n2515, n2047, n2214, n2111, n1989);
xnor g2361 (n2554, n2182, n2168, n2293, n2268);
and  g2362 (n2481, n1870, n2230, n2134, n2255);
xor  g2363 (n2456, n2006, n2160, n2204, n2180);
nand g2364 (n2405, n2215, n2314, n2216, n2284);
xor  g2365 (n2549, n2228, n2157, n2295, n2294);
and  g2366 (n2398, n1896, n2126, n2360, n2075);
xor  g2367 (n2417, n2288, n2218, n2090, n2344);
xnor g2368 (n2499, n1891, n2235, n2145, n2194);
or   g2369 (n2565, n2361, n2356, n1983, n1934);
or   g2370 (n2451, n2128, n1956, n2274, n2163);
nor  g2371 (n2454, n2276, n2107, n2296, n2188);
nor  g2372 (n2513, n2277, n2265, n2186, n1910);
nand g2373 (n2446, n2341, n2265, n2191, n2288);
nor  g2374 (n2489, n2089, n2201, n2254, n2085);
xnor g2375 (n2544, n2312, n2325, n1994, n2327);
xnor g2376 (n2396, n2334, n1841, n2026, n1924);
and  g2377 (n2466, n2173, n1890, n2305, n2055);
nand g2378 (n2505, n1913, n2348, n2116, n2337);
xor  g2379 (n2556, n2034, n2137, n2226, n2328);
and  g2380 (n2385, n2078, n2205, n2190, n2120);
or   g2381 (n2453, n1970, n2202, n2149, n1862);
xor  g2382 (n2403, n2287, n2358, n2255, n1820);
nand g2383 (n2461, n1878, n1980, n2244, n2191);
nor  g2384 (n2529, n2290, n2118, n2147, n2151);
and  g2385 (n2416, n2101, n2269, n1968, n2276);
xor  g2386 (n2412, n2156, n1887, n2100, n2221);
nand g2387 (n2389, n2271, n2308, n2115, n2131);
xor  g2388 (n2437, n2187, n2148, n1986, n1926);
xor  g2389 (n2525, n2110, n2220, n1984, n1822);
xor  g2390 (n2479, n2302, n1837, n2014, n2063);
nor  g2391 (n2474, n2186, n2043, n1908, n1828);
and  g2392 (n2575, n1825, n2246, n2136, n1849);
nor  g2393 (n2587, n2183, n2062, n2230, n2135);
nand g2394 (n2462, n1900, n1819, n2140, n1836);
xor  g2395 (n2573, n2168, n2198, n2227, n2209);
xnor g2396 (n2586, n2263, n2017, n1954, n2097);
nor  g2397 (n2480, n1875, n2133, n2121, n1907);
nor  g2398 (n2563, n2253, n2099, n1960, n1903);
and  g2399 (n2524, n2112, n2155, n2015, n2243);
nand g2400 (n2478, n2259, n2301, n2176, n2125);
xor  g2401 (n2472, n2077, n2005, n2028, n2161);
nor  g2402 (n2557, n1949, n2183, n2358, n2256);
nor  g2403 (n2533, n1917, n1873, n1948, n2101);
xor  g2404 (n2387, n2356, n2152, n1932, n2172);
xor  g2405 (n2476, n1978, n1943, n2088, n2149);
and  g2406 (n2506, n2161, n2221, n2318, n2353);
nor  g2407 (n2568, n2169, n1952, n2263, n2129);
nor  g2408 (n2564, n2162, n1893, n2330, n2136);
xor  g2409 (n2426, n2080, n2106, n2320, n2258);
and  g2410 (n2455, n2289, n1992, n2270, n2122);
or   g2411 (n2503, n2199, n2350, n2339, n2257);
xnor g2412 (n2395, n2319, n2331, n2192, n1827);
and  g2413 (n2532, n2067, n2206, n2158, n1815);
nand g2414 (n2452, n2079, n2133, n2245, n2208);
and  g2415 (n2519, n2317, n2346, n2152, n2351);
or   g2416 (n2578, n2142, n2238, n1976);
and  g2417 (n2439, n1914, n2292, n1920, n2189);
and  g2418 (n2577, n1839, n2329, n2018, n2299);
and  g2419 (n2408, n2347, n2182, n2158, n2035);
nor  g2420 (n2468, n2140, n2210, n2128, n2179);
nand g2421 (n2516, n2181, n1899, n2326, n2156);
nor  g2422 (n2401, n2009, n1911, n1957, n1824);
nor  g2423 (n2580, n2025, n2317, n2138, n2076);
nand g2424 (n2440, n2040, n2195, n2150, n2021);
nor  g2425 (n2393, n2041, n1946, n2159, n2125);
xor  g2426 (n2402, n2096, n1919, n2144, n2245);
nand g2427 (n2407, n1951, n2341, n2170, n2222);
nor  g2428 (n2491, n2258, n1940, n2273, n2131);
and  g2429 (n2507, n2344, n2323, n2081, n2331);
nand g2430 (n2566, n2348, n2298, n1826, n2165);
xor  g2431 (n2435, n2357, n1857, n1889, n2108);
xor  g2432 (n2404, n2240, n2004, n2218, n1982);
or   g2433 (n2444, n2196, n1964, n2316, n1821);
xor  g2434 (n2477, n2173, n2211, n2212, n2209);
nor  g2435 (n2409, n2077, n1996, n2082, n2338);
xnor g2436 (n2588, n2109, n2114, n2307, n2283);
or   g2437 (n2501, n2232, n1999, n2318, n2117);
nor  g2438 (n2482, n1866, n1988, n1835, n1953);
xnor g2439 (n2540, n2180, n2030, n2242, n2144);
nand g2440 (n2530, n1901, n2330, n1955, n2219);
xor  g2441 (n2460, n2162, n2234, n2197, n1981);
nor  g2442 (n2464, n2075, n2112, n1869, n1929);
nor  g2443 (n2422, n2332, n2095, n1925, n1985);
xnor g2444 (n2433, n2281, n2360, n2102, n2118);
nand g2445 (n2441, n2247, n2086, n2165, n2175);
and  g2446 (n2560, n2220, n2107, n2244, n2307);
xnor g2447 (n2527, n1892, n2066, n1856, n2184);
nand g2448 (n2411, n2290, n2332, n2334, n2146);
xor  g2449 (n2486, n2349, n2324, n2248, n2363);
xnor g2450 (n2421, n2325, n2365, n2232, n1833);
xnor g2451 (n2591, n2148, n1977, n2108, n2257);
xor  g2452 (n2518, n2088, n2123, n2310, n2083);
xnor g2453 (n2509, n2203, n1923, n2306, n2011);
nor  g2454 (n2429, n2100, n2294, n2225, n2293);
nand g2455 (n2579, n2003, n2224, n2147, n2177);
and  g2456 (n2448, n1814, n2083, n2189, n1832);
xnor g2457 (n2418, n2187, n1867, n1885, n2116);
xor  g2458 (n2490, n1905, n2250, n2121, n2321);
xor  g2459 (n2553, n2188, n2247, n2104, n1935);
or   g2460 (n2559, n1927, n2207, n2231, n2167);
or   g2461 (n2582, n1939, n2279, n2340, n2145);
or   g2462 (n2457, n2091, n2057, n2051, n2105);
or   g2463 (n2494, n1897, n2184, n1931, n2058);
xor  g2464 (n2425, n2038, n1997, n1854, n1902);
and  g2465 (n2517, n2000, n2216, n2022, n2241);
xor  g2466 (n2526, n2251, n2282, n2027, n2239);
or   g2467 (n2595, n2127, n2124, n2020, n2343);
xor  g2468 (n2465, n2223, n2235, n2090, n2260);
and  g2469 (n2500, n2081, n2286, n2141, n2093);
xnor g2470 (n2423, n2355, n1872, n2319, n2354);
xnor g2471 (n2546, n2142, n2291, n2249, n2141);
xor  g2472 (n2391, n1941, n2217, n2163, n1816);
xor  g2473 (n2576, n2032, n1846, n1962, n2102);
xnor g2474 (n2569, n2060, n2124, n2347, n2266);
and  g2475 (n2543, n2059, n2091, n2335, n2049);
or   g2476 (n2535, n2048, n2069, n1936, n2272);
xnor g2477 (n2434, n1898, n2214, n1906, n1852);
nand g2478 (n2548, n2110, n1847, n2073, n1969);
nor  g2479 (n2400, n2013, n1991, n2164, n2333);
and  g2480 (n2583, n1933, n2267, n1861, n2007);
or   g2481 (n2536, n2178, n2229, n2304, n2119);
nor  g2482 (n2463, n2064, n1883, n2300, n2094);
nor  g2483 (n2534, n2179, n2284, n2260, n2196);
nor  g2484 (n2550, n2302, n2106, n1855, n2076);
xnor g2485 (n2386, n2211, n2084, n2153, n2104);
nand g2486 (n2390, n2251, n2117, n2203, n2252);
and  g2487 (n2510, n1965, n2291, n2315, n2174);
xnor g2488 (n2520, n2237, n2016, n1881, n1882);
nor  g2489 (n2410, n2193, n2310, n2249, n1812);
xor  g2490 (n2485, n2079, n1813, n2243, n2357);
and  g2491 (n2581, n2087, n1918, n2120, n1963);
nor  g2492 (n2470, n2143, n2199, n2008, n2264);
xor  g2493 (n2528, n2233, n2270, n2177, n2364);
xnor g2494 (n2496, n2296, n2217, n2264, n1817);
xor  g2495 (n2431, n1853, n1904, n2099, n2031);
xnor g2496 (n2537, n2335, n2103, n2208, n2150);
nand g2497 (n2572, n1865, n2215, n2213, n2287);
nand g2498 (n2521, n2250, n1930, n2095, n2010);
xor  g2499 (n2450, n2351, n2002, n2153, n2349);
xnor g2500 (n2504, n2139, n2143, n2042, n2023);
xnor g2501 (n2483, n1950, n2001, n2113, n1974);
xnor g2502 (n2512, n2278, n2313, n2098, n1871);
nor  g2503 (n2487, n2070, n2309, n2138, n2224);
and  g2504 (n2399, n2074, n2267, n2024, n2033);
xor  g2505 (n2592, n2094, n2333, n2345, n2092);
xor  g2506 (n2414, n1851, n2313, n2115, n2052);
and  g2507 (n2567, n2363, n2134, n1975, n2213);
xnor g2508 (n2471, n2301, n1928, n2300, n2200);
or   g2509 (n2449, n2322, n2127, n2248, n2185);
and  g2510 (n2397, n2289, n2212, n2241, n2151);
nand g2511 (n2458, n1966, n2114, n2336, n2343);
and  g2512 (n2590, n2337, n2315, n2084, n1947);
xnor g2513 (n2406, n2364, n2266, n1829, n2236);
and  g2514 (n2475, n1834, n2053, n2071, n1868);
nor  g2515 (n2545, n2338, n1967, n2353, n2029);
and  g2516 (n2469, n2275, n2231, n1809, n2253);
and  g2517 (n2547, n2039, n2154, n2362, n2192);
or   g2518 (n2508, n2159, n2297, n2119, n1886);
and  g2519 (n2523, n2303, n2365, n2185, n1848);
nor  g2520 (n2428, n2087, n2272, n2252, n2166);
or   g2521 (n2392, n2036, n1916, n2044, n2103);
and  g2522 (n2413, n2155, n2277, n2197, n1840);
and  g2523 (n2522, n2359, n1915, n1874, n2200);
nor  g2524 (n2570, n2222, n2130, n2061, n2324);
xor  g2525 (n2497, n1850, n2176, n2065, n2135);
nand g2526 (n2555, n2274, n2328, n2164, n2167);
xnor g2527 (n2438, n2236, n1938, n2228, n2195);
or   g2528 (n2430, n2172, n1979, n2194, n2280);
and  g2529 (n2419, n1880, n2154, n2056, n1864);
xnor g2530 (n2467, n2126, n2111, n2352, n2304);
nand g2531 (n2436, n1863, n2242, n2096, n2137);
nand g2532 (n2459, n1860, n2322, n2282, n2285);
nand g2533 (n2384, n1894, n2012, n1858, n1942);
or   g2534 (n2539, n2323, n2285, n2132, n2280);
xnor g2535 (n2571, n1818, n1971, n2093, n1959);
and  g2536 (n2538, n2178, n1884, n2240, n2219);
xnor g2537 (n2442, n2295, n1961, n1859, n2068);
xnor g2538 (n2424, n2097, n1888, n2098, n2246);
or   g2539 (n2473, n2190, n2054, n2362, n2129);
or   g2540 (n2492, n2311, n2340, n2329, n2072);
xnor g2541 (n2589, n2259, n2078, n1993, n2361);
xnor g2542 (n2484, n1879, n2109, n2174, n2201);
and  g2543 (n2552, n2350, n2262, n2019, n2342);
and  g2544 (n2584, n1998, n2354, n2160, n1944);
and  g2545 (n2542, n2298, n2320, n1842, n1921);
nor  g2546 (n2493, n1895, n2261, n2283, n2157);
nor  g2547 (n2511, n2256, n2206, n2286, n1831);
or   g2548 (n2432, n2227, n2303, n2198, n2204);
nand g2549 (n2558, n2089, n2312, n1845, n2352);
nand g2550 (n2502, n2233, n1909, n2092, n2225);
xor  g2551 (n2498, n1958, n1810, n2139, n2237);
nor  g2552 (n2593, n2226, n2234, n1876, n2105);
and  g2553 (n2531, n1877, n1844, n2113, n2130);
nor  g2554 (n2562, n2166, n2327, n2269, n2279);
xor  g2555 (n2594, n1922, n2345, n2205, n1972);
nand g2556 (n2394, n2268, n2299, n2046, n2339);
nor  g2557 (n2447, n2207, n2171, n2132, n2314);
xnor g2558 (n2415, n2271, n2316, n2346, n2239);
nand g2559 (n2551, n1830, n2123, n2297, n2223);
or   g2560 (n2514, n2122, n2273, n2281, n1811);
xnor g2561 (n2574, n1843, n2311, n2305, n2229);
or   g2562 (n2445, n2175, n2193, n2306, n2261);
nor  g2563 (n2608, n2486, n2453, n2415, n2424);
nor  g2564 (n2598, n2500, n2493, n2430, n2487);
and  g2565 (n2612, n2465, n2400, n2483, n2404);
or   g2566 (n2596, n2459, n2452, n2393, n2478);
nand g2567 (n2625, n2392, n2429, n2475, n2451);
xor  g2568 (n2597, n2432, n2388, n2456, n2410);
and  g2569 (n2601, n2420, n2494, n2448, n2398);
nor  g2570 (n2602, n2417, n2394, n2445, n2495);
and  g2571 (n2618, n2454, n2396, n2476, n2403);
nand g2572 (n2609, n2499, n2458, n2413, n2435);
or   g2573 (n2616, n2480, n2431, n2385, n2389);
or   g2574 (n2611, n2390, n2472, n2440, n2473);
or   g2575 (n2617, n2443, n2491, n2479, n2399);
xor  g2576 (n2606, n2488, n2426, n2391, n2497);
xor  g2577 (n2599, n2409, n2384, n2464, n2418);
nand g2578 (n2600, n2484, n2423, n2407, n2433);
or   g2579 (n2622, n2462, n2466, n2455, n2439);
or   g2580 (n2623, n2419, n2470, n2427, n2397);
xnor g2581 (n2607, n2490, n2450, n2469, n2411);
or   g2582 (n2604, n2447, n2401, n2405, n2498);
and  g2583 (n2610, n2428, n2449, n2460, n2422);
xnor g2584 (n2615, n2485, n2461, n2442, n2395);
xor  g2585 (n2624, n2416, n2503, n2437, n2482);
xnor g2586 (n2605, n2434, n2502, n2408, n2444);
nor  g2587 (n2614, n2387, n2406, n2441, n2474);
nand g2588 (n2613, n2438, n2457, n2412, n2468);
or   g2589 (n2621, n2467, n2436, n2481, n2492);
xnor g2590 (n2619, n2425, n2402, n2489, n2446);
xor  g2591 (n2620, n2496, n2386, n2463, n2477);
xnor g2592 (n2603, n2471, n2414, n2421, n2501);
buf  g2593 (n2630, n1299);
buf  g2594 (n2635, n1303);
buf  g2595 (n2632, n2606);
not  g2596 (n2627, n2599);
not  g2597 (n2631, n1298);
buf  g2598 (n2639, n2599);
buf  g2599 (n2626, n2606);
not  g2600 (n2633, n2600);
buf  g2601 (n2628, n1304);
not  g2602 (n2629, n2597);
nand g2603 (n2634, n1310, n1305);
xor  g2604 (n2637, n2596, n2601, n1307, n1300);
xor  g2605 (n2636, n2597, n2601, n2596, n2600);
and  g2606 (n2642, n2602, n2604, n1301, n1308);
xnor g2607 (n2638, n2603, n1302, n2605);
and  g2608 (n2641, n2602, n2603, n2604, n2598);
nor  g2609 (n2640, n1306, n1297, n2598, n1309);
not  g2610 (n2661, n2370);
buf  g2611 (n2650, n2628);
not  g2612 (n2651, n2374);
not  g2613 (n2662, n2630);
buf  g2614 (n2649, n2633);
buf  g2615 (n2669, n2639);
buf  g2616 (n2664, n2627);
buf  g2617 (n2659, n2369);
buf  g2618 (n2652, n2631);
buf  g2619 (n2665, n2373);
buf  g2620 (n2660, n2636);
not  g2621 (n2667, n2368);
buf  g2622 (n2668, n2375);
buf  g2623 (n2671, n2638);
buf  g2624 (n2653, n2631);
not  g2625 (n2656, n2376);
not  g2626 (n2644, n2639);
nand g2627 (n2647, n2381, n2628, n2635);
xor  g2628 (n2658, n2627, n2374, n2634, n2369);
and  g2629 (n2643, n2626, n2383, n2382, n2367);
and  g2630 (n2648, n2378, n2640, n2379, n2634);
or   g2631 (n2663, n2373, n2371, n2368);
nand g2632 (n2666, n2630, n2378, n2629, n2638);
nor  g2633 (n2655, n2626, n2629, n2366, n2632);
xor  g2634 (n2670, n2370, n2372, n2366, n2367);
or   g2635 (n2657, n2377, n2380, n2372, n2636);
xnor g2636 (n2645, n2376, n2379, n2375, n2377);
xnor g2637 (n2654, n2633, n2637, n2632);
nand g2638 (n2646, n2382, n2381, n2635, n2380);
and  g2639 (n2688, n2566, n2576, n2573, n2578);
and  g2640 (n2679, n2648, n2518, n2587, n2519);
nor  g2641 (n2692, n2570, n2582, n2544, n2569);
nand g2642 (n2691, n2555, n2530, n2577, n2644);
nor  g2643 (n2676, n2539, n2564, n2644, n2532);
or   g2644 (n2699, n2552, n2512, n2549, n2560);
xor  g2645 (n2693, n2507, n2643, n2648, n2529);
and  g2646 (n2685, n2551, n2545, n2646);
xor  g2647 (n2694, n2649, n2647, n2583, n2585);
and  g2648 (n2681, n2568, n2649, n2556, n2504);
and  g2649 (n2690, n2575, n2645, n2580, n2584);
nor  g2650 (n2683, n2644, n2557, n2579, n2536);
nand g2651 (n2677, n2644, n2517, n2533, n2506);
xnor g2652 (n2689, n2572, n2565, n2510, n2650);
xnor g2653 (n2680, n2515, n2646, n2521, n2650);
nand g2654 (n2696, n2647, n2561, n2531, n2540);
xor  g2655 (n2672, n2505, n2514, n2527, n2534);
or   g2656 (n2686, n2550, n2535, n2538, n2649);
and  g2657 (n2698, n2523, n2649, n2558, n2516);
nand g2658 (n2678, n2646, n2647, n2548, n2645);
xor  g2659 (n2675, n2547, n2528, n2559, n2525);
and  g2660 (n2684, n2645, n2520, n2542, n2511);
xor  g2661 (n2695, n2522, n2571, n2581, n2537);
xor  g2662 (n2682, n2643, n2567, n2563, n2562);
and  g2663 (n2673, n2543, n2554, n2524, n2648);
or   g2664 (n2687, n2648, n2553, n2574, n2645);
and  g2665 (n2697, n2513, n2509, n2546, n2508);
or   g2666 (n2674, n2541, n2526, n2586, n2647);
not  g2667 (n2701, n2609);
buf  g2668 (n2718, n2675);
not  g2669 (n2710, n2675);
buf  g2670 (n2720, n2676);
not  g2671 (n2714, n2679);
not  g2672 (n2702, n953);
buf  g2673 (n2729, n2617);
buf  g2674 (n2723, n953);
buf  g2675 (n2728, n2678);
not  g2676 (n2713, n954);
not  g2677 (n2700, n2673);
buf  g2678 (n2706, n2675);
buf  g2679 (n2705, n2613);
xor  g2680 (n2704, n2676, n2621, n2607);
or   g2681 (n2707, n954, n2612, n2676, n2614);
xor  g2682 (n2722, n952, n2608, n2624, n2622);
or   g2683 (n2709, n2611, n2619, n2622, n2610);
and  g2684 (n2703, n2608, n2676, n2674, n2625);
and  g2685 (n2727, n2617, n2673, n2677, n2678);
xnor g2686 (n2715, n2672, n2674, n952);
xnor g2687 (n2726, n2672, n2621, n2619, n2674);
xor  g2688 (n2712, n2678, n2677, n2672, n2615);
or   g2689 (n2721, n2610, n2624, n2609, n953);
xor  g2690 (n2724, n2620, n2677, n2613, n953);
nand g2691 (n2711, n2677, n2675, n954, n2673);
xor  g2692 (n2708, n2672, n2611, n2678, n2383);
xnor g2693 (n2725, n2673, n2620, n2679, n2616);
xnor g2694 (n2716, n2625, n2623, n2616, n2615);
xnor g2695 (n2719, n2623, n2607, n954, n2674);
xnor g2696 (n2717, n2618, n2618, n2612, n2614);
nor  g2697 (n2738, n2722, n2714, n2721, n2704);
nor  g2698 (n2742, n2709, n2713, n2710, n2719);
nor  g2699 (n2732, n2722, n2700, n2716, n2706);
xnor g2700 (n2741, n2713, n2718, n2705);
xnor g2701 (n2737, n2716, n2707, n2717, n2703);
nand g2702 (n2731, n2720, n2724, n2721, n2711);
nand g2703 (n2740, n2701, n2706, n2708, n2717);
or   g2704 (n2730, n2724, n2719, n2714, n2704);
nor  g2705 (n2736, n2725, n2725, n2709, n2720);
xnor g2706 (n2735, n2705, n2703, n2701, n2708);
nand g2707 (n2733, n2707, n2700, n2712);
nand g2708 (n2734, n2711, n2715, n2723, n2702);
and  g2709 (n2739, n2715, n2702, n2710, n2723);
xnor g2710 (n2772, n2732, n2651, n2655);
xnor g2711 (n2783, n2731, n2737, n2654);
nor  g2712 (n2762, n2658, n2669, n2662);
and  g2713 (n2775, n2670, n2738, n2737);
xnor g2714 (n2755, n2671, n1443, n2733);
and  g2715 (n2784, n2665, n2663, n2652);
nor  g2716 (n2751, n2728, n2653, n2736);
xor  g2717 (n2753, n2668, n2656, n2732);
or   g2718 (n2757, n2656, n2736, n2671);
nor  g2719 (n2773, n2734, n2728, n1444);
nor  g2720 (n2778, n2660, n2739, n2667);
and  g2721 (n2764, n2662, n2734, n2655);
xnor g2722 (n2766, n2661, n2740, n2659);
nand g2723 (n2779, n2736, n2660);
and  g2724 (n2759, n2661, n2739, n2662);
or   g2725 (n2769, n2664, n2659, n2651, n2655);
xnor g2726 (n2768, n2666, n2742, n1445, n2741);
nand g2727 (n2748, n2657, n2653, n2665, n1314);
xor  g2728 (n2765, n2735, n1311, n2741, n2738);
xnor g2729 (n2756, n2652, n2659, n1316, n2651);
nor  g2730 (n2754, n2738, n2727, n2739);
and  g2731 (n2776, n1313, n2726, n1315, n2730);
xnor g2732 (n2781, n2742, n2731, n2737, n2730);
xnor g2733 (n2770, n2670, n2655, n1312, n1444);
nor  g2734 (n2771, n2740, n2654, n2664, n2662);
and  g2735 (n2782, n2663, n1318, n2669, n2657);
xor  g2736 (n2777, n2670, n2668, n2665, n2666);
xor  g2737 (n2746, n2671, n2651, n2741);
nor  g2738 (n2767, n1444, n2671, n2658, n2668);
nand g2739 (n2745, n2658, n2667, n2738, n2666);
and  g2740 (n2744, n2659, n2661, n2736, n2663);
and  g2741 (n2750, n2664, n2654, n2650, n1319);
xnor g2742 (n2780, n2737, n2661, n2667, n2658);
or   g2743 (n2763, n2657, n2652, n1443, n2656);
xnor g2744 (n2761, n2657, n2652, n2742, n2665);
xnor g2745 (n2743, n2669, n2668, n2650, n2654);
xor  g2746 (n2758, n2726, n2742, n2653, n1317);
xor  g2747 (n2760, n2670, n2728, n2740, n1444);
nor  g2748 (n2749, n1443, n2656, n2660, n2728);
nor  g2749 (n2752, n2740, n2669, n2735, n2664);
nand g2750 (n2774, n2666, n2653, n2735);
xor  g2751 (n2747, n2667, n2739, n2733, n2663);
not  g2752 (n2835, n1461);
buf  g2753 (n2846, n1449);
buf  g2754 (n2898, n2776);
buf  g2755 (n2848, n2764);
not  g2756 (n2852, n1466);
buf  g2757 (n2873, n2754);
not  g2758 (n2795, n2683);
not  g2759 (n2786, n279);
buf  g2760 (n2804, n1457);
not  g2761 (n2794, n1323);
not  g2762 (n2792, n280);
not  g2763 (n2829, n2692);
not  g2764 (n2808, n1465);
not  g2765 (n2904, n2691);
buf  g2766 (n2907, n1459);
buf  g2767 (n2840, n955);
not  g2768 (n2915, n2762);
not  g2769 (n2796, n2745);
buf  g2770 (n2789, n1330);
buf  g2771 (n2924, n1455);
not  g2772 (n2875, n2595);
not  g2773 (n2809, n1334);
not  g2774 (n2903, n1449);
not  g2775 (n2879, n2780);
not  g2776 (n2860, n2695);
buf  g2777 (n2928, n2697);
not  g2778 (n2891, n2699);
not  g2779 (n2830, n2697);
buf  g2780 (n2921, n2684);
buf  g2781 (n2871, n2687);
buf  g2782 (n2837, n1460);
buf  g2783 (n2853, n1333);
buf  g2784 (n2895, n2774);
buf  g2785 (n2888, n2592);
not  g2786 (n2925, n2696);
buf  g2787 (n2920, n2748);
buf  g2788 (n2845, n80);
buf  g2789 (n2843, n1465);
buf  g2790 (n2831, n1445);
buf  g2791 (n2896, n956);
not  g2792 (n2785, n1464);
not  g2793 (n2934, n2753);
buf  g2794 (n2803, n2773);
buf  g2795 (n2890, n2771);
not  g2796 (n2844, n2746);
buf  g2797 (n2828, n2690);
not  g2798 (n2824, n2783);
buf  g2799 (n2936, n2749);
buf  g2800 (n2814, n2745);
buf  g2801 (n2857, n2772);
buf  g2802 (n2894, n1458);
not  g2803 (n2790, n2761);
buf  g2804 (n2869, n2695);
buf  g2805 (n2849, n278);
not  g2806 (n2821, n2589);
not  g2807 (n2932, n2759);
buf  g2808 (n2851, n2688);
buf  g2809 (n2923, n2697);
buf  g2810 (n2867, n1458);
not  g2811 (n2862, n1456);
buf  g2812 (n2842, n2684);
buf  g2813 (n2818, n2777);
not  g2814 (n2900, n1446);
buf  g2815 (n2834, n277);
xnor g2816 (n2820, n2750, n1454, n1464, n277);
xor  g2817 (n2816, n2754, n2779, n2784, n80);
xnor g2818 (n2905, n1451, n1451, n2744, n1448);
or   g2819 (n2791, n2688, n2778, n956, n1455);
xnor g2820 (n2897, n1324, n2691, n2760, n80);
and  g2821 (n2931, n2757, n2692, n2694, n1466);
nor  g2822 (n2918, n2779, n1331, n2640, n2686);
and  g2823 (n2870, n2756, n2782, n957, n2774);
xnor g2824 (n2807, n2767, n2752, n1454, n1456);
nand g2825 (n2832, n1451, n2686, n956, n2757);
nand g2826 (n2910, n276, n2755, n2691);
or   g2827 (n2864, n1446, n2688, n2764, n2689);
or   g2828 (n2926, n2743, n2761, n1366, n1328);
nor  g2829 (n2806, n2641, n2764, n2753, n278);
or   g2830 (n2868, n2766, n2762, n2768, n1320);
or   g2831 (n2911, n2759, n2683, n1464, n1450);
nor  g2832 (n2863, n2777, n2780, n2753, n2771);
xor  g2833 (n2854, n2755, n2593, n1366, n2685);
nand g2834 (n2788, n2683, n2695, n2776, n278);
nand g2835 (n2839, n2768, n2699, n957, n1464);
or   g2836 (n2901, n2698, n2748, n277, n2757);
or   g2837 (n2819, n81, n280, n2751, n2763);
xor  g2838 (n2793, n2749, n2767, n955, n2692);
nand g2839 (n2880, n281, n2681, n2784, n2754);
xnor g2840 (n2865, n1326, n1452, n2679, n2747);
xnor g2841 (n2906, n1459, n2763, n2699, n2783);
xor  g2842 (n2817, n1332, n2686, n2689, n2773);
and  g2843 (n2855, n2755, n2681, n2770, n2747);
and  g2844 (n2833, n1321, n1462, n1446, n2642);
xnor g2845 (n2876, n2760, n2746, n2590, n2745);
xnor g2846 (n2877, n2689, n2775, n2758, n1449);
or   g2847 (n2935, n2763, n1460, n1322, n2744);
xnor g2848 (n2927, n2765, n2680, n2761, n958);
xnor g2849 (n2885, n1463, n82, n2699, n2745);
xnor g2850 (n2799, n2782, n1463, n1446, n2784);
or   g2851 (n2850, n1447, n2766, n1450, n1458);
xnor g2852 (n2827, n2682, n1447, n1366, n2743);
xnor g2853 (n2859, n2778, n958, n2756, n280);
or   g2854 (n2823, n1463, n2693, n2774, n2766);
xor  g2855 (n2914, n1451, n1459, n2750, n2772);
and  g2856 (n2913, n2777, n1457, n2697, n279);
or   g2857 (n2797, n1465, n2780, n2778, n2694);
and  g2858 (n2893, n2747, n2779, n1366, n1462);
or   g2859 (n2919, n2751, n2775, n2750, n2769);
xor  g2860 (n2902, n1452, n1453, n2783, n2758);
nand g2861 (n2882, n279, n2779, n2769, n276);
xnor g2862 (n2922, n958, n2698, n2781, n2690);
xor  g2863 (n2874, n2772, n1450, n2641, n2680);
xor  g2864 (n2802, n2771, n2756, n955, n2744);
and  g2865 (n2841, n1457, n2769, n1455, n2770);
nand g2866 (n2847, n276, n2750, n2759, n1448);
or   g2867 (n2825, n1463, n2696, n1462);
nand g2868 (n2822, n2762, n2692, n2755, n2684);
and  g2869 (n2826, n80, n2758, n2698, n1448);
and  g2870 (n2892, n2681, n1452, n2693, n2680);
xor  g2871 (n2798, n2749, n957, n2751, n1453);
nand g2872 (n2856, n1465, n956, n2694, n2772);
or   g2873 (n2858, n2774, n2743, n1447);
and  g2874 (n2912, n2749, n2758, n1459, n2729);
nand g2875 (n2812, n2679, n2782, n1456, n2698);
nor  g2876 (n2861, n1460, n1457, n2748, n1461);
or   g2877 (n2787, n2767, n2773, n2687, n2680);
xor  g2878 (n2889, n2729, n2770, n1461, n2682);
xor  g2879 (n2930, n280, n2761, n1455, n2773);
nand g2880 (n2933, n2684, n2765, n2759, n1454);
xnor g2881 (n2800, n1325, n1449, n2762, n2696);
nand g2882 (n2884, n958, n2752, n2757, n81);
nor  g2883 (n2916, n81, n277, n1466, n1462);
xor  g2884 (n2838, n2746, n2766, n2771, n2690);
or   g2885 (n2811, n1453, n2687, n2683, n2686);
nor  g2886 (n2908, n2765, n1453, n81, n2770);
and  g2887 (n2866, n2642, n2765, n2694, n2682);
xor  g2888 (n2801, n1456, n2780, n2695, n957);
xnor g2889 (n2929, n2744, n1445, n1447, n2776);
or   g2890 (n2917, n1452, n2775, n2748);
or   g2891 (n2881, n2776, n1461, n2752, n2693);
or   g2892 (n2899, n2781, n2769, n2682, n2688);
and  g2893 (n2815, n2767, n2782, n2756, n1448);
nor  g2894 (n2887, n2746, n2752, n2591, n2693);
nor  g2895 (n2878, n2760, n2687, n1445, n1460);
or   g2896 (n2909, n2754, n2764, n1454, n1450);
xnor g2897 (n2810, n2751, n2690, n2768, n2594);
or   g2898 (n2805, n2781, n2760, n2685, n2763);
xor  g2899 (n2883, n1327, n2689, n2685, n278);
nand g2900 (n2836, n2681, n2588, n1466, n2784);
xnor g2901 (n2886, n279, n2753, n2777, n2781);
xnor g2902 (n2813, n2778, n955, n2685, n2747);
xnor g2903 (n2872, n1458, n2783, n1329, n2768);
xor  g2904 (n2954, n2799, n2813, n2847, n2901);
nor  g2905 (n2943, n2806, n2829, n2885, n2935);
nand g2906 (n2969, n2851, n2830, n2878, n2870);
xnor g2907 (n2952, n2845, n2865, n2869, n2820);
nor  g2908 (n2951, n20, n2906, n2924, n2911);
xor  g2909 (n2947, n17, n2828, n2801, n2922);
xnor g2910 (n2975, n2805, n2825, n2797, n2826);
xor  g2911 (n2966, n2900, n2792, n2863, n2816);
or   g2912 (n2979, n2796, n2929, n2867, n2852);
nor  g2913 (n2978, n2822, n2807, n2888, n2862);
xnor g2914 (n2972, n2894, n2899, n2871, n2932);
xor  g2915 (n2956, n2819, n2927, n2883, n2858);
nor  g2916 (n2942, n2926, n2872, n2884, n2785);
and  g2917 (n2941, n2879, n2896, n2890, n2902);
nand g2918 (n2948, n2930, n2912, n2925, n18);
nor  g2919 (n2959, n2920, n2812, n2895, n21);
xor  g2920 (n2945, n2877, n2892, n2891, n21);
nand g2921 (n2938, n2856, n2860, n2849, n2931);
xnor g2922 (n2939, n2841, n2903, n2889, n2843);
nand g2923 (n2971, n2848, n82, n2803, n2850);
or   g2924 (n2944, n2875, n2793, n2836, n2842);
nand g2925 (n2953, n2923, n2802, n2918, n2853);
xnor g2926 (n2940, n17, n2817, n2789, n2874);
and  g2927 (n2965, n2839, n2790, n20, n2934);
nand g2928 (n2973, n2818, n2897, n2837, n2916);
xor  g2929 (n2960, n2846, n2855, n2913, n2905);
nor  g2930 (n2955, n2919, n2873, n2810, n2834);
xnor g2931 (n2963, n20, n2787, n2910, n2886);
xnor g2932 (n2961, n19, n2887, n21, n18);
or   g2933 (n2976, n2838, n2824, n2811, n2786);
xnor g2934 (n2967, n19, n2880, n2882, n2832);
and  g2935 (n2950, n2933, n2840, n2904, n2808);
nand g2936 (n2968, n2893, n2936, n2833, n2794);
xnor g2937 (n2974, n2791, n2917, n2831, n2914);
or   g2938 (n2949, n18, n2815, n2729, n2876);
nand g2939 (n2937, n2798, n18, n2907, n2835);
or   g2940 (n2958, n2868, n2821, n2844, n2800);
and  g2941 (n2946, n2827, n2729, n19, n2921);
or   g2942 (n2977, n2823, n2864, n2908, n19);
nor  g2943 (n2962, n20, n2909, n2928, n2809);
xor  g2944 (n2964, n2795, n2788, n2814, n2854);
xnor g2945 (n2957, n2881, n2804, n2857, n2861);
xor  g2946 (n2970, n2915, n2898, n2859, n2866);
xnor g2947 (n2981, n2975, n2958, n2968, n2944);
xor  g2948 (n2985, n2963, n2964, n2969, n2962);
xnor g2949 (n2984, n2938, n2959, n2945, n2965);
nor  g2950 (n2983, n2941, n2951, n2947, n2956);
nor  g2951 (n2980, n2967, n2943, n2955, n2960);
or   g2952 (n2986, n2949, n2937, n2950, n2952);
or   g2953 (n2988, n2954, n2948, n2976, n2972);
or   g2954 (n2982, n2961, n2940, n2939, n2953);
xor  g2955 (n2987, n2971, n2970, n2957, n2973);
nor  g2956 (n2989, n2966, n2946, n2942, n2974);
or   g2957 (n2990, n2989, n281);
xor  g2958 (n2992, n961, n960);
nor  g2959 (n2991, n959, n2990, n961);
xnor g2960 (n2994, n2990, n959);
and  g2961 (n2993, n961, n961, n2990, n960);
nand g2962 (n2997, n2992, n27, n2991, n26);
or   g2963 (n2996, n25, n25, n30, n2994);
nor  g2964 (n3000, n29, n28, n27, n2993);
nor  g2965 (n3005, n32, n32, n2994, n2978);
nand g2966 (n3002, n2993, n2994, n2992, n28);
nand g2967 (n3009, n29, n26, n2992);
or   g2968 (n2999, n32, n2993, n26, n31);
or   g2969 (n3004, n2991, n27, n24);
nand g2970 (n2998, n2991, n22, n2994, n26);
and  g2971 (n3007, n32, n28, n30, n23);
xor  g2972 (n2995, n22, n24, n2993, n31);
xor  g2973 (n3010, n21, n23, n24, n22);
or   g2974 (n3003, n2991, n30, n24);
nand g2975 (n3006, n2977, n29, n23, n2979);
xor  g2976 (n3001, n31, n22, n23, n29);
and  g2977 (n3008, n31, n25, n28);
or   g2978 (n3019, n96, n3008, n2995, n86);
xor  g2979 (n3017, n83, n86, n82, n3004);
or   g2980 (n3027, n2996, n93, n83, n92);
xnor g2981 (n3026, n97, n87, n3006, n92);
nor  g2982 (n3025, n3002, n3003, n97, n82);
xor  g2983 (n3012, n2998, n93, n96, n95);
nor  g2984 (n3023, n89, n90, n98, n85);
nor  g2985 (n3015, n96, n94, n3007, n90);
nor  g2986 (n3024, n85, n91, n89, n86);
nand g2987 (n3018, n98, n90, n84, n3006);
and  g2988 (n3011, n83, n3010, n3001, n3007);
and  g2989 (n3028, n93, n84, n3005, n83);
xor  g2990 (n3020, n85, n84, n3008, n3009);
xor  g2991 (n3032, n2999, n92, n90, n84);
nor  g2992 (n3022, n87, n86, n88, n94);
nand g2993 (n3016, n91, n3005, n98, n94);
or   g2994 (n3013, n91, n95);
or   g2995 (n3029, n3010, n3009, n94, n89);
nand g2996 (n3030, n96, n93, n88, n89);
nand g2997 (n3014, n98, n87, n97);
or   g2998 (n3021, n91, n92, n2997, n85);
xnor g2999 (n3031, n3000, n88, n87);
endmodule
