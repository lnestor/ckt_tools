// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_206 written by SynthGen on 2021/04/05 11:23:25
module Stat_2000_206( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n618, n348, n286, n595, n589, n242, n402, n581,
 n428, n537, n426, n171, n433, n311, n337, n329,
 n1918, n1930, n1927, n1946, n1942, n1919, n1923, n1932,
 n1944, n1939, n1938, n1924, n1943, n1948, n1979, n2032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n618, n348, n286, n595, n589, n242, n402, n581,
 n428, n537, n426, n171, n433, n311, n337, n329,
 n1918, n1930, n1927, n1946, n1942, n1919, n1923, n1932,
 n1944, n1939, n1938, n1924, n1943, n1948, n1979, n2032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n287, n288, n289, n290, n291,
 n292, n293, n294, n295, n296, n297, n298, n299,
 n300, n301, n302, n303, n304, n305, n306, n307,
 n308, n309, n310, n312, n313, n314, n315, n316,
 n317, n318, n319, n320, n321, n322, n323, n324,
 n325, n326, n327, n328, n330, n331, n332, n333,
 n334, n335, n336, n338, n339, n340, n341, n342,
 n343, n344, n345, n346, n347, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n427, n429, n430, n431, n432, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n538, n539, n540,
 n541, n542, n543, n544, n545, n546, n547, n548,
 n549, n550, n551, n552, n553, n554, n555, n556,
 n557, n558, n559, n560, n561, n562, n563, n564,
 n565, n566, n567, n568, n569, n570, n571, n572,
 n573, n574, n575, n576, n577, n578, n579, n580,
 n582, n583, n584, n585, n586, n587, n588, n590,
 n591, n592, n593, n594, n596, n597, n598, n599,
 n600, n601, n602, n603, n604, n605, n606, n607,
 n608, n609, n610, n611, n612, n613, n614, n615,
 n616, n617, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
 n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
 n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
 n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
 n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
 n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
 n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
 n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
 n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
 n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
 n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
 n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
 n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
 n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
 n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
 n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
 n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
 n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
 n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
 n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
 n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
 n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
 n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
 n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
 n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
 n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
 n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
 n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
 n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
 n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
 n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
 n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
 n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
 n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
 n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
 n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
 n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
 n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
 n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
 n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
 n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
 n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
 n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
 n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
 n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
 n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
 n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
 n1913, n1914, n1915, n1916, n1917, n1920, n1921, n1922,
 n1925, n1926, n1928, n1929, n1931, n1933, n1934, n1935,
 n1936, n1937, n1940, n1941, n1945, n1947, n1949, n1950,
 n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
 n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
 n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
 n1975, n1976, n1977, n1978, n1980, n1981, n1982, n1983,
 n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
 n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
 n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
 n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
 n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
 n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031;

not  g0 (n44, n22);
not  g1 (n134, n19);
not  g2 (n82, n12);
not  g3 (n72, n32);
buf  g4 (n59, n8);
not  g5 (n156, n20);
not  g6 (n153, n30);
not  g7 (n62, n4);
buf  g8 (n53, n13);
buf  g9 (n151, n7);
buf  g10 (n60, n19);
buf  g11 (n78, n21);
not  g12 (n154, n11);
buf  g13 (n136, n23);
buf  g14 (n51, n19);
not  g15 (n111, n17);
buf  g16 (n104, n24);
buf  g17 (n88, n28);
buf  g18 (n108, n5);
not  g19 (n64, n2);
buf  g20 (n68, n26);
buf  g21 (n140, n7);
buf  g22 (n49, n29);
not  g23 (n145, n27);
buf  g24 (n146, n4);
not  g25 (n147, n2);
buf  g26 (n141, n13);
buf  g27 (n48, n22);
buf  g28 (n61, n18);
buf  g29 (n83, n18);
buf  g30 (n144, n10);
buf  g31 (n152, n9);
buf  g32 (n87, n21);
not  g33 (n159, n15);
not  g34 (n66, n16);
not  g35 (n122, n22);
not  g36 (n132, n3);
not  g37 (n55, n9);
buf  g38 (n69, n14);
not  g39 (n149, n4);
not  g40 (n84, n15);
not  g41 (n105, n3);
buf  g42 (n99, n30);
buf  g43 (n93, n23);
not  g44 (n112, n14);
buf  g45 (n133, n9);
not  g46 (n89, n20);
buf  g47 (n75, n18);
not  g48 (n160, n31);
buf  g49 (n125, n1);
buf  g50 (n142, n17);
not  g51 (n148, n18);
buf  g52 (n115, n2);
not  g53 (n94, n29);
buf  g54 (n98, n27);
not  g55 (n52, n13);
buf  g56 (n63, n24);
not  g57 (n54, n25);
buf  g58 (n85, n12);
buf  g59 (n33, n32);
buf  g60 (n74, n21);
not  g61 (n95, n6);
not  g62 (n114, n24);
buf  g63 (n126, n11);
buf  g64 (n129, n6);
not  g65 (n102, n31);
not  g66 (n91, n26);
buf  g67 (n120, n11);
not  g68 (n65, n8);
not  g69 (n119, n7);
buf  g70 (n41, n5);
not  g71 (n110, n16);
not  g72 (n100, n32);
not  g73 (n70, n6);
not  g74 (n113, n15);
not  g75 (n46, n20);
not  g76 (n101, n31);
buf  g77 (n34, n19);
not  g78 (n39, n1);
not  g79 (n36, n12);
buf  g80 (n155, n25);
not  g81 (n76, n10);
buf  g82 (n73, n29);
not  g83 (n35, n10);
not  g84 (n130, n1);
not  g85 (n127, n27);
not  g86 (n131, n27);
not  g87 (n81, n25);
buf  g88 (n123, n7);
not  g89 (n150, n17);
buf  g90 (n40, n1);
not  g91 (n158, n13);
buf  g92 (n137, n3);
not  g93 (n157, n26);
buf  g94 (n50, n29);
buf  g95 (n47, n30);
buf  g96 (n143, n12);
not  g97 (n71, n2);
buf  g98 (n45, n11);
not  g99 (n109, n24);
not  g100 (n67, n3);
not  g101 (n56, n16);
not  g102 (n97, n17);
buf  g103 (n79, n21);
buf  g104 (n57, n28);
buf  g105 (n80, n6);
not  g106 (n90, n30);
not  g107 (n103, n5);
buf  g108 (n38, n20);
not  g109 (n118, n31);
not  g110 (n92, n8);
buf  g111 (n121, n32);
not  g112 (n58, n22);
not  g113 (n86, n10);
not  g114 (n124, n28);
buf  g115 (n139, n14);
buf  g116 (n117, n9);
buf  g117 (n128, n14);
not  g118 (n43, n26);
not  g119 (n135, n15);
buf  g120 (n77, n5);
buf  g121 (n96, n23);
not  g122 (n138, n25);
buf  g123 (n42, n8);
buf  g124 (n37, n23);
buf  g125 (n116, n4);
buf  g126 (n107, n16);
buf  g127 (n106, n28);
buf  g128 (n618, n159);
buf  g129 (n298, n157);
not  g130 (n539, n58);
not  g131 (n548, n36);
buf  g132 (n313, n141);
buf  g133 (n317, n132);
buf  g134 (n579, n112);
buf  g135 (n216, n115);
buf  g136 (n559, n157);
not  g137 (n401, n125);
buf  g138 (n646, n140);
buf  g139 (n620, n78);
not  g140 (n188, n62);
buf  g141 (n222, n74);
buf  g142 (n501, n69);
not  g143 (n409, n71);
buf  g144 (n277, n35);
not  g145 (n197, n149);
buf  g146 (n275, n142);
not  g147 (n187, n56);
not  g148 (n206, n127);
not  g149 (n638, n136);
not  g150 (n281, n141);
buf  g151 (n371, n52);
not  g152 (n586, n150);
buf  g153 (n498, n73);
not  g154 (n502, n35);
buf  g155 (n219, n61);
buf  g156 (n358, n112);
not  g157 (n417, n84);
buf  g158 (n449, n82);
not  g159 (n228, n106);
not  g160 (n514, n98);
not  g161 (n503, n157);
not  g162 (n563, n98);
not  g163 (n360, n121);
buf  g164 (n648, n138);
not  g165 (n169, n151);
not  g166 (n198, n155);
not  g167 (n565, n111);
buf  g168 (n285, n91);
buf  g169 (n609, n96);
not  g170 (n259, n155);
not  g171 (n348, n53);
buf  g172 (n413, n119);
not  g173 (n301, n80);
buf  g174 (n573, n34);
not  g175 (n430, n68);
buf  g176 (n322, n77);
not  g177 (n634, n102);
buf  g178 (n251, n37);
buf  g179 (n519, n73);
not  g180 (n591, n89);
buf  g181 (n604, n130);
buf  g182 (n584, n122);
not  g183 (n240, n53);
buf  g184 (n201, n84);
buf  g185 (n615, n35);
not  g186 (n581, n75);
not  g187 (n572, n33);
not  g188 (n448, n83);
not  g189 (n438, n123);
not  g190 (n658, n107);
buf  g191 (n276, n55);
buf  g192 (n347, n146);
not  g193 (n661, n75);
buf  g194 (n585, n42);
not  g195 (n459, n77);
not  g196 (n662, n138);
buf  g197 (n190, n66);
buf  g198 (n633, n72);
buf  g199 (n380, n85);
buf  g200 (n659, n71);
buf  g201 (n429, n137);
buf  g202 (n552, n71);
buf  g203 (n587, n92);
buf  g204 (n300, n34);
not  g205 (n555, n132);
not  g206 (n510, n60);
buf  g207 (n506, n86);
buf  g208 (n644, n63);
not  g209 (n230, n56);
not  g210 (n531, n156);
buf  g211 (n242, n48);
not  g212 (n342, n64);
buf  g213 (n299, n67);
not  g214 (n665, n50);
buf  g215 (n370, n122);
buf  g216 (n378, n79);
buf  g217 (n475, n81);
buf  g218 (n522, n43);
buf  g219 (n218, n111);
buf  g220 (n419, n36);
buf  g221 (n428, n158);
not  g222 (n221, n104);
buf  g223 (n214, n125);
not  g224 (n599, n60);
not  g225 (n560, n85);
not  g226 (n390, n92);
not  g227 (n294, n60);
buf  g228 (n166, n125);
buf  g229 (n260, n150);
buf  g230 (n439, n90);
buf  g231 (n177, n114);
not  g232 (n205, n45);
not  g233 (n490, n158);
buf  g234 (n333, n97);
not  g235 (n524, n102);
buf  g236 (n564, n103);
buf  g237 (n554, n39);
buf  g238 (n273, n64);
buf  g239 (n320, n118);
not  g240 (n343, n156);
not  g241 (n422, n116);
not  g242 (n625, n113);
not  g243 (n473, n39);
buf  g244 (n288, n97);
buf  g245 (n469, n115);
buf  g246 (n208, n72);
not  g247 (n264, n36);
not  g248 (n303, n113);
buf  g249 (n639, n129);
buf  g250 (n455, n117);
not  g251 (n279, n140);
not  g252 (n346, n110);
not  g253 (n357, n149);
not  g254 (n404, n115);
not  g255 (n652, n105);
not  g256 (n653, n44);
not  g257 (n189, n70);
buf  g258 (n395, n114);
not  g259 (n664, n49);
buf  g260 (n436, n75);
not  g261 (n593, n54);
buf  g262 (n255, n100);
buf  g263 (n543, n76);
buf  g264 (n534, n103);
not  g265 (n353, n151);
not  g266 (n651, n44);
buf  g267 (n491, n126);
not  g268 (n645, n96);
buf  g269 (n643, n126);
not  g270 (n607, n99);
buf  g271 (n403, n120);
not  g272 (n492, n134);
not  g273 (n266, n106);
buf  g274 (n602, n125);
not  g275 (n306, n78);
not  g276 (n170, n100);
buf  g277 (n537, n131);
buf  g278 (n477, n121);
buf  g279 (n247, n128);
buf  g280 (n258, n130);
buf  g281 (n447, n33);
buf  g282 (n672, n79);
buf  g283 (n296, n72);
buf  g284 (n551, n131);
not  g285 (n458, n68);
not  g286 (n239, n116);
not  g287 (n246, n135);
not  g288 (n619, n144);
buf  g289 (n623, n142);
buf  g290 (n185, n38);
not  g291 (n549, n73);
buf  g292 (n588, n144);
buf  g293 (n257, n121);
buf  g294 (n307, n82);
buf  g295 (n340, n107);
buf  g296 (n364, n100);
buf  g297 (n369, n86);
buf  g298 (n575, n33);
buf  g299 (n457, n110);
buf  g300 (n168, n51);
not  g301 (n541, n33);
buf  g302 (n484, n78);
buf  g303 (n441, n150);
not  g304 (n256, n104);
not  g305 (n666, n123);
buf  g306 (n605, n81);
not  g307 (n546, n77);
not  g308 (n416, n41);
not  g309 (n381, n83);
buf  g310 (n568, n108);
buf  g311 (n411, n58);
not  g312 (n179, n80);
buf  g313 (n305, n143);
buf  g314 (n210, n129);
buf  g315 (n536, n118);
not  g316 (n528, n154);
not  g317 (n224, n83);
not  g318 (n553, n158);
not  g319 (n562, n139);
not  g320 (n284, n91);
buf  g321 (n374, n36);
buf  g322 (n389, n34);
not  g323 (n163, n118);
not  g324 (n345, n51);
not  g325 (n583, n152);
buf  g326 (n194, n80);
not  g327 (n282, n155);
not  g328 (n225, n60);
not  g329 (n407, n154);
buf  g330 (n330, n120);
buf  g331 (n667, n53);
not  g332 (n577, n95);
not  g333 (n570, n152);
not  g334 (n386, n56);
buf  g335 (n200, n49);
buf  g336 (n437, n101);
not  g337 (n377, n100);
not  g338 (n614, n55);
not  g339 (n671, n88);
buf  g340 (n630, n113);
not  g341 (n231, n56);
not  g342 (n452, n90);
buf  g343 (n487, n63);
not  g344 (n505, n41);
buf  g345 (n472, n82);
not  g346 (n649, n57);
buf  g347 (n280, n40);
not  g348 (n592, n57);
not  g349 (n359, n149);
not  g350 (n337, n99);
not  g351 (n451, n94);
buf  g352 (n252, n143);
buf  g353 (n540, n119);
buf  g354 (n466, n65);
not  g355 (n297, n140);
buf  g356 (n654, n76);
not  g357 (n668, n133);
buf  g358 (n557, n88);
buf  g359 (n196, n147);
buf  g360 (n561, n145);
buf  g361 (n464, n159);
buf  g362 (n384, n93);
not  g363 (n178, n47);
not  g364 (n283, n106);
not  g365 (n181, n153);
not  g366 (n408, n59);
not  g367 (n184, n96);
not  g368 (n435, n52);
buf  g369 (n567, n128);
not  g370 (n309, n124);
buf  g371 (n175, n50);
not  g372 (n431, n114);
buf  g373 (n486, n126);
buf  g374 (n631, n41);
not  g375 (n660, n107);
buf  g376 (n215, n149);
buf  g377 (n272, n37);
buf  g378 (n286, n135);
not  g379 (n365, n101);
not  g380 (n456, n94);
not  g381 (n566, n89);
not  g382 (n388, n46);
buf  g383 (n171, n55);
not  g384 (n400, n134);
buf  g385 (n211, n85);
buf  g386 (n292, n50);
buf  g387 (n373, n81);
not  g388 (n350, n134);
buf  g389 (n344, n62);
buf  g390 (n226, n119);
buf  g391 (n293, n43);
buf  g392 (n182, n57);
buf  g393 (n603, n67);
not  g394 (n363, n41);
buf  g395 (n315, n69);
buf  g396 (n589, n48);
not  g397 (n191, n43);
not  g398 (n316, n110);
not  g399 (n600, n70);
not  g400 (n263, n57);
not  g401 (n569, n124);
buf  g402 (n509, n71);
not  g403 (n582, n148);
buf  g404 (n204, n69);
buf  g405 (n445, n122);
not  g406 (n327, n59);
buf  g407 (n596, n122);
not  g408 (n427, n145);
not  g409 (n520, n124);
not  g410 (n499, n153);
buf  g411 (n387, n51);
not  g412 (n328, n101);
not  g413 (n271, n133);
buf  g414 (n595, n47);
buf  g415 (n482, n153);
not  g416 (n249, n133);
not  g417 (n236, n160);
not  g418 (n164, n108);
buf  g419 (n402, n137);
not  g420 (n453, n62);
not  g421 (n287, n37);
not  g422 (n325, n49);
buf  g423 (n629, n136);
buf  g424 (n542, n136);
not  g425 (n202, n156);
buf  g426 (n471, n147);
buf  g427 (n513, n123);
not  g428 (n494, n51);
not  g429 (n248, n142);
buf  g430 (n237, n70);
buf  g431 (n321, n96);
not  g432 (n338, n105);
buf  g433 (n669, n92);
not  g434 (n526, n79);
buf  g435 (n468, n84);
buf  g436 (n580, n58);
buf  g437 (n209, n42);
not  g438 (n594, n145);
buf  g439 (n352, n66);
buf  g440 (n632, n92);
buf  g441 (n335, n54);
buf  g442 (n367, n131);
not  g443 (n311, n99);
buf  g444 (n571, n43);
not  g445 (n176, n109);
not  g446 (n368, n141);
buf  g447 (n545, n130);
buf  g448 (n270, n135);
buf  g449 (n516, n35);
buf  g450 (n462, n151);
buf  g451 (n421, n39);
not  g452 (n324, n136);
not  g453 (n269, n97);
buf  g454 (n418, n145);
not  g455 (n406, n109);
buf  g456 (n642, n160);
not  g457 (n278, n104);
buf  g458 (n465, n93);
buf  g459 (n233, n127);
buf  g460 (n336, n74);
not  g461 (n310, n46);
buf  g462 (n488, n160);
buf  g463 (n597, n142);
buf  g464 (n334, n146);
buf  g465 (n636, n55);
buf  g466 (n532, n98);
not  g467 (n262, n66);
not  g468 (n220, n40);
buf  g469 (n351, n114);
buf  g470 (n254, n45);
buf  g471 (n396, n63);
buf  g472 (n476, n147);
buf  g473 (n504, n47);
buf  g474 (n385, n39);
not  g475 (n195, n160);
not  g476 (n304, n151);
buf  g477 (n641, n109);
buf  g478 (n440, n137);
not  g479 (n393, n112);
not  g480 (n354, n48);
buf  g481 (n394, n139);
not  g482 (n376, n80);
buf  g483 (n574, n158);
not  g484 (n495, n101);
buf  g485 (n601, n95);
not  g486 (n361, n124);
not  g487 (n426, n144);
not  g488 (n606, n67);
not  g489 (n227, n44);
buf  g490 (n339, n141);
not  g491 (n267, n50);
not  g492 (n245, n68);
not  g493 (n234, n45);
buf  g494 (n497, n91);
not  g495 (n640, n90);
not  g496 (n558, n108);
buf  g497 (n443, n144);
not  g498 (n508, n76);
buf  g499 (n444, n61);
buf  g500 (n308, n86);
not  g501 (n479, n147);
buf  g502 (n550, n139);
not  g503 (n663, n120);
buf  g504 (n250, n138);
buf  g505 (n530, n148);
buf  g506 (n523, n65);
not  g507 (n617, n38);
not  g508 (n621, n131);
not  g509 (n538, n129);
buf  g510 (n355, n66);
buf  g511 (n323, n82);
buf  g512 (n332, n48);
not  g513 (n670, n40);
not  g514 (n167, n37);
buf  g515 (n622, n153);
not  g516 (n627, n59);
buf  g517 (n489, n91);
buf  g518 (n397, n159);
buf  g519 (n425, n115);
not  g520 (n511, n120);
not  g521 (n424, n78);
buf  g522 (n527, n111);
buf  g523 (n656, n95);
not  g524 (n392, n64);
buf  g525 (n576, n97);
buf  g526 (n410, n107);
not  g527 (n372, n143);
not  g528 (n474, n76);
not  g529 (n314, n87);
buf  g530 (n405, n62);
buf  g531 (n616, n34);
buf  g532 (n379, n46);
not  g533 (n331, n79);
buf  g534 (n253, n102);
buf  g535 (n493, n128);
buf  g536 (n165, n54);
not  g537 (n478, n42);
not  g538 (n500, n156);
not  g539 (n613, n148);
buf  g540 (n485, n44);
buf  g541 (n268, n143);
buf  g542 (n507, n133);
not  g543 (n173, n106);
buf  g544 (n326, n123);
buf  g545 (n624, n132);
buf  g546 (n243, n94);
not  g547 (n289, n65);
not  g548 (n172, n137);
buf  g549 (n521, n110);
not  g550 (n496, n75);
buf  g551 (n442, n93);
not  g552 (n383, n85);
not  g553 (n415, n134);
not  g554 (n162, n87);
buf  g555 (n290, n87);
not  g556 (n611, n118);
buf  g557 (n512, n95);
buf  g558 (n423, n53);
not  g559 (n341, n77);
not  g560 (n525, n61);
not  g561 (n192, n49);
buf  g562 (n265, n117);
buf  g563 (n657, n154);
buf  g564 (n213, n148);
not  g565 (n318, n140);
buf  g566 (n535, n128);
buf  g567 (n578, n102);
not  g568 (n261, n54);
buf  g569 (n217, n157);
not  g570 (n608, n103);
not  g571 (n650, n74);
not  g572 (n356, n81);
not  g573 (n207, n104);
not  g574 (n635, n59);
buf  g575 (n590, n86);
not  g576 (n362, n45);
buf  g577 (n382, n46);
buf  g578 (n302, n139);
buf  g579 (n432, n61);
not  g580 (n319, n117);
not  g581 (n238, n152);
buf  g582 (n274, n98);
buf  g583 (n463, n138);
not  g584 (n547, n63);
buf  g585 (n626, n117);
buf  g586 (n647, n126);
not  g587 (n349, n65);
buf  g588 (n533, n150);
not  g589 (n180, n109);
not  g590 (n470, n73);
not  g591 (n329, n69);
buf  g592 (n450, n89);
not  g593 (n199, n52);
not  g594 (n366, n146);
not  g595 (n544, n38);
not  g596 (n517, n87);
buf  g597 (n232, n94);
not  g598 (n433, n68);
not  g599 (n412, n52);
not  g600 (n212, n83);
buf  g601 (n446, n116);
buf  g602 (n414, n132);
not  g603 (n183, n40);
buf  g604 (n460, n108);
buf  g605 (n186, n93);
not  g606 (n291, n154);
buf  g607 (n420, n121);
buf  g608 (n399, n111);
not  g609 (n398, n58);
buf  g610 (n461, n84);
not  g611 (n391, n113);
not  g612 (n223, n105);
not  g613 (n454, n90);
not  g614 (n518, n89);
not  g615 (n610, n88);
not  g616 (n481, n67);
not  g617 (n515, n99);
not  g618 (n628, n130);
not  g619 (n312, n159);
buf  g620 (n244, n116);
buf  g621 (n161, n103);
not  g622 (n480, n70);
not  g623 (n235, n152);
buf  g624 (n556, n105);
not  g625 (n295, n88);
not  g626 (n612, n119);
buf  g627 (n229, n64);
buf  g628 (n203, n42);
not  g629 (n529, n38);
not  g630 (n375, n155);
buf  g631 (n655, n112);
buf  g632 (n434, n129);
not  g633 (n637, n127);
buf  g634 (n174, n72);
buf  g635 (n467, n135);
buf  g636 (n483, n127);
buf  g637 (n193, n74);
buf  g638 (n598, n47);
buf  g639 (n241, n146);
not  g640 (n795, n623);
buf  g641 (n804, n509);
not  g642 (n777, n638);
buf  g643 (n764, n643);
buf  g644 (n694, n293);
not  g645 (n832, n640);
not  g646 (n879, n554);
not  g647 (n856, n344);
buf  g648 (n872, n329);
buf  g649 (n805, n636);
not  g650 (n733, n308);
buf  g651 (n867, n651);
not  g652 (n696, n614);
buf  g653 (n893, n457);
buf  g654 (n757, n362);
buf  g655 (n803, n633);
not  g656 (n889, n642);
not  g657 (n870, n470);
buf  g658 (n926, n188);
buf  g659 (n927, n386);
not  g660 (n828, n481);
buf  g661 (n833, n253);
buf  g662 (n880, n173);
buf  g663 (n790, n345);
buf  g664 (n933, n446);
buf  g665 (n682, n527);
not  g666 (n752, n633);
not  g667 (n796, n642);
buf  g668 (n708, n287);
not  g669 (n772, n482);
not  g670 (n836, n609);
not  g671 (n811, n288);
buf  g672 (n944, n197);
buf  g673 (n748, n542);
not  g674 (n892, n654);
not  g675 (n775, n620);
buf  g676 (n865, n621);
not  g677 (n886, n214);
buf  g678 (n746, n597);
buf  g679 (n911, n419);
not  g680 (n849, n629);
not  g681 (n851, n269);
not  g682 (n920, n306);
buf  g683 (n937, n248);
not  g684 (n731, n296);
buf  g685 (n801, n530);
not  g686 (n823, n224);
buf  g687 (n874, n380);
not  g688 (n741, n639);
not  g689 (n825, n409);
not  g690 (n862, n645);
buf  g691 (n739, n366);
not  g692 (n930, n629);
buf  g693 (n939, n373);
not  g694 (n843, n286);
not  g695 (n767, n503);
buf  g696 (n799, n336);
buf  g697 (n840, n353);
buf  g698 (n701, n583);
buf  g699 (n923, n403);
buf  g700 (n759, n593);
not  g701 (n810, n501);
buf  g702 (n830, n648);
not  g703 (n711, n641);
not  g704 (n744, n265);
not  g705 (n773, n580);
buf  g706 (n727, n387);
buf  g707 (n922, n586);
not  g708 (n912, n459);
buf  g709 (n808, n257);
not  g710 (n854, n365);
not  g711 (n848, n604);
buf  g712 (n781, n268);
not  g713 (n783, n210);
not  g714 (n720, n639);
not  g715 (n675, n524);
not  g716 (n863, n515);
buf  g717 (n921, n358);
not  g718 (n765, n635);
buf  g719 (n786, n643);
not  g720 (n941, n557);
not  g721 (n782, n440);
buf  g722 (n894, n543);
not  g723 (n740, n227);
not  g724 (n712, n304);
buf  g725 (n902, n460);
buf  g726 (n705, n472);
buf  g727 (n878, n402);
not  g728 (n692, n385);
not  g729 (n905, n647);
buf  g730 (n932, n600);
buf  g731 (n835, n217);
not  g732 (n850, n444);
buf  g733 (n861, n297);
buf  g734 (n852, n239);
buf  g735 (n907, n652);
buf  g736 (n751, n219);
not  g737 (n895, n312);
buf  g738 (n913, n596);
buf  g739 (n673, n528);
not  g740 (n925, n544);
not  g741 (n723, n479);
not  g742 (n857, n494);
buf  g743 (n837, n627);
buf  g744 (n730, n180);
not  g745 (n877, n626);
not  g746 (n768, n471);
buf  g747 (n871, n536);
buf  g748 (n792, n392);
not  g749 (n859, n454);
buf  g750 (n763, n391);
not  g751 (n858, n251);
buf  g752 (n931, n584);
buf  g753 (n737, n620);
not  g754 (n942, n431);
not  g755 (n706, n653);
not  g756 (n888, n591);
buf  g757 (n690, n637);
buf  g758 (n918, n621);
not  g759 (n697, n311);
not  g760 (n900, n613);
buf  g761 (n695, n480);
buf  g762 (n704, n519);
not  g763 (n735, n327);
not  g764 (n753, n625);
not  g765 (n709, n639);
not  g766 (n684, n437);
not  g767 (n713, n170);
buf  g768 (n940, n649);
buf  g769 (n780, n426);
not  g770 (n891, n178);
buf  g771 (n714, n571);
buf  g772 (n745, n307);
buf  g773 (n917, n207);
buf  g774 (n687, n552);
buf  g775 (n769, n343);
buf  g776 (n758, n309);
not  g777 (n742, n626);
not  g778 (n820, n556);
not  g779 (n732, n521);
not  g780 (n908, n628);
not  g781 (n890, n250);
not  g782 (n928, n526);
buf  g783 (n698, n644);
not  g784 (n729, n242);
not  g785 (n845, n650);
buf  g786 (n699, n175);
buf  g787 (n802, n449);
buf  g788 (n881, n393);
not  g789 (n721, n279);
not  g790 (n770, n379);
buf  g791 (n809, n466);
not  g792 (n869, n201);
buf  g793 (n896, n654);
not  g794 (n674, n619);
buf  g795 (n677, n511);
buf  g796 (n686, n364);
not  g797 (n707, n641);
not  g798 (n813, n598);
not  g799 (n814, n272);
and  g800 (n838, n283, n614, n290, n650);
xnor g801 (n722, n508, n367, n243, n623);
xnor g802 (n778, n588, n360, n314, n216);
or   g803 (n785, n414, n615, n161, n653);
xor  g804 (n885, n640, n602, n334, n498);
nand g805 (n906, n573, n555, n236, n351);
or   g806 (n806, n368, n623, n273, n644);
nand g807 (n882, n421, n356, n432, n410);
nand g808 (n676, n589, n398, n499, n195);
nor  g809 (n734, n291, n168, n648, n585);
xnor g810 (n693, n496, n575, n234, n654);
nor  g811 (n868, n618, n628, n422, n192);
xor  g812 (n816, n164, n189, n274, n319);
nand g813 (n860, n225, n424, n626, n651);
nand g814 (n915, n626, n601, n374, n478);
xor  g815 (n756, n642, n612, n357, n191);
nor  g816 (n824, n282, n247, n448, n442);
and  g817 (n750, n630, n162, n625, n453);
xnor g818 (n685, n537, n605, n644, n637);
and  g819 (n812, n592, n513, n611, n622);
xnor g820 (n728, n635, n220, n622, n633);
or   g821 (n909, n473, n441, n340, n411);
xnor g822 (n821, n324, n474, n627);
or   g823 (n724, n423, n436, n634, n425);
and  g824 (n718, n564, n516, n653, n645);
nor  g825 (n822, n185, n439, n510, n641);
or   g826 (n719, n204, n476, n315, n382);
and  g827 (n943, n464, n649, n622, n491);
or   g828 (n910, n262, n636, n620);
nor  g829 (n754, n255, n233, n539, n559);
and  g830 (n779, n259, n643, n565, n632);
xnor g831 (n680, n485, n582, n384, n203);
or   g832 (n876, n623, n212, n561, n231);
xor  g833 (n797, n632, n369, n415, n627);
xor  g834 (n903, n332, n316, n321, n429);
or   g835 (n817, n427, n545, n570, n645);
nand g836 (n898, n194, n574, n475, n607);
nor  g837 (n855, n167, n462, n375, n241);
nor  g838 (n829, n628, n277, n213, n165);
xor  g839 (n726, n228, n636, n416, n610);
xor  g840 (n929, n244, n634, n456, n560);
nor  g841 (n916, n465, n646, n618, n569);
nor  g842 (n761, n349, n417, n590, n634);
and  g843 (n716, n610, n176, n238, n271);
nand g844 (n717, n443, n323, n337, n451);
nand g845 (n875, n625, n630, n215, n637);
or   g846 (n844, n182, n652, n363, n372);
xnor g847 (n924, n547, n294, n642, n190);
nor  g848 (n897, n330, n594, n579, n370);
or   g849 (n689, n649, n458, n549, n652);
xor  g850 (n794, n518, n184, n587, n646);
nor  g851 (n864, n292, n546, n328, n209);
xor  g852 (n700, n169, n270, n654, n404);
nor  g853 (n743, n650, n647, n377, n620);
nand g854 (n938, n295, n193, n326, n504);
or   g855 (n679, n637, n389, n640, n548);
or   g856 (n789, n396, n299, n383, n278);
or   g857 (n884, n196, n649, n477, n495);
nor  g858 (n873, n260, n468, n625, n240);
and  g859 (n736, n261, n617, n486, n378);
xnor g860 (n683, n407, n651, n608, n435);
xor  g861 (n834, n338, n263, n202, n223);
or   g862 (n826, n581, n333, n445, n399);
xnor g863 (n831, n645, n653, n354, n514);
xor  g864 (n747, n246, n493, n313, n540);
nor  g865 (n819, n531, n381, n434, n232);
or   g866 (n936, n267, n400, n507, n639);
and  g867 (n815, n603, n489, n350, n200);
xor  g868 (n774, n361, n266, n505, n205);
xor  g869 (n688, n611, n631, n452, n487);
xor  g870 (n807, n430, n517, n606, n218);
and  g871 (n846, n635, n303, n461, n355);
or   g872 (n725, n463, n359, n522, n652);
or   g873 (n681, n533, n632, n285, n612);
xnor g874 (n866, n566, n199, n638, n469);
xnor g875 (n787, n226, n621, n211, n648);
xnor g876 (n691, n638, n284, n558, n301);
nand g877 (n853, n624, n567, n289, n406);
or   g878 (n760, n310, n280, n550, n633);
or   g879 (n710, n551, n221, n534, n619);
or   g880 (n899, n438, n245, n252, n655);
xnor g881 (n901, n641, n502, n616, n624);
xnor g882 (n793, n616, n317, n376, n412);
and  g883 (n702, n352, n254, n621, n631);
nor  g884 (n784, n230, n320, n538, n433);
and  g885 (n839, n206, n198, n322, n648);
nor  g886 (n738, n428, n576, n275, n187);
or   g887 (n703, n325, n237, n562, n249);
or   g888 (n749, n346, n629, n395, n331);
nand g889 (n887, n281, n646, n186, n492);
or   g890 (n791, n276, n650, n535, n523);
nor  g891 (n827, n455, n163, n420, n647);
nand g892 (n945, n525, n506, n488, n339);
xnor g893 (n762, n390, n467, n450, n405);
nor  g894 (n771, n408, n520, n563, n512);
nor  g895 (n883, n651, n595, n490, n599);
xnor g896 (n935, n532, n635, n371, n638);
nand g897 (n800, n394, n166, n179, n630);
nand g898 (n755, n348, n640, n529, n335);
xnor g899 (n678, n484, n177, n388, n541);
nand g900 (n818, n342, n171, n572, n229);
nor  g901 (n919, n619, n634, n613, n624);
or   g902 (n766, n483, n318, n500, n644);
nor  g903 (n914, n647, n497, n300, n617);
nand g904 (n934, n629, n632, n298, n553);
xnor g905 (n715, n577, n418, n235, n172);
xnor g906 (n788, n305, n264, n619, n174);
and  g907 (n798, n447, n341, n222, n631);
and  g908 (n841, n643, n347, n302, n397);
nand g909 (n847, n568, n401, n630, n183);
nand g910 (n904, n256, n413, n624, n208);
xor  g911 (n842, n646, n631, n578, n615);
or   g912 (n776, n628, n258, n622, n181);
not  g913 (n948, n865);
not  g914 (n1132, n829);
not  g915 (n1050, n659);
not  g916 (n1059, n702);
buf  g917 (n1109, n827);
not  g918 (n1133, n684);
buf  g919 (n1143, n890);
buf  g920 (n1071, n691);
not  g921 (n981, n918);
not  g922 (n1038, n931);
not  g923 (n1014, n876);
buf  g924 (n1018, n895);
buf  g925 (n975, n746);
buf  g926 (n1099, n792);
not  g927 (n1006, n788);
buf  g928 (n1075, n683);
buf  g929 (n1152, n656);
buf  g930 (n1030, n748);
not  g931 (n1011, n671);
buf  g932 (n1005, n872);
buf  g933 (n966, n806);
not  g934 (n994, n867);
buf  g935 (n953, n833);
buf  g936 (n1022, n810);
buf  g937 (n1141, n738);
not  g938 (n1007, n776);
not  g939 (n998, n658);
not  g940 (n1140, n882);
buf  g941 (n1095, n809);
not  g942 (n967, n662);
not  g943 (n954, n871);
buf  g944 (n1153, n739);
buf  g945 (n950, n716);
buf  g946 (n1097, n828);
not  g947 (n983, n904);
buf  g948 (n1131, n861);
buf  g949 (n1016, n655);
buf  g950 (n1004, n793);
not  g951 (n1128, n759);
buf  g952 (n1103, n846);
not  g953 (n999, n825);
not  g954 (n1126, n857);
buf  g955 (n1151, n710);
buf  g956 (n1015, n780);
not  g957 (n1134, n762);
not  g958 (n1042, n750);
buf  g959 (n988, n718);
buf  g960 (n1025, n903);
not  g961 (n979, n699);
buf  g962 (n1057, n822);
buf  g963 (n1081, n657);
not  g964 (n1149, n929);
buf  g965 (n1056, n933);
buf  g966 (n1105, n930);
not  g967 (n1060, n851);
buf  g968 (n1114, n752);
buf  g969 (n947, n667);
not  g970 (n1062, n832);
not  g971 (n1065, n818);
buf  g972 (n964, n666);
buf  g973 (n1044, n670);
buf  g974 (n1010, n771);
not  g975 (n960, n908);
buf  g976 (n1108, n686);
not  g977 (n1118, n924);
buf  g978 (n1077, n785);
buf  g979 (n970, n720);
not  g980 (n955, n715);
buf  g981 (n996, n880);
not  g982 (n993, n773);
buf  g983 (n1123, n660);
not  g984 (n1063, n919);
not  g985 (n1091, n888);
not  g986 (n1054, n728);
not  g987 (n1098, n664);
not  g988 (n1147, n787);
not  g989 (n1085, n676);
buf  g990 (n1096, n779);
buf  g991 (n958, n915);
not  g992 (n976, n701);
buf  g993 (n1138, n673);
not  g994 (n1080, n875);
buf  g995 (n1031, n671);
not  g996 (n1078, n753);
buf  g997 (n1008, n659);
not  g998 (n1087, n834);
buf  g999 (n1051, n845);
buf  g1000 (n1040, n690);
not  g1001 (n1094, n730);
buf  g1002 (n968, n661);
buf  g1003 (n1032, n669);
not  g1004 (n1124, n669);
not  g1005 (n1017, n841);
not  g1006 (n989, n803);
buf  g1007 (n1090, n657);
not  g1008 (n1034, n923);
not  g1009 (n1041, n693);
not  g1010 (n1089, n782);
not  g1011 (n1021, n911);
buf  g1012 (n1106, n663);
not  g1013 (n1104, n909);
not  g1014 (n1046, n664);
buf  g1015 (n1058, n735);
buf  g1016 (n1073, n751);
not  g1017 (n973, n769);
buf  g1018 (n1100, n835);
not  g1019 (n980, n807);
buf  g1020 (n1111, n749);
buf  g1021 (n1045, n940);
not  g1022 (n1003, n733);
not  g1023 (n1139, n740);
not  g1024 (n986, n860);
buf  g1025 (n1137, n695);
buf  g1026 (n1043, n925);
not  g1027 (n1107, n907);
buf  g1028 (n963, n719);
not  g1029 (n949, n934);
not  g1030 (n1086, n839);
not  g1031 (n946, n665);
buf  g1032 (n1144, n830);
not  g1033 (n1083, n892);
not  g1034 (n1121, n866);
not  g1035 (n978, n671);
not  g1036 (n1142, n714);
buf  g1037 (n1009, n662);
buf  g1038 (n997, n662);
buf  g1039 (n990, n668);
buf  g1040 (n985, n756);
not  g1041 (n1052, n704);
not  g1042 (n1000, n727);
buf  g1043 (n1112, n667);
buf  g1044 (n1125, n667);
not  g1045 (n1033, n801);
not  g1046 (n1013, n850);
not  g1047 (n959, n657);
not  g1048 (n1136, n655);
buf  g1049 (n1129, n886);
buf  g1050 (n1026, n680);
buf  g1051 (n1070, n669);
not  g1052 (n1035, n817);
not  g1053 (n1074, n838);
buf  g1054 (n1066, n795);
buf  g1055 (n1093, n703);
buf  g1056 (n991, n798);
buf  g1057 (n1120, n844);
buf  g1058 (n1150, n900);
buf  g1059 (n1148, n887);
buf  g1060 (n1012, n661);
not  g1061 (n1069, n696);
buf  g1062 (n1072, n778);
not  g1063 (n1146, n672);
buf  g1064 (n1088, n783);
not  g1065 (n961, n898);
not  g1066 (n1119, n913);
buf  g1067 (n956, n662);
buf  g1068 (n952, n758);
buf  g1069 (n1092, n815);
buf  g1070 (n1028, n786);
buf  g1071 (n987, n790);
buf  g1072 (n1001, n687);
not  g1073 (n1115, n698);
not  g1074 (n1102, n799);
not  g1075 (n1036, n939);
and  g1076 (n1110, n734, n883, n840, n781);
or   g1077 (n1122, n935, n858, n881, n712);
and  g1078 (n992, n755, n656, n863, n668);
and  g1079 (n1067, n837, n757, n853, n717);
xor  g1080 (n1127, n668, n666, n692);
or   g1081 (n1064, n681, n760, n794, n893);
and  g1082 (n1113, n889, n685, n766, n942);
and  g1083 (n1020, n705, n774, n660);
nand g1084 (n1116, n700, n663, n669, n665);
and  g1085 (n1061, n679, n884, n873, n894);
or   g1086 (n1053, n697, n777, n808, n658);
xnor g1087 (n1055, n789, n655, n820, n675);
nand g1088 (n1019, n665, n943, n657, n672);
nor  g1089 (n984, n713, n879, n945, n862);
xor  g1090 (n1023, n764, n666, n722, n665);
xnor g1091 (n1082, n896, n723, n660, n656);
and  g1092 (n1101, n842, n906, n688, n732);
or   g1093 (n957, n763, n901, n897, n663);
or   g1094 (n1027, n916, n811, n800, n937);
xor  g1095 (n977, n885, n670, n775, n819);
xor  g1096 (n971, n742, n772, n765, n724);
and  g1097 (n969, n682, n926, n761, n736);
nand g1098 (n1002, n921, n658, n878, n745);
xor  g1099 (n951, n659, n812, n823, n944);
xnor g1100 (n1145, n664, n656, n927, n784);
xor  g1101 (n1029, n726, n864, n874, n928);
xor  g1102 (n972, n744, n813, n741, n848);
or   g1103 (n974, n670, n824, n847, n804);
or   g1104 (n1079, n816, n708, n854, n932);
or   g1105 (n1037, n910, n661, n721, n791);
nand g1106 (n962, n768, n922, n938, n902);
nand g1107 (n1076, n706, n802, n914, n743);
xnor g1108 (n1024, n856, n941, n658, n767);
or   g1109 (n982, n663, n852, n709, n737);
nand g1110 (n1068, n672, n729, n869, n868);
nand g1111 (n965, n670, n843, n912, n689);
or   g1112 (n1047, n711, n877, n826, n661);
and  g1113 (n1084, n659, n936, n668, n667);
nor  g1114 (n995, n796, n855, n707, n836);
xor  g1115 (n1135, n905, n797, n671, n754);
or   g1116 (n1130, n747, n664, n731, n677);
nand g1117 (n1048, n859, n674, n770, n694);
nor  g1118 (n1049, n725, n870, n849, n805);
and  g1119 (n1117, n831, n678, n814, n821);
nor  g1120 (n1039, n899, n920, n891, n917);
not  g1121 (n1163, n967);
not  g1122 (n1174, n1008);
not  g1123 (n1243, n1093);
not  g1124 (n1214, n1094);
not  g1125 (n1208, n1113);
not  g1126 (n1171, n989);
buf  g1127 (n1249, n1029);
not  g1128 (n1239, n1098);
not  g1129 (n1307, n1091);
not  g1130 (n1305, n986);
buf  g1131 (n1312, n974);
not  g1132 (n1184, n1067);
buf  g1133 (n1250, n1071);
buf  g1134 (n1173, n991);
buf  g1135 (n1196, n1077);
buf  g1136 (n1209, n956);
buf  g1137 (n1303, n982);
buf  g1138 (n1298, n971);
buf  g1139 (n1301, n959);
not  g1140 (n1172, n969);
buf  g1141 (n1327, n1003);
buf  g1142 (n1299, n1060);
buf  g1143 (n1289, n947);
buf  g1144 (n1266, n1024);
buf  g1145 (n1178, n962);
not  g1146 (n1186, n1059);
not  g1147 (n1265, n1052);
buf  g1148 (n1260, n976);
buf  g1149 (n1257, n993);
buf  g1150 (n1258, n1013);
not  g1151 (n1245, n1015);
not  g1152 (n1297, n1116);
not  g1153 (n1319, n1105);
not  g1154 (n1204, n952);
buf  g1155 (n1235, n1108);
not  g1156 (n1318, n1085);
buf  g1157 (n1217, n1089);
not  g1158 (n1302, n1112);
buf  g1159 (n1176, n1036);
not  g1160 (n1323, n1072);
buf  g1161 (n1268, n1038);
not  g1162 (n1254, n973);
buf  g1163 (n1255, n1020);
not  g1164 (n1290, n1070);
buf  g1165 (n1213, n1014);
buf  g1166 (n1317, n997);
not  g1167 (n1304, n1106);
buf  g1168 (n1292, n1004);
not  g1169 (n1272, n1055);
buf  g1170 (n1157, n1082);
buf  g1171 (n1169, n1064);
buf  g1172 (n1181, n988);
not  g1173 (n1247, n954);
buf  g1174 (n1237, n1092);
buf  g1175 (n1271, n1007);
not  g1176 (n1241, n1027);
not  g1177 (n1293, n990);
not  g1178 (n1295, n975);
not  g1179 (n1156, n1032);
buf  g1180 (n1309, n1012);
buf  g1181 (n1288, n999);
not  g1182 (n1220, n1066);
not  g1183 (n1286, n966);
buf  g1184 (n1202, n955);
buf  g1185 (n1228, n985);
buf  g1186 (n1324, n1023);
not  g1187 (n1230, n1099);
not  g1188 (n1158, n1058);
buf  g1189 (n1296, n1046);
buf  g1190 (n1308, n1005);
not  g1191 (n1311, n981);
buf  g1192 (n1161, n1006);
buf  g1193 (n1291, n1054);
not  g1194 (n1190, n1031);
buf  g1195 (n1281, n1001);
not  g1196 (n1160, n963);
not  g1197 (n1211, n978);
buf  g1198 (n1183, n972);
not  g1199 (n1270, n1049);
not  g1200 (n1207, n965);
buf  g1201 (n1200, n1068);
buf  g1202 (n1238, n958);
buf  g1203 (n1198, n1076);
not  g1204 (n1216, n1079);
buf  g1205 (n1300, n1065);
not  g1206 (n1267, n1087);
buf  g1207 (n1166, n979);
not  g1208 (n1234, n953);
not  g1209 (n1182, n1056);
buf  g1210 (n1315, n1062);
buf  g1211 (n1306, n980);
not  g1212 (n1180, n1096);
not  g1213 (n1313, n984);
not  g1214 (n1294, n1081);
not  g1215 (n1203, n1073);
buf  g1216 (n1276, n1061);
not  g1217 (n1274, n1034);
not  g1218 (n1251, n1025);
not  g1219 (n1278, n1040);
buf  g1220 (n1229, n1017);
buf  g1221 (n1177, n1115);
not  g1222 (n1310, n1021);
not  g1223 (n1321, n995);
buf  g1224 (n1194, n948);
buf  g1225 (n1154, n992);
buf  g1226 (n1263, n970);
buf  g1227 (n1314, n949);
not  g1228 (n1179, n977);
not  g1229 (n1282, n1018);
not  g1230 (n1259, n1078);
buf  g1231 (n1199, n1084);
not  g1232 (n1215, n1097);
buf  g1233 (n1187, n964);
not  g1234 (n1226, n1118);
buf  g1235 (n1219, n1030);
not  g1236 (n1240, n1104);
buf  g1237 (n1221, n1022);
buf  g1238 (n1188, n1075);
not  g1239 (n1205, n1117);
buf  g1240 (n1231, n987);
buf  g1241 (n1246, n1069);
not  g1242 (n1189, n1047);
buf  g1243 (n1233, n1083);
buf  g1244 (n1283, n961);
buf  g1245 (n1275, n1080);
not  g1246 (n1175, n1101);
buf  g1247 (n1325, n1042);
buf  g1248 (n1192, n1107);
buf  g1249 (n1227, n1111);
not  g1250 (n1256, n1016);
buf  g1251 (n1223, n1000);
not  g1252 (n1222, n983);
not  g1253 (n1164, n1045);
not  g1254 (n1269, n1009);
buf  g1255 (n1248, n1110);
buf  g1256 (n1252, n1100);
buf  g1257 (n1212, n1088);
buf  g1258 (n1159, n1095);
not  g1259 (n1168, n1057);
not  g1260 (n1167, n1028);
buf  g1261 (n1195, n1037);
buf  g1262 (n1210, n1109);
not  g1263 (n1279, n1002);
not  g1264 (n1170, n1119);
not  g1265 (n1185, n1043);
buf  g1266 (n1261, n950);
buf  g1267 (n1201, n1051);
buf  g1268 (n1253, n1011);
not  g1269 (n1287, n1050);
buf  g1270 (n1191, n951);
buf  g1271 (n1273, n998);
buf  g1272 (n1242, n1063);
not  g1273 (n1244, n1039);
buf  g1274 (n1326, n946);
buf  g1275 (n1320, n1090);
buf  g1276 (n1277, n1074);
buf  g1277 (n1316, n1026);
not  g1278 (n1218, n1103);
buf  g1279 (n1193, n1035);
buf  g1280 (n1165, n996);
not  g1281 (n1224, n994);
not  g1282 (n1280, n1114);
buf  g1283 (n1232, n1086);
not  g1284 (n1236, n1010);
not  g1285 (n1162, n1041);
not  g1286 (n1264, n1048);
buf  g1287 (n1206, n1053);
not  g1288 (n1225, n968);
not  g1289 (n1262, n960);
buf  g1290 (n1155, n957);
not  g1291 (n1197, n1033);
not  g1292 (n1322, n1019);
not  g1293 (n1285, n1044);
not  g1294 (n1284, n1102);
not  g1295 (n1351, n1221);
not  g1296 (n1412, n1229);
buf  g1297 (n1355, n1202);
not  g1298 (n1423, n1227);
not  g1299 (n1374, n1159);
buf  g1300 (n1381, n1170);
not  g1301 (n1382, n1230);
buf  g1302 (n1347, n1187);
buf  g1303 (n1372, n1166);
not  g1304 (n1343, n1205);
buf  g1305 (n1334, n1214);
buf  g1306 (n1344, n1230);
not  g1307 (n1389, n1198);
buf  g1308 (n1346, n1172);
not  g1309 (n1333, n1171);
not  g1310 (n1373, n1232);
not  g1311 (n1371, n1186);
buf  g1312 (n1402, n1169);
buf  g1313 (n1364, n1174);
buf  g1314 (n1405, n1230);
buf  g1315 (n1359, n1233);
buf  g1316 (n1362, n1195);
not  g1317 (n1417, n1160);
buf  g1318 (n1366, n1184);
buf  g1319 (n1356, n1196);
buf  g1320 (n1407, n1212);
buf  g1321 (n1406, n1175);
not  g1322 (n1338, n1155);
buf  g1323 (n1397, n1227);
not  g1324 (n1365, n1204);
not  g1325 (n1352, n1193);
not  g1326 (n1378, n1227);
buf  g1327 (n1357, n1200);
buf  g1328 (n1385, n1173);
not  g1329 (n1375, n1223);
not  g1330 (n1369, n1226);
buf  g1331 (n1419, n1197);
buf  g1332 (n1396, n1203);
buf  g1333 (n1349, n1208);
not  g1334 (n1414, n1209);
not  g1335 (n1383, n1231);
not  g1336 (n1330, n1233);
buf  g1337 (n1340, n1224);
not  g1338 (n1350, n1229);
buf  g1339 (n1428, n1215);
buf  g1340 (n1422, n1225);
buf  g1341 (n1360, n1176);
buf  g1342 (n1415, n1220);
not  g1343 (n1413, n1226);
buf  g1344 (n1367, n1192);
buf  g1345 (n1399, n1217);
buf  g1346 (n1410, n1154);
not  g1347 (n1341, n1232);
not  g1348 (n1401, n1232);
buf  g1349 (n1395, n1183);
buf  g1350 (n1411, n1228);
not  g1351 (n1424, n1231);
not  g1352 (n1361, n1167);
buf  g1353 (n1388, n1227);
buf  g1354 (n1426, n1157);
not  g1355 (n1404, n1228);
buf  g1356 (n1408, n1164);
buf  g1357 (n1376, n1230);
not  g1358 (n1329, n1181);
buf  g1359 (n1348, n1194);
buf  g1360 (n1337, n1218);
not  g1361 (n1328, n1213);
not  g1362 (n1392, n1161);
buf  g1363 (n1398, n1216);
buf  g1364 (n1342, n1229);
not  g1365 (n1377, n1191);
not  g1366 (n1386, n1228);
not  g1367 (n1384, n1158);
not  g1368 (n1403, n1177);
not  g1369 (n1394, n1233);
buf  g1370 (n1353, n1210);
buf  g1371 (n1379, n1190);
not  g1372 (n1358, n1201);
buf  g1373 (n1420, n1206);
buf  g1374 (n1363, n1163);
not  g1375 (n1421, n1232);
buf  g1376 (n1370, n1188);
not  g1377 (n1368, n1168);
not  g1378 (n1339, n1229);
not  g1379 (n1380, n1219);
buf  g1380 (n1336, n1180);
not  g1381 (n1387, n1222);
not  g1382 (n1391, n1156);
buf  g1383 (n1345, n1182);
not  g1384 (n1400, n1231);
buf  g1385 (n1416, n1233);
buf  g1386 (n1354, n1162);
not  g1387 (n1331, n1165);
buf  g1388 (n1409, n1185);
buf  g1389 (n1425, n1228);
not  g1390 (n1427, n1179);
buf  g1391 (n1390, n1199);
not  g1392 (n1429, n1178);
buf  g1393 (n1393, n1231);
not  g1394 (n1335, n1207);
not  g1395 (n1332, n1189);
buf  g1396 (n1418, n1211);
not  g1397 (n1435, n1341);
buf  g1398 (n1470, n1346);
buf  g1399 (n1431, n1339);
not  g1400 (n1475, n1334);
not  g1401 (n1472, n1343);
buf  g1402 (n1467, n1338);
not  g1403 (n1494, n1339);
buf  g1404 (n1441, n1336);
buf  g1405 (n1439, n1329);
buf  g1406 (n1442, n1344);
not  g1407 (n1468, n1340);
not  g1408 (n1478, n1333);
not  g1409 (n1469, n1344);
not  g1410 (n1434, n1338);
not  g1411 (n1486, n1334);
buf  g1412 (n1450, n1341);
buf  g1413 (n1471, n1342);
buf  g1414 (n1440, n1330);
not  g1415 (n1430, n1349);
not  g1416 (n1477, n1340);
not  g1417 (n1491, n1334);
buf  g1418 (n1473, n1347);
buf  g1419 (n1455, n1340);
buf  g1420 (n1480, n1333);
buf  g1421 (n1437, n1348);
not  g1422 (n1496, n1337);
buf  g1423 (n1490, n1337);
not  g1424 (n1458, n1333);
not  g1425 (n1445, n1335);
not  g1426 (n1482, n1346);
not  g1427 (n1484, n1350);
buf  g1428 (n1448, n1347);
buf  g1429 (n1464, n1336);
not  g1430 (n1449, n1335);
buf  g1431 (n1451, n1343);
buf  g1432 (n1479, n1345);
buf  g1433 (n1474, n1349);
buf  g1434 (n1495, n1339);
buf  g1435 (n1487, n1342);
not  g1436 (n1499, n1347);
buf  g1437 (n1500, n1337);
not  g1438 (n1433, n1339);
buf  g1439 (n1502, n1336);
buf  g1440 (n1438, n1346);
buf  g1441 (n1465, n1335);
buf  g1442 (n1462, n1338);
not  g1443 (n1483, n1345);
not  g1444 (n1503, n1337);
buf  g1445 (n1459, n1345);
not  g1446 (n1456, n1332);
not  g1447 (n1444, n1348);
buf  g1448 (n1463, n1334);
not  g1449 (n1453, n1348);
not  g1450 (n1498, n1328);
buf  g1451 (n1447, n1336);
buf  g1452 (n1481, n1346);
not  g1453 (n1485, n1341);
not  g1454 (n1460, n1331);
not  g1455 (n1446, n1341);
buf  g1456 (n1493, n1344);
not  g1457 (n1492, n1344);
buf  g1458 (n1457, n1349);
buf  g1459 (n1452, n1338);
buf  g1460 (n1497, n1348);
buf  g1461 (n1489, n1343);
not  g1462 (n1436, n1342);
not  g1463 (n1432, n1345);
not  g1464 (n1501, n1343);
buf  g1465 (n1488, n1333);
buf  g1466 (n1454, n1349);
buf  g1467 (n1476, n1342);
not  g1468 (n1466, n1340);
not  g1469 (n1443, n1347);
not  g1470 (n1461, n1335);
not  g1471 (n1509, n1458);
not  g1472 (n1523, n1456);
not  g1473 (n1512, n1452);
buf  g1474 (n1521, n1451);
not  g1475 (n1513, n1447);
nor  g1476 (n1515, n1440, n1234);
and  g1477 (n1527, n1452, n1235, n1454, n1455);
and  g1478 (n1508, n1452, n1449, n1234, n1455);
xor  g1479 (n1525, n1457, n1459, n1453, n1441);
nand g1480 (n1520, n1447, n1449, n1450, n1234);
or   g1481 (n1510, n1461, n1458, n1443, n1436);
and  g1482 (n1522, n1438, n1459, n1450, n1437);
nor  g1483 (n1506, n1453, n1461, n1430, n1455);
or   g1484 (n1517, n1457, n1460, n1439, n1456);
or   g1485 (n1524, n1235, n1454, n1453, n1451);
xor  g1486 (n1505, n1458, n1456, n1459, n1457);
xor  g1487 (n1519, n1454, n1432, n1450, n1448);
xor  g1488 (n1507, n1451, n1449, n1448, n1444);
nand g1489 (n1526, n1448, n1457, n1235, n1445);
xor  g1490 (n1518, n1435, n1433, n1456, n1431);
xor  g1491 (n1516, n1451, n1434, n1452, n1449);
xor  g1492 (n1514, n1442, n1459, n1448, n1458);
and  g1493 (n1504, n1455, n1446, n1450, n1453);
xor  g1494 (n1511, n1454, n1460);
and  g1495 (n1561, n1237, n1274, n1284, n1267);
or   g1496 (n1595, n1237, n1523, n1242, n1258);
xor  g1497 (n1563, n1241, n1253, n1510, n1505);
xor  g1498 (n1597, n1292, n1267, n1255, n1511);
xnor g1499 (n1570, n1306, n1298, n1303, n1258);
xnor g1500 (n1609, n1295, n1264, n1506, n1254);
and  g1501 (n1602, n1526, n1248, n1302, n1244);
nor  g1502 (n1545, n1304, n1268, n1270, n1525);
xor  g1503 (n1620, n1509, n1245, n1514, n1240);
or   g1504 (n1551, n1284, n1257, n1298, n1256);
or   g1505 (n1538, n1236, n1285, n1514, n1264);
nand g1506 (n1540, n1237, n1302, n1281, n1289);
nor  g1507 (n1608, n1293, n1245, n1285, n1254);
nor  g1508 (n1577, n1265, n1523, n1520, n1261);
nor  g1509 (n1532, n1299, n1277, n1284, n1283);
and  g1510 (n1553, n1237, n1287, n1301, n1521);
nand g1511 (n1548, n1306, n1282, n1285, n1288);
or   g1512 (n1556, n1522, n1296, n1526, n1271);
or   g1513 (n1569, n1270, n1519, n1275, n1246);
nand g1514 (n1610, n1512, n1524, n1516, n1527);
xnor g1515 (n1619, n1238, n1291, n1519, n1239);
nand g1516 (n1539, n1509, n1520, n1511, n1256);
xor  g1517 (n1550, n1250, n1290, n1303, n1305);
nand g1518 (n1566, n1509, n1282, n1280, n1278);
xor  g1519 (n1611, n1249, n1281, n1301, n1297);
nand g1520 (n1592, n1246, n1513, n1303, n1242);
or   g1521 (n1618, n1518, n1297, n1250, n1269);
nand g1522 (n1547, n1274, n1246, n1253, n1507);
nor  g1523 (n1613, n1525, n1292, n1289, n1242);
nand g1524 (n1575, n1517, n1281, n1251, n1265);
and  g1525 (n1591, n1236, n1249, n1513, n1514);
nor  g1526 (n1622, n1516, n1267, n1266);
xnor g1527 (n1586, n1278, n1243, n1513, n1288);
xnor g1528 (n1542, n1507, n1305, n1508, n1253);
and  g1529 (n1603, n1258, n1508, n1262, n1268);
nand g1530 (n1549, n1276, n1515, n1288, n1240);
nor  g1531 (n1546, n1515, n1300, n1270, n1526);
xor  g1532 (n1571, n1239, n1266, n1299, n1506);
xor  g1533 (n1562, n1270, n1291, n1522, n1252);
nand g1534 (n1607, n1516, n1287, n1284, n1291);
nand g1535 (n1541, n1504, n1510, n1293, n1275);
xor  g1536 (n1528, n1276, n1515, n1264, n1517);
xnor g1537 (n1580, n1265, n1246, n1255, n1259);
xor  g1538 (n1587, n1263, n1273, n1257, n1251);
nor  g1539 (n1601, n1504, n1296, n1300, n1299);
nand g1540 (n1579, n1301, n1266, n1241, n1277);
nor  g1541 (n1543, n1505, n1293, n1504, n1271);
xor  g1542 (n1573, n1263, n1307, n1255, n1507);
xnor g1543 (n1584, n1524, n1271, n1294, n1507);
xor  g1544 (n1576, n1514, n1238, n1282, n1526);
or   g1545 (n1554, n1295, n1236, n1260, n1524);
and  g1546 (n1567, n1292, n1295, n1263, n1274);
nand g1547 (n1568, n1522, n1258, n1251, n1240);
nor  g1548 (n1557, n1510, n1261, n1301, n1243);
nor  g1549 (n1552, n1306, n1302, n1298, n1519);
or   g1550 (n1616, n1275, n1518, n1520, n1506);
nand g1551 (n1564, n1512, n1265, n1254, n1518);
xnor g1552 (n1535, n1523, n1241, n1527, n1302);
xor  g1553 (n1593, n1511, n1294, n1292, n1260);
nand g1554 (n1529, n1273, n1300, n1253, n1291);
or   g1555 (n1590, n1260, n1249, n1286, n1513);
and  g1556 (n1581, n1269, n1244, n1286, n1243);
and  g1557 (n1544, n1250, n1283, n1506, n1248);
nand g1558 (n1536, n1243, n1524, n1257, n1242);
nor  g1559 (n1589, n1298, n1269, n1307, n1279);
xor  g1560 (n1558, n1255, n1262, n1304, n1240);
or   g1561 (n1598, n1260, n1282, n1305, n1278);
nor  g1562 (n1588, n1297, n1252, n1286);
xnor g1563 (n1600, n1527, n1273, n1521, n1293);
xnor g1564 (n1594, n1276, n1249, n1290, n1252);
nor  g1565 (n1623, n1286, n1256, n1272, n1280);
xnor g1566 (n1530, n1236, n1262, n1509, n1523);
and  g1567 (n1615, n1272, n1272, n1512, n1248);
nand g1568 (n1604, n1269, n1527, n1277, n1290);
and  g1569 (n1555, n1244, n1508, n1304, n1247);
nor  g1570 (n1621, n1504, n1266, n1275, n1245);
xor  g1571 (n1583, n1283, n1272, n1245, n1261);
and  g1572 (n1578, n1307, n1259, n1522);
nand g1573 (n1617, n1239, n1247, n1288, n1299);
xor  g1574 (n1572, n1515, n1300, n1281, n1248);
xor  g1575 (n1565, n1263, n1295, n1280, n1250);
xor  g1576 (n1596, n1289, n1254, n1510, n1251);
nor  g1577 (n1559, n1505, n1238, n1264, n1304);
or   g1578 (n1560, n1261, n1521, n1274, n1516);
nor  g1579 (n1606, n1279, n1508, n1262, n1287);
or   g1580 (n1582, n1268, n1287, n1289, n1505);
and  g1581 (n1612, n1256, n1277, n1276, n1280);
nor  g1582 (n1614, n1235, n1518, n1247, n1278);
xnor g1583 (n1599, n1285, n1305, n1290, n1279);
nand g1584 (n1534, n1520, n1238, n1511, n1521);
xnor g1585 (n1605, n1294, n1239, n1525, n1296);
nor  g1586 (n1585, n1303, n1517, n1273, n1297);
nor  g1587 (n1537, n1283, n1244, n1519, n1512);
xnor g1588 (n1574, n1294, n1296, n1525, n1241);
nor  g1589 (n1533, n1271, n1259, n1268, n1247);
nand g1590 (n1531, n1517, n1279, n1306, n1257);
not  g1591 (n1665, n1479);
buf  g1592 (n1834, n1359);
buf  g1593 (n1639, n1392);
not  g1594 (n1738, n1570);
buf  g1595 (n1628, n1360);
not  g1596 (n1836, n1602);
not  g1597 (n1864, n1584);
buf  g1598 (n1635, n1572);
not  g1599 (n1658, n1590);
buf  g1600 (n1670, n1574);
not  g1601 (n1809, n1463);
not  g1602 (n1831, n1529);
buf  g1603 (n1739, n1612);
not  g1604 (n1700, n1614);
not  g1605 (n1824, n1480);
buf  g1606 (n1690, n1599);
not  g1607 (n1727, n1403);
not  g1608 (n1710, n1592);
buf  g1609 (n1771, n1616);
buf  g1610 (n1862, n1587);
buf  g1611 (n1755, n1354);
not  g1612 (n1657, n1315);
not  g1613 (n1819, n1583);
not  g1614 (n1741, n1409);
buf  g1615 (n1785, n1534);
buf  g1616 (n1708, n1426);
not  g1617 (n1763, n1600);
not  g1618 (n1797, n1562);
buf  g1619 (n1817, n1566);
buf  g1620 (n1694, n1465);
buf  g1621 (n1717, n1572);
not  g1622 (n1669, n1399);
buf  g1623 (n1861, n1550);
buf  g1624 (n1753, n1308);
buf  g1625 (n1682, n1424);
buf  g1626 (n1769, n1475);
buf  g1627 (n1804, n1536);
buf  g1628 (n1858, n1621);
buf  g1629 (n1656, n1476);
buf  g1630 (n1730, n1350);
not  g1631 (n1848, n1365);
not  g1632 (n1662, n1398);
not  g1633 (n1679, n1480);
buf  g1634 (n1693, n1597);
not  g1635 (n1637, n1592);
not  g1636 (n1788, n1419);
buf  g1637 (n1705, n1594);
buf  g1638 (n1799, n1365);
not  g1639 (n1795, n1609);
not  g1640 (n1641, n1478);
not  g1641 (n1825, n1418);
not  g1642 (n1856, n1611);
buf  g1643 (n1852, n1549);
not  g1644 (n1750, n1356);
not  g1645 (n1860, n1480);
buf  g1646 (n1872, n1563);
buf  g1647 (n1828, n1416);
buf  g1648 (n1719, n1424);
not  g1649 (n1686, n1572);
buf  g1650 (n1840, n1559);
not  g1651 (n1640, n1478);
buf  g1652 (n1666, n1580);
buf  g1653 (n1815, n1426);
not  g1654 (n1777, n1545);
not  g1655 (n1807, n1414);
and  g1656 (n1655, n1557, n1611, n1551, n1559);
nand g1657 (n1742, n1588, n1396, n1571, n1355);
or   g1658 (n1636, n1364, n1312, n1367, n1620);
nor  g1659 (n1781, n1356, n1378, n1595, n1592);
nand g1660 (n1745, n1361, n1409, n1562, n1391);
xnor g1661 (n1849, n1544, n1565, n1528, n1546);
nor  g1662 (n1749, n1353, n1419, n1595, n1589);
nor  g1663 (n1695, n1552, n1587, n1317, n1463);
nand g1664 (n1699, n1354, n1362, n1397, n1382);
and  g1665 (n1687, n1528, n1386, n1363, n1366);
xor  g1666 (n1688, n1312, n1387, n1587, n1405);
xnor g1667 (n1878, n1609, n1403, n1574, n1476);
nor  g1668 (n1761, n1365, n1585, n1601, n1581);
and  g1669 (n1773, n1404, n1426, n1123, n1558);
xor  g1670 (n1783, n1554, n1384, n1125, n1597);
xor  g1671 (n1827, n1318, n1479, n1608, n1555);
or   g1672 (n1629, n1414, n1532, n1559, n1122);
or   g1673 (n1806, n1534, n1407, n1531, n1533);
or   g1674 (n1876, n1318, n1530, n1466, n1415);
and  g1675 (n1627, n1556, n1462, n1473, n1364);
nand g1676 (n1839, n1354, n1564, n1573, n1364);
xor  g1677 (n1718, n1422, n1365, n1468, n1586);
and  g1678 (n1652, n1465, n1590, n1552, n1386);
xor  g1679 (n1835, n1477, n1316, n1580, n1599);
xnor g1680 (n1683, n1568, n1607, n1582, n1609);
and  g1681 (n1638, n1469, n1471, n1551, n1320);
xor  g1682 (n1842, n1586, n1424, n1577, n1391);
xor  g1683 (n1782, n1409, n1568, n1616, n1467);
and  g1684 (n1814, n1405, n1608, n1610, n1535);
xnor g1685 (n1675, n1482, n1551, n1373, n1425);
nor  g1686 (n1855, n1399, n1384, n1355, n1468);
xor  g1687 (n1651, n1360, n1540, n1420, n1619);
xnor g1688 (n1731, n1368, n1418, n1416, n1569);
xor  g1689 (n1674, n1314, n1377, n1545, n1313);
xnor g1690 (n1633, n1623, n1310, n1604, n1359);
or   g1691 (n1676, n1584, n1429, n1360, n1575);
nand g1692 (n1709, n1398, n1475, n1593, n1584);
nand g1693 (n1646, n1597, n1583, n1591, n1354);
and  g1694 (n1768, n1577, n1566, n1376, n1545);
and  g1695 (n1793, n1400, n1604, n1319, n1575);
xnor g1696 (n1701, n1569, n1533, n1543, n1421);
nand g1697 (n1653, n1368, n1311, n1554, n1395);
xor  g1698 (n1772, n1618, n1549, n1368, n1558);
xor  g1699 (n1770, n1617, n1405, n1376, n1373);
or   g1700 (n1830, n1466, n1609, n1576, n1541);
or   g1701 (n1703, n1408, n1400, n1375, n1406);
and  g1702 (n1702, n1558, n1311, n1369, n1466);
xnor g1703 (n1780, n1320, n1622, n1546, n1410);
nand g1704 (n1882, n1385, n1549, n1429, n1586);
nand g1705 (n1845, n1565, n1352, n1578, n1375);
nand g1706 (n1854, n1422, n1309, n1542, n1319);
and  g1707 (n1654, n1316, n1530, n1470, n1557);
or   g1708 (n1649, n1482, n1548, n1413, n1380);
and  g1709 (n1812, n1553, n1531, n1403, n1585);
xor  g1710 (n1645, n1408, n1615, n1390, n1569);
and  g1711 (n1740, n1557, n1370, n1477, n1376);
xor  g1712 (n1767, n1395, n1368, n1394, n1425);
nand g1713 (n1885, n1464, n1470, n1535, n1471);
xor  g1714 (n1714, n1391, n1462, n1351, n1421);
xor  g1715 (n1877, n1562, n1410, n1462, n1579);
and  g1716 (n1648, n1398, n1598, n1587, n1538);
nor  g1717 (n1850, n1567, n1560, n1308, n1614);
nor  g1718 (n1837, n1543, n1566, n1390, n1409);
xnor g1719 (n1796, n1593, n1472, n1376);
nor  g1720 (n1778, n1411, n1623, n1541, n1588);
nand g1721 (n1677, n1411, n1467, n1355, n1316);
xor  g1722 (n1729, n1321, n1621, n1558, n1612);
or   g1723 (n1816, n1617, n1539, n1470, n1538);
and  g1724 (n1692, n1621, n1575, n1422, n1429);
xnor g1725 (n1764, n1320, n1399, n1546, n1581);
nand g1726 (n1671, n1424, n1464, n1372, n1623);
nand g1727 (n1846, n1595, n1571, n1407, n1576);
or   g1728 (n1791, n1483, n1378, n1388, n1537);
or   g1729 (n1681, n1528, n1547, n1573, n1590);
and  g1730 (n1685, n1530, n1538, n1314, n1532);
or   g1731 (n1680, n1374, n1541, n1473, n1355);
and  g1732 (n1863, n1547, n1481, n1402, n1412);
or   g1733 (n1874, n1567, n1540, n1481, n1380);
and  g1734 (n1833, n1591, n1357, n1613, n1367);
xnor g1735 (n1820, n1620, n1475, n1478, n1606);
and  g1736 (n1808, n1422, n1389, n1556, n1375);
xnor g1737 (n1625, n1601, n1381, n1546, n1470);
and  g1738 (n1643, n1552, n1602, n1531, n1564);
xor  g1739 (n1736, n1477, n1604, n1620, n1550);
or   g1740 (n1647, n1384, n1396, n1611, n1416);
xor  g1741 (n1873, n1612, n1359, n1377, n1483);
nand g1742 (n1713, n1529, n1314, n1463, n1420);
xnor g1743 (n1823, n1612, n1608, n1540, n1611);
xor  g1744 (n1841, n1469, n1561, n1351);
xnor g1745 (n1786, n1578, n1352, n1583, n1604);
nor  g1746 (n1821, n1588, n1564, n1465, n1599);
xnor g1747 (n1822, n1401, n1389, n1362, n1474);
xnor g1748 (n1720, n1413, n1322, n1317, n1363);
xor  g1749 (n1765, n1387, n1377, n1425, n1393);
nand g1750 (n1728, n1484, n1623, n1386, n1393);
nor  g1751 (n1744, n1388, n1428, n1610, n1473);
or   g1752 (n1758, n1571, n1351, n1366, n1402);
and  g1753 (n1704, n1381, n1426, n1559, n1532);
xor  g1754 (n1881, n1466, n1580, n1578, n1308);
nor  g1755 (n1724, n1579, n1393, n1577, n1581);
and  g1756 (n1867, n1381, n1383, n1531, n1608);
and  g1757 (n1696, n1565, n1462, n1550, n1321);
and  g1758 (n1868, n1575, n1360, n1555, n1556);
nor  g1759 (n1663, n1483, n1603, n1532, n1586);
nor  g1760 (n1747, n1370, n1423, n1548, n1478);
or   g1761 (n1803, n1400, n1616, n1412, n1469);
and  g1762 (n1829, n1313, n1571, n1362, n1350);
xor  g1763 (n1626, n1402, n1588, n1321, n1124);
xnor g1764 (n1660, n1574, n1483, n1370, n1404);
xor  g1765 (n1673, n1427, n1370, n1555, n1576);
and  g1766 (n1746, n1528, n1309, n1353, n1589);
and  g1767 (n1775, n1417, n1367, n1317, n1411);
or   g1768 (n1698, n1319, n1580, n1615);
xor  g1769 (n1844, n1356, n1534, n1579, n1363);
or   g1770 (n1684, n1382, n1379, n1613, n1384);
and  g1771 (n1801, n1393, n1585, n1390, n1572);
nand g1772 (n1800, n1594, n1315, n1473, n1603);
nand g1773 (n1866, n1394, n1582, n1379, n1351);
nand g1774 (n1659, n1463, n1385, n1421, n1383);
xnor g1775 (n1631, n1554, n1472, n1620, n1366);
or   g1776 (n1784, n1606, n1529, n1534, n1386);
xor  g1777 (n1813, n1569, n1353, n1543, n1392);
or   g1778 (n1787, n1464, n1421, n1621, n1307);
xor  g1779 (n1689, n1598, n1484, n1382, n1394);
xnor g1780 (n1735, n1482, n1544, n1401, n1601);
and  g1781 (n1733, n1361, n1619, n1547, n1467);
or   g1782 (n1805, n1539, n1406, n1591, n1573);
or   g1783 (n1706, n1542, n1357, n1471, n1610);
xor  g1784 (n1774, n1556, n1469, n1598, n1568);
xnor g1785 (n1794, n1120, n1539, n1589, n1364);
xor  g1786 (n1838, n1568, n1387, n1359, n1318);
xnor g1787 (n1756, n1428, n1603, n1385);
or   g1788 (n1650, n1312, n1603, n1318, n1420);
or   g1789 (n1859, n1536, n1613, n1408, n1479);
and  g1790 (n1715, n1406, n1419, n1121, n1540);
nor  g1791 (n1884, n1598, n1464, n1369, n1397);
nor  g1792 (n1678, n1552, n1602, n1581, n1423);
xnor g1793 (n1732, n1417, n1402, n1358, n1363);
or   g1794 (n1697, n1397, n1352, n1311, n1392);
or   g1795 (n1722, n1596, n1415, n1378, n1613);
xor  g1796 (n1726, n1596, n1474, n1388, n1472);
and  g1797 (n1887, n1412, n1563, n1389, n1383);
xnor g1798 (n1752, n1396, n1622, n1413, n1372);
nand g1799 (n1664, n1542, n1371, n1387, n1480);
or   g1800 (n1880, n1560, n1600, n1383, n1427);
nor  g1801 (n1879, n1419, n1405, n1554, n1411);
xnor g1802 (n1751, n1536, n1548, n1400, n1398);
nand g1803 (n1865, n1617, n1536, n1407, n1310);
or   g1804 (n1779, n1321, n1414, n1415, n1616);
nand g1805 (n1883, n1566, n1537, n1310, n1615);
or   g1806 (n1798, n1425, n1594, n1477, n1553);
xnor g1807 (n1851, n1481, n1535, n1563, n1375);
nor  g1808 (n1644, n1350, n1605, n1607, n1589);
and  g1809 (n1672, n1541, n1319, n1361, n1585);
xnor g1810 (n1634, n1372, n1423, n1570, n1427);
nor  g1811 (n1886, n1622, n1380, n1565, n1428);
xor  g1812 (n1630, n1551, n1468, n1369, n1560);
nor  g1813 (n1802, n1417, n1582, n1600, n1310);
and  g1814 (n1871, n1369, n1357, n1570, n1392);
xnor g1815 (n1642, n1371, n1322, n1547, n1394);
xnor g1816 (n1810, n1481, n1371, n1401);
nor  g1817 (n1716, n1395, n1417, n1429, n1555);
xnor g1818 (n1707, n1414, n1308, n1309, n1576);
xnor g1819 (n1754, n1601, n1418, n1361, n1529);
xnor g1820 (n1743, n1377, n1618, n1403, n1390);
nor  g1821 (n1748, n1482, n1408, n1476, n1316);
nand g1822 (n1737, n1600, n1471, n1607, n1476);
or   g1823 (n1760, n1583, n1593, n1557, n1315);
xnor g1824 (n1721, n1549, n1577, n1537, n1374);
xnor g1825 (n1789, n1533, n1597, n1410, n1561);
or   g1826 (n1869, n1605, n1622, n1353, n1320);
and  g1827 (n1632, n1542, n1382, n1607, n1563);
xnor g1828 (n1725, n1545, n1404, n1602, n1538);
and  g1829 (n1826, n1582, n1313, n1389, n1362);
nand g1830 (n1723, n1374, n1605, n1535, n1474);
and  g1831 (n1691, n1315, n1614, n1309, n1619);
nand g1832 (n1762, n1379, n1396, n1366, n1484);
xnor g1833 (n1766, n1617, n1474, n1412, n1605);
xnor g1834 (n1790, n1380, n1567, n1543, n1358);
xor  g1835 (n1759, n1381, n1591, n1420, n1573);
nand g1836 (n1776, n1395, n1567, n1404, n1388);
or   g1837 (n1832, n1606, n1374, n1314, n1311);
xnor g1838 (n1712, n1579, n1592, n1391, n1584);
xnor g1839 (n1853, n1410, n1593, n1461, n1416);
xor  g1840 (n1847, n1427, n1578, n1467, n1367);
nor  g1841 (n1811, n1544, n1356, n1399, n1397);
nor  g1842 (n1734, n1561, n1423, n1574, n1401);
or   g1843 (n1624, n1570, n1407, n1428, n1596);
nand g1844 (n1875, n1413, n1548, n1373, n1465);
and  g1845 (n1667, n1590, n1614, n1479, n1618);
nand g1846 (n1757, n1550, n1539, n1594, n1468);
nor  g1847 (n1870, n1606, n1317, n1564, n1560);
xor  g1848 (n1711, n1619, n1358, n1312, n1599);
xnor g1849 (n1668, n1595, n1415, n1378, n1553);
or   g1850 (n1792, n1313, n1618, n1379, n1537);
nor  g1851 (n1843, n1475, n1544, n1610, n1596);
xor  g1852 (n1661, n1358, n1418, n1357, n1530);
nand g1853 (n1818, n1372, n1533, n1562, n1373);
nand g1854 (n1857, n1461, n1406, n1553, n1352);
or   g1855 (n1899, n1671, n1647, n1733, n1643);
nand g1856 (n1909, n1674, n1633, n1665, n1646);
and  g1857 (n1908, n1635, n1638, n1673, n1737);
nand g1858 (n1890, n1723, n1651, n1712, n1677);
or   g1859 (n1892, n1696, n1714, n1672, n1710);
nor  g1860 (n1904, n1730, n1658, n1653, n1655);
and  g1861 (n1903, n1742, n1705, n1641, n1642);
or   g1862 (n1906, n1703, n1711, n1740, n1729);
xor  g1863 (n1901, n1700, n1727, n1720, n1670);
xnor g1864 (n1900, n1636, n1690, n1676, n1750);
and  g1865 (n1889, n1741, n1666, n1664, n1718);
xnor g1866 (n1894, n1732, n1708, n1744, n1687);
xor  g1867 (n1914, n1688, n1699, n1731, n1650);
nor  g1868 (n1898, n1660, n1656, n1679, n1663);
nor  g1869 (n1913, n1667, n1686, n1652, n1697);
nor  g1870 (n1907, n1748, n1702, n1725, n1685);
or   g1871 (n1915, n1715, n1644, n1639, n1648);
and  g1872 (n1888, n1735, n1689, n1661, n1722);
xor  g1873 (n1891, n1649, n1717, n1706, n1728);
or   g1874 (n1911, n1675, n1657, n1747, n1640);
nand g1875 (n1905, n1694, n1745, n1743, n1707);
nor  g1876 (n1902, n1716, n1726, n1701, n1662);
nor  g1877 (n1917, n1682, n1669, n1746, n1724);
nand g1878 (n1893, n1738, n1637, n1634, n1698);
xnor g1879 (n1895, n1739, n1692, n1645, n1654);
nand g1880 (n1916, n1704, n1693, n1751, n1736);
xor  g1881 (n1910, n1749, n1668, n1719, n1659);
xor  g1882 (n1897, n1691, n1695, n1734, n1713);
and  g1883 (n1912, n1681, n1752, n1721, n1684);
and  g1884 (n1896, n1683, n1709, n1678, n1680);
nand g1885 (n1941, n1837, n1817, n1900, n1916);
xor  g1886 (n1939, n1812, n1763, n1901, n1899);
nor  g1887 (n1926, n1775, n1807, n1907, n1903);
or   g1888 (n1944, n1829, n1799, n1801, n1784);
or   g1889 (n1933, n1766, n1781, n1838, n1791);
and  g1890 (n1945, n1841, n1805, n1811, n1789);
or   g1891 (n1942, n1843, n1814, n1760, n1764);
nand g1892 (n1946, n1772, n1754, n1792, n1819);
nand g1893 (n1948, n1800, n1910, n1902, n1757);
xor  g1894 (n1931, n1786, n1828, n1777, n1911);
and  g1895 (n1918, n1787, n1780, n1844, n1771);
nor  g1896 (n1929, n1917, n1822, n1768, n1836);
nand g1897 (n1927, n1826, n1906, n1794, n1904);
and  g1898 (n1936, n1897, n1840, n1825, n1783);
xnor g1899 (n1935, n1773, n1815, n1898, n1782);
or   g1900 (n1938, n1917, n1821, n1756, n1761);
and  g1901 (n1940, n1788, n1755, n1830, n1809);
nor  g1902 (n1937, n1824, n1758, n1767, n1917);
or   g1903 (n1947, n1895, n1804, n1833, n1823);
nor  g1904 (n1922, n1802, n1842, n1806, n1916);
or   g1905 (n1924, n1776, n1762, n1896, n1891);
xor  g1906 (n1925, n1914, n1778, n1915, n1779);
nor  g1907 (n1932, n1795, n1913, n1892, n1905);
xor  g1908 (n1920, n1816, n1810, n1835, n1818);
and  g1909 (n1921, n1793, n1909, n1831, n1894);
nand g1910 (n1934, n1839, n1845, n1797, n1759);
nor  g1911 (n1923, n1820, n1834, n1893, n1832);
nand g1912 (n1928, n1790, n1803, n1753, n1769);
or   g1913 (n1943, n1796, n1785, n1917, n1908);
and  g1914 (n1919, n1770, n1808, n1798, n1813);
and  g1915 (n1930, n1765, n1827, n1774, n1912);
nor  g1916 (n1951, n1323, n1938, n1128, n1134);
nor  g1917 (n1949, n1940, n1324, n1937, n1846);
nor  g1918 (n1952, n1323, n1136, n1935, n1133);
xor  g1919 (n1955, n1323, n1324, n1130, n1932);
and  g1920 (n1956, n1324, n1126, n1934, n1936);
xnor g1921 (n1954, n1135, n1939, n1933, n1131);
and  g1922 (n1953, n1323, n1942, n1322);
xor  g1923 (n1950, n1127, n1132, n1129, n1941);
nand g1924 (n1960, n1325, n1325, n1951, n1852);
nand g1925 (n1958, n1847, n1851, n1853, n1850);
or   g1926 (n1959, n1950, n1324, n1855, n1848);
nor  g1927 (n1961, n1949, n1849, n1854, n1857);
nor  g1928 (n1957, n1325, n1952, n1953, n1856);
not  g1929 (n1962, n1957);
buf  g1930 (n1965, n1958);
buf  g1931 (n1964, n1959);
not  g1932 (n1963, n1960);
xor  g1933 (n1967, n1964, n1965);
nand g1934 (n1977, n1870, n1869);
and  g1935 (n1972, n1866, n1963, n1326);
xnor g1936 (n1968, n1963, n1964, n1945);
nand g1937 (n1970, n1943, n1965, n1865);
xor  g1938 (n1966, n1871, n1864, n1862);
or   g1939 (n1969, n1962, n1860, n1963);
xnor g1940 (n1973, n1962, n1326, n1863);
and  g1941 (n1979, n1868, n1948, n1961);
and  g1942 (n1978, n1867, n1325, n1965);
nand g1943 (n1975, n1965, n1944, n1963);
and  g1944 (n1976, n1861, n1946, n1947);
nor  g1945 (n1974, n1872, n1326, n1858);
nor  g1946 (n1971, n1859, n1964);
xnor g1947 (n1980, n1978, n1487, n1976, n1977);
xnor g1948 (n1982, n1503, n1881, n1495, n1488);
and  g1949 (n2012, n1878, n1873, n1492, n1979);
or   g1950 (n1991, n1974, n1977, n1485, n1490);
xnor g1951 (n2003, n1486, n1503, n1489, n1954);
xnor g1952 (n1998, n1495, n1494, n1882, n1883);
xor  g1953 (n1995, n1876, n1489, n1497, n1972);
xnor g1954 (n1999, n1977, n1491, n1971, n1500);
xnor g1955 (n1986, n1491, n1499, n1882, n1976);
xnor g1956 (n1989, n1501, n1979, n1489, n1975);
nor  g1957 (n2011, n1877, n1974, n1485, n1973);
or   g1958 (n1994, n1488, n1975, n1487, n1979);
xnor g1959 (n1990, n1486, n1498, n1492, n1497);
nor  g1960 (n2009, n1884, n1137, n1487, n1503);
xnor g1961 (n2004, n1502, n1972, n1491, n1490);
xnor g1962 (n1992, n1979, n1497, n1485, n1491);
nand g1963 (n2001, n1486, n1502, n1975, n1495);
and  g1964 (n2007, n1492, n1503, n1972, n1489);
and  g1965 (n1984, n1487, n1973, n1500, n1497);
nor  g1966 (n1985, n1138, n1875, n1485, n1883);
xor  g1967 (n1981, n1973, n1493, n1502);
or   g1968 (n2005, n1879, n1496, n1498, n1493);
xor  g1969 (n1987, n1499, n1493, n1139, n1492);
nand g1970 (n1993, n1486, n1502, n1973, n1495);
and  g1971 (n1988, n1499, n1498, n1976, n1956);
nor  g1972 (n2010, n1496, n1484, n1881, n1490);
and  g1973 (n2008, n1874, n1496, n1494, n1500);
nand g1974 (n2002, n1490, n1501, n1955, n1884);
nand g1975 (n1997, n1500, n1974, n1972, n1498);
nand g1976 (n2000, n1488, n1978, n1501);
xnor g1977 (n2006, n1880, n1974, n1499, n1978);
nand g1978 (n1983, n1978, n1488, n1494);
nand g1979 (n1996, n1976, n1496, n1975, n1977);
xor  g1980 (n2016, n1327, n1987, n1986, n2003);
nand g1981 (n2013, n1992, n1145, n1990, n1983);
xnor g1982 (n2021, n672, n1887, n1144);
or   g1983 (n2025, n2005, n1150, n1885, n1998);
nand g1984 (n2024, n1143, n1326, n1989, n2009);
nor  g1985 (n2020, n1146, n1981, n1886, n1887);
nand g1986 (n2023, n1151, n1153, n1152, n1140);
and  g1987 (n2019, n1980, n2002, n1885, n2012);
xnor g1988 (n2027, n1327, n2006, n1996, n1995);
or   g1989 (n2014, n1985, n1994, n1993, n2008);
xor  g1990 (n2022, n2004, n1327, n2010, n2000);
nor  g1991 (n2015, n1142, n1997, n2007, n1141);
nand g1992 (n2017, n2001, n1147, n1149, n1988);
and  g1993 (n2026, n1984, n1999, n1886, n1982);
nor  g1994 (n2018, n1148, n1327, n2011, n1991);
nand g1995 (n2031, n2026, n2023, n2027, n2014);
or   g1996 (n2029, n2024, n2021, n2018, n2016);
nand g1997 (n2028, n2020, n2015, n1887, n2017);
and  g1998 (n2030, n2022, n2025, n2013, n2019);
xor  g1999 (n2032, n2031, n2028, n2029, n2030);
endmodule
