

module Stat_1027_28_12
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n769,
  n767,
  n762,
  n815,
  n819,
  n822,
  n821,
  n811,
  n814,
  n817,
  n823,
  n824,
  n816,
  n810,
  n830,
  n1060,
  n1051,
  n1063,
  n1064,
  n1061,
  n1054,
  n1062,
  n1050,
  n1056,
  n1066,
  n1059,
  n1058,
  n1053,
  n1057,
  n1065,
  n1052,
  n1055
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n769;output n767;output n762;output n815;output n819;output n822;output n821;output n811;output n814;output n817;output n823;output n824;output n816;output n810;output n830;output n1060;output n1051;output n1063;output n1064;output n1061;output n1054;output n1062;output n1050;output n1056;output n1066;output n1059;output n1058;output n1053;output n1057;output n1065;output n1052;output n1055;
  wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n763;wire n764;wire n765;wire n766;wire n768;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n812;wire n813;wire n818;wire n820;wire n825;wire n826;wire n827;wire n828;wire n829;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  buf
  g0
  (
    n41,
    n12
  );


  not
  g1
  (
    n59,
    n1
  );


  not
  g2
  (
    n68,
    n5
  );


  buf
  g3
  (
    n67,
    n10
  );


  not
  g4
  (
    n52,
    n6
  );


  not
  g5
  (
    n47,
    n4
  );


  not
  g6
  (
    n48,
    n10
  );


  buf
  g7
  (
    n50,
    n7
  );


  buf
  g8
  (
    n40,
    n1
  );


  buf
  g9
  (
    n56,
    n13
  );


  not
  g10
  (
    n66,
    n9
  );


  buf
  g11
  (
    n43,
    n13
  );


  buf
  g12
  (
    n58,
    n15
  );


  buf
  g13
  (
    n63,
    n8
  );


  not
  g14
  (
    n45,
    n3
  );


  buf
  g15
  (
    n49,
    n7
  );


  buf
  g16
  (
    n53,
    n9
  );


  buf
  g17
  (
    n54,
    n14
  );


  buf
  g18
  (
    n55,
    n6
  );


  buf
  g19
  (
    n42,
    n5
  );


  not
  g20
  (
    n44,
    n2
  );


  buf
  g21
  (
    n65,
    n4
  );


  not
  g22
  (
    KeyWire_0_1,
    n12
  );


  buf
  g23
  (
    n64,
    n2
  );


  not
  g24
  (
    n57,
    n8
  );


  not
  g25
  (
    n51,
    n14
  );


  buf
  g26
  (
    n46,
    n15
  );


  buf
  g27
  (
    n69,
    n11
  );


  buf
  g28
  (
    n61,
    n11
  );


  buf
  g29
  (
    n62,
    n3
  );


  buf
  g30
  (
    n88,
    n62
  );


  not
  g31
  (
    n103,
    n54
  );


  not
  g32
  (
    n140,
    n49
  );


  buf
  g33
  (
    n131,
    n45
  );


  not
  g34
  (
    KeyWire_0_2,
    n57
  );


  not
  g35
  (
    n137,
    n48
  );


  not
  g36
  (
    n159,
    n42
  );


  not
  g37
  (
    n76,
    n64
  );


  buf
  g38
  (
    n177,
    n43
  );


  not
  g39
  (
    n115,
    n43
  );


  not
  g40
  (
    n119,
    n57
  );


  not
  g41
  (
    n87,
    n42
  );


  not
  g42
  (
    n124,
    n44
  );


  buf
  g43
  (
    n164,
    n58
  );


  not
  g44
  (
    n166,
    n66
  );


  not
  g45
  (
    n171,
    n51
  );


  not
  g46
  (
    n114,
    n66
  );


  buf
  g47
  (
    n134,
    n67
  );


  not
  g48
  (
    n121,
    n60
  );


  not
  g49
  (
    n75,
    n58
  );


  buf
  g50
  (
    n150,
    n45
  );


  not
  g51
  (
    n71,
    n66
  );


  not
  g52
  (
    n130,
    n50
  );


  buf
  g53
  (
    KeyWire_0_11,
    n46
  );


  not
  g54
  (
    n145,
    n41
  );


  buf
  g55
  (
    n162,
    n52
  );


  not
  g56
  (
    n123,
    n16
  );


  not
  g57
  (
    n111,
    n52
  );


  not
  g58
  (
    n94,
    n63
  );


  not
  g59
  (
    n156,
    n50
  );


  buf
  g60
  (
    n73,
    n48
  );


  buf
  g61
  (
    n174,
    n41
  );


  buf
  g62
  (
    n92,
    n59
  );


  not
  g63
  (
    n81,
    n67
  );


  not
  g64
  (
    n95,
    n53
  );


  buf
  g65
  (
    n146,
    n52
  );


  buf
  g66
  (
    n90,
    n56
  );


  buf
  g67
  (
    n169,
    n60
  );


  buf
  g68
  (
    n70,
    n50
  );


  buf
  g69
  (
    n147,
    n42
  );


  buf
  g70
  (
    n112,
    n52
  );


  not
  g71
  (
    n93,
    n42
  );


  buf
  g72
  (
    n125,
    n16
  );


  buf
  g73
  (
    n126,
    n63
  );


  buf
  g74
  (
    n89,
    n55
  );


  not
  g75
  (
    n101,
    n55
  );


  not
  g76
  (
    n98,
    n47
  );


  buf
  g77
  (
    n182,
    n46
  );


  buf
  g78
  (
    n136,
    n48
  );


  buf
  g79
  (
    n108,
    n59
  );


  not
  g80
  (
    n122,
    n49
  );


  buf
  g81
  (
    n77,
    n64
  );


  buf
  g82
  (
    n173,
    n41
  );


  not
  g83
  (
    n82,
    n40
  );


  not
  g84
  (
    n152,
    n46
  );


  buf
  g85
  (
    n99,
    n62
  );


  not
  g86
  (
    n167,
    n62
  );


  buf
  g87
  (
    n72,
    n57
  );


  buf
  g88
  (
    n165,
    n51
  );


  not
  g89
  (
    n153,
    n67
  );


  buf
  g90
  (
    n109,
    n49
  );


  not
  g91
  (
    n151,
    n63
  );


  buf
  g92
  (
    n179,
    n50
  );


  not
  g93
  (
    n170,
    n57
  );


  not
  g94
  (
    n163,
    n66
  );


  not
  g95
  (
    n102,
    n55
  );


  buf
  g96
  (
    n138,
    n61
  );


  buf
  g97
  (
    n157,
    n62
  );


  not
  g98
  (
    n158,
    n63
  );


  not
  g99
  (
    n100,
    n53
  );


  not
  g100
  (
    n149,
    n61
  );


  buf
  g101
  (
    n113,
    n65
  );


  buf
  g102
  (
    n116,
    n65
  );


  not
  g103
  (
    n106,
    n44
  );


  buf
  g104
  (
    n154,
    n53
  );


  not
  g105
  (
    n78,
    n65
  );


  not
  g106
  (
    n83,
    n53
  );


  not
  g107
  (
    n161,
    n58
  );


  not
  g108
  (
    n117,
    n40
  );


  buf
  g109
  (
    n104,
    n40
  );


  not
  g110
  (
    n180,
    n67
  );


  buf
  g111
  (
    n80,
    n47
  );


  buf
  g112
  (
    n178,
    n56
  );


  buf
  g113
  (
    n175,
    n17
  );


  not
  g114
  (
    n144,
    n54
  );


  not
  g115
  (
    n181,
    n51
  );


  buf
  g116
  (
    n84,
    n59
  );


  buf
  g117
  (
    n155,
    n51
  );


  not
  g118
  (
    n74,
    n56
  );


  buf
  g119
  (
    n91,
    n64
  );


  not
  g120
  (
    n86,
    n61
  );


  not
  g121
  (
    n139,
    n46
  );


  buf
  g122
  (
    n160,
    n17
  );


  buf
  g123
  (
    n105,
    n44
  );


  not
  g124
  (
    n176,
    n45
  );


  not
  g125
  (
    n168,
    n49
  );


  buf
  g126
  (
    n142,
    n48
  );


  buf
  g127
  (
    n110,
    n41
  );


  not
  g128
  (
    n148,
    n43
  );


  not
  g129
  (
    n143,
    n68
  );


  not
  g130
  (
    n127,
    n45
  );


  not
  g131
  (
    n172,
    n54
  );


  buf
  g132
  (
    n133,
    n65
  );


  buf
  g133
  (
    KeyWire_0_13,
    n55
  );


  buf
  g134
  (
    n141,
    n59
  );


  buf
  g135
  (
    n129,
    n60
  );


  not
  g136
  (
    n85,
    n43
  );


  buf
  g137
  (
    n79,
    n54
  );


  xor
  g138
  (
    n132,
    n56,
    n58
  );


  not
  g139
  (
    n97,
    n47
  );


  nor
  g140
  (
    n128,
    n64,
    n40
  );


  and
  g141
  (
    n135,
    n61,
    n18
  );


  and
  g142
  (
    n120,
    n44,
    n60
  );


  buf
  g143
  (
    n264,
    n77
  );


  buf
  g144
  (
    n218,
    n71
  );


  not
  g145
  (
    n255,
    n116
  );


  not
  g146
  (
    n402,
    n22
  );


  buf
  g147
  (
    n195,
    n74
  );


  not
  g148
  (
    n288,
    n73
  );


  not
  g149
  (
    n366,
    n123
  );


  not
  g150
  (
    n368,
    n20
  );


  not
  g151
  (
    n290,
    n104
  );


  buf
  g152
  (
    n370,
    n76
  );


  not
  g153
  (
    n381,
    n93
  );


  buf
  g154
  (
    n231,
    n113
  );


  not
  g155
  (
    n353,
    n114
  );


  buf
  g156
  (
    n286,
    n95
  );


  buf
  g157
  (
    n317,
    n121
  );


  not
  g158
  (
    n310,
    n68
  );


  not
  g159
  (
    n365,
    n123
  );


  not
  g160
  (
    n320,
    n121
  );


  buf
  g161
  (
    n340,
    n26
  );


  not
  g162
  (
    n240,
    n111
  );


  not
  g163
  (
    n394,
    n106
  );


  buf
  g164
  (
    n335,
    n30
  );


  buf
  g165
  (
    n345,
    n103
  );


  not
  g166
  (
    n208,
    n69
  );


  buf
  g167
  (
    n346,
    n84
  );


  buf
  g168
  (
    n247,
    n110
  );


  buf
  g169
  (
    n197,
    n101
  );


  buf
  g170
  (
    n200,
    n76
  );


  not
  g171
  (
    n403,
    n126
  );


  buf
  g172
  (
    n262,
    n84
  );


  buf
  g173
  (
    n324,
    n99
  );


  not
  g174
  (
    n216,
    n83
  );


  buf
  g175
  (
    n242,
    n19
  );


  buf
  g176
  (
    n331,
    n117
  );


  buf
  g177
  (
    n246,
    n78
  );


  buf
  g178
  (
    n226,
    n77
  );


  buf
  g179
  (
    n248,
    n88
  );


  not
  g180
  (
    n251,
    n94
  );


  buf
  g181
  (
    n260,
    n91
  );


  buf
  g182
  (
    n296,
    n23
  );


  buf
  g183
  (
    n308,
    n109
  );


  not
  g184
  (
    n285,
    n124
  );


  buf
  g185
  (
    n322,
    n89
  );


  buf
  g186
  (
    n344,
    n118
  );


  buf
  g187
  (
    n342,
    n113
  );


  not
  g188
  (
    n193,
    n126
  );


  buf
  g189
  (
    n404,
    n117
  );


  buf
  g190
  (
    n333,
    n114
  );


  buf
  g191
  (
    n327,
    n100
  );


  not
  g192
  (
    n241,
    n96
  );


  not
  g193
  (
    n228,
    n82
  );


  buf
  g194
  (
    n237,
    n74
  );


  not
  g195
  (
    n258,
    n122
  );


  not
  g196
  (
    n371,
    n85
  );


  not
  g197
  (
    n254,
    n25
  );


  not
  g198
  (
    n232,
    n92
  );


  buf
  g199
  (
    n294,
    n71
  );


  not
  g200
  (
    n211,
    n90
  );


  not
  g201
  (
    n406,
    n102
  );


  not
  g202
  (
    n362,
    n69
  );


  buf
  g203
  (
    n321,
    n72
  );


  not
  g204
  (
    n385,
    n78
  );


  not
  g205
  (
    n401,
    n115
  );


  buf
  g206
  (
    n309,
    n98
  );


  buf
  g207
  (
    n319,
    n71
  );


  buf
  g208
  (
    n348,
    n115
  );


  buf
  g209
  (
    n313,
    n68
  );


  not
  g210
  (
    n206,
    n73
  );


  buf
  g211
  (
    n379,
    n79
  );


  not
  g212
  (
    KeyWire_0_6,
    n123
  );


  buf
  g213
  (
    n257,
    n108
  );


  not
  g214
  (
    n374,
    n107
  );


  not
  g215
  (
    n358,
    n111
  );


  buf
  g216
  (
    n219,
    n24
  );


  not
  g217
  (
    n350,
    n125
  );


  not
  g218
  (
    n210,
    n106
  );


  not
  g219
  (
    n217,
    n85
  );


  not
  g220
  (
    n187,
    n103
  );


  buf
  g221
  (
    n375,
    n94
  );


  buf
  g222
  (
    n279,
    n84
  );


  not
  g223
  (
    n407,
    n102
  );


  buf
  g224
  (
    n227,
    n19
  );


  buf
  g225
  (
    n273,
    n75
  );


  buf
  g226
  (
    n334,
    n95
  );


  buf
  g227
  (
    n305,
    n81
  );


  not
  g228
  (
    n389,
    n118
  );


  not
  g229
  (
    n192,
    n110
  );


  buf
  g230
  (
    n399,
    n76
  );


  not
  g231
  (
    n220,
    n101
  );


  buf
  g232
  (
    n300,
    n112
  );


  not
  g233
  (
    n269,
    n88
  );


  buf
  g234
  (
    n297,
    n111
  );


  buf
  g235
  (
    n198,
    n77
  );


  buf
  g236
  (
    n222,
    n104
  );


  not
  g237
  (
    n304,
    n92
  );


  not
  g238
  (
    n386,
    n109
  );


  buf
  g239
  (
    n225,
    n72
  );


  buf
  g240
  (
    n337,
    n102
  );


  not
  g241
  (
    n359,
    n99
  );


  not
  g242
  (
    n190,
    n115
  );


  buf
  g243
  (
    n376,
    n124
  );


  buf
  g244
  (
    n214,
    n105
  );


  buf
  g245
  (
    n265,
    n115
  );


  not
  g246
  (
    KeyWire_0_9,
    n78
  );


  buf
  g247
  (
    n189,
    n108
  );


  buf
  g248
  (
    n291,
    n120
  );


  buf
  g249
  (
    n382,
    n73
  );


  not
  g250
  (
    n377,
    n24
  );


  not
  g251
  (
    n356,
    n94
  );


  buf
  g252
  (
    n184,
    n18
  );


  buf
  g253
  (
    n263,
    n110
  );


  buf
  g254
  (
    n280,
    n77
  );


  not
  g255
  (
    n328,
    n74
  );


  buf
  g256
  (
    n292,
    n97
  );


  not
  g257
  (
    n205,
    n86
  );


  not
  g258
  (
    n229,
    n87
  );


  buf
  g259
  (
    n405,
    n70
  );


  not
  g260
  (
    n387,
    n119
  );


  not
  g261
  (
    n398,
    n111
  );


  not
  g262
  (
    n277,
    n72
  );


  not
  g263
  (
    n278,
    n72
  );


  not
  g264
  (
    n256,
    n121
  );


  buf
  g265
  (
    n338,
    n68
  );


  buf
  g266
  (
    n349,
    n118
  );


  not
  g267
  (
    n325,
    n71
  );


  not
  g268
  (
    n261,
    n100
  );


  buf
  g269
  (
    n276,
    n114
  );


  not
  g270
  (
    n303,
    n75
  );


  buf
  g271
  (
    n293,
    n98
  );


  buf
  g272
  (
    n185,
    n27
  );


  not
  g273
  (
    n207,
    n87
  );


  buf
  g274
  (
    n196,
    n105
  );


  buf
  g275
  (
    n272,
    n116
  );


  buf
  g276
  (
    n253,
    n106
  );


  buf
  g277
  (
    n336,
    n80
  );


  buf
  g278
  (
    n239,
    n112
  );


  not
  g279
  (
    n312,
    n121
  );


  buf
  g280
  (
    n224,
    n85
  );


  not
  g281
  (
    n383,
    n110
  );


  not
  g282
  (
    n183,
    n70
  );


  not
  g283
  (
    n400,
    n122
  );


  buf
  g284
  (
    n347,
    n123
  );


  not
  g285
  (
    n364,
    n81
  );


  not
  g286
  (
    n409,
    n105
  );


  not
  g287
  (
    n318,
    n76
  );


  not
  g288
  (
    n270,
    n98
  );


  not
  g289
  (
    n281,
    n80
  );


  buf
  g290
  (
    n355,
    n70
  );


  not
  g291
  (
    n212,
    n87
  );


  not
  g292
  (
    n289,
    n28
  );


  buf
  g293
  (
    n373,
    n122
  );


  not
  g294
  (
    n267,
    n88
  );


  buf
  g295
  (
    n250,
    n100
  );


  buf
  g296
  (
    n343,
    n105
  );


  buf
  g297
  (
    n384,
    n124
  );


  not
  g298
  (
    n213,
    n109
  );


  buf
  g299
  (
    n266,
    n97
  );


  buf
  g300
  (
    n245,
    n101
  );


  buf
  g301
  (
    n298,
    n119
  );


  buf
  g302
  (
    n369,
    n113
  );


  buf
  g303
  (
    n352,
    n83
  );


  not
  g304
  (
    n186,
    n83
  );


  buf
  g305
  (
    n363,
    n126
  );


  not
  g306
  (
    n307,
    n118
  );


  buf
  g307
  (
    n282,
    n93
  );


  buf
  g308
  (
    n188,
    n106
  );


  buf
  g309
  (
    n199,
    n75
  );


  not
  g310
  (
    n203,
    n80
  );


  buf
  g311
  (
    n271,
    n116
  );


  not
  g312
  (
    n194,
    n116
  );


  not
  g313
  (
    n259,
    n79
  );


  buf
  g314
  (
    n249,
    n83
  );


  not
  g315
  (
    n341,
    n120
  );


  buf
  g316
  (
    n299,
    n21
  );


  not
  g317
  (
    n332,
    n109
  );


  not
  g318
  (
    n201,
    n27
  );


  buf
  g319
  (
    n380,
    n95
  );


  buf
  g320
  (
    n360,
    n79
  );


  buf
  g321
  (
    n390,
    n90
  );


  not
  g322
  (
    n388,
    n96
  );


  not
  g323
  (
    n230,
    n120
  );


  buf
  g324
  (
    n215,
    n112
  );


  buf
  g325
  (
    n223,
    n96
  );


  not
  g326
  (
    n396,
    n93
  );


  not
  g327
  (
    n354,
    n89
  );


  not
  g328
  (
    n316,
    n84
  );


  buf
  g329
  (
    n284,
    n82
  );


  not
  g330
  (
    n287,
    n125
  );


  not
  g331
  (
    n392,
    n86
  );


  buf
  g332
  (
    n372,
    n92
  );


  buf
  g333
  (
    n391,
    n23
  );


  buf
  g334
  (
    KeyWire_0_5,
    n91
  );


  buf
  g335
  (
    n339,
    n86
  );


  buf
  g336
  (
    n393,
    n73
  );


  not
  g337
  (
    n314,
    n85
  );


  not
  g338
  (
    n302,
    n28
  );


  not
  g339
  (
    n315,
    n20
  );


  not
  g340
  (
    n351,
    n96
  );


  not
  g341
  (
    n235,
    n29
  );


  buf
  g342
  (
    n191,
    n82
  );


  not
  g343
  (
    n283,
    n108
  );


  not
  g344
  (
    n252,
    n122
  );


  not
  g345
  (
    n268,
    n107
  );


  not
  g346
  (
    n397,
    n125
  );


  not
  g347
  (
    n244,
    n92
  );


  buf
  g348
  (
    KeyWire_0_7,
    n108
  );


  not
  g349
  (
    KeyWire_0_10,
    n117
  );


  not
  g350
  (
    n243,
    n103
  );


  not
  g351
  (
    n378,
    n89
  );


  buf
  g352
  (
    n330,
    n86
  );


  buf
  g353
  (
    n221,
    n107
  );


  not
  g354
  (
    n209,
    n113
  );


  not
  g355
  (
    n275,
    n94
  );


  not
  g356
  (
    n234,
    n89
  );


  not
  g357
  (
    n295,
    n119
  );


  not
  g358
  (
    n236,
    n75
  );


  not
  g359
  (
    n311,
    n99
  );


  nor
  g360
  (
    n202,
    n103,
    n95,
    n93
  );


  xor
  g361
  (
    n238,
    n74,
    n21,
    n22,
    n104
  );


  xor
  g362
  (
    n326,
    n125,
    n100,
    n91
  );


  xnor
  g363
  (
    n274,
    n81,
    n78,
    n120,
    n25
  );


  or
  g364
  (
    n233,
    n119,
    n81,
    n80,
    n88
  );


  nor
  g365
  (
    n323,
    n112,
    n82,
    n98,
    n104
  );


  xnor
  g366
  (
    n301,
    n114,
    n70,
    n97,
    n29
  );


  and
  g367
  (
    n367,
    n117,
    n79,
    n90,
    n97
  );


  xor
  g368
  (
    n361,
    n107,
    n90,
    n87,
    n102
  );


  or
  g369
  (
    n408,
    n101,
    n124,
    n99,
    n26
  );


  buf
  g370
  (
    n459,
    n35
  );


  buf
  g371
  (
    n421,
    n192
  );


  buf
  g372
  (
    n589,
    n197
  );


  not
  g373
  (
    n578,
    n161
  );


  not
  g374
  (
    n604,
    n133
  );


  not
  g375
  (
    n422,
    n256
  );


  not
  g376
  (
    n591,
    n146
  );


  buf
  g377
  (
    n609,
    n141
  );


  buf
  g378
  (
    n460,
    n269
  );


  buf
  g379
  (
    n575,
    n221
  );


  nor
  g380
  (
    n512,
    n313,
    n335,
    n243
  );


  or
  g381
  (
    n440,
    n211,
    n379,
    n144,
    n152
  );


  xor
  g382
  (
    n583,
    n130,
    n316,
    n348,
    n222
  );


  and
  g383
  (
    n630,
    n366,
    n387,
    n234,
    n142
  );


  and
  g384
  (
    n449,
    n322,
    n230,
    n360,
    n138
  );


  nand
  g385
  (
    n484,
    n149,
    n187,
    n346,
    n126
  );


  xnor
  g386
  (
    n542,
    n186,
    n352,
    n164,
    n259
  );


  xor
  g387
  (
    n553,
    n155,
    n345,
    n309,
    n282
  );


  xor
  g388
  (
    n615,
    n194,
    n170,
    n268,
    n196
  );


  nor
  g389
  (
    n534,
    n326,
    n163,
    n370,
    n388
  );


  nand
  g390
  (
    n446,
    n238,
    n373,
    n198
  );


  xor
  g391
  (
    n582,
    n309,
    n158,
    n142,
    n393
  );


  xor
  g392
  (
    n586,
    n318,
    n359,
    n136,
    n233
  );


  nand
  g393
  (
    n562,
    n226,
    n262,
    n132,
    n342
  );


  and
  g394
  (
    n419,
    n264,
    n283,
    n284,
    n241
  );


  xnor
  g395
  (
    n445,
    n336,
    n385,
    n168,
    n192
  );


  and
  g396
  (
    n528,
    n208,
    n142,
    n205,
    n311
  );


  nand
  g397
  (
    n550,
    n205,
    n368,
    n310,
    n374
  );


  xor
  g398
  (
    KeyWire_0_12,
    n223,
    n188,
    n153,
    n345
  );


  nor
  g399
  (
    n631,
    n387,
    n189,
    n359,
    n212
  );


  xnor
  g400
  (
    n437,
    n383,
    n274,
    n218,
    n393
  );


  nand
  g401
  (
    n577,
    n352,
    n321,
    n364,
    n250
  );


  or
  g402
  (
    n442,
    n135,
    n148,
    n145,
    n32
  );


  xnor
  g403
  (
    n557,
    n132,
    n273,
    n269,
    n212
  );


  xor
  g404
  (
    n545,
    n236,
    n284,
    n135,
    n308
  );


  xor
  g405
  (
    n639,
    n136,
    n371,
    n265,
    n242
  );


  nor
  g406
  (
    n593,
    n340,
    n324,
    n330,
    n325
  );


  or
  g407
  (
    n555,
    n314,
    n247,
    n289,
    n347
  );


  nand
  g408
  (
    n510,
    n215,
    n305,
    n355,
    n386
  );


  nand
  g409
  (
    n447,
    n148,
    n275,
    n340,
    n258
  );


  or
  g410
  (
    n611,
    n129,
    n191,
    n319,
    n357
  );


  nand
  g411
  (
    n569,
    n369,
    n384,
    n151,
    n144
  );


  xor
  g412
  (
    n413,
    n170,
    n210,
    n253,
    n169
  );


  xor
  g413
  (
    n482,
    n327,
    n379,
    n391,
    n232
  );


  nand
  g414
  (
    n415,
    n357,
    n363,
    n350,
    n220
  );


  or
  g415
  (
    n548,
    n173,
    n356,
    n354,
    n323
  );


  or
  g416
  (
    n666,
    n223,
    n382,
    n141,
    n200
  );


  nand
  g417
  (
    n636,
    n36,
    n223,
    n291,
    n320
  );


  xnor
  g418
  (
    n535,
    n154,
    n194,
    n381,
    n171
  );


  and
  g419
  (
    n461,
    n165,
    n158,
    n299,
    n294
  );


  or
  g420
  (
    n595,
    n153,
    n388,
    n264,
    n347
  );


  xnor
  g421
  (
    n602,
    n265,
    n128,
    n366,
    n188
  );


  nor
  g422
  (
    n477,
    n311,
    n302,
    n217,
    n325
  );


  and
  g423
  (
    n652,
    n163,
    n358,
    n140,
    n374
  );


  or
  g424
  (
    n521,
    n298,
    n255,
    n273,
    n140
  );


  xnor
  g425
  (
    n601,
    n330,
    n190,
    n270,
    n135
  );


  or
  g426
  (
    n585,
    n257,
    n184,
    n262,
    n218
  );


  nor
  g427
  (
    n468,
    n249,
    n340,
    n145,
    n200
  );


  nor
  g428
  (
    n464,
    n260,
    n156,
    n148,
    n146
  );


  nor
  g429
  (
    n450,
    n213,
    n167,
    n234,
    n246
  );


  or
  g430
  (
    n662,
    n350,
    n382,
    n189,
    n321
  );


  and
  g431
  (
    n470,
    n156,
    n141,
    n261,
    n334
  );


  xnor
  g432
  (
    n489,
    n302,
    n285,
    n343,
    n231
  );


  nor
  g433
  (
    n412,
    n325,
    n390,
    n270,
    n217
  );


  nand
  g434
  (
    n570,
    n143,
    n209,
    n225,
    n206
  );


  xnor
  g435
  (
    n527,
    n168,
    n337,
    n161,
    n173
  );


  nand
  g436
  (
    n645,
    n241,
    n378,
    n202
  );


  nand
  g437
  (
    n655,
    n127,
    n235,
    n287,
    n240
  );


  xnor
  g438
  (
    n499,
    n368,
    n316,
    n276,
    n219
  );


  and
  g439
  (
    n566,
    n201,
    n295,
    n190,
    n221
  );


  or
  g440
  (
    n597,
    n313,
    n267,
    n247,
    n266
  );


  nand
  g441
  (
    n531,
    n305,
    n242,
    n276,
    n216
  );


  xor
  g442
  (
    n678,
    n312,
    n270,
    n298,
    n252
  );


  nand
  g443
  (
    n669,
    n150,
    n349,
    n341,
    n384
  );


  nand
  g444
  (
    n659,
    n229,
    n307,
    n379,
    n345
  );


  xor
  g445
  (
    n504,
    n277,
    n312,
    n243,
    n387
  );


  and
  g446
  (
    n568,
    n335,
    n151,
    n361,
    n313
  );


  nand
  g447
  (
    n519,
    n38,
    n229,
    n292,
    n219
  );


  xnor
  g448
  (
    n665,
    n358,
    n364,
    n189,
    n321
  );


  xnor
  g449
  (
    n670,
    n240,
    n344,
    n195
  );


  nand
  g450
  (
    n634,
    n155,
    n158,
    n347,
    n352
  );


  xnor
  g451
  (
    n410,
    n216,
    n275,
    n267,
    n192
  );


  nor
  g452
  (
    n536,
    n361,
    n210,
    n197,
    n339
  );


  xnor
  g453
  (
    n514,
    n225,
    n378,
    n343,
    n288
  );


  or
  g454
  (
    n674,
    n257,
    n150,
    n336,
    n356
  );


  or
  g455
  (
    n476,
    n367,
    n127,
    n318,
    n263
  );


  and
  g456
  (
    n560,
    n300,
    n267,
    n368,
    n157
  );


  xor
  g457
  (
    n603,
    n308,
    n359,
    n289,
    n193
  );


  nand
  g458
  (
    n642,
    n210,
    n214,
    n227,
    n203
  );


  or
  g459
  (
    n438,
    n162,
    n266,
    n145,
    n317
  );


  or
  g460
  (
    n456,
    n378,
    n295,
    n145,
    n202
  );


  or
  g461
  (
    n506,
    n272,
    n364,
    n329,
    n149
  );


  nor
  g462
  (
    n623,
    n276,
    n387,
    n226,
    n311
  );


  xor
  g463
  (
    n508,
    n310,
    n342,
    n331,
    n337
  );


  xor
  g464
  (
    n605,
    n266,
    n344,
    n274,
    n245
  );


  nor
  g465
  (
    n500,
    n197,
    n339,
    n162,
    n244
  );


  nor
  g466
  (
    n418,
    n139,
    n389,
    n318,
    n360
  );


  xor
  g467
  (
    n430,
    n226,
    n167,
    n372,
    n269
  );


  xnor
  g468
  (
    n607,
    n362,
    n316,
    n367,
    n160
  );


  and
  g469
  (
    n651,
    n253,
    n311,
    n128,
    n147
  );


  nand
  g470
  (
    n474,
    n324,
    n223,
    n264,
    n204
  );


  or
  g471
  (
    n495,
    n346,
    n343,
    n293,
    n149
  );


  and
  g472
  (
    n511,
    n351,
    n196,
    n218,
    n152
  );


  xor
  g473
  (
    n587,
    n265,
    n159,
    n388,
    n203
  );


  nor
  g474
  (
    n620,
    n165,
    n130,
    n274,
    n281
  );


  xnor
  g475
  (
    n600,
    n200,
    n131,
    n353,
    n332
  );


  and
  g476
  (
    n592,
    n258,
    n357,
    n390,
    n303
  );


  nand
  g477
  (
    n572,
    n300,
    n225,
    n391,
    n170
  );


  xor
  g478
  (
    n416,
    n308,
    n248,
    n326,
    n164
  );


  nor
  g479
  (
    n457,
    n263,
    n238,
    n144,
    n206
  );


  nor
  g480
  (
    n580,
    n308,
    n257,
    n310,
    n128
  );


  xor
  g481
  (
    n417,
    n361,
    n365,
    n199,
    n348
  );


  xor
  g482
  (
    n453,
    n320,
    n204,
    n32,
    n263
  );


  nand
  g483
  (
    n565,
    n383,
    n207,
    n245,
    n265
  );


  xor
  g484
  (
    n539,
    n284,
    n389,
    n254,
    n304
  );


  and
  g485
  (
    n455,
    n164,
    n195,
    n310,
    n264
  );


  nor
  g486
  (
    n516,
    n293,
    n374,
    n219,
    n254
  );


  nor
  g487
  (
    n626,
    n249,
    n366,
    n326,
    n34
  );


  or
  g488
  (
    n584,
    n271,
    n342,
    n350,
    n312
  );


  and
  g489
  (
    n530,
    n156,
    n362,
    n162,
    n147
  );


  nand
  g490
  (
    n646,
    n196,
    n363,
    n186,
    n184
  );


  xnor
  g491
  (
    n661,
    n245,
    n152,
    n134,
    n329
  );


  xnor
  g492
  (
    n428,
    n202,
    n184,
    n200,
    n360
  );


  nor
  g493
  (
    n648,
    n135,
    n244
  );


  nand
  g494
  (
    n679,
    n384,
    n306,
    n383,
    n334
  );


  or
  g495
  (
    n571,
    n187,
    n386,
    n221,
    n292
  );


  xor
  g496
  (
    n491,
    n322,
    n143,
    n323,
    n307
  );


  xor
  g497
  (
    n478,
    n377,
    n355,
    n380,
    n278
  );


  xor
  g498
  (
    n481,
    n390,
    n166,
    n309,
    n130
  );


  xnor
  g499
  (
    n411,
    n231,
    n185,
    n209,
    n377
  );


  xor
  g500
  (
    n547,
    n222,
    n280,
    n163,
    n320
  );


  or
  g501
  (
    n518,
    n33,
    n319,
    n137,
    n353
  );


  and
  g502
  (
    n434,
    n259,
    n369,
    n393,
    n362
  );


  xnor
  g503
  (
    n673,
    n338,
    n213,
    n323,
    n330
  );


  xnor
  g504
  (
    n501,
    n375,
    n286,
    n185,
    n370
  );


  or
  g505
  (
    n473,
    n144,
    n204,
    n274,
    n220
  );


  or
  g506
  (
    n554,
    n152,
    n267,
    n291,
    n332
  );


  xnor
  g507
  (
    n629,
    n183,
    n143,
    n154,
    n307
  );


  and
  g508
  (
    n452,
    n382,
    n174,
    n353,
    n235
  );


  or
  g509
  (
    n425,
    n304,
    n260,
    n381,
    n328
  );


  xnor
  g510
  (
    n640,
    n256,
    n295,
    n242,
    n240
  );


  and
  g511
  (
    n641,
    n232,
    n338,
    n336,
    n218
  );


  xor
  g512
  (
    n596,
    n351,
    n166,
    n327,
    n127
  );


  nand
  g513
  (
    n599,
    n167,
    n228,
    n306,
    n301
  );


  nor
  g514
  (
    n479,
    n328,
    n231,
    n280,
    n164
  );


  nand
  g515
  (
    n574,
    n138,
    n233,
    n131,
    n369
  );


  xor
  g516
  (
    n541,
    n227,
    n168,
    n140,
    n371
  );


  nor
  g517
  (
    n458,
    n389,
    n277,
    n230,
    n213
  );


  or
  g518
  (
    n469,
    n331,
    n339,
    n377,
    n304
  );


  or
  g519
  (
    n656,
    n369,
    n333,
    n157,
    n288
  );


  or
  g520
  (
    n448,
    n210,
    n235,
    n283,
    n324
  );


  or
  g521
  (
    n497,
    n187,
    n313,
    n258,
    n203
  );


  nor
  g522
  (
    n588,
    n296,
    n360,
    n290,
    n262
  );


  xnor
  g523
  (
    n617,
    n288,
    n306,
    n150,
    n294
  );


  nor
  g524
  (
    n664,
    n314,
    n385,
    n332,
    n186
  );


  nor
  g525
  (
    n524,
    n303,
    n297,
    n220,
    n208
  );


  and
  g526
  (
    n618,
    n169,
    n173,
    n255,
    n336
  );


  nand
  g527
  (
    n668,
    n249,
    n165,
    n139,
    n155
  );


  nand
  g528
  (
    n515,
    n260,
    n196,
    n385,
    n356
  );


  xnor
  g529
  (
    n653,
    n185,
    n31,
    n228,
    n256
  );


  nor
  g530
  (
    n567,
    n272,
    n163,
    n215,
    n290
  );


  nor
  g531
  (
    n467,
    n153,
    n240,
    n322,
    n370
  );


  nor
  g532
  (
    n431,
    n248,
    n241,
    n138,
    n33
  );


  xnor
  g533
  (
    n672,
    n285,
    n297,
    n236,
    n235
  );


  nor
  g534
  (
    n635,
    n334,
    n224,
    n253,
    n380
  );


  nor
  g535
  (
    n429,
    n257,
    n351,
    n317,
    n247
  );


  or
  g536
  (
    n624,
    n341,
    n286,
    n224,
    n172
  );


  xnor
  g537
  (
    n676,
    n129,
    n375,
    n185,
    n136
  );


  nor
  g538
  (
    n426,
    n349,
    n198,
    n283,
    n337
  );


  or
  g539
  (
    n598,
    n329,
    n159,
    n165,
    n250
  );


  nor
  g540
  (
    n544,
    n146,
    n213,
    n239,
    n224
  );


  and
  g541
  (
    n680,
    n282,
    n166,
    n193,
    n214
  );


  and
  g542
  (
    n488,
    n389,
    n262,
    n258,
    n316
  );


  xnor
  g543
  (
    n414,
    n295,
    n302,
    n296,
    n243
  );


  and
  g544
  (
    n543,
    n368,
    n385,
    n209,
    n251
  );


  xor
  g545
  (
    n493,
    n349,
    n228,
    n193,
    n227
  );


  xnor
  g546
  (
    n613,
    n207,
    n211,
    n278,
    n149
  );


  nand
  g547
  (
    n654,
    n306,
    n259,
    n378,
    n151
  );


  or
  g548
  (
    n487,
    n341,
    n322,
    n194,
    n315
  );


  xor
  g549
  (
    n509,
    n340,
    n161,
    n151,
    n354
  );


  xor
  g550
  (
    n667,
    n359,
    n323,
    n188,
    n349
  );


  nand
  g551
  (
    KeyWire_0_14,
    n199,
    n228,
    n365,
    n328
  );


  nor
  g552
  (
    n427,
    n365,
    n160,
    n327,
    n351
  );


  nand
  g553
  (
    n537,
    n269,
    n217,
    n318,
    n201
  );


  or
  g554
  (
    n507,
    n285,
    n159,
    n364,
    n292
  );


  xnor
  g555
  (
    n671,
    n143,
    n314,
    n171,
    n261
  );


  xor
  g556
  (
    n522,
    n146,
    n246,
    n291,
    n137
  );


  nand
  g557
  (
    n619,
    n300,
    n272,
    n133,
    n246
  );


  xnor
  g558
  (
    n533,
    n233,
    n293,
    n128,
    n358
  );


  xor
  g559
  (
    n525,
    n242,
    n384,
    n127,
    n38
  );


  nand
  g560
  (
    n551,
    n216,
    n365,
    n372,
    n333
  );


  nor
  g561
  (
    n505,
    n217,
    n192,
    n270,
    n376
  );


  or
  g562
  (
    n556,
    n380,
    n277,
    n314
  );


  and
  g563
  (
    n564,
    n191,
    n372,
    n35,
    n391
  );


  xnor
  g564
  (
    n643,
    n191,
    n190,
    n250,
    n215
  );


  xor
  g565
  (
    n540,
    n331,
    n285,
    n197,
    n159
  );


  nor
  g566
  (
    n675,
    n279,
    n317,
    n332,
    n221
  );


  nand
  g567
  (
    n513,
    n261,
    n392,
    n312,
    n220
  );


  nor
  g568
  (
    n443,
    n297,
    n288,
    n172,
    n239
  );


  xor
  g569
  (
    n644,
    n238,
    n231,
    n195,
    n279
  );


  xor
  g570
  (
    n594,
    n237,
    n157,
    n211,
    n254
  );


  nand
  g571
  (
    n621,
    n160,
    n261,
    n133,
    n183
  );


  nand
  g572
  (
    n463,
    n230,
    n132,
    n191,
    n303
  );


  and
  g573
  (
    n490,
    n236,
    n355,
    n246,
    n232
  );


  nand
  g574
  (
    n546,
    n251,
    n150,
    n272,
    n190
  );


  xnor
  g575
  (
    n423,
    n206,
    n169,
    n222,
    n250
  );


  nand
  g576
  (
    n638,
    n204,
    n286,
    n307,
    n370
  );


  xnor
  g577
  (
    n420,
    n294,
    n138,
    n142,
    n320
  );


  nor
  g578
  (
    n432,
    n229,
    n134,
    n315,
    n195
  );


  xnor
  g579
  (
    n454,
    n376,
    n289,
    n281,
    n325
  );


  nor
  g580
  (
    n494,
    n199,
    n225,
    n329,
    n304
  );


  nand
  g581
  (
    n558,
    n208,
    n345,
    n187,
    n381
  );


  xnor
  g582
  (
    n502,
    n362,
    n234,
    n278,
    n393
  );


  nor
  g583
  (
    n451,
    n346,
    n157,
    n172,
    n130
  );


  nor
  g584
  (
    n462,
    n184,
    n154,
    n36,
    n339
  );


  nand
  g585
  (
    n538,
    n348,
    n134,
    n170,
    n188
  );


  nand
  g586
  (
    n559,
    n317,
    n245,
    n183,
    n254
  );


  nand
  g587
  (
    n677,
    n342,
    n309,
    n305,
    n361
  );


  nor
  g588
  (
    n465,
    n222,
    n209,
    n199,
    n347
  );


  nor
  g589
  (
    n529,
    n275,
    n282,
    n294,
    n373
  );


  and
  g590
  (
    n658,
    n214,
    n287,
    n132,
    n241
  );


  or
  g591
  (
    n627,
    n171,
    n154,
    n215,
    n198
  );


  and
  g592
  (
    n616,
    n248,
    n252,
    n377,
    n205
  );


  nand
  g593
  (
    n444,
    n315,
    n319,
    n352,
    n303
  );


  and
  g594
  (
    n435,
    n355,
    n168,
    n301,
    n271
  );


  xnor
  g595
  (
    n485,
    n203,
    n367,
    n375,
    n238
  );


  nand
  g596
  (
    n650,
    n374,
    n208,
    n381,
    n30
  );


  xnor
  g597
  (
    n472,
    n344,
    n333,
    n367,
    n328
  );


  and
  g598
  (
    n625,
    n379,
    n287,
    n376,
    n219
  );


  xor
  g599
  (
    n614,
    n34,
    n148,
    n296,
    n259
  );


  and
  g600
  (
    n436,
    n354,
    n189,
    n346,
    n319
  );


  nor
  g601
  (
    n498,
    n302,
    n249,
    n252,
    n153
  );


  or
  g602
  (
    n576,
    n233,
    n280,
    n212,
    n292
  );


  nand
  g603
  (
    n496,
    n207,
    n253,
    n324,
    n386
  );


  or
  g604
  (
    n608,
    n299,
    n139,
    n263,
    n194
  );


  nor
  g605
  (
    n649,
    n237,
    n214,
    n239,
    n388
  );


  xor
  g606
  (
    n663,
    n358,
    n206,
    n391,
    n160
  );


  and
  g607
  (
    n441,
    n158,
    n207,
    n330,
    n354
  );


  nor
  g608
  (
    n424,
    n281,
    n372,
    n133,
    n380
  );


  xnor
  g609
  (
    n660,
    n234,
    n290,
    n266,
    n230
  );


  nand
  g610
  (
    n503,
    n299,
    n147,
    n273,
    n275
  );


  xnor
  g611
  (
    n573,
    n205,
    n137,
    n247,
    n287
  );


  and
  g612
  (
    n483,
    n356,
    n390,
    n140,
    n237
  );


  and
  g613
  (
    n579,
    n37,
    n392,
    n268,
    n371
  );


  nor
  g614
  (
    n606,
    n279,
    n315,
    n301,
    n69
  );


  xnor
  g615
  (
    n647,
    n300,
    n363,
    n293,
    n284
  );


  and
  g616
  (
    n480,
    n290,
    n129,
    n232,
    n386
  );


  nand
  g617
  (
    n628,
    n348,
    n392,
    n299,
    n350
  );


  or
  g618
  (
    n561,
    n260,
    n251,
    n371,
    n268
  );


  and
  g619
  (
    n622,
    n251,
    n376,
    n327,
    n273
  );


  xnor
  g620
  (
    n633,
    n136,
    n282,
    n224,
    n297
  );


  xnor
  g621
  (
    n517,
    n286,
    n276,
    n183,
    n193
  );


  xnor
  g622
  (
    n475,
    n162,
    n375,
    n141,
    n296
  );


  nand
  g623
  (
    n612,
    n298,
    n37,
    n171,
    n335
  );


  xnor
  g624
  (
    n590,
    n382,
    n291,
    n331,
    n201
  );


  xnor
  g625
  (
    n439,
    n278,
    n161,
    n341,
    n39
  );


  and
  g626
  (
    n552,
    n186,
    n283,
    n243,
    n301
  );


  or
  g627
  (
    n563,
    n131,
    n289,
    n169,
    n252
  );


  nand
  g628
  (
    n520,
    n174,
    n255,
    n226,
    n236
  );


  nand
  g629
  (
    n486,
    n212,
    n268,
    n333,
    n337
  );


  nand
  g630
  (
    n632,
    n201,
    n366,
    n353,
    n131
  );


  nand
  g631
  (
    n549,
    n357,
    n305,
    n255,
    n298
  );


  nor
  g632
  (
    n657,
    n237,
    n343,
    n326,
    n173
  );


  nor
  g633
  (
    n581,
    n281,
    n334,
    n248,
    n383
  );


  nand
  g634
  (
    n637,
    n338,
    n155,
    n280,
    n279
  );


  and
  g635
  (
    n526,
    n167,
    n271,
    n229,
    n147
  );


  xnor
  g636
  (
    n466,
    n139,
    n198,
    n363,
    n216
  );


  xor
  g637
  (
    n492,
    n129,
    n166,
    n134,
    n239
  );


  xor
  g638
  (
    n471,
    n31,
    n392,
    n271,
    n172
  );


  nand
  g639
  (
    n532,
    n321,
    n156,
    n338,
    n373
  );


  and
  g640
  (
    n433,
    n137,
    n227,
    n211,
    n256
  );


  and
  g641
  (
    n681,
    n424,
    n411,
    n421
  );


  xor
  g642
  (
    n686,
    n414,
    n412,
    n410,
    n420
  );


  or
  g643
  (
    n682,
    n420,
    n425,
    n423,
    n417
  );


  xnor
  g644
  (
    n685,
    n413,
    n410,
    n423,
    n418
  );


  nor
  g645
  (
    n687,
    n421,
    n417,
    n416,
    n413
  );


  nor
  g646
  (
    n688,
    n422,
    n415,
    n416,
    n419
  );


  nor
  g647
  (
    n683,
    n412,
    n424,
    n415,
    n414
  );


  nor
  g648
  (
    n684,
    n425,
    n422,
    n419,
    n418
  );


  xnor
  g649
  (
    n691,
    n426,
    n431,
    n427,
    n683
  );


  xnor
  g650
  (
    n690,
    n430,
    n432,
    n429,
    n685
  );


  and
  g651
  (
    n693,
    n428,
    n684,
    n432,
    n431
  );


  xnor
  g652
  (
    n692,
    n430,
    n428,
    n681,
    n426
  );


  xor
  g653
  (
    n689,
    n682,
    n429,
    n427,
    n433
  );


  and
  g654
  (
    n702,
    n693,
    n446,
    n690
  );


  xnor
  g655
  (
    n697,
    n691,
    n442,
    n438
  );


  nand
  g656
  (
    n698,
    n438,
    n444,
    n448,
    n692
  );


  nand
  g657
  (
    n701,
    n440,
    n441,
    n435,
    n445
  );


  xnor
  g658
  (
    n703,
    n437,
    n435,
    n444,
    n691
  );


  and
  g659
  (
    n696,
    n441,
    n437,
    n447
  );


  or
  g660
  (
    n695,
    n689,
    n690,
    n443,
    n434
  );


  nor
  g661
  (
    n700,
    n439,
    n436,
    n693,
    n434
  );


  or
  g662
  (
    n694,
    n436,
    n443,
    n439,
    n692
  );


  or
  g663
  (
    n699,
    n440,
    n689,
    n433,
    n445
  );


  xnor
  g664
  (
    n708,
    n395,
    n394
  );


  or
  g665
  (
    n704,
    n694,
    n394
  );


  xnor
  g666
  (
    n707,
    n395,
    n396,
    n694,
    n394
  );


  nand
  g667
  (
    n705,
    n396,
    n694,
    n395
  );


  nand
  g668
  (
    n706,
    n395,
    n394,
    n695,
    n396
  );


  not
  g669
  (
    n710,
    n704
  );


  not
  g670
  (
    n709,
    n704
  );


  buf
  g671
  (
    n711,
    n704
  );


  buf
  g672
  (
    n712,
    n704
  );


  not
  g673
  (
    n720,
    n710
  );


  not
  g674
  (
    n725,
    n686
  );


  buf
  g675
  (
    n714,
    n695
  );


  buf
  g676
  (
    n723,
    n710
  );


  buf
  g677
  (
    n722,
    n687
  );


  not
  g678
  (
    n721,
    n712
  );


  not
  g679
  (
    n719,
    n687
  );


  buf
  g680
  (
    n728,
    n710
  );


  buf
  g681
  (
    n718,
    n695
  );


  not
  g682
  (
    n713,
    n712
  );


  buf
  g683
  (
    n727,
    n710
  );


  not
  g684
  (
    n724,
    n711
  );


  not
  g685
  (
    n716,
    n709
  );


  xor
  g686
  (
    n715,
    n712,
    n709
  );


  and
  g687
  (
    n726,
    n688,
    n448,
    n711,
    n712
  );


  xor
  g688
  (
    n717,
    n709,
    n711,
    n688
  );


  nand
  g689
  (
    n753,
    n399,
    n450,
    n449,
    n708
  );


  nor
  g690
  (
    n755,
    n717,
    n697,
    n716,
    n459
  );


  xor
  g691
  (
    n729,
    n177,
    n713,
    n706
  );


  nor
  g692
  (
    n747,
    n455,
    n715,
    n174
  );


  xor
  g693
  (
    n743,
    n696,
    n697,
    n698,
    n451
  );


  and
  g694
  (
    n736,
    n698,
    n698,
    n696,
    n452
  );


  nand
  g695
  (
    n746,
    n720,
    n717,
    n177,
    n716
  );


  xnor
  g696
  (
    n758,
    n454,
    n398,
    n461,
    n176
  );


  xnor
  g697
  (
    n738,
    n399,
    n719,
    n401
  );


  xnor
  g698
  (
    n745,
    n718,
    n397,
    n696,
    n461
  );


  xnor
  g699
  (
    n751,
    n399,
    n396,
    n454,
    n715
  );


  and
  g700
  (
    n732,
    n453,
    n177,
    n706,
    n175
  );


  xnor
  g701
  (
    n759,
    n175,
    n713,
    n397,
    n705
  );


  nand
  g702
  (
    n740,
    n397,
    n463,
    n719,
    n457
  );


  and
  g703
  (
    n757,
    n697,
    n707,
    n705
  );


  xnor
  g704
  (
    n737,
    n707,
    n720,
    n708,
    n457
  );


  xnor
  g705
  (
    n730,
    n456,
    n705,
    n718,
    n717
  );


  nor
  g706
  (
    n735,
    n397,
    n714,
    n400,
    n176
  );


  and
  g707
  (
    n741,
    n453,
    n450,
    n714,
    n715
  );


  or
  g708
  (
    n752,
    n706,
    n716,
    n713,
    n720
  );


  xnor
  g709
  (
    KeyWire_0_4,
    n452,
    n69,
    n462,
    n714
  );


  xor
  g710
  (
    n754,
    n174,
    n714,
    n718,
    n458
  );


  nor
  g711
  (
    n756,
    n460,
    n705,
    n449,
    n463
  );


  xnor
  g712
  (
    n760,
    n460,
    n451,
    n399,
    n698
  );


  and
  g713
  (
    n734,
    n696,
    n464,
    n175,
    n720
  );


  and
  g714
  (
    n750,
    n398,
    n718,
    n697,
    n400
  );


  nand
  g715
  (
    n749,
    n175,
    n717,
    n719,
    n400
  );


  or
  g716
  (
    n739,
    n398,
    n462,
    n176,
    n708
  );


  and
  g717
  (
    n742,
    n695,
    n398,
    n456,
    n716
  );


  and
  g718
  (
    n733,
    n400,
    n458,
    n176,
    n464
  );


  xor
  g719
  (
    n744,
    n708,
    n713,
    n707,
    n719
  );


  or
  g720
  (
    n731,
    n459,
    n455,
    n699,
    n177
  );


  nor
  g721
  (
    n761,
    n402,
    n701,
    n465,
    n700
  );


  nand
  g722
  (
    n766,
    n470,
    n401,
    n402,
    n701
  );


  xor
  g723
  (
    n763,
    n702,
    n733,
    n736,
    n468
  );


  nor
  g724
  (
    n764,
    n467,
    n732,
    n735,
    n466
  );


  xnor
  g725
  (
    n770,
    n730,
    n465,
    n701,
    n699
  );


  xnor
  g726
  (
    n762,
    n731,
    n738,
    n702,
    n401
  );


  nand
  g727
  (
    n765,
    n699,
    n469,
    n700
  );


  and
  g728
  (
    n767,
    n466,
    n702,
    n467,
    n699
  );


  xor
  g729
  (
    n768,
    n737,
    n701,
    n734,
    n468
  );


  xor
  g730
  (
    n769,
    n702,
    n700,
    n729,
    n469
  );


  xor
  g731
  (
    n777,
    n475,
    n765,
    n766,
    n769
  );


  xor
  g732
  (
    n776,
    n479,
    n471,
    n767
  );


  nand
  g733
  (
    n772,
    n472,
    n478,
    n770,
    n764
  );


  or
  g734
  (
    n773,
    n479,
    n478,
    n477
  );


  or
  g735
  (
    n775,
    n473,
    n474,
    n480
  );


  nand
  g736
  (
    n771,
    n480,
    n472,
    n476
  );


  xor
  g737
  (
    n774,
    n475,
    n470,
    n473,
    n768
  );


  not
  g738
  (
    n782,
    n771
  );


  not
  g739
  (
    n778,
    n772
  );


  buf
  g740
  (
    n783,
    n481
  );


  buf
  g741
  (
    n779,
    n772
  );


  not
  g742
  (
    n780,
    n771
  );


  xor
  g743
  (
    n781,
    n481,
    n771
  );


  xor
  g744
  (
    n785,
    n740,
    n482,
    n778
  );


  and
  g745
  (
    n784,
    n739,
    n772,
    n779
  );


  nor
  g746
  (
    n786,
    n784,
    n741
  );


  or
  g747
  (
    n787,
    n786,
    n773
  );


  or
  g748
  (
    n788,
    n774,
    n786,
    n773
  );


  buf
  g749
  (
    n792,
    n787
  );


  buf
  g750
  (
    n791,
    n774
  );


  xor
  g751
  (
    n789,
    n787,
    n775
  );


  xnor
  g752
  (
    n790,
    n774,
    n788
  );


  nor
  g753
  (
    n796,
    n181,
    n181,
    n791,
    n782
  );


  xnor
  g754
  (
    n800,
    n791,
    n721,
    n745,
    n780
  );


  and
  g755
  (
    n801,
    n182,
    n785,
    n722,
    n180
  );


  xnor
  g756
  (
    n804,
    n180,
    n179,
    n790
  );


  or
  g757
  (
    n797,
    n178,
    n178,
    n721,
    n179
  );


  xor
  g758
  (
    n799,
    n178,
    n721,
    n792,
    n789
  );


  and
  g759
  (
    n802,
    n181,
    n182,
    n789,
    n180
  );


  nand
  g760
  (
    n798,
    n791,
    n783,
    n722,
    n746
  );


  or
  g761
  (
    n793,
    n722,
    n744,
    n179,
    n791
  );


  or
  g762
  (
    n803,
    n721,
    n182,
    n781
  );


  and
  g763
  (
    n795,
    n790,
    n786,
    n789
  );


  xor
  g764
  (
    n794,
    n181,
    n180,
    n743,
    n790
  );


  xor
  g765
  (
    n805,
    n742,
    n178,
    n789,
    n790
  );


  xnor
  g766
  (
    n807,
    n754,
    n756,
    n757,
    n796
  );


  nand
  g767
  (
    n808,
    n795,
    n755,
    n757,
    n748
  );


  or
  g768
  (
    n806,
    n749,
    n793,
    n750,
    n751
  );


  or
  g769
  (
    n809,
    n747,
    n753,
    n794,
    n752
  );


  xor
  g770
  (
    n818,
    n498,
    n487,
    n807,
    n505
  );


  and
  g771
  (
    n820,
    n485,
    n501,
    n492,
    n808
  );


  nor
  g772
  (
    n814,
    n495,
    n489,
    n494,
    n488
  );


  and
  g773
  (
    n811,
    n492,
    n499,
    n502,
    n497
  );


  xnor
  g774
  (
    n810,
    n491,
    n502,
    n484,
    n506
  );


  or
  g775
  (
    n813,
    n496,
    n503,
    n486,
    n497
  );


  or
  g776
  (
    n825,
    n489,
    n487,
    n501,
    n809
  );


  nor
  g777
  (
    n819,
    n496,
    n495,
    n807,
    n488
  );


  and
  g778
  (
    n815,
    n506,
    n504,
    n503,
    n499
  );


  or
  g779
  (
    n816,
    n808,
    n494,
    n491,
    n809
  );


  xnor
  g780
  (
    n822,
    n484,
    n490,
    n808,
    n498
  );


  xor
  g781
  (
    n812,
    n808,
    n486,
    n483,
    n809
  );


  and
  g782
  (
    n823,
    n490,
    n500,
    n806
  );


  xnor
  g783
  (
    n824,
    n806,
    n807,
    n505
  );


  and
  g784
  (
    n821,
    n483,
    n493,
    n806,
    n504
  );


  and
  g785
  (
    n817,
    n809,
    n485,
    n806,
    n493
  );


  not
  g786
  (
    n828,
    n823
  );


  buf
  g787
  (
    n826,
    n821
  );


  buf
  g788
  (
    n827,
    n822
  );


  buf
  g789
  (
    n831,
    n798
  );


  nand
  g790
  (
    n834,
    n826,
    n512,
    n511
  );


  nand
  g791
  (
    n833,
    n510,
    n775,
    n826,
    n797
  );


  nor
  g792
  (
    n830,
    n799,
    n510,
    n509,
    n827
  );


  and
  g793
  (
    n836,
    n507,
    n827,
    n775,
    n792
  );


  xnor
  g794
  (
    n835,
    n512,
    n508,
    n827,
    n826
  );


  and
  g795
  (
    n832,
    n826,
    n775,
    n800,
    n509
  );


  xor
  g796
  (
    n829,
    n507,
    n508,
    n511,
    n827
  );


  nor
  g797
  (
    n838,
    n513,
    n517,
    n805,
    n514
  );


  xor
  g798
  (
    n839,
    n833,
    n804,
    n834,
    n519
  );


  or
  g799
  (
    n842,
    n520,
    n836,
    n518,
    n517
  );


  nor
  g800
  (
    n841,
    n516,
    n515,
    n802,
    n520
  );


  and
  g801
  (
    n843,
    n832,
    n515,
    n835,
    n830
  );


  nor
  g802
  (
    n837,
    n518,
    n516,
    n831,
    n803
  );


  xor
  g803
  (
    n840,
    n513,
    n801,
    n514,
    n519
  );


  buf
  g804
  (
    n866,
    n758
  );


  not
  g805
  (
    n850,
    n405
  );


  nand
  g806
  (
    n844,
    n522,
    n404,
    n406,
    n837
  );


  xor
  g807
  (
    n856,
    n406,
    n703,
    n404,
    n407
  );


  xnor
  g808
  (
    n854,
    n404,
    n842,
    n405,
    n521
  );


  or
  g809
  (
    n849,
    n408,
    n535,
    n703,
    n842
  );


  or
  g810
  (
    n871,
    n532,
    n841,
    n839,
    n408
  );


  and
  g811
  (
    n868,
    n406,
    n525,
    n824,
    n405
  );


  and
  g812
  (
    n845,
    n536,
    n409,
    n406,
    n402
  );


  or
  g813
  (
    n847,
    n521,
    n528,
    n408,
    n404
  );


  xor
  g814
  (
    n865,
    n403,
    n405,
    n531,
    n842
  );


  nand
  g815
  (
    n859,
    n530,
    n703,
    n537,
    n837
  );


  xor
  g816
  (
    n863,
    n534,
    n535,
    n524,
    n538
  );


  or
  g817
  (
    KeyWire_0_15,
    n703,
    n838,
    n837,
    n409
  );


  nor
  g818
  (
    n861,
    n841,
    n523,
    n403,
    n843
  );


  or
  g819
  (
    n848,
    n527,
    n838,
    n534,
    n407
  );


  and
  g820
  (
    n846,
    n530,
    n760,
    n841,
    n840
  );


  xnor
  g821
  (
    n867,
    n408,
    n526,
    n529,
    n536
  );


  nor
  g822
  (
    n864,
    n843,
    n538,
    n523,
    n402
  );


  xor
  g823
  (
    n852,
    n837,
    n843,
    n533
  );


  nand
  g824
  (
    n855,
    n760,
    n527,
    n403,
    n407
  );


  and
  g825
  (
    n860,
    n840,
    n522,
    n531,
    n403
  );


  nand
  g826
  (
    n858,
    n758,
    n407,
    n528,
    n839
  );


  nor
  g827
  (
    n857,
    n839,
    n839,
    n838,
    n529
  );


  and
  g828
  (
    n862,
    n825,
    n759,
    n838
  );


  nand
  g829
  (
    n870,
    n842,
    n409,
    n526,
    n533
  );


  nor
  g830
  (
    n869,
    n524,
    n409,
    n537,
    n525
  );


  xor
  g831
  (
    n853,
    n841,
    n840,
    n532
  );


  xor
  g832
  (
    n918,
    n855,
    n871,
    n860,
    n858
  );


  xor
  g833
  (
    n976,
    n569,
    n573,
    n850,
    n648
  );


  xor
  g834
  (
    n919,
    n586,
    n675,
    n866,
    n616
  );


  and
  g835
  (
    n969,
    n654,
    n651,
    n859,
    n676
  );


  and
  g836
  (
    n940,
    n865,
    n848,
    n673,
    n605
  );


  xor
  g837
  (
    n934,
    n599,
    n655,
    n870,
    n614
  );


  xnor
  g838
  (
    n951,
    n649,
    n857,
    n542,
    n593
  );


  nor
  g839
  (
    n909,
    n656,
    n606,
    n637,
    n599
  );


  or
  g840
  (
    n872,
    n671,
    n564,
    n850,
    n590
  );


  xnor
  g841
  (
    n927,
    n595,
    n610,
    n661,
    n628
  );


  xor
  g842
  (
    n899,
    n668,
    n861,
    n657,
    n846
  );


  xor
  g843
  (
    n935,
    n583,
    n857,
    n662,
    n639
  );


  or
  g844
  (
    n973,
    n630,
    n666,
    n548,
    n871
  );


  nor
  g845
  (
    n968,
    n652,
    n669,
    n675,
    n863
  );


  or
  g846
  (
    n895,
    n661,
    n620,
    n651,
    n854
  );


  xor
  g847
  (
    n876,
    n676,
    n856,
    n870,
    n669
  );


  xnor
  g848
  (
    n936,
    n578,
    n590,
    n629,
    n604
  );


  xor
  g849
  (
    n942,
    n605,
    n549,
    n568,
    n857
  );


  nor
  g850
  (
    n930,
    n586,
    n562,
    n849,
    n543
  );


  or
  g851
  (
    n894,
    n672,
    n675,
    n634,
    n567
  );


  nand
  g852
  (
    n924,
    n847,
    n626,
    n851,
    n610
  );


  and
  g853
  (
    n944,
    n859,
    n600,
    n563,
    n643
  );


  xor
  g854
  (
    n981,
    n539,
    n844,
    n646,
    n665
  );


  and
  g855
  (
    n974,
    n660,
    n673,
    n661,
    n554
  );


  and
  g856
  (
    n911,
    n858,
    n553,
    n661,
    n847
  );


  nand
  g857
  (
    n938,
    n556,
    n653,
    n664,
    n596
  );


  or
  g858
  (
    n896,
    n642,
    n608,
    n656,
    n553
  );


  nand
  g859
  (
    n960,
    n598,
    n626,
    n640,
    n607
  );


  xor
  g860
  (
    n910,
    n867,
    n637,
    n576,
    n555
  );


  nand
  g861
  (
    n879,
    n667,
    n566,
    n663,
    n662
  );


  or
  g862
  (
    n933,
    n647,
    n613,
    n864,
    n555
  );


  or
  g863
  (
    n954,
    n667,
    n648,
    n859,
    n635
  );


  xnor
  g864
  (
    n945,
    n552,
    n870,
    n543,
    n672
  );


  xor
  g865
  (
    n982,
    n663,
    n854,
    n849,
    n561
  );


  and
  g866
  (
    n941,
    n865,
    n572,
    n667,
    n582
  );


  and
  g867
  (
    n939,
    n660,
    n551,
    n860,
    n861
  );


  and
  g868
  (
    n901,
    n650,
    n672,
    n853,
    n611
  );


  and
  g869
  (
    n975,
    n663,
    n592,
    n585,
    n674
  );


  and
  g870
  (
    n950,
    n587,
    n665,
    n636,
    n670
  );


  xor
  g871
  (
    n878,
    n560,
    n654,
    n618
  );


  and
  g872
  (
    n965,
    n588,
    n624,
    n869,
    n602
  );


  xor
  g873
  (
    n972,
    n846,
    n860,
    n559,
    n674
  );


  nor
  g874
  (
    n885,
    n852,
    n854,
    n670,
    n615
  );


  and
  g875
  (
    n953,
    n570,
    n578,
    n865,
    n565
  );


  nand
  g876
  (
    n964,
    n544,
    n39,
    n863,
    n613
  );


  and
  g877
  (
    n912,
    n673,
    n622,
    n862,
    n868
  );


  or
  g878
  (
    n977,
    n858,
    n546,
    n591,
    n606
  );


  nor
  g879
  (
    n883,
    n862,
    n659,
    n547,
    n570
  );


  nor
  g880
  (
    n886,
    n557,
    n653,
    n587,
    n615
  );


  nand
  g881
  (
    n923,
    n646,
    n647,
    n612,
    n847
  );


  xor
  g882
  (
    n949,
    n633,
    n653,
    n564,
    n561
  );


  and
  g883
  (
    n908,
    n868,
    n649,
    n552,
    n851
  );


  nand
  g884
  (
    n931,
    n647,
    n636,
    n581,
    n642
  );


  or
  g885
  (
    n880,
    n655,
    n849,
    n847,
    n556
  );


  nand
  g886
  (
    n943,
    n623,
    n871,
    n583,
    n562
  );


  nor
  g887
  (
    n915,
    n569,
    n848,
    n594,
    n625
  );


  xnor
  g888
  (
    n900,
    n567,
    n669,
    n663,
    n632
  );


  nand
  g889
  (
    n979,
    n650,
    n573,
    n674,
    n593
  );


  and
  g890
  (
    n897,
    n603,
    n855,
    n651,
    n671
  );


  xnor
  g891
  (
    n921,
    n609,
    n617,
    n643,
    n545
  );


  or
  g892
  (
    n891,
    n545,
    n664,
    n860,
    n589
  );


  nor
  g893
  (
    n905,
    n635,
    n659,
    n575,
    n609
  );


  xor
  g894
  (
    n873,
    n619,
    n868,
    n853,
    n604
  );


  or
  g895
  (
    n884,
    n670,
    n865,
    n598,
    n550
  );


  or
  g896
  (
    n937,
    n666,
    n676,
    n541,
    n596
  );


  xnor
  g897
  (
    n932,
    n644,
    n601,
    n568,
    n845
  );


  and
  g898
  (
    n881,
    n614,
    n857,
    n579,
    n858
  );


  or
  g899
  (
    n928,
    n577,
    n657,
    n844,
    n592
  );


  xnor
  g900
  (
    n882,
    n634,
    n576,
    n655,
    n851
  );


  or
  g901
  (
    n963,
    n584,
    n584,
    n852,
    n577
  );


  xor
  g902
  (
    n875,
    n601,
    n670,
    n565,
    n600
  );


  xor
  g903
  (
    n890,
    n866,
    n861,
    n668,
    n627
  );


  or
  g904
  (
    n898,
    n862,
    n668,
    n660,
    n616
  );


  xor
  g905
  (
    n952,
    n867,
    n856,
    n547,
    n656
  );


  xnor
  g906
  (
    n889,
    n621,
    n868,
    n859,
    n867
  );


  and
  g907
  (
    n893,
    n845,
    n659,
    n658,
    n563
  );


  nor
  g908
  (
    n929,
    n665,
    n648,
    n658,
    n585
  );


  xor
  g909
  (
    n948,
    n594,
    n632,
    n628,
    n645
  );


  and
  g910
  (
    n926,
    n645,
    n588,
    n673,
    n657
  );


  xor
  g911
  (
    n917,
    n627,
    n623,
    n558,
    n668
  );


  and
  g912
  (
    n903,
    n639,
    n864,
    n652,
    n617
  );


  nand
  g913
  (
    n966,
    n638,
    n853,
    n620,
    n602
  );


  nor
  g914
  (
    n957,
    n652,
    n618,
    n665,
    n574
  );


  or
  g915
  (
    n947,
    n846,
    n539,
    n581,
    n548
  );


  and
  g916
  (
    n904,
    n624,
    n861,
    n852,
    n580
  );


  or
  g917
  (
    n956,
    n651,
    n867,
    n579,
    n549
  );


  xor
  g918
  (
    n971,
    n671,
    n644,
    n844,
    n647
  );


  and
  g919
  (
    n888,
    n844,
    n851,
    n855,
    n629
  );


  nor
  g920
  (
    n978,
    n597,
    n660,
    n559,
    n870
  );


  xor
  g921
  (
    n887,
    n630,
    n641,
    n845,
    n657
  );


  xor
  g922
  (
    n906,
    n658,
    n664,
    n648,
    n846
  );


  and
  g923
  (
    n962,
    n560,
    n850,
    n649,
    n582
  );


  and
  g924
  (
    n967,
    n654,
    n869,
    n864,
    n667
  );


  xor
  g925
  (
    n925,
    n608,
    n633,
    n557,
    n669
  );


  and
  g926
  (
    n892,
    n546,
    n671,
    n674,
    n591
  );


  and
  g927
  (
    n907,
    n855,
    n848,
    n863,
    n856
  );


  xor
  g928
  (
    n874,
    n849,
    n672,
    n653,
    n554
  );


  xor
  g929
  (
    n983,
    n848,
    n659,
    n580,
    n864
  );


  or
  g930
  (
    n913,
    n866,
    n641,
    n572,
    n856
  );


  nand
  g931
  (
    n920,
    n542,
    n650,
    n854,
    n655
  );


  xnor
  g932
  (
    n946,
    n571,
    n607,
    n574,
    n550
  );


  nor
  g933
  (
    n980,
    n621,
    n869,
    n652,
    n871
  );


  and
  g934
  (
    n959,
    n597,
    n853,
    n622,
    n850
  );


  nand
  g935
  (
    n916,
    n675,
    n658,
    n640,
    n664
  );


  nor
  g936
  (
    n958,
    n650,
    n666,
    n619,
    n625
  );


  xor
  g937
  (
    n902,
    n638,
    n649,
    n666,
    n575
  );


  nor
  g938
  (
    n914,
    n852,
    n558,
    n662,
    n866
  );


  xnor
  g939
  (
    n922,
    n541,
    n589,
    n603,
    n862
  );


  xnor
  g940
  (
    n955,
    n611,
    n612,
    n544,
    n595
  );


  xor
  g941
  (
    n970,
    n540,
    n551,
    n631,
    n656
  );


  nand
  g942
  (
    n877,
    n662,
    n571,
    n540,
    n863
  );


  xor
  g943
  (
    n961,
    n869,
    n631,
    n566,
    n845
  );


  or
  g944
  (
    n1016,
    n725,
    n980,
    n726,
    n777
  );


  nor
  g945
  (
    n1029,
    n878,
    n925,
    n968,
    n906
  );


  xor
  g946
  (
    n1002,
    n938,
    n950,
    n723,
    n966
  );


  xor
  g947
  (
    n1043,
    n728,
    n981,
    n945
  );


  nor
  g948
  (
    n1012,
    n939,
    n728,
    n892,
    n964
  );


  nor
  g949
  (
    n1023,
    n920,
    n935,
    n960,
    n724
  );


  xor
  g950
  (
    n992,
    n978,
    n900,
    n953,
    n942
  );


  xnor
  g951
  (
    n1007,
    n939,
    n887,
    n970,
    n944
  );


  or
  g952
  (
    n1046,
    n943,
    n727,
    n879,
    n677
  );


  and
  g953
  (
    n1044,
    n776,
    n911,
    n723,
    n947
  );


  xnor
  g954
  (
    n1039,
    n967,
    n726,
    n926,
    n902
  );


  and
  g955
  (
    n1042,
    n972,
    n958,
    n975,
    n941
  );


  nand
  g956
  (
    n1040,
    n676,
    n932,
    n896,
    n916
  );


  nor
  g957
  (
    n1037,
    n955,
    n971,
    n931,
    n977
  );


  and
  g958
  (
    n996,
    n962,
    n979,
    n967,
    n908
  );


  nor
  g959
  (
    n1028,
    n959,
    n898,
    n896,
    n900
  );


  xnor
  g960
  (
    n987,
    n901,
    n969,
    n924,
    n828
  );


  nand
  g961
  (
    n986,
    n895,
    n951,
    n929,
    n945
  );


  and
  g962
  (
    n1030,
    n919,
    n828,
    n725,
    n907
  );


  xor
  g963
  (
    n1020,
    n918,
    n941,
    n927,
    n679
  );


  xnor
  g964
  (
    n1000,
    n952,
    n876,
    n956,
    n921
  );


  nand
  g965
  (
    n1004,
    n883,
    n919,
    n678,
    n909
  );


  nor
  g966
  (
    n1034,
    n920,
    n723,
    n899,
    n892
  );


  or
  g967
  (
    n1021,
    n724,
    n908,
    n961,
    n39
  );


  nor
  g968
  (
    n998,
    n909,
    n950,
    n937,
    n928
  );


  or
  g969
  (
    n1045,
    n952,
    n961,
    n777,
    n917
  );


  nor
  g970
  (
    n984,
    n902,
    n973,
    n777,
    n679
  );


  nand
  g971
  (
    n999,
    n935,
    n898,
    n936,
    n888
  );


  or
  g972
  (
    n1026,
    n922,
    n901,
    n903,
    n983
  );


  xnor
  g973
  (
    n1025,
    n872,
    n680,
    n956,
    n905
  );


  nand
  g974
  (
    n988,
    n979,
    n885,
    n726,
    n940
  );


  xor
  g975
  (
    n1018,
    n873,
    n954,
    n894,
    n891
  );


  and
  g976
  (
    n1011,
    n947,
    n891,
    n910,
    n915
  );


  nor
  g977
  (
    n1031,
    n776,
    n959,
    n971,
    n972
  );


  nand
  g978
  (
    n1048,
    n946,
    n677,
    n728,
    n679
  );


  nand
  g979
  (
    KeyWire_0_3,
    n934,
    n678,
    n726,
    n976
  );


  and
  g980
  (
    n1036,
    n966,
    n882,
    n970,
    n936
  );


  and
  g981
  (
    n1001,
    n969,
    n727,
    n923,
    n680
  );


  nor
  g982
  (
    KeyWire_0_0,
    n924,
    n792,
    n903,
    n932
  );


  or
  g983
  (
    n1032,
    n968,
    n962,
    n725,
    n722
  );


  nand
  g984
  (
    n991,
    n897,
    n914,
    n982,
    n907
  );


  nor
  g985
  (
    n989,
    n965,
    n728,
    n890,
    n949
  );


  xor
  g986
  (
    n1003,
    n889,
    n938,
    n888,
    n978
  );


  xnor
  g987
  (
    n1013,
    n976,
    n777,
    n899,
    n881
  );


  nor
  g988
  (
    n1005,
    n977,
    n916,
    n937,
    n725
  );


  xnor
  g989
  (
    n985,
    n677,
    n957,
    n946,
    n960
  );


  nor
  g990
  (
    n1010,
    n955,
    n929,
    n724,
    n982
  );


  nand
  g991
  (
    n993,
    n875,
    n983,
    n905,
    n930
  );


  or
  g992
  (
    n990,
    n894,
    n678,
    n923,
    n943
  );


  xnor
  g993
  (
    n1047,
    n890,
    n957,
    n963,
    n724
  );


  xor
  g994
  (
    n1033,
    n897,
    n874,
    n828,
    n776
  );


  xnor
  g995
  (
    n1019,
    n931,
    n926,
    n913,
    n963
  );


  xor
  g996
  (
    n1022,
    n928,
    n973,
    n679,
    n39
  );


  xor
  g997
  (
    n1027,
    n895,
    n911,
    n953,
    n958
  );


  nand
  g998
  (
    n1017,
    n880,
    n910,
    n904,
    n886
  );


  xnor
  g999
  (
    n1049,
    n904,
    n948,
    n934
  );


  xor
  g1000
  (
    n1006,
    n917,
    n918,
    n942,
    n949
  );


  xor
  g1001
  (
    n1008,
    n974,
    n974,
    n913,
    n927
  );


  nor
  g1002
  (
    n1038,
    n980,
    n921,
    n914,
    n975
  );


  or
  g1003
  (
    n1024,
    n915,
    n828,
    n965,
    n930
  );


  and
  g1004
  (
    n1035,
    n944,
    n677,
    n893,
    n884
  );


  xnor
  g1005
  (
    n1014,
    n877,
    n951,
    n933
  );


  xor
  g1006
  (
    n995,
    n889,
    n727,
    n723,
    n925
  );


  nor
  g1007
  (
    n994,
    n912,
    n776,
    n906,
    n727
  );


  nor
  g1008
  (
    n1041,
    n792,
    n954,
    n922,
    n893
  );


  or
  g1009
  (
    n1009,
    n940,
    n964,
    n678,
    n912
  );


  or
  g1010
  (
    n1061,
    n987,
    n996,
    n1034,
    n1008
  );


  nand
  g1011
  (
    n1065,
    n1023,
    n1040,
    n989,
    n1009
  );


  xnor
  g1012
  (
    n1050,
    n1035,
    n997,
    n994,
    n986
  );


  or
  g1013
  (
    KeyWire_0_8,
    n1003,
    n1047,
    n680,
    n1005
  );


  xnor
  g1014
  (
    n1052,
    n1017,
    n1037,
    n1000,
    n1031
  );


  nor
  g1015
  (
    n1064,
    n1013,
    n1001,
    n1026,
    n990
  );


  nor
  g1016
  (
    n1059,
    n1020,
    n993,
    n1028,
    n1024
  );


  nand
  g1017
  (
    n1051,
    n1043,
    n1044,
    n1045,
    n1036
  );


  xor
  g1018
  (
    n1063,
    n1042,
    n1006,
    n1048,
    n1046
  );


  xnor
  g1019
  (
    n1062,
    n1015,
    n1027,
    n1030,
    n1032
  );


  xor
  g1020
  (
    n1057,
    n1039,
    n1014,
    n1019,
    n1007
  );


  nor
  g1021
  (
    n1056,
    n1010,
    n1029,
    n1041,
    n1016
  );


  nand
  g1022
  (
    n1055,
    n985,
    n1011,
    n999,
    n1018
  );


  xor
  g1023
  (
    n1060,
    n1025,
    n1002,
    n1004,
    n1038
  );


  nand
  g1024
  (
    n1058,
    n1012,
    n991,
    n992,
    n984
  );


  nor
  g1025
  (
    n1066,
    n998,
    n1022,
    n1033,
    n988
  );


  nor
  g1026
  (
    n1054,
    n995,
    n680,
    n1021,
    n1049
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1015,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n60,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n96,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n997,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n748,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n329,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n395,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n306,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1053,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n204,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n357,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n107,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n523,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n118,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n610,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n851,
    KeyNOTWire_0_15
  );


endmodule


