

module Stat_1648_36_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n1465,
  n1461,
  n1457,
  n1463,
  n1464,
  n1517,
  n1520,
  n1512,
  n1515,
  n1522,
  n1507,
  n1514,
  n1519,
  n1620,
  n1619,
  n1616,
  n1613,
  n1612,
  n1611,
  n1610,
  n1622,
  n1615,
  n1670,
  n1672,
  n1671,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n1465;
  output n1461;
  output n1457;
  output n1463;
  output n1464;
  output n1517;
  output n1520;
  output n1512;
  output n1515;
  output n1522;
  output n1507;
  output n1514;
  output n1519;
  output n1620;
  output n1619;
  output n1616;
  output n1613;
  output n1612;
  output n1611;
  output n1610;
  output n1622;
  output n1615;
  output n1670;
  output n1672;
  output n1671;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1462;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1513;
  wire n1516;
  wire n1518;
  wire n1521;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1614;
  wire n1617;
  wire n1618;
  wire n1621;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n71,
    n9
  );


  buf
  g1
  (
    n60,
    n17
  );


  not
  g2
  (
    n96,
    n23
  );


  not
  g3
  (
    n85,
    n14
  );


  buf
  g4
  (
    n75,
    n17
  );


  buf
  g5
  (
    n47,
    n18
  );


  buf
  g6
  (
    n77,
    n19
  );


  not
  g7
  (
    n119,
    n10
  );


  buf
  g8
  (
    n101,
    n7
  );


  not
  g9
  (
    n40,
    n24
  );


  buf
  g10
  (
    n45,
    n7
  );


  not
  g11
  (
    n62,
    n22
  );


  not
  g12
  (
    n42,
    n8
  );


  not
  g13
  (
    n98,
    n16
  );


  not
  g14
  (
    n68,
    n18
  );


  buf
  g15
  (
    n25,
    n11
  );


  not
  g16
  (
    n104,
    n4
  );


  buf
  g17
  (
    n81,
    n20
  );


  buf
  g18
  (
    n66,
    n3
  );


  buf
  g19
  (
    n107,
    n6
  );


  buf
  g20
  (
    n103,
    n9
  );


  not
  g21
  (
    n43,
    n7
  );


  buf
  g22
  (
    n110,
    n16
  );


  buf
  g23
  (
    n30,
    n12
  );


  not
  g24
  (
    n111,
    n22
  );


  not
  g25
  (
    n72,
    n5
  );


  not
  g26
  (
    n76,
    n10
  );


  buf
  g27
  (
    n65,
    n18
  );


  buf
  g28
  (
    n33,
    n10
  );


  not
  g29
  (
    n79,
    n4
  );


  not
  g30
  (
    n88,
    n15
  );


  buf
  g31
  (
    n93,
    n16
  );


  buf
  g32
  (
    n97,
    n19
  );


  not
  g33
  (
    n69,
    n12
  );


  not
  g34
  (
    n27,
    n5
  );


  not
  g35
  (
    n31,
    n13
  );


  not
  g36
  (
    n36,
    n22
  );


  not
  g37
  (
    n78,
    n20
  );


  not
  g38
  (
    n92,
    n19
  );


  not
  g39
  (
    n74,
    n1
  );


  buf
  g40
  (
    n99,
    n15
  );


  buf
  g41
  (
    n37,
    n23
  );


  not
  g42
  (
    n114,
    n24
  );


  buf
  g43
  (
    n61,
    n19
  );


  not
  g44
  (
    n34,
    n2
  );


  buf
  g45
  (
    n38,
    n15
  );


  buf
  g46
  (
    n82,
    n7
  );


  not
  g47
  (
    n115,
    n17
  );


  not
  g48
  (
    n113,
    n17
  );


  buf
  g49
  (
    n52,
    n24
  );


  buf
  g50
  (
    n39,
    n23
  );


  not
  g51
  (
    n64,
    n20
  );


  buf
  g52
  (
    n46,
    n21
  );


  not
  g53
  (
    n84,
    n11
  );


  buf
  g54
  (
    n109,
    n3
  );


  buf
  g55
  (
    n80,
    n20
  );


  buf
  g56
  (
    n63,
    n6
  );


  buf
  g57
  (
    n117,
    n21
  );


  not
  g58
  (
    n116,
    n1
  );


  not
  g59
  (
    n95,
    n6
  );


  buf
  g60
  (
    n53,
    n9
  );


  not
  g61
  (
    n83,
    n13
  );


  buf
  g62
  (
    n54,
    n18
  );


  buf
  g63
  (
    n118,
    n2
  );


  not
  g64
  (
    n48,
    n1
  );


  buf
  g65
  (
    n86,
    n12
  );


  not
  g66
  (
    n100,
    n3
  );


  not
  g67
  (
    n51,
    n13
  );


  not
  g68
  (
    n32,
    n14
  );


  buf
  g69
  (
    n91,
    n5
  );


  buf
  g70
  (
    n49,
    n8
  );


  buf
  g71
  (
    KeyWire_0_5,
    n5
  );


  buf
  g72
  (
    n108,
    n6
  );


  buf
  g73
  (
    n26,
    n8
  );


  not
  g74
  (
    n58,
    n21
  );


  not
  g75
  (
    n59,
    n3
  );


  buf
  g76
  (
    n112,
    n12
  );


  not
  g77
  (
    n29,
    n23
  );


  buf
  g78
  (
    n90,
    n14
  );


  buf
  g79
  (
    n50,
    n2
  );


  buf
  g80
  (
    n106,
    n9
  );


  buf
  g81
  (
    n67,
    n24
  );


  buf
  g82
  (
    n73,
    n11
  );


  buf
  g83
  (
    n55,
    n2
  );


  not
  g84
  (
    n44,
    n21
  );


  not
  g85
  (
    n87,
    n14
  );


  not
  g86
  (
    n102,
    n22
  );


  buf
  g87
  (
    n28,
    n11
  );


  not
  g88
  (
    n105,
    n15
  );


  buf
  g89
  (
    n89,
    n4
  );


  buf
  g90
  (
    n120,
    n4
  );


  not
  g91
  (
    n41,
    n1
  );


  not
  g92
  (
    n70,
    n8
  );


  buf
  g93
  (
    n56,
    n16
  );


  not
  g94
  (
    n57,
    n13
  );


  not
  g95
  (
    n94,
    n10
  );


  not
  g96
  (
    n299,
    n60
  );


  not
  g97
  (
    n419,
    n71
  );


  buf
  g98
  (
    n329,
    n60
  );


  buf
  g99
  (
    n246,
    n93
  );


  buf
  g100
  (
    n418,
    n93
  );


  buf
  g101
  (
    n214,
    n73
  );


  buf
  g102
  (
    n307,
    n34
  );


  not
  g103
  (
    n305,
    n96
  );


  buf
  g104
  (
    n279,
    n100
  );


  not
  g105
  (
    n163,
    n47
  );


  not
  g106
  (
    n421,
    n92
  );


  buf
  g107
  (
    n232,
    n76
  );


  buf
  g108
  (
    n170,
    n102
  );


  not
  g109
  (
    n455,
    n43
  );


  buf
  g110
  (
    n258,
    n46
  );


  buf
  g111
  (
    n426,
    n97
  );


  not
  g112
  (
    n260,
    n39
  );


  not
  g113
  (
    n135,
    n33
  );


  not
  g114
  (
    n159,
    n70
  );


  buf
  g115
  (
    n193,
    n29
  );


  not
  g116
  (
    n189,
    n46
  );


  buf
  g117
  (
    n321,
    n70
  );


  not
  g118
  (
    n318,
    n67
  );


  not
  g119
  (
    n282,
    n101
  );


  not
  g120
  (
    n177,
    n87
  );


  buf
  g121
  (
    n148,
    n74
  );


  not
  g122
  (
    n197,
    n55
  );


  not
  g123
  (
    n451,
    n104
  );


  buf
  g124
  (
    n306,
    n108
  );


  buf
  g125
  (
    n141,
    n53
  );


  not
  g126
  (
    KeyWire_0_13,
    n34
  );


  not
  g127
  (
    n338,
    n42
  );


  not
  g128
  (
    n179,
    n86
  );


  not
  g129
  (
    n295,
    n46
  );


  not
  g130
  (
    n291,
    n102
  );


  buf
  g131
  (
    n406,
    n47
  );


  not
  g132
  (
    n132,
    n85
  );


  buf
  g133
  (
    n427,
    n50
  );


  buf
  g134
  (
    n263,
    n77
  );


  buf
  g135
  (
    n371,
    n82
  );


  not
  g136
  (
    n271,
    n37
  );


  not
  g137
  (
    n350,
    n90
  );


  buf
  g138
  (
    n269,
    n51
  );


  buf
  g139
  (
    n182,
    n57
  );


  buf
  g140
  (
    n396,
    n79
  );


  buf
  g141
  (
    n278,
    n82
  );


  buf
  g142
  (
    n274,
    n37
  );


  not
  g143
  (
    n340,
    n86
  );


  buf
  g144
  (
    n326,
    n62
  );


  not
  g145
  (
    n313,
    n49
  );


  buf
  g146
  (
    n252,
    n62
  );


  buf
  g147
  (
    n443,
    n94
  );


  buf
  g148
  (
    n411,
    n96
  );


  not
  g149
  (
    n225,
    n66
  );


  buf
  g150
  (
    n178,
    n101
  );


  buf
  g151
  (
    n454,
    n28
  );


  buf
  g152
  (
    n367,
    n80
  );


  buf
  g153
  (
    n127,
    n41
  );


  not
  g154
  (
    n211,
    n95
  );


  buf
  g155
  (
    n123,
    n39
  );


  buf
  g156
  (
    n188,
    n56
  );


  buf
  g157
  (
    n283,
    n99
  );


  not
  g158
  (
    n156,
    n76
  );


  not
  g159
  (
    n288,
    n36
  );


  buf
  g160
  (
    n187,
    n40
  );


  buf
  g161
  (
    n137,
    n104
  );


  not
  g162
  (
    n139,
    n63
  );


  buf
  g163
  (
    n292,
    n58
  );


  not
  g164
  (
    n361,
    n30
  );


  not
  g165
  (
    n368,
    n59
  );


  not
  g166
  (
    n277,
    n105
  );


  not
  g167
  (
    n234,
    n84
  );


  not
  g168
  (
    n233,
    n25
  );


  buf
  g169
  (
    n324,
    n44
  );


  not
  g170
  (
    n248,
    n43
  );


  not
  g171
  (
    n147,
    n58
  );


  not
  g172
  (
    n357,
    n69
  );


  not
  g173
  (
    n390,
    n54
  );


  not
  g174
  (
    n124,
    n32
  );


  not
  g175
  (
    n227,
    n52
  );


  not
  g176
  (
    n181,
    n33
  );


  not
  g177
  (
    n237,
    n107
  );


  buf
  g178
  (
    n374,
    n36
  );


  not
  g179
  (
    n265,
    n35
  );


  not
  g180
  (
    n304,
    n26
  );


  buf
  g181
  (
    n398,
    n85
  );


  buf
  g182
  (
    n196,
    n97
  );


  not
  g183
  (
    n360,
    n27
  );


  not
  g184
  (
    n228,
    n106
  );


  buf
  g185
  (
    n138,
    n94
  );


  not
  g186
  (
    n449,
    n89
  );


  buf
  g187
  (
    n180,
    n108
  );


  not
  g188
  (
    n164,
    n91
  );


  not
  g189
  (
    n207,
    n54
  );


  not
  g190
  (
    n273,
    n71
  );


  not
  g191
  (
    n302,
    n54
  );


  not
  g192
  (
    n199,
    n68
  );


  buf
  g193
  (
    n257,
    n88
  );


  buf
  g194
  (
    n134,
    n86
  );


  buf
  g195
  (
    n221,
    n52
  );


  buf
  g196
  (
    n422,
    n40
  );


  not
  g197
  (
    n415,
    n41
  );


  not
  g198
  (
    n363,
    n50
  );


  not
  g199
  (
    n145,
    n74
  );


  buf
  g200
  (
    n190,
    n48
  );


  buf
  g201
  (
    n369,
    n52
  );


  not
  g202
  (
    n408,
    n51
  );


  not
  g203
  (
    n131,
    n65
  );


  not
  g204
  (
    n430,
    n75
  );


  buf
  g205
  (
    n158,
    n102
  );


  buf
  g206
  (
    n401,
    n42
  );


  not
  g207
  (
    KeyWire_0_9,
    n75
  );


  not
  g208
  (
    n143,
    n59
  );


  not
  g209
  (
    n250,
    n45
  );


  not
  g210
  (
    n424,
    n38
  );


  not
  g211
  (
    n373,
    n49
  );


  not
  g212
  (
    n389,
    n95
  );


  buf
  g213
  (
    n121,
    n75
  );


  buf
  g214
  (
    n384,
    n105
  );


  not
  g215
  (
    n375,
    n49
  );


  not
  g216
  (
    n416,
    n100
  );


  not
  g217
  (
    n270,
    n58
  );


  not
  g218
  (
    n383,
    n105
  );


  not
  g219
  (
    n376,
    n35
  );


  not
  g220
  (
    n428,
    n47
  );


  buf
  g221
  (
    n312,
    n72
  );


  buf
  g222
  (
    n323,
    n39
  );


  buf
  g223
  (
    n447,
    n82
  );


  buf
  g224
  (
    n267,
    n96
  );


  buf
  g225
  (
    n414,
    n92
  );


  buf
  g226
  (
    n412,
    n44
  );


  buf
  g227
  (
    n290,
    n71
  );


  buf
  g228
  (
    n315,
    n108
  );


  buf
  g229
  (
    n355,
    n35
  );


  buf
  g230
  (
    n325,
    n104
  );


  buf
  g231
  (
    n186,
    n100
  );


  buf
  g232
  (
    n435,
    n26
  );


  buf
  g233
  (
    n423,
    n96
  );


  buf
  g234
  (
    n378,
    n79
  );


  not
  g235
  (
    n438,
    n78
  );


  not
  g236
  (
    n266,
    n62
  );


  buf
  g237
  (
    n217,
    n75
  );


  not
  g238
  (
    n169,
    n83
  );


  not
  g239
  (
    n393,
    n60
  );


  not
  g240
  (
    n388,
    n66
  );


  not
  g241
  (
    n289,
    n34
  );


  not
  g242
  (
    n236,
    n90
  );


  not
  g243
  (
    n184,
    n55
  );


  buf
  g244
  (
    n446,
    n69
  );


  not
  g245
  (
    n353,
    n87
  );


  not
  g246
  (
    n351,
    n57
  );


  buf
  g247
  (
    n344,
    n32
  );


  not
  g248
  (
    n404,
    n89
  );


  not
  g249
  (
    n151,
    n25
  );


  buf
  g250
  (
    n339,
    n78
  );


  buf
  g251
  (
    n162,
    n108
  );


  not
  g252
  (
    n173,
    n63
  );


  buf
  g253
  (
    n335,
    n98
  );


  not
  g254
  (
    n294,
    n101
  );


  not
  g255
  (
    n209,
    n33
  );


  not
  g256
  (
    n342,
    n77
  );


  buf
  g257
  (
    n429,
    n68
  );


  buf
  g258
  (
    n439,
    n48
  );


  buf
  g259
  (
    n198,
    n77
  );


  buf
  g260
  (
    n372,
    n68
  );


  buf
  g261
  (
    n166,
    n36
  );


  buf
  g262
  (
    n285,
    n80
  );


  buf
  g263
  (
    n358,
    n83
  );


  not
  g264
  (
    n402,
    n66
  );


  buf
  g265
  (
    n347,
    n101
  );


  not
  g266
  (
    n433,
    n28
  );


  buf
  g267
  (
    n276,
    n102
  );


  buf
  g268
  (
    n334,
    n94
  );


  buf
  g269
  (
    n224,
    n37
  );


  buf
  g270
  (
    n332,
    n30
  );


  buf
  g271
  (
    n275,
    n62
  );


  buf
  g272
  (
    n254,
    n55
  );


  not
  g273
  (
    n249,
    n81
  );


  not
  g274
  (
    n385,
    n27
  );


  buf
  g275
  (
    n168,
    n76
  );


  buf
  g276
  (
    n204,
    n79
  );


  buf
  g277
  (
    n440,
    n59
  );


  not
  g278
  (
    n327,
    n36
  );


  not
  g279
  (
    n153,
    n60
  );


  buf
  g280
  (
    n434,
    n88
  );


  not
  g281
  (
    n400,
    n48
  );


  buf
  g282
  (
    n301,
    n44
  );


  buf
  g283
  (
    n210,
    n63
  );


  not
  g284
  (
    n136,
    n72
  );


  not
  g285
  (
    n235,
    n71
  );


  buf
  g286
  (
    n175,
    n67
  );


  not
  g287
  (
    n296,
    n69
  );


  buf
  g288
  (
    n413,
    n25
  );


  not
  g289
  (
    n392,
    n95
  );


  buf
  g290
  (
    n445,
    n86
  );


  buf
  g291
  (
    n195,
    n70
  );


  not
  g292
  (
    n231,
    n35
  );


  not
  g293
  (
    n394,
    n32
  );


  not
  g294
  (
    n407,
    n80
  );


  buf
  g295
  (
    n280,
    n64
  );


  buf
  g296
  (
    n300,
    n40
  );


  not
  g297
  (
    n432,
    n43
  );


  buf
  g298
  (
    n441,
    n107
  );


  not
  g299
  (
    n238,
    n34
  );


  buf
  g300
  (
    n262,
    n106
  );


  not
  g301
  (
    n208,
    n29
  );


  buf
  g302
  (
    n382,
    n103
  );


  not
  g303
  (
    n272,
    n90
  );


  buf
  g304
  (
    n409,
    n38
  );


  not
  g305
  (
    n160,
    n74
  );


  not
  g306
  (
    n205,
    n47
  );


  not
  g307
  (
    n444,
    n78
  );


  buf
  g308
  (
    n442,
    n100
  );


  not
  g309
  (
    n206,
    n61
  );


  not
  g310
  (
    n377,
    n26
  );


  buf
  g311
  (
    n259,
    n74
  );


  buf
  g312
  (
    n330,
    n33
  );


  not
  g313
  (
    n176,
    n38
  );


  buf
  g314
  (
    n144,
    n53
  );


  not
  g315
  (
    n133,
    n85
  );


  buf
  g316
  (
    n171,
    n107
  );


  not
  g317
  (
    n352,
    n50
  );


  not
  g318
  (
    n391,
    n93
  );


  not
  g319
  (
    n146,
    n84
  );


  not
  g320
  (
    n431,
    n54
  );


  buf
  g321
  (
    n345,
    n67
  );


  not
  g322
  (
    n436,
    n56
  );


  buf
  g323
  (
    n129,
    n81
  );


  not
  g324
  (
    n310,
    n89
  );


  not
  g325
  (
    n229,
    n61
  );


  not
  g326
  (
    n161,
    n40
  );


  buf
  g327
  (
    n216,
    n83
  );


  buf
  g328
  (
    n215,
    n43
  );


  buf
  g329
  (
    n309,
    n95
  );


  buf
  g330
  (
    n450,
    n73
  );


  not
  g331
  (
    n245,
    n52
  );


  buf
  g332
  (
    n341,
    n104
  );


  not
  g333
  (
    n150,
    n53
  );


  buf
  g334
  (
    n255,
    n50
  );


  not
  g335
  (
    n316,
    n92
  );


  not
  g336
  (
    n319,
    n30
  );


  buf
  g337
  (
    n293,
    n51
  );


  not
  g338
  (
    n303,
    n97
  );


  buf
  g339
  (
    n356,
    n69
  );


  buf
  g340
  (
    n247,
    n80
  );


  not
  g341
  (
    n240,
    n31
  );


  not
  g342
  (
    n379,
    n97
  );


  buf
  g343
  (
    n425,
    n37
  );


  buf
  g344
  (
    n222,
    n88
  );


  buf
  g345
  (
    n328,
    n82
  );


  buf
  g346
  (
    n452,
    n57
  );


  not
  g347
  (
    n241,
    n94
  );


  not
  g348
  (
    n268,
    n51
  );


  buf
  g349
  (
    n314,
    n63
  );


  not
  g350
  (
    n251,
    n42
  );


  buf
  g351
  (
    n410,
    n98
  );


  buf
  g352
  (
    n287,
    n83
  );


  not
  g353
  (
    n362,
    n99
  );


  not
  g354
  (
    n337,
    n67
  );


  not
  g355
  (
    n218,
    n53
  );


  buf
  g356
  (
    n308,
    n41
  );


  buf
  g357
  (
    n167,
    n91
  );


  not
  g358
  (
    n261,
    n31
  );


  not
  g359
  (
    n243,
    n91
  );


  buf
  g360
  (
    n380,
    n49
  );


  not
  g361
  (
    n405,
    n32
  );


  buf
  g362
  (
    n122,
    n30
  );


  buf
  g363
  (
    n201,
    n55
  );


  buf
  g364
  (
    n183,
    n65
  );


  not
  g365
  (
    n343,
    n31
  );


  buf
  g366
  (
    n399,
    n28
  );


  buf
  g367
  (
    n253,
    n99
  );


  buf
  g368
  (
    n298,
    n103
  );


  not
  g369
  (
    n165,
    n84
  );


  not
  g370
  (
    n320,
    n29
  );


  buf
  g371
  (
    n157,
    n39
  );


  not
  g372
  (
    n230,
    n78
  );


  not
  g373
  (
    n403,
    n84
  );


  buf
  g374
  (
    n456,
    n64
  );


  buf
  g375
  (
    n223,
    n87
  );


  buf
  g376
  (
    n366,
    n64
  );


  not
  g377
  (
    n155,
    n76
  );


  not
  g378
  (
    n212,
    n38
  );


  not
  g379
  (
    n364,
    n103
  );


  buf
  g380
  (
    n354,
    n90
  );


  buf
  g381
  (
    n317,
    n88
  );


  not
  g382
  (
    n386,
    n56
  );


  not
  g383
  (
    n281,
    n31
  );


  not
  g384
  (
    n346,
    n25
  );


  buf
  g385
  (
    n128,
    n107
  );


  not
  g386
  (
    n311,
    n99
  );


  buf
  g387
  (
    n239,
    n81
  );


  not
  g388
  (
    n203,
    n27
  );


  not
  g389
  (
    n125,
    n70
  );


  not
  g390
  (
    n220,
    n59
  );


  buf
  g391
  (
    n286,
    n106
  );


  not
  g392
  (
    n370,
    n89
  );


  not
  g393
  (
    n126,
    n72
  );


  not
  g394
  (
    n152,
    n26
  );


  buf
  g395
  (
    n149,
    n46
  );


  buf
  g396
  (
    n172,
    n66
  );


  buf
  g397
  (
    n264,
    n28
  );


  buf
  g398
  (
    n417,
    n57
  );


  not
  g399
  (
    n244,
    n93
  );


  not
  g400
  (
    n395,
    n81
  );


  not
  g401
  (
    n365,
    n29
  );


  not
  g402
  (
    n381,
    n98
  );


  buf
  g403
  (
    n256,
    n106
  );


  buf
  g404
  (
    n242,
    n61
  );


  not
  g405
  (
    n336,
    n61
  );


  not
  g406
  (
    n331,
    n72
  );


  not
  g407
  (
    n348,
    n98
  );


  not
  g408
  (
    n387,
    n42
  );


  not
  g409
  (
    n448,
    n44
  );


  buf
  g410
  (
    n349,
    n105
  );


  not
  g411
  (
    n453,
    n41
  );


  buf
  g412
  (
    n333,
    n73
  );


  buf
  g413
  (
    n322,
    n103
  );


  buf
  g414
  (
    n142,
    n56
  );


  buf
  g415
  (
    n185,
    n87
  );


  not
  g416
  (
    n284,
    n48
  );


  buf
  g417
  (
    n200,
    n45
  );


  not
  g418
  (
    n213,
    n73
  );


  buf
  g419
  (
    n297,
    n68
  );


  buf
  g420
  (
    n154,
    n85
  );


  not
  g421
  (
    n191,
    n77
  );


  buf
  g422
  (
    n202,
    n65
  );


  buf
  g423
  (
    n140,
    n58
  );


  not
  g424
  (
    n359,
    n92
  );


  not
  g425
  (
    n420,
    n45
  );


  not
  g426
  (
    n174,
    n91
  );


  buf
  g427
  (
    n194,
    n45
  );


  not
  g428
  (
    n397,
    n79
  );


  not
  g429
  (
    n130,
    n65
  );


  not
  g430
  (
    n192,
    n27
  );


  buf
  g431
  (
    n226,
    n64
  );


  not
  g432
  (
    n968,
    n325
  );


  buf
  g433
  (
    n876,
    n136
  );


  buf
  g434
  (
    n911,
    n342
  );


  buf
  g435
  (
    n465,
    n236
  );


  buf
  g436
  (
    n841,
    n237
  );


  not
  g437
  (
    n637,
    n297
  );


  not
  g438
  (
    n551,
    n259
  );


  not
  g439
  (
    KeyWire_0_24,
    n310
  );


  not
  g440
  (
    n684,
    n311
  );


  buf
  g441
  (
    KeyWire_0_10,
    n154
  );


  not
  g442
  (
    n1085,
    n354
  );


  not
  g443
  (
    n902,
    n200
  );


  not
  g444
  (
    n622,
    n274
  );


  buf
  g445
  (
    n807,
    n397
  );


  not
  g446
  (
    n895,
    n294
  );


  buf
  g447
  (
    n910,
    n229
  );


  buf
  g448
  (
    n1090,
    n370
  );


  buf
  g449
  (
    n963,
    n308
  );


  buf
  g450
  (
    n1045,
    n242
  );


  buf
  g451
  (
    n692,
    n135
  );


  buf
  g452
  (
    n881,
    n281
  );


  not
  g453
  (
    n512,
    n182
  );


  not
  g454
  (
    n998,
    n201
  );


  buf
  g455
  (
    n765,
    n329
  );


  buf
  g456
  (
    n974,
    n313
  );


  not
  g457
  (
    n562,
    n270
  );


  not
  g458
  (
    n888,
    n202
  );


  buf
  g459
  (
    n492,
    n341
  );


  buf
  g460
  (
    n1030,
    n132
  );


  buf
  g461
  (
    n1081,
    n260
  );


  not
  g462
  (
    n935,
    n360
  );


  buf
  g463
  (
    n697,
    n196
  );


  buf
  g464
  (
    n770,
    n194
  );


  buf
  g465
  (
    n750,
    n333
  );


  not
  g466
  (
    n889,
    n181
  );


  buf
  g467
  (
    n972,
    n127
  );


  not
  g468
  (
    n698,
    n302
  );


  buf
  g469
  (
    n548,
    n123
  );


  not
  g470
  (
    n1067,
    n227
  );


  not
  g471
  (
    n952,
    n195
  );


  not
  g472
  (
    n913,
    n138
  );


  not
  g473
  (
    n555,
    n275
  );


  buf
  g474
  (
    n1040,
    n276
  );


  buf
  g475
  (
    n604,
    n380
  );


  buf
  g476
  (
    n1051,
    n363
  );


  buf
  g477
  (
    n489,
    n299
  );


  not
  g478
  (
    n701,
    n194
  );


  buf
  g479
  (
    n494,
    n346
  );


  not
  g480
  (
    n845,
    n369
  );


  not
  g481
  (
    n740,
    n149
  );


  not
  g482
  (
    n1025,
    n222
  );


  not
  g483
  (
    n606,
    n165
  );


  not
  g484
  (
    n837,
    n305
  );


  not
  g485
  (
    n679,
    n265
  );


  not
  g486
  (
    n655,
    n249
  );


  buf
  g487
  (
    n703,
    n186
  );


  buf
  g488
  (
    n1003,
    n284
  );


  buf
  g489
  (
    n1041,
    n328
  );


  buf
  g490
  (
    n1075,
    n374
  );


  not
  g491
  (
    n1064,
    n124
  );


  buf
  g492
  (
    n839,
    n249
  );


  not
  g493
  (
    n651,
    n132
  );


  buf
  g494
  (
    n771,
    n273
  );


  not
  g495
  (
    n941,
    n366
  );


  not
  g496
  (
    KeyWire_0_11,
    n214
  );


  buf
  g497
  (
    KeyWire_0_17,
    n273
  );


  buf
  g498
  (
    n868,
    n182
  );


  buf
  g499
  (
    n857,
    n374
  );


  buf
  g500
  (
    n626,
    n160
  );


  not
  g501
  (
    n472,
    n336
  );


  buf
  g502
  (
    n653,
    n265
  );


  buf
  g503
  (
    n970,
    n201
  );


  not
  g504
  (
    n973,
    n348
  );


  buf
  g505
  (
    n783,
    n366
  );


  buf
  g506
  (
    n1046,
    n168
  );


  not
  g507
  (
    n619,
    n349
  );


  not
  g508
  (
    n930,
    n262
  );


  not
  g509
  (
    n519,
    n288
  );


  buf
  g510
  (
    n775,
    n171
  );


  buf
  g511
  (
    n798,
    n291
  );


  not
  g512
  (
    n744,
    n351
  );


  not
  g513
  (
    n938,
    n175
  );


  buf
  g514
  (
    n1019,
    n122
  );


  not
  g515
  (
    n909,
    n290
  );


  buf
  g516
  (
    n931,
    n269
  );


  not
  g517
  (
    n578,
    n125
  );


  not
  g518
  (
    n991,
    n133
  );


  not
  g519
  (
    n939,
    n404
  );


  not
  g520
  (
    n590,
    n156
  );


  buf
  g521
  (
    n797,
    n276
  );


  buf
  g522
  (
    n733,
    n286
  );


  not
  g523
  (
    n975,
    n328
  );


  not
  g524
  (
    n836,
    n398
  );


  not
  g525
  (
    n460,
    n230
  );


  buf
  g526
  (
    n721,
    n341
  );


  buf
  g527
  (
    n708,
    n153
  );


  buf
  g528
  (
    n936,
    n202
  );


  not
  g529
  (
    n649,
    n394
  );


  not
  g530
  (
    n793,
    n367
  );


  buf
  g531
  (
    n1035,
    n244
  );


  not
  g532
  (
    n746,
    n357
  );


  not
  g533
  (
    n745,
    n255
  );


  not
  g534
  (
    n874,
    n342
  );


  buf
  g535
  (
    n865,
    n240
  );


  not
  g536
  (
    n903,
    n403
  );


  not
  g537
  (
    n675,
    n165
  );


  not
  g538
  (
    n1071,
    n255
  );


  not
  g539
  (
    n628,
    n396
  );


  buf
  g540
  (
    n470,
    n199
  );


  buf
  g541
  (
    n1082,
    n300
  );


  not
  g542
  (
    n769,
    n206
  );


  buf
  g543
  (
    n802,
    n329
  );


  not
  g544
  (
    n486,
    n271
  );


  buf
  g545
  (
    n751,
    n161
  );


  not
  g546
  (
    n831,
    n326
  );


  buf
  g547
  (
    n550,
    n237
  );


  buf
  g548
  (
    n464,
    n131
  );


  not
  g549
  (
    KeyWire_0_4,
    n160
  );


  not
  g550
  (
    n468,
    n121
  );


  buf
  g551
  (
    n695,
    n309
  );


  buf
  g552
  (
    n988,
    n351
  );


  buf
  g553
  (
    n912,
    n397
  );


  not
  g554
  (
    n875,
    n304
  );


  not
  g555
  (
    n821,
    n128
  );


  buf
  g556
  (
    n672,
    n383
  );


  buf
  g557
  (
    n761,
    n338
  );


  buf
  g558
  (
    n1055,
    n307
  );


  buf
  g559
  (
    n537,
    n338
  );


  not
  g560
  (
    n525,
    n369
  );


  not
  g561
  (
    n820,
    n394
  );


  buf
  g562
  (
    n1006,
    n355
  );


  not
  g563
  (
    n789,
    n388
  );


  buf
  g564
  (
    n914,
    n213
  );


  buf
  g565
  (
    n849,
    n206
  );


  not
  g566
  (
    n1066,
    n124
  );


  buf
  g567
  (
    n869,
    n172
  );


  buf
  g568
  (
    n995,
    n340
  );


  not
  g569
  (
    n908,
    n325
  );


  not
  g570
  (
    n459,
    n371
  );


  not
  g571
  (
    n710,
    n213
  );


  not
  g572
  (
    n905,
    n268
  );


  buf
  g573
  (
    n1094,
    n270
  );


  buf
  g574
  (
    n728,
    n221
  );


  buf
  g575
  (
    n843,
    n357
  );


  buf
  g576
  (
    n917,
    n384
  );


  not
  g577
  (
    n508,
    n159
  );


  not
  g578
  (
    n530,
    n188
  );


  buf
  g579
  (
    n884,
    n360
  );


  not
  g580
  (
    n1037,
    n389
  );


  not
  g581
  (
    n906,
    n290
  );


  buf
  g582
  (
    n501,
    n173
  );


  buf
  g583
  (
    n536,
    n217
  );


  not
  g584
  (
    n561,
    n287
  );


  not
  g585
  (
    n483,
    n207
  );


  not
  g586
  (
    n1088,
    n141
  );


  not
  g587
  (
    n682,
    n208
  );


  not
  g588
  (
    n620,
    n297
  );


  buf
  g589
  (
    n481,
    n281
  );


  buf
  g590
  (
    n907,
    n303
  );


  not
  g591
  (
    n773,
    n373
  );


  not
  g592
  (
    n947,
    n220
  );


  buf
  g593
  (
    n829,
    n243
  );


  not
  g594
  (
    n623,
    n138
  );


  not
  g595
  (
    n986,
    n300
  );


  buf
  g596
  (
    n864,
    n305
  );


  not
  g597
  (
    n593,
    n296
  );


  buf
  g598
  (
    n523,
    n241
  );


  not
  g599
  (
    n899,
    n336
  );


  not
  g600
  (
    n702,
    n164
  );


  not
  g601
  (
    n1059,
    n309
  );


  buf
  g602
  (
    n654,
    n387
  );


  not
  g603
  (
    n861,
    n137
  );


  buf
  g604
  (
    n810,
    n193
  );


  buf
  g605
  (
    n630,
    n201
  );


  buf
  g606
  (
    n473,
    n390
  );


  not
  g607
  (
    n602,
    n387
  );


  not
  g608
  (
    n854,
    n221
  );


  buf
  g609
  (
    n663,
    n384
  );


  not
  g610
  (
    n573,
    n121
  );


  not
  g611
  (
    n475,
    n307
  );


  buf
  g612
  (
    n560,
    n143
  );


  not
  g613
  (
    n502,
    n173
  );


  not
  g614
  (
    n648,
    n333
  );


  buf
  g615
  (
    n923,
    n129
  );


  not
  g616
  (
    n642,
    n225
  );


  buf
  g617
  (
    n901,
    n401
  );


  not
  g618
  (
    n785,
    n289
  );


  buf
  g619
  (
    n940,
    n376
  );


  not
  g620
  (
    n1038,
    n365
  );


  buf
  g621
  (
    n982,
    n247
  );


  not
  g622
  (
    n535,
    n323
  );


  buf
  g623
  (
    n678,
    n219
  );


  not
  g624
  (
    n656,
    n307
  );


  buf
  g625
  (
    n925,
    n398
  );


  not
  g626
  (
    n597,
    n128
  );


  buf
  g627
  (
    n600,
    n347
  );


  buf
  g628
  (
    n801,
    n258
  );


  buf
  g629
  (
    n463,
    n202
  );


  buf
  g630
  (
    n474,
    n159
  );


  not
  g631
  (
    n981,
    n295
  );


  buf
  g632
  (
    KeyWire_0_0,
    n326
  );


  not
  g633
  (
    n687,
    n145
  );


  buf
  g634
  (
    n738,
    n339
  );


  buf
  g635
  (
    n513,
    n380
  );


  not
  g636
  (
    n873,
    n181
  );


  buf
  g637
  (
    n815,
    n373
  );


  buf
  g638
  (
    n499,
    n127
  );


  not
  g639
  (
    n599,
    n278
  );


  not
  g640
  (
    n476,
    n133
  );


  buf
  g641
  (
    n497,
    n314
  );


  buf
  g642
  (
    n929,
    n270
  );


  not
  g643
  (
    n894,
    n241
  );


  not
  g644
  (
    n479,
    n337
  );


  not
  g645
  (
    n457,
    n364
  );


  buf
  g646
  (
    n1073,
    n391
  );


  not
  g647
  (
    n595,
    n176
  );


  not
  g648
  (
    n953,
    n340
  );


  buf
  g649
  (
    n987,
    n306
  );


  not
  g650
  (
    n1086,
    n330
  );


  buf
  g651
  (
    n670,
    n286
  );


  not
  g652
  (
    n778,
    n207
  );


  buf
  g653
  (
    KeyWire_0_16,
    n375
  );


  not
  g654
  (
    n661,
    n257
  );


  not
  g655
  (
    n541,
    n281
  );


  buf
  g656
  (
    n976,
    n350
  );


  not
  g657
  (
    n1016,
    n167
  );


  not
  g658
  (
    n824,
    n324
  );


  not
  g659
  (
    n503,
    n308
  );


  not
  g660
  (
    n830,
    n388
  );


  not
  g661
  (
    n961,
    n129
  );


  not
  g662
  (
    n633,
    n330
  );


  buf
  g663
  (
    n1023,
    n158
  );


  buf
  g664
  (
    n927,
    n241
  );


  buf
  g665
  (
    n847,
    n172
  );


  buf
  g666
  (
    n786,
    n150
  );


  buf
  g667
  (
    n956,
    n167
  );


  not
  g668
  (
    n747,
    n354
  );


  buf
  g669
  (
    n488,
    n329
  );


  buf
  g670
  (
    n724,
    n321
  );


  not
  g671
  (
    n531,
    n337
  );


  not
  g672
  (
    n552,
    n356
  );


  buf
  g673
  (
    n646,
    n125
  );


  not
  g674
  (
    n681,
    n122
  );


  not
  g675
  (
    n1028,
    n277
  );


  buf
  g676
  (
    n569,
    n370
  );


  not
  g677
  (
    n493,
    n403
  );


  not
  g678
  (
    n683,
    n222
  );


  not
  g679
  (
    n496,
    n373
  );


  not
  g680
  (
    n916,
    n232
  );


  buf
  g681
  (
    n962,
    n302
  );


  not
  g682
  (
    n856,
    n344
  );


  not
  g683
  (
    n618,
    n190
  );


  not
  g684
  (
    n583,
    n197
  );


  buf
  g685
  (
    n858,
    n385
  );


  buf
  g686
  (
    n559,
    n198
  );


  buf
  g687
  (
    n674,
    n169
  );


  buf
  g688
  (
    n992,
    n287
  );


  buf
  g689
  (
    n652,
    n127
  );


  not
  g690
  (
    n641,
    n193
  );


  not
  g691
  (
    n1049,
    n154
  );


  buf
  g692
  (
    n877,
    n196
  );


  not
  g693
  (
    n1009,
    n304
  );


  not
  g694
  (
    n870,
    n285
  );


  buf
  g695
  (
    n669,
    n231
  );


  buf
  g696
  (
    n983,
    n225
  );


  not
  g697
  (
    n645,
    n124
  );


  buf
  g698
  (
    n546,
    n169
  );


  not
  g699
  (
    n896,
    n350
  );


  not
  g700
  (
    n926,
    n404
  );


  buf
  g701
  (
    n1018,
    n395
  );


  not
  g702
  (
    n885,
    n239
  );


  buf
  g703
  (
    n671,
    n247
  );


  not
  g704
  (
    n514,
    n374
  );


  not
  g705
  (
    n693,
    n284
  );


  not
  g706
  (
    n589,
    n252
  );


  not
  g707
  (
    n601,
    n199
  );


  not
  g708
  (
    n577,
    n228
  );


  buf
  g709
  (
    n631,
    n317
  );


  not
  g710
  (
    n462,
    n145
  );


  not
  g711
  (
    n580,
    n159
  );


  buf
  g712
  (
    n774,
    n243
  );


  not
  g713
  (
    n752,
    n259
  );


  buf
  g714
  (
    n491,
    n232
  );


  buf
  g715
  (
    n521,
    n369
  );


  not
  g716
  (
    n1061,
    n320
  );


  not
  g717
  (
    n900,
    n285
  );


  buf
  g718
  (
    n760,
    n226
  );


  buf
  g719
  (
    n504,
    n313
  );


  not
  g720
  (
    n754,
    n151
  );


  buf
  g721
  (
    n755,
    n153
  );


  not
  g722
  (
    n598,
    n312
  );


  not
  g723
  (
    n1010,
    n130
  );


  not
  g724
  (
    n1057,
    n240
  );


  buf
  g725
  (
    n1031,
    n303
  );


  not
  g726
  (
    n1027,
    n375
  );


  buf
  g727
  (
    n1033,
    n399
  );


  buf
  g728
  (
    n461,
    n279
  );


  buf
  g729
  (
    n1074,
    n388
  );


  not
  g730
  (
    n964,
    n396
  );


  not
  g731
  (
    n542,
    n310
  );


  buf
  g732
  (
    n629,
    n402
  );


  buf
  g733
  (
    n1000,
    n303
  );


  not
  g734
  (
    n706,
    n144
  );


  not
  g735
  (
    n634,
    n335
  );


  not
  g736
  (
    n920,
    n350
  );


  buf
  g737
  (
    n759,
    n195
  );


  not
  g738
  (
    n776,
    n343
  );


  buf
  g739
  (
    n1052,
    n284
  );


  not
  g740
  (
    n731,
    n151
  );


  buf
  g741
  (
    n665,
    n283
  );


  buf
  g742
  (
    KeyWire_0_23,
    n212
  );


  buf
  g743
  (
    n1079,
    n321
  );


  buf
  g744
  (
    n607,
    n298
  );


  not
  g745
  (
    n1062,
    n334
  );


  not
  g746
  (
    n781,
    n244
  );


  not
  g747
  (
    n640,
    n336
  );


  buf
  g748
  (
    n539,
    n394
  );


  not
  g749
  (
    n919,
    n249
  );


  buf
  g750
  (
    n1092,
    n283
  );


  not
  g751
  (
    n758,
    n174
  );


  buf
  g752
  (
    n534,
    n244
  );


  not
  g753
  (
    n570,
    n389
  );


  buf
  g754
  (
    KeyWire_0_19,
    n136
  );


  not
  g755
  (
    n526,
    n251
  );


  not
  g756
  (
    n804,
    n266
  );


  buf
  g757
  (
    n532,
    n242
  );


  not
  g758
  (
    n588,
    n332
  );


  not
  g759
  (
    n1087,
    n400
  );


  not
  g760
  (
    n689,
    n171
  );


  buf
  g761
  (
    n712,
    n210
  );


  buf
  g762
  (
    n835,
    n140
  );


  not
  g763
  (
    n500,
    n275
  );


  buf
  g764
  (
    n1015,
    n403
  );


  not
  g765
  (
    n848,
    n358
  );


  not
  g766
  (
    n587,
    n196
  );


  not
  g767
  (
    n887,
    n378
  );


  not
  g768
  (
    n667,
    n147
  );


  not
  g769
  (
    n891,
    n185
  );


  buf
  g770
  (
    n796,
    n132
  );


  not
  g771
  (
    n517,
    n223
  );


  not
  g772
  (
    n959,
    n238
  );


  buf
  g773
  (
    n568,
    n129
  );


  buf
  g774
  (
    n734,
    n138
  );


  not
  g775
  (
    n1043,
    n263
  );


  buf
  g776
  (
    n719,
    n355
  );


  buf
  g777
  (
    n784,
    n393
  );


  not
  g778
  (
    n709,
    n172
  );


  buf
  g779
  (
    n1007,
    n256
  );


  buf
  g780
  (
    n522,
    n377
  );


  buf
  g781
  (
    n613,
    n290
  );


  buf
  g782
  (
    n699,
    n168
  );


  not
  g783
  (
    n647,
    n262
  );


  not
  g784
  (
    n490,
    n187
  );


  buf
  g785
  (
    n495,
    n225
  );


  not
  g786
  (
    n1072,
    n355
  );


  buf
  g787
  (
    n768,
    n211
  );


  not
  g788
  (
    n715,
    n233
  );


  buf
  g789
  (
    n1017,
    n313
  );


  buf
  g790
  (
    n965,
    n204
  );


  not
  g791
  (
    n777,
    n348
  );


  buf
  g792
  (
    n605,
    n363
  );


  buf
  g793
  (
    n720,
    n139
  );


  not
  g794
  (
    n766,
    n179
  );


  not
  g795
  (
    n1091,
    n251
  );


  buf
  g796
  (
    n487,
    n176
  );


  not
  g797
  (
    n883,
    n309
  );


  not
  g798
  (
    n694,
    n256
  );


  not
  g799
  (
    n934,
    n202
  );


  buf
  g800
  (
    n680,
    n327
  );


  buf
  g801
  (
    n586,
    n133
  );


  not
  g802
  (
    n557,
    n280
  );


  not
  g803
  (
    n800,
    n292
  );


  not
  g804
  (
    n825,
    n387
  );


  not
  g805
  (
    n932,
    n275
  );


  buf
  g806
  (
    n458,
    n322
  );


  not
  g807
  (
    n538,
    n146
  );


  buf
  g808
  (
    n677,
    n281
  );


  buf
  g809
  (
    n612,
    n360
  );


  buf
  g810
  (
    n608,
    n178
  );


  not
  g811
  (
    n817,
    n242
  );


  not
  g812
  (
    n632,
    n371
  );


  not
  g813
  (
    n749,
    n292
  );


  buf
  g814
  (
    n1005,
    n386
  );


  buf
  g815
  (
    n544,
    n279
  );


  buf
  g816
  (
    n1044,
    n246
  );


  buf
  g817
  (
    n897,
    n289
  );


  not
  g818
  (
    n506,
    n184
  );


  buf
  g819
  (
    n918,
    n135
  );


  not
  g820
  (
    n753,
    n301
  );


  buf
  g821
  (
    n624,
    n126
  );


  buf
  g822
  (
    n466,
    n334
  );


  buf
  g823
  (
    n928,
    n198
  );


  not
  g824
  (
    n756,
    n204
  );


  not
  g825
  (
    n809,
    n136
  );


  buf
  g826
  (
    n871,
    n344
  );


  buf
  g827
  (
    n478,
    n167
  );


  buf
  g828
  (
    n772,
    n177
  );


  buf
  g829
  (
    KeyWire_0_25,
    n174
  );


  buf
  g830
  (
    n921,
    n386
  );


  not
  g831
  (
    n558,
    n273
  );


  not
  g832
  (
    n924,
    n263
  );


  not
  g833
  (
    n611,
    n211
  );


  not
  g834
  (
    n567,
    n297
  );


  not
  g835
  (
    n575,
    n157
  );


  buf
  g836
  (
    n549,
    n333
  );


  not
  g837
  (
    n615,
    n400
  );


  buf
  g838
  (
    n1026,
    n218
  );


  buf
  g839
  (
    n650,
    n166
  );


  buf
  g840
  (
    n1070,
    n339
  );


  buf
  g841
  (
    n997,
    n261
  );


  not
  g842
  (
    n566,
    n142
  );


  buf
  g843
  (
    n859,
    n361
  );


  buf
  g844
  (
    n516,
    n162
  );


  buf
  g845
  (
    n945,
    n322
  );


  not
  g846
  (
    n886,
    n207
  );


  buf
  g847
  (
    n882,
    n200
  );


  not
  g848
  (
    n554,
    n191
  );


  not
  g849
  (
    n993,
    n300
  );


  buf
  g850
  (
    n862,
    n382
  );


  buf
  g851
  (
    n565,
    n214
  );


  buf
  g852
  (
    n563,
    n164
  );


  buf
  g853
  (
    n617,
    n321
  );


  buf
  g854
  (
    n545,
    n204
  );


  buf
  g855
  (
    n950,
    n276
  );


  buf
  g856
  (
    n676,
    n141
  );


  buf
  g857
  (
    n943,
    n230
  );


  buf
  g858
  (
    n507,
    n279
  );


  buf
  g859
  (
    n937,
    n399
  );


  not
  g860
  (
    n949,
    n161
  );


  buf
  g861
  (
    n511,
    n384
  );


  not
  g862
  (
    n994,
    n259
  );


  not
  g863
  (
    KeyWire_0_28,
    n256
  );


  buf
  g864
  (
    n644,
    n158
  );


  buf
  g865
  (
    n716,
    n388
  );


  buf
  g866
  (
    n571,
    n293
  );


  not
  g867
  (
    n543,
    n262
  );


  buf
  g868
  (
    n527,
    n174
  );


  buf
  g869
  (
    n805,
    n228
  );


  not
  g870
  (
    n584,
    n272
  );


  not
  g871
  (
    n1065,
    n196
  );


  not
  g872
  (
    n1054,
    n362
  );


  not
  g873
  (
    n795,
    n234
  );


  buf
  g874
  (
    n579,
    n170
  );


  buf
  g875
  (
    n1034,
    n132
  );


  not
  g876
  (
    n1077,
    n130
  );


  not
  g877
  (
    n814,
    n296
  );


  not
  g878
  (
    n515,
    n179
  );


  not
  g879
  (
    n572,
    n311
  );


  buf
  g880
  (
    n610,
    n343
  );


  buf
  g881
  (
    n614,
    n309
  );


  not
  g882
  (
    n625,
    n146
  );


  buf
  g883
  (
    n529,
    n138
  );


  buf
  g884
  (
    n1013,
    n208
  );


  not
  g885
  (
    n658,
    n358
  );


  not
  g886
  (
    n985,
    n175
  );


  buf
  g887
  (
    n700,
    n331
  );


  not
  g888
  (
    n484,
    n379
  );


  not
  g889
  (
    n627,
    n404
  );


  buf
  g890
  (
    n971,
    n233
  );


  not
  g891
  (
    n743,
    n166
  );


  buf
  g892
  (
    n1053,
    n335
  );


  buf
  g893
  (
    n838,
    n124
  );


  buf
  g894
  (
    n1048,
    n288
  );


  buf
  g895
  (
    n840,
    n368
  );


  not
  g896
  (
    n828,
    n342
  );


  not
  g897
  (
    n1014,
    n170
  );


  not
  g898
  (
    n764,
    n228
  );


  buf
  g899
  (
    n1024,
    n125
  );


  not
  g900
  (
    n853,
    n191
  );


  not
  g901
  (
    n748,
    n319
  );


  not
  g902
  (
    n790,
    n301
  );


  buf
  g903
  (
    n482,
    n322
  );


  not
  g904
  (
    KeyWire_0_20,
    n327
  );


  nand
  g905
  (
    n788,
    n143,
    n126,
    n277
  );


  xor
  g906
  (
    n946,
    n376,
    n376,
    n316,
    n157
  );


  or
  g907
  (
    n585,
    n299,
    n391,
    n302
  );


  nor
  g908
  (
    n1078,
    n314,
    n121,
    n123,
    n130
  );


  xor
  g909
  (
    n969,
    n177,
    n122,
    n367,
    n158
  );


  or
  g910
  (
    n1029,
    n268,
    n283,
    n231,
    n240
  );


  xnor
  g911
  (
    n855,
    n165,
    n398,
    n192,
    n324
  );


  and
  g912
  (
    n803,
    n338,
    n122,
    n395,
    n334
  );


  xor
  g913
  (
    n851,
    n162,
    n327,
    n221,
    n323
  );


  xor
  g914
  (
    n999,
    n156,
    n384,
    n277,
    n206
  );


  nor
  g915
  (
    n852,
    n250,
    n317,
    n379,
    n365
  );


  and
  g916
  (
    n933,
    n382,
    n293,
    n188,
    n294
  );


  nand
  g917
  (
    n603,
    n177,
    n169,
    n334,
    n387
  );


  nor
  g918
  (
    n948,
    n297,
    n218,
    n318,
    n222
  );


  xor
  g919
  (
    n966,
    n348,
    n152,
    n180,
    n342
  );


  xnor
  g920
  (
    n685,
    n362,
    n150,
    n261,
    n279
  );


  xor
  g921
  (
    n833,
    n344,
    n137,
    n237,
    n129
  );


  xnor
  g922
  (
    n711,
    n250,
    n335,
    n183,
    n240
  );


  and
  g923
  (
    n621,
    n352,
    n142,
    n339,
    n227
  );


  xor
  g924
  (
    n915,
    n134,
    n318,
    n254,
    n381
  );


  and
  g925
  (
    n505,
    n361,
    n146,
    n184,
    n402
  );


  xnor
  g926
  (
    n872,
    n285,
    n348,
    n298,
    n347
  );


  xnor
  g927
  (
    n942,
    n359,
    n378,
    n167,
    n247
  );


  xnor
  g928
  (
    n705,
    n209,
    n292,
    n148,
    n267
  );


  xor
  g929
  (
    n1069,
    n170,
    n178,
    n152,
    n197
  );


  nor
  g930
  (
    n844,
    n185,
    n404,
    n378,
    n241
  );


  or
  g931
  (
    n832,
    n157,
    n231,
    n171,
    n263
  );


  nor
  g932
  (
    n890,
    n382,
    n197,
    n326,
    n343
  );


  nor
  g933
  (
    n860,
    n187,
    n274,
    n245,
    n148
  );


  xor
  g934
  (
    n659,
    n189,
    n305,
    n390,
    n235
  );


  and
  g935
  (
    n850,
    n216,
    n153,
    n353,
    n135
  );


  xor
  g936
  (
    n739,
    n345,
    n218,
    n263,
    n308
  );


  and
  g937
  (
    n1056,
    n352,
    n372,
    n264,
    n338
  );


  xnor
  g938
  (
    n666,
    n189,
    n308,
    n194,
    n280
  );


  xor
  g939
  (
    n967,
    n150,
    n294,
    n248,
    n211
  );


  and
  g940
  (
    n1036,
    n381,
    n340,
    n402,
    n255
  );


  or
  g941
  (
    n581,
    n272,
    n320,
    n291,
    n315
  );


  nand
  g942
  (
    n707,
    n146,
    n368,
    n400,
    n140
  );


  and
  g943
  (
    n791,
    n319,
    n231,
    n229,
    n162
  );


  nand
  g944
  (
    n979,
    n359,
    n271,
    n335,
    n225
  );


  or
  g945
  (
    n528,
    n380,
    n262,
    n347,
    n366
  );


  xor
  g946
  (
    n547,
    n214,
    n275,
    n186,
    n242
  );


  and
  g947
  (
    n480,
    n284,
    n253,
    n361,
    n299
  );


  and
  g948
  (
    n811,
    n220,
    n217,
    n266,
    n195
  );


  and
  g949
  (
    n727,
    n175,
    n312,
    n126,
    n212
  );


  and
  g950
  (
    n1002,
    n180,
    n173,
    n217,
    n254
  );


  xnor
  g951
  (
    n984,
    n220,
    n392,
    n178,
    n156
  );


  and
  g952
  (
    n1032,
    n254,
    n216,
    n350,
    n316
  );


  xnor
  g953
  (
    n737,
    n269,
    n188,
    n251,
    n212
  );


  or
  g954
  (
    n763,
    n299,
    n223,
    n185,
    n228
  );


  nor
  g955
  (
    n989,
    n316,
    n227,
    n339,
    n327
  );


  xnor
  g956
  (
    n725,
    n367,
    n180,
    n318,
    n216
  );


  or
  g957
  (
    n673,
    n304,
    n291,
    n361,
    n176
  );


  xor
  g958
  (
    n518,
    n184,
    n389,
    n251,
    n187
  );


  or
  g959
  (
    n1068,
    n311,
    n160,
    n294,
    n253
  );


  nor
  g960
  (
    n638,
    n197,
    n137,
    n346,
    n199
  );


  or
  g961
  (
    n980,
    n278,
    n219,
    n330,
    n161
  );


  xor
  g962
  (
    n616,
    n224,
    n155,
    n364,
    n398
  );


  nand
  g963
  (
    n713,
    n154,
    n250,
    n349,
    n229
  );


  xnor
  g964
  (
    n813,
    n357,
    n374,
    n267,
    n223
  );


  xnor
  g965
  (
    n664,
    n271,
    n325,
    n166,
    n131
  );


  xor
  g966
  (
    n990,
    n311,
    n246,
    n230,
    n265
  );


  xor
  g967
  (
    n510,
    n337,
    n301,
    n252,
    n312
  );


  xor
  g968
  (
    n582,
    n383,
    n362,
    n292,
    n190
  );


  nor
  g969
  (
    KeyWire_0_2,
    n238,
    n218,
    n375,
    n168
  );


  nor
  g970
  (
    n736,
    n343,
    n368,
    n286,
    n315
  );


  nor
  g971
  (
    n826,
    n226,
    n219,
    n333,
    n237
  );


  nor
  g972
  (
    n1039,
    n359,
    n346,
    n216,
    n212
  );


  xnor
  g973
  (
    n1022,
    n187,
    n331,
    n205,
    n246
  );


  nand
  g974
  (
    n686,
    n382,
    n219,
    n134,
    n385
  );


  xor
  g975
  (
    n867,
    n203,
    n230,
    n385,
    n127
  );


  nor
  g976
  (
    n696,
    n234,
    n286,
    n141,
    n372
  );


  nand
  g977
  (
    n1076,
    n405,
    n295,
    n345,
    n289
  );


  and
  g978
  (
    n757,
    n236,
    n296,
    n268
  );


  nor
  g979
  (
    n730,
    n390,
    n226,
    n371,
    n375
  );


  xor
  g980
  (
    n842,
    n365,
    n363,
    n140,
    n236
  );


  nor
  g981
  (
    n792,
    n192,
    n328,
    n293,
    n377
  );


  or
  g982
  (
    n735,
    n315,
    n357,
    n215,
    n145
  );


  nor
  g983
  (
    n1020,
    n220,
    n288,
    n395,
    n142
  );


  nand
  g984
  (
    n892,
    n211,
    n149,
    n249
  );


  and
  g985
  (
    n574,
    n204,
    n224,
    n165,
    n168
  );


  nand
  g986
  (
    n996,
    n314,
    n247,
    n258,
    n269
  );


  nand
  g987
  (
    n958,
    n381,
    n182,
    n163,
    n235
  );


  xor
  g988
  (
    n893,
    n221,
    n386,
    n401
  );


  xnor
  g989
  (
    n767,
    n215,
    n353,
    n283,
    n194
  );


  and
  g990
  (
    n477,
    n215,
    n200,
    n224,
    n186
  );


  nand
  g991
  (
    n1021,
    n390,
    n155,
    n352,
    n145
  );


  xnor
  g992
  (
    n726,
    n393,
    n189,
    n389,
    n368
  );


  xnor
  g993
  (
    n660,
    n278,
    n295,
    n261,
    n143
  );


  or
  g994
  (
    n704,
    n356,
    n171,
    n351,
    n369
  );


  xnor
  g995
  (
    n1093,
    n224,
    n300,
    n152,
    n229
  );


  xnor
  g996
  (
    n823,
    n192,
    n144,
    n270,
    n155
  );


  xnor
  g997
  (
    n957,
    n355,
    n322,
    n341,
    n188
  );


  xor
  g998
  (
    n799,
    n266,
    n233,
    n125,
    n301
  );


  nor
  g999
  (
    n553,
    n181,
    n253,
    n235,
    n314
  );


  and
  g1000
  (
    n564,
    n190,
    n269,
    n298,
    n257
  );


  or
  g1001
  (
    n808,
    n159,
    n205,
    n213,
    n372
  );


  xor
  g1002
  (
    n819,
    n280,
    n252,
    n260,
    n287
  );


  and
  g1003
  (
    n904,
    n207,
    n376,
    n400,
    n163
  );


  xor
  g1004
  (
    n880,
    n373,
    n130,
    n177,
    n282
  );


  xor
  g1005
  (
    n556,
    n193,
    n319,
    n245,
    n273
  );


  or
  g1006
  (
    n485,
    n257,
    n358,
    n136,
    n250
  );


  or
  g1007
  (
    n1004,
    n307,
    n366,
    n201,
    n134
  );


  nor
  g1008
  (
    n955,
    n399,
    n319,
    n179,
    n392
  );


  and
  g1009
  (
    n732,
    n397,
    n143,
    n248,
    n148
  );


  nor
  g1010
  (
    n846,
    n278,
    n131,
    n320,
    n217
  );


  xor
  g1011
  (
    n818,
    n174,
    n175,
    n393,
    n379
  );


  nand
  g1012
  (
    n834,
    n244,
    n182,
    n399,
    n260
  );


  nor
  g1013
  (
    n729,
    n203,
    n139,
    n205,
    n150
  );


  xor
  g1014
  (
    n520,
    n123,
    n312,
    n403,
    n172
  );


  nor
  g1015
  (
    n794,
    n363,
    n209,
    n282,
    n144
  );


  and
  g1016
  (
    n762,
    n285,
    n318,
    n134,
    n298
  );


  xnor
  g1017
  (
    n596,
    n226,
    n257,
    n155,
    n290
  );


  and
  g1018
  (
    n1080,
    n253,
    n209,
    n317,
    n239
  );


  and
  g1019
  (
    n812,
    n128,
    n323,
    n183,
    n264
  );


  or
  g1020
  (
    n467,
    n372,
    n364,
    n392,
    n356
  );


  or
  g1021
  (
    n951,
    n296,
    n176,
    n149,
    n401
  );


  xor
  g1022
  (
    n722,
    n289,
    n246,
    n227,
    n340
  );


  and
  g1023
  (
    n668,
    n169,
    n325,
    n282,
    n192
  );


  or
  g1024
  (
    n592,
    n324,
    n179,
    n267,
    n397
  );


  nor
  g1025
  (
    n690,
    n256,
    n328,
    n181,
    n293
  );


  or
  g1026
  (
    n742,
    n208,
    n255,
    n198,
    n393
  );


  and
  g1027
  (
    n866,
    n248,
    n123,
    n385,
    n203
  );


  xnor
  g1028
  (
    n1063,
    n364,
    n236,
    n383,
    n261
  );


  or
  g1029
  (
    n576,
    n140,
    n164,
    n203,
    n233
  );


  xor
  g1030
  (
    n636,
    n133,
    n354,
    n391,
    n258
  );


  or
  g1031
  (
    n1011,
    n213,
    n239,
    n252,
    n178
  );


  nor
  g1032
  (
    n782,
    n232,
    n137,
    n379,
    n323
  );


  xor
  g1033
  (
    n1089,
    n154,
    n265,
    n248,
    n210
  );


  xnor
  g1034
  (
    n827,
    n362,
    n238,
    n234,
    n184
  );


  nor
  g1035
  (
    n978,
    n164,
    n356,
    n332,
    n346
  );


  xnor
  g1036
  (
    n591,
    n259,
    n332,
    n239,
    n222
  );


  and
  g1037
  (
    n1042,
    n147,
    n258,
    n148,
    n391
  );


  xor
  g1038
  (
    n863,
    n321,
    n317,
    n271,
    n324
  );


  xor
  g1039
  (
    n960,
    n180,
    n267,
    n190,
    n232
  );


  nor
  g1040
  (
    KeyWire_0_7,
    n210,
    n245,
    n353,
    n354
  );


  xnor
  g1041
  (
    n471,
    n352,
    n235,
    n153,
    n287
  );


  or
  g1042
  (
    n779,
    n185,
    n147,
    n156,
    n336
  );


  nand
  g1043
  (
    n533,
    n288,
    n378,
    n131,
    n396
  );


  nand
  g1044
  (
    n609,
    n206,
    n310,
    n349,
    n245
  );


  and
  g1045
  (
    n780,
    n272,
    n191,
    n310,
    n282
  );


  nand
  g1046
  (
    n714,
    n331,
    n392,
    n359,
    n186
  );


  xor
  g1047
  (
    n806,
    n349,
    n320,
    n243,
    n329
  );


  and
  g1048
  (
    n977,
    n147,
    n365,
    n160,
    n272
  );


  nand
  g1049
  (
    n540,
    n306,
    n306,
    n345,
    n341
  );


  xor
  g1050
  (
    n717,
    n276,
    n280,
    n144,
    n199
  );


  or
  g1051
  (
    n944,
    n223,
    n158,
    n163,
    n396
  );


  xor
  g1052
  (
    n635,
    n209,
    n254,
    n377,
    n260
  );


  nor
  g1053
  (
    n1083,
    n128,
    n313,
    n198,
    n170
  );


  and
  g1054
  (
    n498,
    n210,
    n173,
    n166,
    n360
  );


  or
  g1055
  (
    n1012,
    n139,
    n291,
    n234,
    n347
  );


  or
  g1056
  (
    n878,
    n121,
    n274,
    n191,
    n331
  );


  nor
  g1057
  (
    n691,
    n353,
    n304,
    n316,
    n208
  );


  nand
  g1058
  (
    n787,
    n395,
    n371,
    n386,
    n351
  );


  xor
  g1059
  (
    n822,
    n238,
    n135,
    n193,
    n142
  );


  nor
  g1060
  (
    n922,
    n306,
    n189,
    n381,
    n183
  );


  xnor
  g1061
  (
    n524,
    n264,
    n337,
    n151,
    n139
  );


  xnor
  g1062
  (
    n662,
    n274,
    n332,
    n157,
    n394
  );


  xor
  g1063
  (
    n657,
    n380,
    n200,
    n266,
    n264
  );


  nand
  g1064
  (
    n509,
    n305,
    n195,
    n370,
    n330
  );


  and
  g1065
  (
    n1050,
    n163,
    n326,
    n383,
    n315
  );


  nand
  g1066
  (
    n723,
    n141,
    n214,
    n277,
    n161
  );


  and
  g1067
  (
    n1058,
    n303,
    n215,
    n183,
    n367
  );


  xnor
  g1068
  (
    n954,
    n205,
    n162,
    n152,
    n151
  );


  nand
  g1069
  (
    n816,
    n358,
    n344,
    n243,
    n377
  );


  xnor
  g1070
  (
    n1060,
    n370,
    n295,
    n402,
    n345
  );


  nor
  g1071
  (
    n1112,
    n887,
    n1056,
    n811,
    n518
  );


  nand
  g1072
  (
    n1246,
    n601,
    n1007,
    n889,
    n1028
  );


  or
  g1073
  (
    n1182,
    n700,
    n791,
    n538,
    n1036
  );


  and
  g1074
  (
    n1291,
    n1035,
    n637,
    n875,
    n505
  );


  or
  g1075
  (
    n1268,
    n837,
    n999,
    n486,
    n1037
  );


  nand
  g1076
  (
    n1128,
    n789,
    n1017,
    n583,
    n733
  );


  and
  g1077
  (
    n1265,
    n1002,
    n1045,
    n1025,
    n673
  );


  xor
  g1078
  (
    n1152,
    n592,
    n1016,
    n737,
    n540
  );


  nand
  g1079
  (
    n1193,
    n1001,
    n479,
    n1057,
    n1056
  );


  nand
  g1080
  (
    n1274,
    n993,
    n892,
    n1053,
    n1024
  );


  xor
  g1081
  (
    n1174,
    n1058,
    n618,
    n516,
    n463
  );


  and
  g1082
  (
    n1191,
    n406,
    n690,
    n1024,
    n968
  );


  xnor
  g1083
  (
    n1187,
    n807,
    n748,
    n405,
    n1028
  );


  and
  g1084
  (
    n1264,
    n1023,
    n669,
    n965,
    n955
  );


  nand
  g1085
  (
    n1203,
    n903,
    n407,
    n406,
    n469
  );


  and
  g1086
  (
    n1284,
    n653,
    n1005,
    n823,
    n1010
  );


  or
  g1087
  (
    n1277,
    n487,
    n899,
    n512,
    n1038
  );


  xnor
  g1088
  (
    n1161,
    n1011,
    n747,
    n997,
    n490
  );


  nor
  g1089
  (
    n1287,
    n1008,
    n740,
    n991,
    n1004
  );


  and
  g1090
  (
    n1101,
    n913,
    n559,
    n483,
    n942
  );


  nand
  g1091
  (
    n1189,
    n982,
    n876,
    n974,
    n783
  );


  xor
  g1092
  (
    n1097,
    n1058,
    n621,
    n1051,
    n663
  );


  xnor
  g1093
  (
    n1146,
    n666,
    n1020,
    n860,
    n711
  );


  xor
  g1094
  (
    n1144,
    n704,
    n1047,
    n808,
    n523
  );


  xor
  g1095
  (
    n1202,
    n667,
    n588,
    n1009,
    n616
  );


  xor
  g1096
  (
    n1234,
    n1007,
    n950,
    n987,
    n554
  );


  nand
  g1097
  (
    n1273,
    n477,
    n785,
    n992,
    n1044
  );


  xnor
  g1098
  (
    n1185,
    n932,
    n629,
    n1025,
    n741
  );


  or
  g1099
  (
    n1233,
    n956,
    n951,
    n1028,
    n794
  );


  nand
  g1100
  (
    n1210,
    n833,
    n976,
    n739,
    n979
  );


  nand
  g1101
  (
    n1109,
    n934,
    n1058,
    n914,
    n575
  );


  nand
  g1102
  (
    n1239,
    n1035,
    n746,
    n983,
    n765
  );


  xor
  g1103
  (
    n1281,
    n639,
    n688,
    n874,
    n574
  );


  nand
  g1104
  (
    n1134,
    n1059,
    n978,
    n752,
    n775
  );


  nand
  g1105
  (
    n1117,
    n727,
    n846,
    n865,
    n933
  );


  and
  g1106
  (
    n1290,
    n1057,
    n1055,
    n524,
    n936
  );


  or
  g1107
  (
    n1242,
    n743,
    n541,
    n1036,
    n949
  );


  nor
  g1108
  (
    n1236,
    n1004,
    n569,
    n1005,
    n1033
  );


  and
  g1109
  (
    n1288,
    n707,
    n1046,
    n548,
    n953
  );


  nor
  g1110
  (
    n1098,
    n528,
    n1025,
    n1015,
    n696
  );


  nor
  g1111
  (
    n1299,
    n894,
    n814,
    n879,
    n826
  );


  and
  g1112
  (
    n1162,
    n1029,
    n1034,
    n898,
    n1049
  );


  xnor
  g1113
  (
    n1119,
    n972,
    n992,
    n937,
    n582
  );


  nor
  g1114
  (
    n1296,
    n705,
    n1041,
    n999,
    n687
  );


  nor
  g1115
  (
    KeyWire_0_30,
    n699,
    n986,
    n702,
    n732
  );


  nor
  g1116
  (
    n1186,
    n1027,
    n864,
    n1039,
    n810
  );


  and
  g1117
  (
    n1136,
    n407,
    n1006,
    n646,
    n661
  );


  nand
  g1118
  (
    n1137,
    n499,
    n1042,
    n551,
    n1022
  );


  xor
  g1119
  (
    n1244,
    n763,
    n905,
    n944,
    n797
  );


  nor
  g1120
  (
    n1169,
    n710,
    n780,
    n1056,
    n1045
  );


  and
  g1121
  (
    n1200,
    n1041,
    n1050,
    n935,
    n605
  );


  and
  g1122
  (
    n1212,
    n468,
    n1037,
    n1001,
    n1021
  );


  xor
  g1123
  (
    n1141,
    n1049,
    n1020,
    n586,
    n466
  );


  xor
  g1124
  (
    n1197,
    n542,
    n1039,
    n1006,
    n973
  );


  and
  g1125
  (
    n1165,
    n851,
    n536,
    n1011,
    n754
  );


  xor
  g1126
  (
    n1159,
    n585,
    n604,
    n614,
    n762
  );


  and
  g1127
  (
    n1139,
    n998,
    n553,
    n990,
    n838
  );


  xor
  g1128
  (
    n1209,
    n994,
    n579,
    n1037,
    n460
  );


  nand
  g1129
  (
    n1247,
    n720,
    n886,
    n990,
    n1053
  );


  xnor
  g1130
  (
    n1215,
    n723,
    n495,
    n996,
    n910
  );


  xnor
  g1131
  (
    n1104,
    n576,
    n897,
    n929,
    n578
  );


  and
  g1132
  (
    n1132,
    n709,
    n1026,
    n482,
    n835
  );


  nand
  g1133
  (
    n1131,
    n842,
    n1027,
    n1000,
    n960
  );


  and
  g1134
  (
    n1301,
    n1039,
    n868,
    n654,
    n547
  );


  nand
  g1135
  (
    n1278,
    n729,
    n680,
    n921,
    n924
  );


  and
  g1136
  (
    n1107,
    n1027,
    n1032,
    n990,
    n1052
  );


  and
  g1137
  (
    n1181,
    n861,
    n781,
    n461,
    n917
  );


  nor
  g1138
  (
    n1108,
    n721,
    n497,
    n545,
    n992
  );


  and
  g1139
  (
    n1173,
    n764,
    n1040,
    n790,
    n1054
  );


  and
  g1140
  (
    n1275,
    n947,
    n1016,
    n817,
    n1030
  );


  nand
  g1141
  (
    n1262,
    n698,
    n855,
    n850,
    n788
  );


  nor
  g1142
  (
    n1178,
    n703,
    n985,
    n624,
    n757
  );


  or
  g1143
  (
    n1195,
    n776,
    n1049,
    n1031,
    n626
  );


  or
  g1144
  (
    n1280,
    n1018,
    n594,
    n1006,
    n513
  );


  xnor
  g1145
  (
    n1143,
    n907,
    n471,
    n692,
    n954
  );


  xnor
  g1146
  (
    n1164,
    n640,
    n1011,
    n844,
    n971
  );


  nor
  g1147
  (
    n1263,
    n631,
    n537,
    n1012,
    n572
  );


  xnor
  g1148
  (
    n1255,
    n465,
    n693,
    n590,
    n1043
  );


  xnor
  g1149
  (
    KeyWire_0_21,
    n998,
    n1014,
    n724,
    n676
  );


  or
  g1150
  (
    n1285,
    n1021,
    n1015,
    n1020,
    n1017
  );


  nand
  g1151
  (
    n1167,
    n577,
    n493,
    n563,
    n406
  );


  and
  g1152
  (
    n1192,
    n997,
    n1047,
    n602,
    n1014
  );


  or
  g1153
  (
    n1283,
    n998,
    n625,
    n975,
    n997
  );


  xnor
  g1154
  (
    n1116,
    n1038,
    n1053,
    n503,
    n964
  );


  xor
  g1155
  (
    n1267,
    n558,
    n1008,
    n726,
    n1057
  );


  xnor
  g1156
  (
    n1150,
    n1032,
    n830,
    n596,
    n651
  );


  xor
  g1157
  (
    n1163,
    n464,
    n501,
    n1019,
    n531
  );


  xnor
  g1158
  (
    n1276,
    n1025,
    n405,
    n925,
    n525
  );


  xnor
  g1159
  (
    n1175,
    n750,
    n598,
    n589,
    n519
  );


  nor
  g1160
  (
    n1292,
    n580,
    n535,
    n928,
    n1026
  );


  and
  g1161
  (
    n1251,
    n526,
    n694,
    n1050,
    n856
  );


  xor
  g1162
  (
    n1133,
    n1055,
    n675,
    n1037,
    n802
  );


  and
  g1163
  (
    n1124,
    n1042,
    n1013,
    n896,
    n557
  );


  xor
  g1164
  (
    n1138,
    n992,
    n859,
    n565,
    n664
  );


  nor
  g1165
  (
    n1135,
    n1045,
    n931,
    n824,
    n885
  );


  nor
  g1166
  (
    n1241,
    n866,
    n1052,
    n407,
    n1003
  );


  nor
  g1167
  (
    n1257,
    n806,
    n990,
    n970,
    n1022
  );


  xnor
  g1168
  (
    n1145,
    n660,
    n840,
    n591,
    n1023
  );


  xor
  g1169
  (
    n1240,
    n1018,
    n641,
    n803,
    n570
  );


  nand
  g1170
  (
    n1130,
    n828,
    n948,
    n995,
    n532
  );


  nand
  g1171
  (
    n1270,
    n1029,
    n561,
    n991,
    n1052
  );


  nand
  g1172
  (
    n1204,
    n798,
    n734,
    n584,
    n1015
  );


  xor
  g1173
  (
    n1170,
    n507,
    n717,
    n731,
    n800
  );


  or
  g1174
  (
    n1120,
    n945,
    n1044,
    n510,
    n1019
  );


  xor
  g1175
  (
    n1129,
    n1013,
    n728,
    n1041,
    n686
  );


  or
  g1176
  (
    n1232,
    n777,
    n478,
    n989,
    n527
  );


  and
  g1177
  (
    n1171,
    n792,
    n611,
    n782,
    n1030
  );


  or
  g1178
  (
    n1157,
    n888,
    n556,
    n1047,
    n1021
  );


  xnor
  g1179
  (
    n1252,
    n636,
    n1051,
    n595,
    n1011
  );


  xnor
  g1180
  (
    n1188,
    n679,
    n681,
    n1017,
    n890
  );


  nand
  g1181
  (
    n1211,
    n751,
    n829,
    n1008,
    n1041
  );


  nor
  g1182
  (
    n1148,
    n701,
    n564,
    n943,
    n517
  );


  and
  g1183
  (
    n1190,
    n995,
    n1029,
    n1050,
    n1047
  );


  nand
  g1184
  (
    n1103,
    n1014,
    n993,
    n984,
    n511
  );


  nand
  g1185
  (
    KeyWire_0_18,
    n994,
    n647,
    n670,
    n665
  );


  xnor
  g1186
  (
    n1219,
    n1045,
    n902,
    n714,
    n996
  );


  xnor
  g1187
  (
    n1220,
    n612,
    n650,
    n1046,
    n961
  );


  xor
  g1188
  (
    n1147,
    n1026,
    n645,
    n508,
    n1008
  );


  nor
  g1189
  (
    n1230,
    n857,
    n1043,
    n995,
    n1034
  );


  nand
  g1190
  (
    n1207,
    n1056,
    n918,
    n767,
    n996
  );


  and
  g1191
  (
    n1295,
    n927,
    n847,
    n546,
    n597
  );


  nor
  g1192
  (
    n1166,
    n1010,
    n522,
    n820,
    n539
  );


  nor
  g1193
  (
    n1260,
    n642,
    n1055,
    n1052,
    n735
  );


  xor
  g1194
  (
    n1243,
    n716,
    n843,
    n533,
    n768
  );


  xor
  g1195
  (
    n1121,
    n1007,
    n1009,
    n870,
    n1035
  );


  xor
  g1196
  (
    n1223,
    n689,
    n1042,
    n652,
    n1004
  );


  or
  g1197
  (
    n1258,
    n919,
    n872,
    n1046,
    n562
  );


  xnor
  g1198
  (
    n1127,
    n836,
    n488,
    n515,
    n644
  );


  or
  g1199
  (
    n1156,
    n869,
    n749,
    n1002,
    n656
  );


  nor
  g1200
  (
    n1229,
    n1054,
    n1048,
    n549,
    n793
  );


  xor
  g1201
  (
    n1096,
    n922,
    n1033,
    n832,
    n481
  );


  xnor
  g1202
  (
    n1153,
    n1059,
    n609,
    n1027,
    n685
  );


  and
  g1203
  (
    n1100,
    n472,
    n809,
    n1016,
    n697
  );


  or
  g1204
  (
    n1102,
    n476,
    n801,
    n957,
    n1058
  );


  nand
  g1205
  (
    n1269,
    n655,
    n1024,
    n1005,
    n755
  );


  nor
  g1206
  (
    n1125,
    n1026,
    n643,
    n1003,
    n962
  );


  nand
  g1207
  (
    n1254,
    n1001,
    n995,
    n1033,
    n1036
  );


  xor
  g1208
  (
    n1106,
    n502,
    n1022,
    n520,
    n719
  );


  xor
  g1209
  (
    n1149,
    n738,
    n952,
    n991,
    n407
  );


  and
  g1210
  (
    n1155,
    n1059,
    n881,
    n758,
    n1043
  );


  xor
  g1211
  (
    n1279,
    n993,
    n1030,
    n509,
    n635
  );


  xor
  g1212
  (
    n1261,
    n852,
    n969,
    n1020,
    n834
  );


  or
  g1213
  (
    n1235,
    n683,
    n682,
    n587,
    n462
  );


  and
  g1214
  (
    n1208,
    n930,
    n1022,
    n470,
    n786
  );


  xnor
  g1215
  (
    n1259,
    n1044,
    n1039,
    n1048,
    n867
  );


  xnor
  g1216
  (
    n1253,
    n459,
    n911,
    n713,
    n893
  );


  nor
  g1217
  (
    n1231,
    n1012,
    n521,
    n494,
    n825
  );


  and
  g1218
  (
    n1218,
    n779,
    n671,
    n759,
    n1050
  );


  or
  g1219
  (
    n1272,
    n993,
    n940,
    n648,
    n994
  );


  xnor
  g1220
  (
    n1216,
    n496,
    n606,
    n1051,
    n610
  );


  nor
  g1221
  (
    n1194,
    n678,
    n853,
    n467,
    n958
  );


  nand
  g1222
  (
    n1199,
    n1001,
    n1029,
    n1017,
    n1038
  );


  nor
  g1223
  (
    n1176,
    n492,
    n550,
    n1023,
    n573
  );


  and
  g1224
  (
    n1184,
    n1006,
    n506,
    n725,
    n1019
  );


  nor
  g1225
  (
    n1172,
    n1032,
    n848,
    n849,
    n630
  );


  nor
  g1226
  (
    n1266,
    n555,
    n474,
    n884,
    n996
  );


  xnor
  g1227
  (
    n1154,
    n514,
    n963,
    n1036,
    n674
  );


  and
  g1228
  (
    n1110,
    n581,
    n772,
    n1034,
    n1053
  );


  xor
  g1229
  (
    n1217,
    n858,
    n1040,
    n926,
    n668
  );


  nand
  g1230
  (
    n1168,
    n988,
    n742,
    n566,
    n649
  );


  and
  g1231
  (
    n1115,
    n500,
    n672,
    n1040,
    n1021
  );


  xor
  g1232
  (
    n1198,
    n760,
    n839,
    n920,
    n1019
  );


  nand
  g1233
  (
    n1228,
    n1057,
    n708,
    n1031,
    n981
  );


  xor
  g1234
  (
    n1293,
    n753,
    n534,
    n882,
    n977
  );


  and
  g1235
  (
    n1298,
    n871,
    n608,
    n900,
    n819
  );


  and
  g1236
  (
    n1140,
    n895,
    n1000,
    n543,
    n544
  );


  nand
  g1237
  (
    n1237,
    n530,
    n1002,
    n1042,
    n622
  );


  nor
  g1238
  (
    n1300,
    n1013,
    n1004,
    n1010,
    n863
  );


  nand
  g1239
  (
    n1226,
    n916,
    n1024,
    n659,
    n473
  );


  xnor
  g1240
  (
    n1179,
    n405,
    n1014,
    n706,
    n1015
  );


  nand
  g1241
  (
    n1142,
    n998,
    n770,
    n552,
    n745
  );


  xnor
  g1242
  (
    n1213,
    n1002,
    n458,
    n1031,
    n769
  );


  nor
  g1243
  (
    KeyWire_0_6,
    n923,
    n778,
    n1013,
    n796
  );


  nor
  g1244
  (
    n1126,
    n818,
    n1012,
    n1010,
    n662
  );


  xor
  g1245
  (
    n1221,
    n1054,
    n1000,
    n891,
    n633
  );


  and
  g1246
  (
    n1214,
    n912,
    n600,
    n638,
    n634
  );


  and
  g1247
  (
    n1114,
    n877,
    n1007,
    n980,
    n736
  );


  and
  g1248
  (
    n1289,
    n1043,
    n1009,
    n1038,
    n489
  );


  and
  g1249
  (
    n1206,
    n862,
    n722,
    n878,
    n677
  );


  xor
  g1250
  (
    n1205,
    n593,
    n568,
    n784,
    n1033
  );


  xor
  g1251
  (
    n1294,
    n1018,
    n915,
    n816,
    n938
  );


  xor
  g1252
  (
    n1099,
    n787,
    n504,
    n567,
    n774
  );


  nor
  g1253
  (
    n1225,
    n1005,
    n560,
    n491,
    n1054
  );


  or
  g1254
  (
    n1297,
    n408,
    n999,
    n822,
    n991
  );


  or
  g1255
  (
    n1113,
    n1003,
    n1012,
    n744,
    n997
  );


  nor
  g1256
  (
    n1227,
    n632,
    n1028,
    n946,
    n756
  );


  and
  g1257
  (
    n1249,
    n627,
    n909,
    n1018,
    n827
  );


  nor
  g1258
  (
    n1238,
    n880,
    n959,
    n715,
    n620
  );


  nand
  g1259
  (
    n1122,
    n607,
    n718,
    n712,
    n841
  );


  nand
  g1260
  (
    n1183,
    n813,
    n966,
    n831,
    n773
  );


  xor
  g1261
  (
    n1245,
    n730,
    n1051,
    n571,
    n1035
  );


  nand
  g1262
  (
    n1160,
    n480,
    n1003,
    n1048,
    n617
  );


  xor
  g1263
  (
    n1286,
    n603,
    n812,
    n805,
    n967
  );


  xnor
  g1264
  (
    n1282,
    n1023,
    n799,
    n1009,
    n1000
  );


  or
  g1265
  (
    n1224,
    n845,
    n1030,
    n761,
    n1046
  );


  nand
  g1266
  (
    n1256,
    n475,
    n766,
    n771,
    n684
  );


  nand
  g1267
  (
    n1271,
    n1032,
    n1040,
    n457,
    n599
  );


  nor
  g1268
  (
    n1118,
    n821,
    n901,
    n994,
    n1034
  );


  xnor
  g1269
  (
    n1222,
    n815,
    n695,
    n498,
    n883
  );


  and
  g1270
  (
    n1151,
    n619,
    n795,
    n999,
    n1016
  );


  nand
  g1271
  (
    n1123,
    n804,
    n485,
    n908,
    n628
  );


  and
  g1272
  (
    n1180,
    n1049,
    n1031,
    n613,
    n1044
  );


  xor
  g1273
  (
    n1111,
    n854,
    n657,
    n1048,
    n939
  );


  and
  g1274
  (
    n1250,
    n658,
    n691,
    n873,
    n1055
  );


  xor
  g1275
  (
    n1177,
    n406,
    n529,
    n615,
    n904
  );


  nor
  g1276
  (
    n1105,
    n623,
    n941,
    n484,
    n906
  );


  buf
  g1277
  (
    n1305,
    n1097
  );


  buf
  g1278
  (
    n1311,
    n1109
  );


  not
  g1279
  (
    n1314,
    n1107
  );


  not
  g1280
  (
    n1319,
    n1113
  );


  buf
  g1281
  (
    n1313,
    n1104
  );


  not
  g1282
  (
    n1303,
    n1099
  );


  buf
  g1283
  (
    n1317,
    n1098
  );


  not
  g1284
  (
    n1304,
    n1096
  );


  buf
  g1285
  (
    KeyWire_0_27,
    n1112
  );


  not
  g1286
  (
    n1318,
    n1106
  );


  not
  g1287
  (
    n1312,
    n1115
  );


  buf
  g1288
  (
    n1309,
    n1108
  );


  not
  g1289
  (
    n1306,
    n1101
  );


  buf
  g1290
  (
    n1321,
    n1103
  );


  not
  g1291
  (
    n1315,
    n1105
  );


  buf
  g1292
  (
    n1316,
    n1100
  );


  not
  g1293
  (
    n1308,
    n1114
  );


  buf
  g1294
  (
    n1307,
    n1110
  );


  buf
  g1295
  (
    n1310,
    n1102
  );


  not
  g1296
  (
    n1302,
    n1111
  );


  xor
  g1297
  (
    n1334,
    n425,
    n411,
    n417,
    n1070
  );


  xor
  g1298
  (
    n1356,
    n1302,
    n1064,
    n1304,
    n1303
  );


  xor
  g1299
  (
    n1377,
    n1316,
    n423,
    n429,
    n413
  );


  or
  g1300
  (
    n1347,
    n1061,
    n410,
    n1073,
    n1067
  );


  or
  g1301
  (
    n1381,
    n1302,
    n1303,
    n409,
    n416
  );


  xor
  g1302
  (
    n1333,
    n1061,
    n418,
    n1309,
    n1062
  );


  nor
  g1303
  (
    n1370,
    n410,
    n1308,
    n425,
    n1060
  );


  nand
  g1304
  (
    n1332,
    n1309,
    n431,
    n424,
    n1075
  );


  xnor
  g1305
  (
    n1369,
    n1315,
    n431,
    n1077,
    n1078
  );


  xor
  g1306
  (
    n1338,
    n1071,
    n411,
    n1062,
    n1312
  );


  xnor
  g1307
  (
    n1345,
    n408,
    n1305,
    n1306,
    n421
  );


  or
  g1308
  (
    n1366,
    n1072,
    n1067,
    n422,
    n417
  );


  xnor
  g1309
  (
    n1353,
    n1306,
    n414,
    n415,
    n1067
  );


  xnor
  g1310
  (
    n1348,
    n1066,
    n1061,
    n413,
    n425
  );


  xnor
  g1311
  (
    n1325,
    n1311,
    n427,
    n426,
    n1065
  );


  nand
  g1312
  (
    n1326,
    n1309,
    n1080,
    n1305,
    n418
  );


  nand
  g1313
  (
    n1355,
    n425,
    n1077,
    n1070,
    n1310
  );


  nor
  g1314
  (
    n1371,
    n1310,
    n1075,
    n426,
    n1313
  );


  xor
  g1315
  (
    n1351,
    n1309,
    n1314,
    n1313,
    n427
  );


  or
  g1316
  (
    n1349,
    n1314,
    n1059,
    n423,
    n1079
  );


  xnor
  g1317
  (
    n1358,
    n1305,
    n1310,
    n428,
    n1066
  );


  or
  g1318
  (
    n1374,
    n1080,
    n1078,
    n426
  );


  or
  g1319
  (
    n1373,
    n422,
    n409,
    n1307,
    n416
  );


  nand
  g1320
  (
    n1375,
    n430,
    n1316,
    n1313,
    n420
  );


  or
  g1321
  (
    n1341,
    n1063,
    n1074,
    n1079,
    n1075
  );


  nand
  g1322
  (
    n1368,
    n412,
    n429,
    n420,
    n419
  );


  xor
  g1323
  (
    n1346,
    n1308,
    n1315,
    n1067,
    n1071
  );


  or
  g1324
  (
    n1359,
    n1314,
    n1081,
    n421,
    n1311
  );


  xor
  g1325
  (
    n1336,
    n1314,
    n429,
    n413,
    n1306
  );


  nand
  g1326
  (
    n1378,
    n1066,
    n1315,
    n1303,
    n1074
  );


  xnor
  g1327
  (
    n1367,
    n419,
    n1062,
    n415,
    n426
  );


  xor
  g1328
  (
    n1339,
    n1065,
    n1076,
    n1063,
    n414
  );


  nor
  g1329
  (
    n1364,
    n428,
    n420,
    n1080,
    n415
  );


  or
  g1330
  (
    n1329,
    n422,
    n1063,
    n1069,
    n430
  );


  or
  g1331
  (
    n1342,
    n1062,
    n1312,
    n1071,
    n1079
  );


  or
  g1332
  (
    n1324,
    n414,
    n414,
    n1060,
    n1068
  );


  and
  g1333
  (
    KeyWire_0_29,
    n1064,
    n428,
    n1063,
    n1068
  );


  and
  g1334
  (
    n1328,
    n1065,
    n1307,
    n1073,
    n1060
  );


  nand
  g1335
  (
    n1344,
    n1070,
    n419,
    n1064,
    n431
  );


  xor
  g1336
  (
    n1327,
    n418,
    n412,
    n1069,
    n1068
  );


  and
  g1337
  (
    n1322,
    n412,
    n416,
    n1074,
    n1316
  );


  xnor
  g1338
  (
    n1363,
    n1305,
    n422,
    n410,
    n409
  );


  nand
  g1339
  (
    n1360,
    n1079,
    n419,
    n1072,
    n416
  );


  xnor
  g1340
  (
    n1335,
    n1308,
    n1302,
    n424,
    n1311
  );


  xnor
  g1341
  (
    n1372,
    n1315,
    n415,
    n1303,
    n1312
  );


  xor
  g1342
  (
    n1380,
    n430,
    n1073,
    n1080,
    n1061
  );


  xor
  g1343
  (
    n1376,
    n1078,
    n1308,
    n1065,
    n1072
  );


  nor
  g1344
  (
    n1362,
    n1069,
    n1074,
    n421,
    n427
  );


  xnor
  g1345
  (
    n1382,
    n1071,
    n418,
    n1076,
    n408
  );


  and
  g1346
  (
    KeyWire_0_31,
    n1312,
    n1310,
    n412,
    n429
  );


  nor
  g1347
  (
    n1352,
    n1081,
    n411,
    n1313,
    n1068
  );


  xor
  g1348
  (
    n1323,
    n1311,
    n1304,
    n1072,
    n420
  );


  nand
  g1349
  (
    n1340,
    n409,
    n408,
    n424,
    n1081
  );


  nor
  g1350
  (
    n1354,
    n1064,
    n1316,
    n1304,
    n417
  );


  xor
  g1351
  (
    n1337,
    n1081,
    n1317,
    n1066,
    n423
  );


  or
  g1352
  (
    n1365,
    n423,
    n1077,
    n1307,
    n427
  );


  and
  g1353
  (
    n1343,
    n411,
    n1075,
    n1304,
    n1069
  );


  or
  g1354
  (
    n1331,
    n1077,
    n410,
    n1306,
    n421
  );


  xor
  g1355
  (
    n1330,
    n1070,
    n1060,
    n1076,
    n424
  );


  nor
  g1356
  (
    n1350,
    n413,
    n1073,
    n428,
    n1307
  );


  and
  g1357
  (
    n1379,
    n1302,
    n430,
    n417,
    n1076
  );


  nand
  g1358
  (
    n1384,
    n1335,
    n1155,
    n1332,
    n1152
  );


  xor
  g1359
  (
    n1391,
    n1133,
    n1325,
    n1118,
    n1127
  );


  or
  g1360
  (
    n1398,
    n1336,
    n1324,
    n1151,
    n1141
  );


  and
  g1361
  (
    n1397,
    n1126,
    n1138,
    n1140,
    n1135
  );


  nand
  g1362
  (
    n1392,
    n1160,
    n1123,
    n1124,
    n1329
  );


  xnor
  g1363
  (
    n1386,
    n1322,
    n1158,
    n1129,
    n1163
  );


  nor
  g1364
  (
    n1383,
    n1120,
    n1117,
    n1161,
    n1147
  );


  nand
  g1365
  (
    n1387,
    n1331,
    n1137,
    n1136,
    n1330
  );


  or
  g1366
  (
    n1395,
    n1333,
    n1328,
    n1122,
    n1159
  );


  or
  g1367
  (
    n1389,
    n1156,
    n1327,
    n1153,
    n1131
  );


  xor
  g1368
  (
    n1393,
    n1119,
    n1134,
    n1337,
    n1128
  );


  xor
  g1369
  (
    n1396,
    n1125,
    n1146,
    n1143,
    n1145
  );


  and
  g1370
  (
    n1388,
    n1323,
    n1132,
    n1157,
    n1148
  );


  nand
  g1371
  (
    n1390,
    n1154,
    n1130,
    n1121,
    n1139
  );


  nor
  g1372
  (
    n1385,
    n1162,
    n1116,
    n1149,
    n1150
  );


  and
  g1373
  (
    n1394,
    n1142,
    n1326,
    n1334,
    n1144
  );


  and
  g1374
  (
    n1410,
    n1390,
    n1082,
    n1083,
    n1172
  );


  nor
  g1375
  (
    n1402,
    n1183,
    n1202,
    n1084,
    n1187
  );


  nand
  g1376
  (
    n1407,
    n1177,
    n1188,
    n1389,
    n1169
  );


  or
  g1377
  (
    n1399,
    n1383,
    n1190,
    n1168,
    n1388
  );


  nor
  g1378
  (
    n1406,
    n1388,
    n1171,
    n1082,
    n1195
  );


  nor
  g1379
  (
    n1412,
    n1192,
    n1186,
    n1083,
    n1391
  );


  nor
  g1380
  (
    n1405,
    n1083,
    n1389,
    n1173,
    n1200
  );


  xor
  g1381
  (
    n1401,
    n1181,
    n1082,
    n1385,
    n1084
  );


  xor
  g1382
  (
    n1408,
    n1179,
    n1387,
    n1205,
    n1203
  );


  xor
  g1383
  (
    n1403,
    n1196,
    n1390,
    n1191,
    n1197
  );


  xnor
  g1384
  (
    n1400,
    n1189,
    n1182,
    n1198,
    n1388
  );


  and
  g1385
  (
    n1415,
    n1180,
    n1389,
    n1175,
    n1199
  );


  or
  g1386
  (
    n1416,
    n1390,
    n1174,
    n1185,
    n1166
  );


  nand
  g1387
  (
    n1413,
    n1167,
    n1384,
    n1184,
    n1389
  );


  xor
  g1388
  (
    n1404,
    n1170,
    n1084,
    n1164,
    n1386
  );


  nand
  g1389
  (
    n1409,
    n1193,
    n1165,
    n1390,
    n1204
  );


  or
  g1390
  (
    n1414,
    n1178,
    n1391,
    n1083,
    n1201
  );


  or
  g1391
  (
    n1411,
    n1084,
    n1082,
    n1176,
    n1194
  );


  xnor
  g1392
  (
    n1417,
    n1208,
    n1206,
    n1399,
    n1207
  );


  xnor
  g1393
  (
    n1418,
    n1209,
    n1215,
    n1417,
    n1210
  );


  xnor
  g1394
  (
    n1420,
    n1211,
    n1212,
    n1417,
    n1214
  );


  xnor
  g1395
  (
    n1419,
    n1417,
    n1216,
    n1217,
    n1213
  );


  xnor
  g1396
  (
    n1428,
    n1218,
    n1226,
    n1339,
    n1419
  );


  nor
  g1397
  (
    n1421,
    n1420,
    n1229,
    n1338,
    n1340
  );


  xnor
  g1398
  (
    n1424,
    n1228,
    n1419,
    n1341
  );


  nand
  g1399
  (
    n1422,
    n1221,
    n1418,
    n1085
  );


  nor
  g1400
  (
    n1429,
    n1087,
    n1086,
    n1085
  );


  xnor
  g1401
  (
    n1430,
    n1220,
    n1418,
    n1222,
    n1342
  );


  xor
  g1402
  (
    n1426,
    n1227,
    n1420,
    n1219,
    n1317
  );


  nor
  g1403
  (
    n1425,
    n1085,
    n1086,
    n1230,
    n1418
  );


  and
  g1404
  (
    n1423,
    n1317,
    n1419,
    n1224,
    n1085
  );


  nand
  g1405
  (
    n1427,
    n1223,
    n1317,
    n1086,
    n1225
  );


  buf
  g1406
  (
    n1431,
    n1423
  );


  not
  g1407
  (
    n1433,
    n1421
  );


  not
  g1408
  (
    n1434,
    n1424
  );


  buf
  g1409
  (
    n1432,
    n1422
  );


  nand
  g1410
  (
    n1442,
    n1432,
    n1431,
    n1411
  );


  nand
  g1411
  (
    n1440,
    n1318,
    n1403,
    n1432,
    n1431
  );


  or
  g1412
  (
    n1438,
    n1319,
    n1320,
    n1410
  );


  xor
  g1413
  (
    n1444,
    n1406,
    n1402,
    n1318,
    n1414
  );


  and
  g1414
  (
    n1439,
    n1432,
    n1391,
    n1319
  );


  and
  g1415
  (
    n1437,
    n1432,
    n1318,
    n1405,
    n1407
  );


  xnor
  g1416
  (
    n1435,
    n1318,
    n1401,
    n1433,
    n1319
  );


  and
  g1417
  (
    n1443,
    n1431,
    n1413,
    n1412,
    n1404
  );


  nand
  g1418
  (
    n1441,
    n1409,
    n1415,
    n1408,
    n1416
  );


  nand
  g1419
  (
    n1436,
    n1433,
    n1391,
    n1320,
    n1400
  );


  buf
  g1420
  (
    n1448,
    n1437
  );


  buf
  g1421
  (
    n1453,
    n1439
  );


  not
  g1422
  (
    n1452,
    n1440
  );


  buf
  g1423
  (
    n1446,
    n1442
  );


  buf
  g1424
  (
    n1445,
    n1441
  );


  buf
  g1425
  (
    n1449,
    n1438
  );


  xnor
  g1426
  (
    n1447,
    n1233,
    n1425,
    n1443,
    n1426
  );


  nor
  g1427
  (
    n1451,
    n1426,
    n1232,
    n1435,
    n1436
  );


  or
  g1428
  (
    n1450,
    n1231,
    n1234,
    n1425
  );


  nor
  g1429
  (
    n1464,
    n1427,
    n1447,
    n1430,
    n1446
  );


  and
  g1430
  (
    n1465,
    n1448,
    n1428,
    n1429,
    n1088
  );


  nor
  g1431
  (
    n1462,
    n1420,
    n1087,
    n1427
  );


  and
  g1432
  (
    n1454,
    n1448,
    n1235,
    n432,
    n1428
  );


  nand
  g1433
  (
    n1458,
    n1433,
    n1420,
    n1237,
    n1447
  );


  or
  g1434
  (
    n1460,
    n1426,
    n1087,
    n1446
  );


  xor
  g1435
  (
    n1461,
    n1429,
    n1446,
    n1447,
    n1427
  );


  xor
  g1436
  (
    n1459,
    n1448,
    n1238,
    n1089,
    n431
  );


  xnor
  g1437
  (
    n1466,
    n1445,
    n1429,
    n1088,
    n432
  );


  nand
  g1438
  (
    n1457,
    n432,
    n1434,
    n1428
  );


  nor
  g1439
  (
    n1467,
    n1430,
    n1445,
    n1088,
    n1434
  );


  and
  g1440
  (
    n1455,
    n1434,
    n1429,
    n1428,
    n1446
  );


  nand
  g1441
  (
    n1463,
    n1089,
    n1430,
    n1445
  );


  xnor
  g1442
  (
    n1456,
    n1447,
    n1236,
    n1433,
    n1088
  );


  not
  g1443
  (
    n1469,
    n1460
  );


  buf
  g1444
  (
    n1470,
    n1459
  );


  not
  g1445
  (
    n1471,
    n1461
  );


  not
  g1446
  (
    n1468,
    n1462
  );


  or
  g1447
  (
    n1480,
    n1464,
    n1467,
    n1450,
    n1452
  );


  nand
  g1448
  (
    n1484,
    n1469,
    n1453,
    n1450,
    n1243
  );


  nand
  g1449
  (
    n1482,
    n1453,
    n1453,
    n1452,
    n1449
  );


  xor
  g1450
  (
    n1478,
    n1449,
    n1449,
    n1089,
    n1444
  );


  nand
  g1451
  (
    n1476,
    n1470,
    n1451,
    n1090,
    n1471
  );


  xor
  g1452
  (
    n1474,
    n1469,
    n1451,
    n1468,
    n1090
  );


  and
  g1453
  (
    n1472,
    n1090,
    n1465,
    n1450,
    n1468
  );


  nor
  g1454
  (
    n1485,
    n1241,
    n1091,
    n1470,
    n1471
  );


  xor
  g1455
  (
    n1481,
    n1471,
    n1449,
    n1448,
    n1453
  );


  xor
  g1456
  (
    n1475,
    n1470,
    n1091,
    n1463,
    n1451
  );


  nand
  g1457
  (
    n1473,
    n1242,
    n1444,
    n1452,
    n1466
  );


  xnor
  g1458
  (
    n1479,
    n1469,
    n1444,
    n1091,
    n1090
  );


  and
  g1459
  (
    n1477,
    n433,
    n1089,
    n1470,
    n1240
  );


  xnor
  g1460
  (
    n1486,
    n1471,
    n1469,
    n432,
    n1468
  );


  or
  g1461
  (
    n1483,
    n1239,
    n1451,
    n1450,
    n1452
  );


  nor
  g1462
  (
    n1495,
    n1480,
    n1472,
    n1476,
    n1479
  );


  nor
  g1463
  (
    n1493,
    n1477,
    n1476,
    n1480,
    n1473
  );


  nor
  g1464
  (
    n1488,
    n1476,
    n1478,
    n1475
  );


  nor
  g1465
  (
    n1490,
    n1477,
    n1474,
    n1478
  );


  xnor
  g1466
  (
    n1491,
    n1472,
    n1477,
    n1476
  );


  xor
  g1467
  (
    n1487,
    n1474,
    n1473,
    n1478,
    n1472
  );


  xor
  g1468
  (
    n1489,
    n1480,
    n1475,
    n1478
  );


  nor
  g1469
  (
    n1494,
    n1472,
    n1479,
    n1480
  );


  xnor
  g1470
  (
    n1492,
    n1479,
    n1474,
    n1473
  );


  not
  g1471
  (
    n1502,
    n1482
  );


  not
  g1472
  (
    n1498,
    n1482
  );


  buf
  g1473
  (
    n1501,
    n433
  );


  buf
  g1474
  (
    KeyWire_0_3,
    n1493
  );


  not
  g1475
  (
    n1503,
    n1495
  );


  not
  g1476
  (
    n1499,
    n1494
  );


  nor
  g1477
  (
    n1500,
    n1482,
    n1489,
    n1487
  );


  and
  g1478
  (
    n1496,
    n1490,
    n1481,
    n1091,
    n1482
  );


  or
  g1479
  (
    n1497,
    n1495,
    n1481
  );


  nor
  g1480
  (
    n1504,
    n1481,
    n1483,
    n1495
  );


  and
  g1481
  (
    n1505,
    n1492,
    n433,
    n1488,
    n1491
  );


  xnor
  g1482
  (
    KeyWire_0_14,
    n1499,
    n1483,
    n1496,
    n1486
  );


  nand
  g1483
  (
    n1511,
    n440,
    n1498,
    n1484
  );


  and
  g1484
  (
    n1515,
    n436,
    n1498,
    n438,
    n1496
  );


  xor
  g1485
  (
    n1514,
    n1498,
    n439
  );


  or
  g1486
  (
    n1509,
    n1497,
    n1496,
    n437,
    n440
  );


  and
  g1487
  (
    n1516,
    n1486,
    n441,
    n1497,
    n434
  );


  or
  g1488
  (
    n1510,
    n441,
    n1497,
    n1483,
    n438
  );


  xnor
  g1489
  (
    n1521,
    n1484,
    n441,
    n1496,
    n1499
  );


  and
  g1490
  (
    n1517,
    n442,
    n433,
    n1498,
    n1485
  );


  nand
  g1491
  (
    n1519,
    n437,
    n434,
    n440,
    n1499
  );


  xnor
  g1492
  (
    n1520,
    n440,
    n1485,
    n438,
    n1497
  );


  and
  g1493
  (
    n1507,
    n436,
    n437,
    n1485
  );


  nand
  g1494
  (
    n1512,
    n1486,
    n435,
    n439
  );


  xor
  g1495
  (
    n1508,
    n436,
    n435,
    n1486,
    n441
  );


  nor
  g1496
  (
    n1522,
    n436,
    n1485,
    n1499,
    n438
  );


  nand
  g1497
  (
    n1513,
    n434,
    n434,
    n1484,
    n435
  );


  and
  g1498
  (
    n1525,
    n1500,
    n1520,
    n444,
    n1092
  );


  xnor
  g1499
  (
    n1530,
    n446,
    n445,
    n1519
  );


  nor
  g1500
  (
    n1524,
    n1500,
    n1092,
    n445,
    n1522
  );


  nor
  g1501
  (
    n1528,
    n1516,
    n1515,
    n444,
    n1092
  );


  xor
  g1502
  (
    n1526,
    n1518,
    n442,
    n1500,
    n443
  );


  xor
  g1503
  (
    n1523,
    n443,
    n444
  );


  nand
  g1504
  (
    n1529,
    n446,
    n443,
    n1521,
    n1517
  );


  or
  g1505
  (
    n1527,
    n1500,
    n445,
    n442
  );


  xor
  g1506
  (
    n1535,
    n1528,
    n1529,
    n116,
    n1246
  );


  xor
  g1507
  (
    n1544,
    n1524,
    n1501,
    n447,
    n115
  );


  nand
  g1508
  (
    n1545,
    n1523,
    n1530,
    n1261,
    n1525
  );


  nor
  g1509
  (
    n1552,
    n110,
    n113,
    n114,
    n1273
  );


  xnor
  g1510
  (
    n1536,
    n113,
    n1258,
    n1530,
    n1504
  );


  or
  g1511
  (
    n1561,
    n1525,
    n1505,
    n1501,
    n1502
  );


  or
  g1512
  (
    n1557,
    n1502,
    n1528,
    n114,
    n110
  );


  nor
  g1513
  (
    n1531,
    n1272,
    n447,
    n1506,
    n1527
  );


  nand
  g1514
  (
    n1541,
    n112,
    n110,
    n1506,
    n1248
  );


  and
  g1515
  (
    n1559,
    n1503,
    n109,
    n1249,
    n447
  );


  xor
  g1516
  (
    n1534,
    n1504,
    n1251,
    n1267,
    n1501
  );


  nor
  g1517
  (
    KeyWire_0_22,
    n1262,
    n448,
    n1530,
    n1255
  );


  xnor
  g1518
  (
    n1547,
    n112,
    n446,
    n1524,
    n1260
  );


  nand
  g1519
  (
    n1549,
    n1266,
    n1526,
    n1506,
    n1529
  );


  nor
  g1520
  (
    n1558,
    n1257,
    n110,
    n1504,
    n1524
  );


  nor
  g1521
  (
    n1538,
    n1526,
    n112,
    n109,
    n114
  );


  and
  g1522
  (
    n1556,
    n1525,
    n1501,
    n1528,
    n1529
  );


  xnor
  g1523
  (
    n1548,
    n1529,
    n1523,
    n111,
    n1259
  );


  xor
  g1524
  (
    n1553,
    n109,
    n1504,
    n1530,
    n1524
  );


  xnor
  g1525
  (
    n1540,
    n1523,
    n1244,
    n109,
    n1502
  );


  or
  g1526
  (
    n1543,
    n1506,
    n1527,
    n116,
    n1503
  );


  nor
  g1527
  (
    n1532,
    n1503,
    n117,
    n1250,
    n1264
  );


  or
  g1528
  (
    n1554,
    n1526,
    n1505,
    n111,
    n1254
  );


  or
  g1529
  (
    n1560,
    n113,
    n1527,
    n116,
    n448
  );


  xor
  g1530
  (
    n1542,
    n446,
    n1270,
    n1263,
    n1528
  );


  or
  g1531
  (
    n1537,
    n1523,
    n111,
    n114,
    n1271
  );


  xnor
  g1532
  (
    n1550,
    n115,
    n1527,
    n1526,
    n1268
  );


  nand
  g1533
  (
    n1551,
    n1265,
    n117,
    n1502,
    n1505
  );


  and
  g1534
  (
    n1562,
    n113,
    n1252,
    n112,
    n115
  );


  xor
  g1535
  (
    n1539,
    n115,
    n1245,
    n1269,
    n1247
  );


  xnor
  g1536
  (
    n1555,
    n447,
    n1503,
    n1505,
    n1253
  );


  nor
  g1537
  (
    n1546,
    n1525,
    n116,
    n111,
    n1256
  );


  nor
  g1538
  (
    n1563,
    n450,
    n449,
    n1538,
    n452
  );


  xor
  g1539
  (
    n1565,
    n448,
    n452,
    n450,
    n449
  );


  nand
  g1540
  (
    n1569,
    n1533,
    n1531,
    n451,
    n1539
  );


  xor
  g1541
  (
    KeyWire_0_8,
    n448,
    n451,
    n1535,
    n449
  );


  and
  g1542
  (
    n1566,
    n452,
    n453,
    n451,
    n450
  );


  nor
  g1543
  (
    n1568,
    n1536,
    n449,
    n450,
    n452
  );


  xnor
  g1544
  (
    n1567,
    n1532,
    n1534,
    n1537,
    n451
  );


  xor
  g1545
  (
    n1570,
    n454,
    n455
  );


  xnor
  g1546
  (
    n1574,
    n1565,
    n456,
    n453
  );


  and
  g1547
  (
    n1572,
    n453,
    n454,
    n1567,
    n1564
  );


  nor
  g1548
  (
    n1571,
    n454,
    n454,
    n453,
    n1563
  );


  nand
  g1549
  (
    n1573,
    n1566,
    n455,
    n456
  );


  not
  g1550
  (
    n1576,
    n1572
  );


  buf
  g1551
  (
    n1578,
    n1570
  );


  buf
  g1552
  (
    n1577,
    n1573
  );


  not
  g1553
  (
    n1575,
    n1571
  );


  nor
  g1554
  (
    n1588,
    n1575,
    n1277,
    n1552,
    n1549
  );


  xnor
  g1555
  (
    n1582,
    n1542,
    n1094,
    n1276,
    n1553
  );


  or
  g1556
  (
    n1587,
    n1577,
    n1093,
    n1554
  );


  and
  g1557
  (
    n1580,
    n1094,
    n1576,
    n1092,
    n1275
  );


  nand
  g1558
  (
    n1584,
    n1095,
    n1550,
    n1545,
    n1548
  );


  nor
  g1559
  (
    n1586,
    n1093,
    n1577,
    n1547,
    n1551
  );


  and
  g1560
  (
    n1583,
    n1544,
    n1575,
    n1541,
    n1543
  );


  xor
  g1561
  (
    n1585,
    n1094,
    n1576,
    n1278,
    n1274
  );


  nand
  g1562
  (
    n1579,
    n1575,
    n1576,
    n1540,
    n1094
  );


  nand
  g1563
  (
    n1581,
    n1576,
    n1546,
    n1093,
    n1575
  );


  buf
  g1564
  (
    n1591,
    n1580
  );


  buf
  g1565
  (
    n1589,
    n1580
  );


  not
  g1566
  (
    n1590,
    n1579
  );


  not
  g1567
  (
    n1592,
    n1580
  );


  nand
  g1568
  (
    n1603,
    n1291,
    n1589,
    n1590,
    n1288
  );


  xor
  g1569
  (
    n1608,
    n1556,
    n1577,
    n1289,
    n1591
  );


  and
  g1570
  (
    n1606,
    n1294,
    n1569,
    n1562,
    n1282
  );


  nor
  g1571
  (
    n1597,
    n1284,
    n1321,
    n1568,
    n1561
  );


  xnor
  g1572
  (
    n1602,
    n1589,
    n1562,
    n1560,
    n1592
  );


  nor
  g1573
  (
    n1593,
    n1562,
    n1560,
    n1591,
    n1286
  );


  nor
  g1574
  (
    n1596,
    n1577,
    n1590,
    n1280,
    n1320
  );


  or
  g1575
  (
    n1604,
    n1590,
    n1559,
    n1292
  );


  and
  g1576
  (
    n1601,
    n1561,
    n1592,
    n1321
  );


  and
  g1577
  (
    n1605,
    n1591,
    n1558,
    n1560
  );


  xnor
  g1578
  (
    KeyWire_0_15,
    n1321,
    n1290,
    n1578,
    n1555
  );


  xnor
  g1579
  (
    n1594,
    n1293,
    n1578,
    n1561,
    n1558
  );


  xor
  g1580
  (
    n1598,
    n1321,
    n1287,
    n1558,
    n1557
  );


  nor
  g1581
  (
    n1599,
    n1279,
    n1589,
    n1591
  );


  and
  g1582
  (
    n1600,
    n1590,
    n1281,
    n1559,
    n1283
  );


  xor
  g1583
  (
    n1607,
    n1285,
    n1562,
    n1561,
    n1592
  );


  nand
  g1584
  (
    n1615,
    n1585,
    n120,
    n1597,
    n1593
  );


  nand
  g1585
  (
    n1613,
    n120,
    n1584,
    n1588,
    n1582
  );


  nand
  g1586
  (
    n1619,
    n1601,
    n119,
    n118,
    n1587
  );


  or
  g1587
  (
    n1617,
    n1583,
    n1578,
    n1596,
    n1587
  );


  xor
  g1588
  (
    n1614,
    n1587,
    n1588,
    n1603,
    n117
  );


  xnor
  g1589
  (
    KeyWire_0_26,
    n1585,
    n1602,
    n1578,
    n1584
  );


  and
  g1590
  (
    n1618,
    n119,
    n1582,
    n1585,
    n1594
  );


  and
  g1591
  (
    n1609,
    n1599,
    n1583,
    n1582,
    n1602
  );


  and
  g1592
  (
    n1621,
    n1602,
    n1586,
    n1584
  );


  and
  g1593
  (
    n1624,
    n1581,
    n118,
    n1583,
    n117
  );


  nor
  g1594
  (
    n1610,
    n1588,
    n119,
    n120
  );


  or
  g1595
  (
    n1622,
    n1595,
    n1581,
    n1600,
    n1588
  );


  xnor
  g1596
  (
    n1623,
    n1581,
    n118,
    n1602
  );


  nand
  g1597
  (
    n1620,
    n1582,
    n1586,
    n1583,
    n1603
  );


  xnor
  g1598
  (
    n1616,
    n119,
    n1585,
    n1584,
    n1587
  );


  xor
  g1599
  (
    n1612,
    n1574,
    n1603,
    n1598,
    n1586
  );


  not
  g1600
  (
    n1629,
    n1619
  );


  buf
  g1601
  (
    n1627,
    n1622
  );


  not
  g1602
  (
    n1626,
    n1618
  );


  not
  g1603
  (
    n1625,
    n1620
  );


  buf
  g1604
  (
    n1628,
    n1621
  );


  nand
  g1605
  (
    n1630,
    n1625,
    n1095
  );


  xor
  g1606
  (
    n1631,
    n1300,
    n1296,
    n1630,
    n1299
  );


  and
  g1607
  (
    n1632,
    n1630,
    n1298,
    n1295,
    n1297
  );


  xnor
  g1608
  (
    n1634,
    n1632,
    n1604,
    n1605
  );


  or
  g1609
  (
    n1636,
    n1606,
    n1605,
    n1607
  );


  xnor
  g1610
  (
    n1633,
    n1605,
    n1607,
    n1604
  );


  and
  g1611
  (
    n1635,
    n1603,
    n1632,
    n1631
  );


  nand
  g1612
  (
    n1637,
    n1632,
    n1606
  );


  nor
  g1613
  (
    n1647,
    n1379,
    n1361,
    n1627,
    n1355
  );


  and
  g1614
  (
    n1649,
    n1633,
    n1637,
    n1353,
    n1381
  );


  xor
  g1615
  (
    n1648,
    n1354,
    n1358,
    n1608,
    n1637
  );


  xnor
  g1616
  (
    n1642,
    n1370,
    n1345,
    n1377,
    n1343
  );


  xor
  g1617
  (
    n1638,
    n1628,
    n1624,
    n1351,
    n1347
  );


  xnor
  g1618
  (
    n1653,
    n1635,
    n1365,
    n1637,
    n1608
  );


  xor
  g1619
  (
    n1645,
    n1367,
    n1629,
    n1372,
    n1607
  );


  xor
  g1620
  (
    n1641,
    n1356,
    n1627,
    n1359,
    n1607
  );


  xnor
  g1621
  (
    n1643,
    n1637,
    n1608,
    n1362,
    n1629
  );


  and
  g1622
  (
    n1650,
    n1629,
    n1636,
    n1346,
    n1371
  );


  nand
  g1623
  (
    KeyWire_0_1,
    n1623,
    n1378,
    n1357,
    n1349
  );


  nor
  g1624
  (
    n1646,
    n1633,
    n1626,
    n1369,
    n1350
  );


  or
  g1625
  (
    n1639,
    n1634,
    n1635,
    n1363
  );


  xor
  g1626
  (
    n1651,
    n1360,
    n1628,
    n1635,
    n1608
  );


  xor
  g1627
  (
    n1644,
    n1368,
    n1636,
    n1633,
    n1352
  );


  or
  g1628
  (
    n1656,
    n1628,
    n1634,
    n1633,
    n1344
  );


  or
  g1629
  (
    n1655,
    n1376,
    n1382,
    n1366,
    n1636
  );


  and
  g1630
  (
    n1640,
    n1634,
    n1636,
    n1364,
    n1301
  );


  nand
  g1631
  (
    n1654,
    n1348,
    n1374,
    n1375,
    n1634
  );


  xor
  g1632
  (
    n1652,
    n1628,
    n1629,
    n1373,
    n1380
  );


  nor
  g1633
  (
    n1658,
    n1397,
    n1396,
    n1398,
    n1394
  );


  xnor
  g1634
  (
    n1668,
    n1396,
    n1395,
    n1648,
    n1394
  );


  and
  g1635
  (
    n1664,
    n1652,
    n1393,
    n1646,
    n1638
  );


  and
  g1636
  (
    KeyWire_0_12,
    n1397,
    n1654,
    n1650,
    n1644
  );


  nor
  g1637
  (
    n1666,
    n1651,
    n1397,
    n1640,
    n1396
  );


  or
  g1638
  (
    n1662,
    n1393,
    n1393,
    n1392,
    n1639
  );


  xnor
  g1639
  (
    n1659,
    n1655,
    n1397,
    n1398,
    n1642
  );


  nand
  g1640
  (
    n1661,
    n1398,
    n1395,
    n1656
  );


  xor
  g1641
  (
    n1669,
    n1392,
    n1394,
    n1653,
    n1647
  );


  xor
  g1642
  (
    n1667,
    n1395,
    n1396,
    n1398,
    n1394
  );


  or
  g1643
  (
    n1660,
    n1392,
    n1649,
    n1643,
    n1645
  );


  nand
  g1644
  (
    n1665,
    n1392,
    n1393,
    n1657,
    n1641
  );


  xnor
  g1645
  (
    n1670,
    n1659,
    n1668,
    n1666,
    n1667
  );


  xnor
  g1646
  (
    n1672,
    n1664,
    n1660,
    n1669,
    n1662
  );


  or
  g1647
  (
    n1671,
    n1665,
    n1663,
    n1658,
    n1661
  );


  xor
  KeyGate_0_0
  (
    n688,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1657,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1084,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1506,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n639,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n35,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1248,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n643,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1564,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n219,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n741,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1047,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1663,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n437,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1518,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n1595,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n718,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1095,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1158,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n594,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1008,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1196,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n1533,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1001,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n879,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n469,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1611,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1320,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n898,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n1361,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1201,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1357,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

