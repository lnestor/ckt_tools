

module Stat_1046_20_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n1020,
  n1014,
  n1015,
  n1016,
  n1018,
  n1049,
  n1042,
  n1047,
  n1043,
  n1053,
  n1051,
  n1033,
  n1040,
  n1034,
  n1044,
  n1032,
  n1050,
  n1048,
  n1046,
  n1038,
  n1071,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1020;output n1014;output n1015;output n1016;output n1018;output n1049;output n1042;output n1047;output n1043;output n1053;output n1051;output n1033;output n1040;output n1034;output n1044;output n1032;output n1050;output n1048;output n1046;output n1038;output n1071;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1017;wire n1019;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1035;wire n1036;wire n1037;wire n1039;wire n1041;wire n1045;wire n1052;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n59,
    n25
  );


  buf
  g1
  (
    n35,
    n22
  );


  not
  g2
  (
    n32,
    n11
  );


  buf
  g3
  (
    n112,
    n20
  );


  buf
  g4
  (
    n92,
    n16
  );


  not
  g5
  (
    n42,
    n11
  );


  buf
  g6
  (
    n62,
    n22
  );


  buf
  g7
  (
    n115,
    n13
  );


  not
  g8
  (
    n36,
    n12
  );


  not
  g9
  (
    n77,
    n10
  );


  buf
  g10
  (
    n29,
    n19
  );


  buf
  g11
  (
    n110,
    n1
  );


  buf
  g12
  (
    n71,
    n13
  );


  buf
  g13
  (
    n124,
    n2
  );


  not
  g14
  (
    n44,
    n24
  );


  not
  g15
  (
    n96,
    n5
  );


  buf
  g16
  (
    n83,
    n17
  );


  not
  g17
  (
    n63,
    n15
  );


  buf
  g18
  (
    n57,
    n20
  );


  buf
  g19
  (
    n38,
    n6
  );


  not
  g20
  (
    n40,
    n14
  );


  buf
  g21
  (
    n27,
    n4
  );


  not
  g22
  (
    n94,
    n17
  );


  buf
  g23
  (
    n108,
    n18
  );


  not
  g24
  (
    n50,
    n14
  );


  not
  g25
  (
    n75,
    n7
  );


  not
  g26
  (
    n87,
    n25
  );


  buf
  g27
  (
    n54,
    n14
  );


  buf
  g28
  (
    n118,
    n3
  );


  not
  g29
  (
    n49,
    n21
  );


  not
  g30
  (
    n56,
    n15
  );


  buf
  g31
  (
    n122,
    n22
  );


  buf
  g32
  (
    n66,
    n19
  );


  buf
  g33
  (
    n123,
    n6
  );


  not
  g34
  (
    n72,
    n16
  );


  buf
  g35
  (
    n125,
    n17
  );


  not
  g36
  (
    n116,
    n2
  );


  not
  g37
  (
    n89,
    n5
  );


  not
  g38
  (
    n98,
    n10
  );


  buf
  g39
  (
    n41,
    n16
  );


  not
  g40
  (
    n101,
    n10
  );


  not
  g41
  (
    n119,
    n12
  );


  not
  g42
  (
    n74,
    n9
  );


  not
  g43
  (
    n82,
    n10
  );


  buf
  g44
  (
    n104,
    n25
  );


  not
  g45
  (
    n47,
    n2
  );


  not
  g46
  (
    n46,
    n5
  );


  buf
  g47
  (
    n73,
    n23
  );


  buf
  g48
  (
    n97,
    n16
  );


  not
  g49
  (
    n111,
    n13
  );


  buf
  g50
  (
    n88,
    n20
  );


  not
  g51
  (
    n65,
    n1
  );


  not
  g52
  (
    n106,
    n9
  );


  buf
  g53
  (
    n90,
    n12
  );


  buf
  g54
  (
    n30,
    n8
  );


  not
  g55
  (
    n51,
    n8
  );


  not
  g56
  (
    n113,
    n21
  );


  buf
  g57
  (
    n76,
    n3
  );


  not
  g58
  (
    n79,
    n21
  );


  not
  g59
  (
    n69,
    n15
  );


  not
  g60
  (
    n60,
    n11
  );


  buf
  g61
  (
    n80,
    n13
  );


  not
  g62
  (
    n53,
    n6
  );


  not
  g63
  (
    n95,
    n12
  );


  buf
  g64
  (
    n67,
    n18
  );


  not
  g65
  (
    n99,
    n23
  );


  not
  g66
  (
    n34,
    n11
  );


  buf
  g67
  (
    n91,
    n2
  );


  not
  g68
  (
    n81,
    n3
  );


  buf
  g69
  (
    n58,
    n23
  );


  buf
  g70
  (
    n45,
    n19
  );


  buf
  g71
  (
    n33,
    n18
  );


  buf
  g72
  (
    n26,
    n21
  );


  not
  g73
  (
    n31,
    n1
  );


  not
  g74
  (
    n78,
    n7
  );


  not
  g75
  (
    n48,
    n9
  );


  not
  g76
  (
    n28,
    n14
  );


  buf
  g77
  (
    n55,
    n8
  );


  not
  g78
  (
    n68,
    n5
  );


  not
  g79
  (
    n107,
    n17
  );


  not
  g80
  (
    n109,
    n22
  );


  not
  g81
  (
    n70,
    n25
  );


  buf
  g82
  (
    n102,
    n24
  );


  not
  g83
  (
    n114,
    n4
  );


  not
  g84
  (
    n84,
    n8
  );


  buf
  g85
  (
    n100,
    n20
  );


  buf
  g86
  (
    n86,
    n6
  );


  buf
  g87
  (
    n61,
    n7
  );


  buf
  g88
  (
    n93,
    n4
  );


  buf
  g89
  (
    n103,
    n7
  );


  not
  g90
  (
    n120,
    n1
  );


  not
  g91
  (
    n85,
    n19
  );


  not
  g92
  (
    n105,
    n24
  );


  not
  g93
  (
    n117,
    n24
  );


  buf
  g94
  (
    KeyWire_0_2,
    n18
  );


  not
  g95
  (
    n52,
    n23
  );


  not
  g96
  (
    n64,
    n9
  );


  buf
  g97
  (
    n39,
    n3
  );


  buf
  g98
  (
    n37,
    n4
  );


  not
  g99
  (
    n43,
    n15
  );


  buf
  g100
  (
    n328,
    n44
  );


  buf
  g101
  (
    n389,
    n111
  );


  buf
  g102
  (
    n268,
    n104
  );


  not
  g103
  (
    n145,
    n114
  );


  buf
  g104
  (
    n164,
    n90
  );


  buf
  g105
  (
    n150,
    n79
  );


  not
  g106
  (
    n421,
    n33
  );


  buf
  g107
  (
    n146,
    n40
  );


  not
  g108
  (
    n376,
    n96
  );


  not
  g109
  (
    n281,
    n32
  );


  buf
  g110
  (
    KeyWire_0_25,
    n75
  );


  buf
  g111
  (
    KeyWire_0_9,
    n48
  );


  not
  g112
  (
    n353,
    n118
  );


  not
  g113
  (
    n235,
    n81
  );


  buf
  g114
  (
    n203,
    n42
  );


  buf
  g115
  (
    n149,
    n82
  );


  buf
  g116
  (
    n296,
    n52
  );


  not
  g117
  (
    n291,
    n87
  );


  not
  g118
  (
    n129,
    n113
  );


  not
  g119
  (
    n357,
    n40
  );


  buf
  g120
  (
    n254,
    n106
  );


  not
  g121
  (
    n229,
    n108
  );


  buf
  g122
  (
    n304,
    n66
  );


  not
  g123
  (
    n356,
    n81
  );


  not
  g124
  (
    n209,
    n83
  );


  not
  g125
  (
    n270,
    n52
  );


  buf
  g126
  (
    n190,
    n114
  );


  not
  g127
  (
    n211,
    n63
  );


  not
  g128
  (
    n132,
    n98
  );


  not
  g129
  (
    n240,
    n106
  );


  not
  g130
  (
    n228,
    n108
  );


  buf
  g131
  (
    n382,
    n92
  );


  not
  g132
  (
    n162,
    n111
  );


  not
  g133
  (
    n364,
    n115
  );


  not
  g134
  (
    n180,
    n109
  );


  buf
  g135
  (
    n276,
    n75
  );


  not
  g136
  (
    n323,
    n38
  );


  not
  g137
  (
    n142,
    n101
  );


  not
  g138
  (
    n166,
    n71
  );


  buf
  g139
  (
    n206,
    n91
  );


  not
  g140
  (
    n222,
    n117
  );


  not
  g141
  (
    n322,
    n55
  );


  buf
  g142
  (
    n195,
    n31
  );


  buf
  g143
  (
    n255,
    n88
  );


  not
  g144
  (
    n262,
    n37
  );


  not
  g145
  (
    n163,
    n37
  );


  not
  g146
  (
    n422,
    n117
  );


  not
  g147
  (
    n303,
    n94
  );


  not
  g148
  (
    n175,
    n35
  );


  buf
  g149
  (
    n143,
    n29
  );


  not
  g150
  (
    n367,
    n54
  );


  buf
  g151
  (
    n196,
    n92
  );


  not
  g152
  (
    n324,
    n62
  );


  buf
  g153
  (
    n212,
    n104
  );


  not
  g154
  (
    n371,
    n68
  );


  not
  g155
  (
    n340,
    n117
  );


  not
  g156
  (
    n373,
    n96
  );


  not
  g157
  (
    n370,
    n55
  );


  buf
  g158
  (
    n266,
    n44
  );


  not
  g159
  (
    n396,
    n72
  );


  buf
  g160
  (
    n297,
    n121
  );


  not
  g161
  (
    n401,
    n109
  );


  not
  g162
  (
    n326,
    n76
  );


  buf
  g163
  (
    n273,
    n93
  );


  not
  g164
  (
    n147,
    n63
  );


  buf
  g165
  (
    KeyWire_0_4,
    n105
  );


  not
  g166
  (
    n365,
    n39
  );


  buf
  g167
  (
    n137,
    n80
  );


  buf
  g168
  (
    n355,
    n102
  );


  not
  g169
  (
    n290,
    n59
  );


  not
  g170
  (
    n127,
    n84
  );


  not
  g171
  (
    n295,
    n93
  );


  buf
  g172
  (
    n408,
    n77
  );


  buf
  g173
  (
    n292,
    n39
  );


  buf
  g174
  (
    n413,
    n58
  );


  buf
  g175
  (
    n181,
    n35
  );


  buf
  g176
  (
    n378,
    n72
  );


  buf
  g177
  (
    n397,
    n109
  );


  buf
  g178
  (
    n253,
    n35
  );


  not
  g179
  (
    n139,
    n119
  );


  not
  g180
  (
    n243,
    n48
  );


  not
  g181
  (
    n360,
    n60
  );


  not
  g182
  (
    n199,
    n54
  );


  buf
  g183
  (
    n411,
    n70
  );


  buf
  g184
  (
    n284,
    n49
  );


  buf
  g185
  (
    n395,
    n67
  );


  not
  g186
  (
    n171,
    n42
  );


  not
  g187
  (
    n403,
    n97
  );


  not
  g188
  (
    n272,
    n113
  );


  not
  g189
  (
    KeyWire_0_6,
    n105
  );


  buf
  g190
  (
    n156,
    n101
  );


  not
  g191
  (
    n423,
    n96
  );


  buf
  g192
  (
    n336,
    n65
  );


  not
  g193
  (
    n305,
    n98
  );


  not
  g194
  (
    n242,
    n117
  );


  buf
  g195
  (
    KeyWire_0_1,
    n36
  );


  not
  g196
  (
    n309,
    n74
  );


  buf
  g197
  (
    n167,
    n54
  );


  not
  g198
  (
    n264,
    n83
  );


  not
  g199
  (
    n354,
    n58
  );


  not
  g200
  (
    n289,
    n38
  );


  buf
  g201
  (
    n213,
    n52
  );


  not
  g202
  (
    n398,
    n39
  );


  buf
  g203
  (
    n417,
    n111
  );


  not
  g204
  (
    n188,
    n86
  );


  buf
  g205
  (
    n249,
    n109
  );


  not
  g206
  (
    n241,
    n114
  );


  not
  g207
  (
    n218,
    n99
  );


  buf
  g208
  (
    n148,
    n77
  );


  not
  g209
  (
    n233,
    n39
  );


  buf
  g210
  (
    KeyWire_0_16,
    n46
  );


  buf
  g211
  (
    n133,
    n71
  );


  buf
  g212
  (
    n221,
    n100
  );


  not
  g213
  (
    n252,
    n32
  );


  buf
  g214
  (
    n178,
    n84
  );


  not
  g215
  (
    n189,
    n40
  );


  buf
  g216
  (
    n332,
    n33
  );


  not
  g217
  (
    n329,
    n54
  );


  not
  g218
  (
    n191,
    n116
  );


  buf
  g219
  (
    n311,
    n98
  );


  buf
  g220
  (
    n391,
    n62
  );


  not
  g221
  (
    n394,
    n26
  );


  not
  g222
  (
    KeyWire_0_17,
    n80
  );


  not
  g223
  (
    n339,
    n27
  );


  not
  g224
  (
    n186,
    n67
  );


  buf
  g225
  (
    n207,
    n118
  );


  not
  g226
  (
    n239,
    n74
  );


  not
  g227
  (
    n414,
    n76
  );


  buf
  g228
  (
    n280,
    n82
  );


  buf
  g229
  (
    n306,
    n75
  );


  not
  g230
  (
    n138,
    n100
  );


  buf
  g231
  (
    n251,
    n105
  );


  buf
  g232
  (
    n381,
    n34
  );


  buf
  g233
  (
    n154,
    n113
  );


  not
  g234
  (
    n232,
    n62
  );


  buf
  g235
  (
    n294,
    n68
  );


  not
  g236
  (
    n317,
    n89
  );


  not
  g237
  (
    n351,
    n41
  );


  not
  g238
  (
    n177,
    n51
  );


  not
  g239
  (
    KeyWire_0_20,
    n38
  );


  not
  g240
  (
    n275,
    n118
  );


  not
  g241
  (
    n410,
    n112
  );


  buf
  g242
  (
    n238,
    n51
  );


  buf
  g243
  (
    n141,
    n27
  );


  not
  g244
  (
    n308,
    n53
  );


  not
  g245
  (
    n214,
    n78
  );


  not
  g246
  (
    n227,
    n106
  );


  buf
  g247
  (
    n259,
    n31
  );


  not
  g248
  (
    n344,
    n61
  );


  not
  g249
  (
    n318,
    n46
  );


  not
  g250
  (
    n205,
    n29
  );


  not
  g251
  (
    n346,
    n67
  );


  buf
  g252
  (
    n320,
    n48
  );


  not
  g253
  (
    n247,
    n41
  );


  buf
  g254
  (
    n193,
    n50
  );


  buf
  g255
  (
    n299,
    n45
  );


  buf
  g256
  (
    n341,
    n103
  );


  not
  g257
  (
    n271,
    n28
  );


  not
  g258
  (
    n237,
    n26
  );


  not
  g259
  (
    n263,
    n107
  );


  not
  g260
  (
    n159,
    n115
  );


  buf
  g261
  (
    n361,
    n61
  );


  not
  g262
  (
    n377,
    n110
  );


  buf
  g263
  (
    n334,
    n73
  );


  not
  g264
  (
    n282,
    n80
  );


  buf
  g265
  (
    n165,
    n72
  );


  buf
  g266
  (
    n220,
    n82
  );


  buf
  g267
  (
    n316,
    n83
  );


  buf
  g268
  (
    n315,
    n80
  );


  not
  g269
  (
    n134,
    n99
  );


  buf
  g270
  (
    n170,
    n120
  );


  not
  g271
  (
    n173,
    n31
  );


  buf
  g272
  (
    n285,
    n85
  );


  buf
  g273
  (
    n256,
    n99
  );


  not
  g274
  (
    n385,
    n120
  );


  not
  g275
  (
    n368,
    n32
  );


  buf
  g276
  (
    n418,
    n86
  );


  buf
  g277
  (
    n161,
    n113
  );


  not
  g278
  (
    n404,
    n38
  );


  buf
  g279
  (
    n380,
    n116
  );


  buf
  g280
  (
    n208,
    n42
  );


  buf
  g281
  (
    KeyWire_0_21,
    n61
  );


  not
  g282
  (
    n257,
    n75
  );


  buf
  g283
  (
    n302,
    n85
  );


  not
  g284
  (
    n277,
    n110
  );


  not
  g285
  (
    n183,
    n64
  );


  buf
  g286
  (
    n347,
    n36
  );


  not
  g287
  (
    n325,
    n36
  );


  buf
  g288
  (
    KeyWire_0_7,
    n84
  );


  not
  g289
  (
    n250,
    n92
  );


  buf
  g290
  (
    n168,
    n72
  );


  buf
  g291
  (
    n331,
    n96
  );


  buf
  g292
  (
    n374,
    n30
  );


  not
  g293
  (
    n261,
    n69
  );


  not
  g294
  (
    n187,
    n79
  );


  buf
  g295
  (
    n210,
    n45
  );


  buf
  g296
  (
    n388,
    n71
  );


  buf
  g297
  (
    n293,
    n103
  );


  not
  g298
  (
    n267,
    n94
  );


  buf
  g299
  (
    n269,
    n46
  );


  not
  g300
  (
    n307,
    n34
  );


  not
  g301
  (
    n366,
    n53
  );


  not
  g302
  (
    n202,
    n64
  );


  not
  g303
  (
    n384,
    n62
  );


  not
  g304
  (
    n260,
    n65
  );


  not
  g305
  (
    n246,
    n34
  );


  buf
  g306
  (
    n225,
    n49
  );


  not
  g307
  (
    n416,
    n118
  );


  buf
  g308
  (
    n258,
    n100
  );


  not
  g309
  (
    n185,
    n93
  );


  buf
  g310
  (
    n363,
    n34
  );


  buf
  g311
  (
    n409,
    n63
  );


  buf
  g312
  (
    n279,
    n91
  );


  not
  g313
  (
    n359,
    n94
  );


  buf
  g314
  (
    n201,
    n97
  );


  buf
  g315
  (
    n330,
    n74
  );


  buf
  g316
  (
    n224,
    n119
  );


  buf
  g317
  (
    n400,
    n115
  );


  buf
  g318
  (
    n236,
    n66
  );


  buf
  g319
  (
    n379,
    n43
  );


  not
  g320
  (
    n230,
    n33
  );


  not
  g321
  (
    n226,
    n28
  );


  buf
  g322
  (
    n152,
    n45
  );


  buf
  g323
  (
    n349,
    n63
  );


  buf
  g324
  (
    n198,
    n74
  );


  buf
  g325
  (
    n223,
    n49
  );


  buf
  g326
  (
    n286,
    n120
  );


  not
  g327
  (
    n415,
    n29
  );


  buf
  g328
  (
    n372,
    n30
  );


  buf
  g329
  (
    n406,
    n60
  );


  not
  g330
  (
    n369,
    n43
  );


  not
  g331
  (
    n265,
    n55
  );


  not
  g332
  (
    n300,
    n66
  );


  buf
  g333
  (
    n169,
    n85
  );


  buf
  g334
  (
    n153,
    n70
  );


  buf
  g335
  (
    n128,
    n59
  );


  buf
  g336
  (
    n200,
    n64
  );


  not
  g337
  (
    n287,
    n27
  );


  buf
  g338
  (
    n362,
    n98
  );


  not
  g339
  (
    n350,
    n82
  );


  buf
  g340
  (
    n278,
    n51
  );


  not
  g341
  (
    n126,
    n104
  );


  not
  g342
  (
    n197,
    n102
  );


  not
  g343
  (
    n245,
    n77
  );


  buf
  g344
  (
    n312,
    n110
  );


  buf
  g345
  (
    n182,
    n69
  );


  buf
  g346
  (
    n321,
    n49
  );


  buf
  g347
  (
    n313,
    n108
  );


  not
  g348
  (
    n131,
    n86
  );


  not
  g349
  (
    n335,
    n120
  );


  not
  g350
  (
    n219,
    n47
  );


  buf
  g351
  (
    n244,
    n40
  );


  not
  g352
  (
    n338,
    n30
  );


  buf
  g353
  (
    n283,
    n90
  );


  buf
  g354
  (
    n160,
    n58
  );


  not
  g355
  (
    n402,
    n89
  );


  not
  g356
  (
    n342,
    n30
  );


  buf
  g357
  (
    n343,
    n101
  );


  buf
  g358
  (
    n204,
    n47
  );


  not
  g359
  (
    n194,
    n28
  );


  buf
  g360
  (
    n135,
    n100
  );


  buf
  g361
  (
    n319,
    n119
  );


  buf
  g362
  (
    n176,
    n32
  );


  buf
  g363
  (
    n298,
    n45
  );


  buf
  g364
  (
    n174,
    n53
  );


  not
  g365
  (
    n333,
    n55
  );


  not
  g366
  (
    n157,
    n26
  );


  not
  g367
  (
    n387,
    n95
  );


  not
  g368
  (
    n231,
    n104
  );


  buf
  g369
  (
    n412,
    n107
  );


  xor
  g370
  (
    n144,
    n57,
    n43,
    n88,
    n91
  );


  nor
  g371
  (
    n216,
    n102,
    n105,
    n110,
    n65
  );


  nor
  g372
  (
    n337,
    n37,
    n88,
    n27,
    n101
  );


  or
  g373
  (
    n419,
    n50,
    n106,
    n116,
    n69
  );


  or
  g374
  (
    n288,
    n73,
    n112,
    n70,
    n37
  );


  and
  g375
  (
    n155,
    n26,
    n51,
    n50,
    n78
  );


  and
  g376
  (
    n215,
    n44,
    n57,
    n70,
    n73
  );


  xnor
  g377
  (
    n248,
    n56,
    n47,
    n35,
    n97
  );


  nand
  g378
  (
    n301,
    n33,
    n56,
    n61
  );


  nor
  g379
  (
    n348,
    n60,
    n103,
    n71,
    n58
  );


  and
  g380
  (
    n420,
    n78,
    n67,
    n59
  );


  xnor
  g381
  (
    n130,
    n87,
    n114,
    n89,
    n91
  );


  and
  g382
  (
    n310,
    n93,
    n48,
    n52,
    n81
  );


  or
  g383
  (
    n392,
    n85,
    n57,
    n79
  );


  and
  g384
  (
    n172,
    n41,
    n84,
    n90,
    n87
  );


  nor
  g385
  (
    KeyWire_0_29,
    n95,
    n115,
    n43,
    n97
  );


  nand
  g386
  (
    n192,
    n121,
    n112,
    n56,
    n44
  );


  nand
  g387
  (
    n352,
    n50,
    n66,
    n29,
    n42
  );


  and
  g388
  (
    n136,
    n95,
    n103,
    n68,
    n65
  );


  xor
  g389
  (
    n184,
    n36,
    n28,
    n90,
    n60
  );


  nor
  g390
  (
    n158,
    n107,
    n99,
    n77,
    n68
  );


  nand
  g391
  (
    n399,
    n94,
    n47,
    n53,
    n116
  );


  xor
  g392
  (
    n234,
    n87,
    n31,
    n46,
    n111
  );


  nand
  g393
  (
    n405,
    n81,
    n88,
    n41,
    n119
  );


  or
  g394
  (
    n390,
    n83,
    n64,
    n107,
    n92
  );


  xor
  g395
  (
    n140,
    n73,
    n69,
    n102,
    n89
  );


  nor
  g396
  (
    n358,
    n78,
    n95,
    n112,
    n86
  );


  xnor
  g397
  (
    n393,
    n108,
    n76,
    n57
  );


  buf
  g398
  (
    n559,
    n401
  );


  buf
  g399
  (
    n501,
    n137
  );


  not
  g400
  (
    n462,
    n405
  );


  not
  g401
  (
    KeyWire_0_18,
    n199
  );


  not
  g402
  (
    n449,
    n416
  );


  not
  g403
  (
    n620,
    n140
  );


  buf
  g404
  (
    n459,
    n239
  );


  not
  g405
  (
    n483,
    n225
  );


  buf
  g406
  (
    KeyWire_0_5,
    n417
  );


  buf
  g407
  (
    n496,
    n310
  );


  not
  g408
  (
    n486,
    n262
  );


  buf
  g409
  (
    n550,
    n254
  );


  not
  g410
  (
    n546,
    n409
  );


  not
  g411
  (
    n468,
    n155
  );


  not
  g412
  (
    n473,
    n211
  );


  buf
  g413
  (
    n520,
    n298
  );


  buf
  g414
  (
    n553,
    n419
  );


  buf
  g415
  (
    n564,
    n388
  );


  not
  g416
  (
    n622,
    n381
  );


  not
  g417
  (
    n545,
    n332
  );


  not
  g418
  (
    n528,
    n404
  );


  buf
  g419
  (
    n603,
    n361
  );


  buf
  g420
  (
    n600,
    n409
  );


  not
  g421
  (
    n508,
    n385
  );


  buf
  g422
  (
    n618,
    n218
  );


  buf
  g423
  (
    n482,
    n313
  );


  buf
  g424
  (
    n605,
    n148
  );


  not
  g425
  (
    n439,
    n127
  );


  buf
  g426
  (
    n525,
    n191
  );


  buf
  g427
  (
    n594,
    n166
  );


  buf
  g428
  (
    n572,
    n280
  );


  not
  g429
  (
    n437,
    n412
  );


  buf
  g430
  (
    n460,
    n221
  );


  not
  g431
  (
    n441,
    n349
  );


  buf
  g432
  (
    n587,
    n295
  );


  buf
  g433
  (
    n596,
    n245
  );


  not
  g434
  (
    n613,
    n241
  );


  buf
  g435
  (
    n498,
    n227
  );


  not
  g436
  (
    n466,
    n357
  );


  not
  g437
  (
    n476,
    n396
  );


  buf
  g438
  (
    n591,
    n244
  );


  not
  g439
  (
    n541,
    n371
  );


  not
  g440
  (
    n563,
    n407
  );


  not
  g441
  (
    n532,
    n350
  );


  buf
  g442
  (
    n581,
    n418
  );


  buf
  g443
  (
    n531,
    n272
  );


  not
  g444
  (
    n509,
    n412
  );


  buf
  g445
  (
    n542,
    n387
  );


  buf
  g446
  (
    n503,
    n401
  );


  not
  g447
  (
    n457,
    n405
  );


  buf
  g448
  (
    n555,
    n392
  );


  not
  g449
  (
    n463,
    n356
  );


  buf
  g450
  (
    n454,
    n268
  );


  buf
  g451
  (
    n526,
    n216
  );


  buf
  g452
  (
    n608,
    n267
  );


  not
  g453
  (
    n464,
    n386
  );


  not
  g454
  (
    n538,
    n233
  );


  not
  g455
  (
    n616,
    n173
  );


  not
  g456
  (
    n549,
    n365
  );


  buf
  g457
  (
    n442,
    n418
  );


  buf
  g458
  (
    n495,
    n215
  );


  not
  g459
  (
    n478,
    n286
  );


  buf
  g460
  (
    n604,
    n398
  );


  not
  g461
  (
    n621,
    n396
  );


  buf
  g462
  (
    n598,
    n400
  );


  buf
  g463
  (
    n443,
    n399
  );


  buf
  g464
  (
    KeyWire_0_24,
    n184
  );


  not
  g465
  (
    n534,
    n383
  );


  not
  g466
  (
    n516,
    n144
  );


  buf
  g467
  (
    n585,
    n407
  );


  not
  g468
  (
    n456,
    n395
  );


  not
  g469
  (
    n461,
    n327
  );


  not
  g470
  (
    n433,
    n150
  );


  not
  g471
  (
    n432,
    n346
  );


  buf
  g472
  (
    n446,
    n400
  );


  not
  g473
  (
    n584,
    n419
  );


  buf
  g474
  (
    n597,
    n415
  );


  buf
  g475
  (
    n575,
    n411
  );


  not
  g476
  (
    n610,
    n279
  );


  not
  g477
  (
    n448,
    n305
  );


  buf
  g478
  (
    n440,
    n414
  );


  not
  g479
  (
    n588,
    n408
  );


  buf
  g480
  (
    n609,
    n402
  );


  not
  g481
  (
    n434,
    n275
  );


  not
  g482
  (
    n453,
    n354
  );


  not
  g483
  (
    n519,
    n363
  );


  not
  g484
  (
    n494,
    n363
  );


  not
  g485
  (
    n576,
    n281
  );


  buf
  g486
  (
    n471,
    n384
  );


  not
  g487
  (
    n429,
    n373
  );


  buf
  g488
  (
    n497,
    n411
  );


  buf
  g489
  (
    n565,
    n260
  );


  not
  g490
  (
    n615,
    n371
  );


  not
  g491
  (
    n580,
    n415
  );


  buf
  g492
  (
    n424,
    n373
  );


  buf
  g493
  (
    n554,
    n196
  );


  not
  g494
  (
    KeyWire_0_11,
    n256
  );


  buf
  g495
  (
    n537,
    n374
  );


  not
  g496
  (
    n477,
    n186
  );


  not
  g497
  (
    n493,
    n394
  );


  buf
  g498
  (
    n571,
    n364
  );


  not
  g499
  (
    n527,
    n389
  );


  not
  g500
  (
    n578,
    n419
  );


  buf
  g501
  (
    n570,
    n315
  );


  not
  g502
  (
    n548,
    n230
  );


  buf
  g503
  (
    n522,
    n179
  );


  buf
  g504
  (
    n436,
    n405
  );


  buf
  g505
  (
    n487,
    n338
  );


  not
  g506
  (
    n540,
    n365
  );


  buf
  g507
  (
    n518,
    n171
  );


  buf
  g508
  (
    n427,
    n377
  );


  not
  g509
  (
    n455,
    n183
  );


  not
  g510
  (
    n491,
    n367
  );


  buf
  g511
  (
    n517,
    n362
  );


  not
  g512
  (
    n558,
    n253
  );


  not
  g513
  (
    n617,
    n217
  );


  not
  g514
  (
    n595,
    n167
  );


  buf
  g515
  (
    n511,
    n411
  );


  not
  g516
  (
    n623,
    n379
  );


  buf
  g517
  (
    n474,
    n408
  );


  buf
  g518
  (
    n431,
    n411
  );


  not
  g519
  (
    n438,
    n231
  );


  buf
  g520
  (
    n450,
    n282
  );


  buf
  g521
  (
    n430,
    n247
  );


  not
  g522
  (
    n592,
    n158
  );


  buf
  g523
  (
    n512,
    n135
  );


  buf
  g524
  (
    n467,
    n188
  );


  not
  g525
  (
    KeyWire_0_22,
    n406
  );


  buf
  g526
  (
    n606,
    n401
  );


  buf
  g527
  (
    n561,
    n169
  );


  not
  g528
  (
    n586,
    n293
  );


  buf
  g529
  (
    n485,
    n278
  );


  not
  g530
  (
    n614,
    n403
  );


  xnor
  g531
  (
    n544,
    n415,
    n388,
    n270
  );


  xnor
  g532
  (
    n490,
    n189,
    n136,
    n399,
    n202
  );


  nand
  g533
  (
    n529,
    n381,
    n416,
    n408,
    n157
  );


  nor
  g534
  (
    n515,
    n128,
    n328,
    n333,
    n208
  );


  xnor
  g535
  (
    n547,
    n403,
    n406,
    n318,
    n133
  );


  xnor
  g536
  (
    n472,
    n257,
    n214,
    n154,
    n190
  );


  and
  g537
  (
    n480,
    n251,
    n405,
    n391,
    n366
  );


  xnor
  g538
  (
    n444,
    n141,
    n300,
    n409,
    n417
  );


  xnor
  g539
  (
    n543,
    n307,
    n395,
    n209,
    n134
  );


  and
  g540
  (
    n425,
    n195,
    n416,
    n240,
    n370
  );


  or
  g541
  (
    n452,
    n403,
    n410,
    n418,
    n250
  );


  xnor
  g542
  (
    n577,
    n398,
    n414,
    n314,
    n368
  );


  and
  g543
  (
    n451,
    n168,
    n376,
    n418,
    n229
  );


  and
  g544
  (
    n602,
    n283,
    n181,
    n413,
    n206
  );


  and
  g545
  (
    n513,
    n159,
    n263,
    n362,
    n163
  );


  xor
  g546
  (
    n500,
    n384,
    n367,
    n355,
    n242
  );


  and
  g547
  (
    n539,
    n324,
    n406,
    n311,
    n330
  );


  xnor
  g548
  (
    n445,
    n285,
    n175,
    n419,
    n265
  );


  xnor
  g549
  (
    n562,
    n177,
    n224,
    n308,
    n336
  );


  or
  g550
  (
    n524,
    n347,
    n234,
    n129,
    n248
  );


  xor
  g551
  (
    n568,
    n382,
    n397,
    n152,
    n200
  );


  and
  g552
  (
    n514,
    n370,
    n301,
    n413,
    n299
  );


  or
  g553
  (
    n612,
    n219,
    n326,
    n138,
    n126
  );


  or
  g554
  (
    n533,
    n376,
    n352,
    n397,
    n404
  );


  nor
  g555
  (
    n574,
    n382,
    n412,
    n383,
    n296
  );


  xnor
  g556
  (
    n428,
    n368,
    n403,
    n372,
    n304
  );


  xnor
  g557
  (
    n535,
    n130,
    n153,
    n243,
    n390
  );


  and
  g558
  (
    n489,
    n170,
    n359,
    n412,
    n132
  );


  and
  g559
  (
    n510,
    n297,
    n402,
    n249,
    n415
  );


  and
  g560
  (
    n479,
    n151,
    n303,
    n386,
    n145
  );


  xor
  g561
  (
    n492,
    n409,
    n162,
    n187,
    n391
  );


  xor
  g562
  (
    n536,
    n342,
    n156,
    n287,
    n372
  );


  or
  g563
  (
    n569,
    n407,
    n406,
    n420,
    n400
  );


  xor
  g564
  (
    n573,
    n174,
    n139,
    n237,
    n316
  );


  or
  g565
  (
    n601,
    n178,
    n198,
    n375,
    n417
  );


  or
  g566
  (
    n582,
    n292,
    n399,
    n176,
    n375
  );


  and
  g567
  (
    n560,
    n374,
    n402,
    n320,
    n369
  );


  xnor
  g568
  (
    n607,
    n213,
    n259,
    n197,
    n274
  );


  or
  g569
  (
    n469,
    n339,
    n389,
    n193,
    n341
  );


  nor
  g570
  (
    n499,
    n210,
    n345,
    n393,
    n390
  );


  or
  g571
  (
    n593,
    n204,
    n246,
    n331,
    n238
  );


  xnor
  g572
  (
    n481,
    n325,
    n322,
    n165,
    n414
  );


  xnor
  g573
  (
    n556,
    n266,
    n416,
    n340,
    n261
  );


  and
  g574
  (
    n521,
    n258,
    n172,
    n402,
    n398
  );


  or
  g575
  (
    n551,
    n321,
    n401,
    n180,
    n417
  );


  or
  g576
  (
    n523,
    n410,
    n410,
    n212,
    n407
  );


  xnor
  g577
  (
    KeyWire_0_19,
    n205,
    n353,
    n379,
    n276
  );


  xnor
  g578
  (
    n447,
    n378,
    n226,
    n413,
    n164
  );


  xor
  g579
  (
    n619,
    n392,
    n397,
    n264,
    n400
  );


  and
  g580
  (
    n599,
    n337,
    n236,
    n147,
    n377
  );


  xnor
  g581
  (
    n484,
    n410,
    n142,
    n358,
    n387
  );


  xor
  g582
  (
    n589,
    n323,
    n161,
    n220,
    n317
  );


  or
  g583
  (
    n458,
    n420,
    n291,
    n334,
    n306
  );


  nand
  g584
  (
    n435,
    n273,
    n309,
    n344,
    n329
  );


  or
  g585
  (
    n567,
    n394,
    n351,
    n223,
    n290
  );


  and
  g586
  (
    n507,
    n194,
    n203,
    n271,
    n319
  );


  nor
  g587
  (
    n557,
    n185,
    n207,
    n277,
    n131
  );


  xnor
  g588
  (
    KeyWire_0_12,
    n143,
    n289,
    n414,
    n232
  );


  nand
  g589
  (
    n426,
    n360,
    n201,
    n404,
    n149
  );


  or
  g590
  (
    n505,
    n408,
    n399,
    n192,
    n335
  );


  nand
  g591
  (
    n506,
    n284,
    n222,
    n182,
    n413
  );


  and
  g592
  (
    n504,
    n294,
    n255,
    n380,
    n235
  );


  nand
  g593
  (
    n611,
    n404,
    n343,
    n378,
    n288
  );


  nor
  g594
  (
    n465,
    n366,
    n228,
    n369,
    n302
  );


  or
  g595
  (
    n470,
    n380,
    n312,
    n385,
    n146
  );


  nand
  g596
  (
    n488,
    n397,
    n393,
    n364,
    n348
  );


  and
  g597
  (
    KeyWire_0_27,
    n252,
    n160,
    n398,
    n269
  );


  buf
  g598
  (
    KeyWire_0_3,
    n611
  );


  buf
  g599
  (
    n783,
    n588
  );


  not
  g600
  (
    n729,
    n497
  );


  not
  g601
  (
    n692,
    n454
  );


  not
  g602
  (
    n708,
    n530
  );


  not
  g603
  (
    n716,
    n503
  );


  not
  g604
  (
    n733,
    n504
  );


  not
  g605
  (
    n720,
    n528
  );


  not
  g606
  (
    n706,
    n523
  );


  buf
  g607
  (
    n719,
    n510
  );


  not
  g608
  (
    n661,
    n531
  );


  buf
  g609
  (
    n786,
    n576
  );


  not
  g610
  (
    n691,
    n426
  );


  buf
  g611
  (
    n656,
    n519
  );


  buf
  g612
  (
    n637,
    n606
  );


  buf
  g613
  (
    n702,
    n458
  );


  buf
  g614
  (
    n646,
    n478
  );


  not
  g615
  (
    n684,
    n490
  );


  not
  g616
  (
    n703,
    n509
  );


  buf
  g617
  (
    n765,
    n442
  );


  not
  g618
  (
    n794,
    n500
  );


  buf
  g619
  (
    n690,
    n592
  );


  buf
  g620
  (
    n739,
    n494
  );


  not
  g621
  (
    KeyWire_0_26,
    n595
  );


  buf
  g622
  (
    n761,
    n526
  );


  buf
  g623
  (
    n774,
    n566
  );


  buf
  g624
  (
    n798,
    n541
  );


  buf
  g625
  (
    n705,
    n506
  );


  not
  g626
  (
    n704,
    n601
  );


  buf
  g627
  (
    n649,
    n425
  );


  buf
  g628
  (
    n693,
    n584
  );


  not
  g629
  (
    n662,
    n420
  );


  not
  g630
  (
    n771,
    n618
  );


  not
  g631
  (
    n689,
    n439
  );


  not
  g632
  (
    n767,
    n533
  );


  not
  g633
  (
    n773,
    n456
  );


  not
  g634
  (
    n743,
    n433
  );


  not
  g635
  (
    n792,
    n483
  );


  not
  g636
  (
    n759,
    n516
  );


  buf
  g637
  (
    n751,
    n556
  );


  buf
  g638
  (
    n632,
    n448
  );


  not
  g639
  (
    n781,
    n596
  );


  buf
  g640
  (
    n640,
    n515
  );


  not
  g641
  (
    n747,
    n590
  );


  not
  g642
  (
    n688,
    n614
  );


  not
  g643
  (
    KeyWire_0_15,
    n571
  );


  buf
  g644
  (
    n659,
    n473
  );


  not
  g645
  (
    n731,
    n543
  );


  not
  g646
  (
    n666,
    n492
  );


  not
  g647
  (
    n727,
    n451
  );


  not
  g648
  (
    n777,
    n487
  );


  buf
  g649
  (
    n757,
    n529
  );


  buf
  g650
  (
    n707,
    n455
  );


  not
  g651
  (
    n634,
    n466
  );


  not
  g652
  (
    n764,
    n517
  );


  buf
  g653
  (
    n795,
    n615
  );


  not
  g654
  (
    n698,
    n482
  );


  buf
  g655
  (
    n700,
    n604
  );


  not
  g656
  (
    n676,
    n430
  );


  buf
  g657
  (
    n658,
    n484
  );


  buf
  g658
  (
    n709,
    n472
  );


  buf
  g659
  (
    n730,
    n598
  );


  buf
  g660
  (
    n726,
    n512
  );


  not
  g661
  (
    n626,
    n432
  );


  buf
  g662
  (
    n636,
    n508
  );


  buf
  g663
  (
    n741,
    n498
  );


  buf
  g664
  (
    n769,
    n612
  );


  buf
  g665
  (
    n799,
    n438
  );


  buf
  g666
  (
    n647,
    n593
  );


  not
  g667
  (
    n744,
    n513
  );


  buf
  g668
  (
    n724,
    n546
  );


  buf
  g669
  (
    n665,
    n552
  );


  buf
  g670
  (
    n776,
    n514
  );


  buf
  g671
  (
    n701,
    n469
  );


  not
  g672
  (
    n748,
    n549
  );


  buf
  g673
  (
    n770,
    n610
  );


  not
  g674
  (
    n674,
    n501
  );


  not
  g675
  (
    n740,
    n561
  );


  not
  g676
  (
    n775,
    n603
  );


  not
  g677
  (
    n790,
    n585
  );


  not
  g678
  (
    n742,
    n580
  );


  buf
  g679
  (
    n663,
    n538
  );


  buf
  g680
  (
    n660,
    n445
  );


  not
  g681
  (
    n627,
    n461
  );


  buf
  g682
  (
    n746,
    n511
  );


  buf
  g683
  (
    n717,
    n579
  );


  not
  g684
  (
    n749,
    n560
  );


  not
  g685
  (
    n756,
    n496
  );


  buf
  g686
  (
    n687,
    n547
  );


  buf
  g687
  (
    n657,
    n479
  );


  buf
  g688
  (
    n673,
    n453
  );


  not
  g689
  (
    n758,
    n577
  );


  buf
  g690
  (
    n778,
    n518
  );


  not
  g691
  (
    KeyWire_0_10,
    n481
  );


  not
  g692
  (
    n734,
    n440
  );


  not
  g693
  (
    n679,
    n465
  );


  buf
  g694
  (
    n737,
    n502
  );


  not
  g695
  (
    n655,
    n617
  );


  not
  g696
  (
    n639,
    n565
  );


  buf
  g697
  (
    n686,
    n477
  );


  not
  g698
  (
    n654,
    n608
  );


  not
  g699
  (
    n683,
    n486
  );


  buf
  g700
  (
    n682,
    n551
  );


  buf
  g701
  (
    n788,
    n540
  );


  not
  g702
  (
    n644,
    n476
  );


  buf
  g703
  (
    n735,
    n535
  );


  buf
  g704
  (
    n642,
    n605
  );


  buf
  g705
  (
    n750,
    n475
  );


  buf
  g706
  (
    n768,
    n505
  );


  buf
  g707
  (
    n784,
    n429
  );


  not
  g708
  (
    n723,
    n493
  );


  buf
  g709
  (
    n711,
    n539
  );


  buf
  g710
  (
    n696,
    n545
  );


  not
  g711
  (
    n712,
    n499
  );


  not
  g712
  (
    n680,
    n441
  );


  buf
  g713
  (
    n685,
    n573
  );


  buf
  g714
  (
    n793,
    n587
  );


  not
  g715
  (
    n641,
    n589
  );


  not
  g716
  (
    n787,
    n452
  );


  not
  g717
  (
    n650,
    n420
  );


  not
  g718
  (
    n668,
    n431
  );


  buf
  g719
  (
    n772,
    n447
  );


  buf
  g720
  (
    n667,
    n544
  );


  buf
  g721
  (
    n633,
    n443
  );


  not
  g722
  (
    n728,
    n474
  );


  not
  g723
  (
    n736,
    n488
  );


  not
  g724
  (
    n766,
    n428
  );


  buf
  g725
  (
    n752,
    n525
  );


  buf
  g726
  (
    n753,
    n436
  );


  not
  g727
  (
    n678,
    n567
  );


  not
  g728
  (
    KeyWire_0_28,
    n434
  );


  not
  g729
  (
    n670,
    n507
  );


  not
  g730
  (
    n635,
    n557
  );


  buf
  g731
  (
    n629,
    n572
  );


  buf
  g732
  (
    n715,
    n532
  );


  buf
  g733
  (
    n710,
    n424
  );


  not
  g734
  (
    n648,
    n489
  );


  buf
  g735
  (
    n681,
    n559
  );


  buf
  g736
  (
    n738,
    n520
  );


  buf
  g737
  (
    n722,
    n460
  );


  buf
  g738
  (
    n779,
    n568
  );


  not
  g739
  (
    n714,
    n575
  );


  not
  g740
  (
    n651,
    n542
  );


  not
  g741
  (
    n785,
    n597
  );


  buf
  g742
  (
    n652,
    n537
  );


  buf
  g743
  (
    n625,
    n459
  );


  buf
  g744
  (
    n782,
    n521
  );


  buf
  g745
  (
    n669,
    n527
  );


  not
  g746
  (
    n762,
    n427
  );


  buf
  g747
  (
    n628,
    n574
  );


  buf
  g748
  (
    n713,
    n449
  );


  buf
  g749
  (
    n638,
    n554
  );


  buf
  g750
  (
    n675,
    n491
  );


  buf
  g751
  (
    n789,
    n600
  );


  buf
  g752
  (
    n631,
    n446
  );


  buf
  g753
  (
    n725,
    n609
  );


  not
  g754
  (
    n677,
    n586
  );


  buf
  g755
  (
    n645,
    n534
  );


  not
  g756
  (
    n745,
    n564
  );


  buf
  g757
  (
    n664,
    n548
  );


  buf
  g758
  (
    n796,
    n570
  );


  not
  g759
  (
    n755,
    n536
  );


  not
  g760
  (
    n630,
    n578
  );


  buf
  g761
  (
    n732,
    n562
  );


  not
  g762
  (
    n760,
    n444
  );


  buf
  g763
  (
    KeyWire_0_0,
    n581
  );


  not
  g764
  (
    n653,
    n550
  );


  not
  g765
  (
    n672,
    n599
  );


  or
  g766
  (
    n780,
    n582,
    n467
  );


  nand
  g767
  (
    n694,
    n583,
    n558,
    n591,
    n607
  );


  nand
  g768
  (
    n671,
    n618,
    n613,
    n464,
    n435
  );


  and
  g769
  (
    n718,
    n485,
    n555,
    n616,
    n468
  );


  nand
  g770
  (
    n643,
    n524,
    n594,
    n522,
    n462
  );


  nand
  g771
  (
    n791,
    n569,
    n463,
    n553,
    n471
  );


  nor
  g772
  (
    n697,
    n602,
    n563,
    n495,
    n437
  );


  xnor
  g773
  (
    n624,
    n480,
    n457,
    n470,
    n450
  );


  or
  g774
  (
    n965,
    n628,
    n752,
    n680,
    n677
  );


  or
  g775
  (
    n899,
    n655,
    n737,
    n675,
    n744
  );


  nand
  g776
  (
    n900,
    n681,
    n769,
    n678,
    n659
  );


  xor
  g777
  (
    n809,
    n705,
    n744,
    n694,
    n714
  );


  and
  g778
  (
    n847,
    n631,
    n713,
    n705,
    n731
  );


  and
  g779
  (
    n910,
    n703,
    n728,
    n738,
    n671
  );


  nor
  g780
  (
    n914,
    n773,
    n710,
    n792,
    n704
  );


  or
  g781
  (
    n868,
    n784,
    n729,
    n777,
    n691
  );


  or
  g782
  (
    n969,
    n649,
    n643,
    n627,
    n745
  );


  or
  g783
  (
    n820,
    n641,
    n642,
    n678,
    n625
  );


  xor
  g784
  (
    n951,
    n640,
    n672,
    n663,
    n756
  );


  nand
  g785
  (
    KeyWire_0_23,
    n747,
    n657,
    n646,
    n641
  );


  and
  g786
  (
    n913,
    n654,
    n786,
    n690,
    n723
  );


  nor
  g787
  (
    n814,
    n759,
    n683,
    n788,
    n709
  );


  nand
  g788
  (
    n954,
    n789,
    n651,
    n763,
    n701
  );


  xor
  g789
  (
    n828,
    n672,
    n688,
    n742,
    n698
  );


  nor
  g790
  (
    n879,
    n626,
    n670,
    n777,
    n754
  );


  and
  g791
  (
    n829,
    n732,
    n700,
    n703,
    n733
  );


  and
  g792
  (
    n906,
    n629,
    n757,
    n736,
    n624
  );


  or
  g793
  (
    n819,
    n658,
    n642,
    n627,
    n759
  );


  nor
  g794
  (
    n804,
    n683,
    n650,
    n627,
    n758
  );


  xnor
  g795
  (
    n855,
    n775,
    n728,
    n749,
    n647
  );


  xor
  g796
  (
    n810,
    n769,
    n699,
    n739,
    n675
  );


  nor
  g797
  (
    n834,
    n749,
    n749,
    n767,
    n653
  );


  xor
  g798
  (
    n926,
    n732,
    n755,
    n719,
    n757
  );


  nand
  g799
  (
    n864,
    n752,
    n725,
    n751,
    n687
  );


  nor
  g800
  (
    n953,
    n643,
    n730,
    n725,
    n708
  );


  and
  g801
  (
    n904,
    n756,
    n790,
    n724,
    n658
  );


  nand
  g802
  (
    n805,
    n651,
    n780,
    n770,
    n741
  );


  xor
  g803
  (
    n883,
    n677,
    n784,
    n662,
    n716
  );


  nor
  g804
  (
    n872,
    n699,
    n662,
    n642,
    n717
  );


  xnor
  g805
  (
    n958,
    n721,
    n758,
    n785,
    n779
  );


  nand
  g806
  (
    n932,
    n639,
    n790,
    n748,
    n698
  );


  nand
  g807
  (
    n806,
    n676,
    n775,
    n733,
    n673
  );


  xor
  g808
  (
    n860,
    n762,
    n774,
    n734,
    n765
  );


  nand
  g809
  (
    n970,
    n708,
    n738,
    n739,
    n636
  );


  nand
  g810
  (
    n947,
    n771,
    n763,
    n791,
    n754
  );


  xnor
  g811
  (
    n896,
    n734,
    n742,
    n652,
    n705
  );


  xnor
  g812
  (
    n858,
    n686,
    n669,
    n765,
    n764
  );


  xor
  g813
  (
    n939,
    n732,
    n695,
    n785,
    n652
  );


  and
  g814
  (
    n842,
    n725,
    n682,
    n761,
    n712
  );


  xnor
  g815
  (
    n917,
    n685,
    n739,
    n667,
    n716
  );


  xor
  g816
  (
    n826,
    n661,
    n646,
    n730,
    n776
  );


  or
  g817
  (
    n833,
    n779,
    n791,
    n696,
    n692
  );


  and
  g818
  (
    n801,
    n773,
    n711,
    n674,
    n696
  );


  nand
  g819
  (
    n830,
    n676,
    n793,
    n694,
    n691
  );


  xnor
  g820
  (
    n807,
    n668,
    n778,
    n709,
    n670
  );


  xor
  g821
  (
    n895,
    n660,
    n631,
    n774,
    n747
  );


  xor
  g822
  (
    n835,
    n781,
    n789,
    n795,
    n635
  );


  nand
  g823
  (
    n870,
    n770,
    n722,
    n772,
    n710
  );


  or
  g824
  (
    n822,
    n740,
    n638,
    n751,
    n720
  );


  nor
  g825
  (
    n946,
    n648,
    n703,
    n629,
    n765
  );


  or
  g826
  (
    n878,
    n628,
    n726,
    n660,
    n734
  );


  xor
  g827
  (
    n941,
    n779,
    n659,
    n654,
    n755
  );


  xor
  g828
  (
    n825,
    n632,
    n660,
    n727,
    n647
  );


  xnor
  g829
  (
    KeyWire_0_13,
    n689,
    n704,
    n724,
    n766
  );


  nand
  g830
  (
    n902,
    n757,
    n620,
    n698,
    n771
  );


  nor
  g831
  (
    n854,
    n632,
    n736,
    n759,
    n645
  );


  nor
  g832
  (
    n943,
    n644,
    n747,
    n656,
    n743
  );


  or
  g833
  (
    n903,
    n625,
    n683,
    n632,
    n743
  );


  xor
  g834
  (
    n890,
    n771,
    n691,
    n717,
    n732
  );


  or
  g835
  (
    n874,
    n703,
    n766,
    n633,
    n783
  );


  or
  g836
  (
    n856,
    n723,
    n786,
    n738,
    n648
  );


  nand
  g837
  (
    n861,
    n766,
    n758,
    n656,
    n772
  );


  or
  g838
  (
    n885,
    n692,
    n788,
    n721,
    n727
  );


  xor
  g839
  (
    n869,
    n650,
    n740,
    n701,
    n785
  );


  nand
  g840
  (
    n840,
    n715,
    n652,
    n707,
    n653
  );


  or
  g841
  (
    n891,
    n783,
    n664,
    n712,
    n654
  );


  nand
  g842
  (
    n931,
    n667,
    n630,
    n752,
    n625
  );


  and
  g843
  (
    n876,
    n643,
    n634,
    n644
  );


  nand
  g844
  (
    n887,
    n775,
    n693,
    n771,
    n637
  );


  nand
  g845
  (
    n905,
    n746,
    n733,
    n680,
    n663
  );


  and
  g846
  (
    n909,
    n702,
    n695,
    n698,
    n789
  );


  or
  g847
  (
    n884,
    n684,
    n764,
    n658,
    n782
  );


  xnor
  g848
  (
    n873,
    n646,
    n750,
    n645,
    n776
  );


  nand
  g849
  (
    n892,
    n629,
    n630,
    n697,
    n666
  );


  xor
  g850
  (
    n908,
    n750,
    n696,
    n787,
    n645
  );


  and
  g851
  (
    n960,
    n688,
    n671,
    n638,
    n637
  );


  nand
  g852
  (
    n928,
    n671,
    n708,
    n626,
    n686
  );


  and
  g853
  (
    n837,
    n690,
    n717,
    n760,
    n790
  );


  xnor
  g854
  (
    n816,
    n648,
    n768,
    n744,
    n740
  );


  xnor
  g855
  (
    n881,
    n633,
    n649,
    n674,
    n713
  );


  and
  g856
  (
    n924,
    n640,
    n639,
    n661,
    n761
  );


  or
  g857
  (
    n929,
    n742,
    n746,
    n726,
    n668
  );


  xor
  g858
  (
    n849,
    n678,
    n633,
    n685,
    n787
  );


  xor
  g859
  (
    n934,
    n769,
    n721,
    n739
  );


  xnor
  g860
  (
    n952,
    n761,
    n772,
    n794,
    n746
  );


  nand
  g861
  (
    n919,
    n679,
    n692,
    n741,
    n772
  );


  xor
  g862
  (
    n967,
    n737,
    n729,
    n664,
    n643
  );


  or
  g863
  (
    n831,
    n662,
    n750,
    n684,
    n753
  );


  and
  g864
  (
    n894,
    n778,
    n657,
    n716,
    n755
  );


  xor
  g865
  (
    n927,
    n719,
    n729,
    n743,
    n696
  );


  nand
  g866
  (
    n907,
    n659,
    n781,
    n651,
    n767
  );


  and
  g867
  (
    n957,
    n641,
    n786,
    n636,
    n701
  );


  nor
  g868
  (
    n959,
    n761,
    n738,
    n791,
    n760
  );


  and
  g869
  (
    n824,
    n634,
    n668,
    n651,
    n718
  );


  or
  g870
  (
    n803,
    n680,
    n709,
    n692,
    n712
  );


  or
  g871
  (
    n838,
    n688,
    n722,
    n650,
    n760
  );


  and
  g872
  (
    n916,
    n655,
    n713,
    n788,
    n682
  );


  nor
  g873
  (
    n938,
    n684,
    n789,
    n723,
    n666
  );


  nand
  g874
  (
    n933,
    n675,
    n768,
    n707,
    n624
  );


  or
  g875
  (
    n920,
    n690,
    n654,
    n763,
    n748
  );


  and
  g876
  (
    n821,
    n619,
    n635,
    n706,
    n727
  );


  and
  g877
  (
    n877,
    n762,
    n730,
    n628,
    n648
  );


  nor
  g878
  (
    n882,
    n619,
    n730,
    n741,
    n649
  );


  xnor
  g879
  (
    n937,
    n774,
    n724,
    n718,
    n791
  );


  or
  g880
  (
    n968,
    n624,
    n631,
    n672,
    n702
  );


  xor
  g881
  (
    n918,
    n733,
    n687,
    n745,
    n787
  );


  xor
  g882
  (
    n966,
    n725,
    n670,
    n674,
    n719
  );


  nand
  g883
  (
    n961,
    n763,
    n704,
    n783,
    n735
  );


  xnor
  g884
  (
    n922,
    n637,
    n635,
    n784,
    n627
  );


  or
  g885
  (
    n930,
    n677,
    n628,
    n759,
    n686
  );


  or
  g886
  (
    n962,
    n655,
    n645,
    n764,
    n737
  );


  nand
  g887
  (
    n808,
    n782,
    n778,
    n716,
    n672
  );


  xor
  g888
  (
    n846,
    n762,
    n664,
    n767,
    n713
  );


  or
  g889
  (
    n898,
    n709,
    n793,
    n768,
    n710
  );


  xor
  g890
  (
    KeyWire_0_30,
    n686,
    n676,
    n770,
    n681
  );


  or
  g891
  (
    n911,
    n669,
    n720,
    n636,
    n694
  );


  nor
  g892
  (
    n818,
    n794,
    n647,
    n650,
    n677
  );


  xor
  g893
  (
    n923,
    n773,
    n776,
    n634,
    n704
  );


  nor
  g894
  (
    n871,
    n750,
    n736,
    n777,
    n752
  );


  xnor
  g895
  (
    n850,
    n694,
    n679,
    n661,
    n722
  );


  and
  g896
  (
    n880,
    n794,
    n719,
    n637,
    n640
  );


  or
  g897
  (
    n921,
    n665,
    n681,
    n724,
    n707
  );


  nand
  g898
  (
    n851,
    n728,
    n667,
    n758,
    n711
  );


  xnor
  g899
  (
    n811,
    n699,
    n775,
    n734,
    n679
  );


  xnor
  g900
  (
    n945,
    n737,
    n700,
    n680,
    n714
  );


  xor
  g901
  (
    n815,
    n673,
    n711,
    n665,
    n668
  );


  xor
  g902
  (
    n844,
    n699,
    n715,
    n678,
    n770
  );


  xnor
  g903
  (
    n949,
    n718,
    n787,
    n736,
    n726
  );


  xor
  g904
  (
    n863,
    n691,
    n685,
    n706,
    n700
  );


  xor
  g905
  (
    n836,
    n639,
    n640,
    n792,
    n708
  );


  xnor
  g906
  (
    n956,
    n782,
    n697,
    n717,
    n769
  );


  nand
  g907
  (
    n823,
    n655,
    n741,
    n777,
    n652
  );


  and
  g908
  (
    n875,
    n665,
    n753,
    n731,
    n774
  );


  nor
  g909
  (
    n817,
    n629,
    n638,
    n751,
    n641
  );


  nor
  g910
  (
    n853,
    n673,
    n679,
    n712,
    n706
  );


  xor
  g911
  (
    n893,
    n682,
    n667,
    n702,
    n690
  );


  nand
  g912
  (
    n859,
    n665,
    n659,
    n657,
    n673
  );


  nand
  g913
  (
    n827,
    n745,
    n657,
    n674,
    n735
  );


  nor
  g914
  (
    n942,
    n780,
    n745,
    n671,
    n751
  );


  and
  g915
  (
    n901,
    n765,
    n676,
    n785,
    n747
  );


  and
  g916
  (
    n888,
    n754,
    n779,
    n731,
    n664
  );


  nor
  g917
  (
    n886,
    n710,
    n748,
    n780,
    n653
  );


  and
  g918
  (
    n862,
    n723,
    n669,
    n756,
    n660
  );


  xor
  g919
  (
    n812,
    n661,
    n735,
    n695,
    n663
  );


  nor
  g920
  (
    n915,
    n626,
    n633,
    n666,
    n682
  );


  xnor
  g921
  (
    KeyWire_0_31,
    n702,
    n687,
    n635,
    n689
  );


  and
  g922
  (
    n936,
    n764,
    n762,
    n647,
    n722
  );


  or
  g923
  (
    n841,
    n644,
    n663,
    n743,
    n705
  );


  and
  g924
  (
    n800,
    n776,
    n631,
    n624,
    n697
  );


  xnor
  g925
  (
    n925,
    n634,
    n656,
    n684,
    n630
  );


  nor
  g926
  (
    n971,
    n649,
    n669,
    n753,
    n793
  );


  or
  g927
  (
    n865,
    n766,
    n720,
    n781,
    n783
  );


  xor
  g928
  (
    n963,
    n768,
    n742,
    n683,
    n715
  );


  nand
  g929
  (
    n843,
    n639,
    n706,
    n662,
    n792
  );


  and
  g930
  (
    n802,
    n697,
    n715,
    n784,
    n693
  );


  xor
  g931
  (
    n940,
    n731,
    n658,
    n670,
    n760
  );


  or
  g932
  (
    n889,
    n632,
    n689,
    n707,
    n675
  );


  xor
  g933
  (
    n935,
    n748,
    n792,
    n718,
    n656
  );


  and
  g934
  (
    n948,
    n689,
    n778,
    n638,
    n642
  );


  nand
  g935
  (
    n857,
    n685,
    n795,
    n695
  );


  or
  g936
  (
    n972,
    n754,
    n773,
    n749,
    n720
  );


  nor
  g937
  (
    n912,
    n729,
    n740,
    n728,
    n794
  );


  xnor
  g938
  (
    n832,
    n781,
    n653,
    n714,
    n746
  );


  and
  g939
  (
    n813,
    n701,
    n711,
    n693,
    n625
  );


  xnor
  g940
  (
    n867,
    n767,
    n636,
    n700,
    n630
  );


  nand
  g941
  (
    n950,
    n790,
    n646,
    n693,
    n788
  );


  xor
  g942
  (
    KeyWire_0_14,
    n626,
    n681,
    n753,
    n755
  );


  nand
  g943
  (
    n848,
    n793,
    n786,
    n796,
    n757
  );


  or
  g944
  (
    n866,
    n687,
    n795,
    n780,
    n744
  );


  and
  g945
  (
    n845,
    n714,
    n735,
    n726,
    n727
  );


  nor
  g946
  (
    n964,
    n666,
    n782,
    n688,
    n756
  );


  xor
  g947
  (
    n995,
    n813,
    n825,
    n824,
    n829
  );


  nor
  g948
  (
    n986,
    n871,
    n802,
    n867,
    n883
  );


  nand
  g949
  (
    n983,
    n872,
    n820,
    n830,
    n854
  );


  nand
  g950
  (
    n988,
    n827,
    n819,
    n814,
    n821
  );


  and
  g951
  (
    n973,
    n891,
    n897,
    n880,
    n902
  );


  nand
  g952
  (
    n980,
    n808,
    n889,
    n855,
    n899
  );


  xor
  g953
  (
    n976,
    n905,
    n847,
    n870,
    n822
  );


  xnor
  g954
  (
    n987,
    n809,
    n841,
    n896,
    n810
  );


  xnor
  g955
  (
    n978,
    n906,
    n888,
    n823,
    n816
  );


  nor
  g956
  (
    n979,
    n904,
    n832,
    n877,
    n853
  );


  and
  g957
  (
    n998,
    n859,
    n845,
    n878,
    n887
  );


  xor
  g958
  (
    n989,
    n834,
    n831,
    n884,
    n826
  );


  nor
  g959
  (
    n991,
    n869,
    n876,
    n811,
    n839
  );


  nand
  g960
  (
    n992,
    n858,
    n907,
    n806,
    n894
  );


  nor
  g961
  (
    n974,
    n836,
    n833,
    n842,
    n849
  );


  xnor
  g962
  (
    KeyWire_0_8,
    n850,
    n801,
    n893,
    n840
  );


  nor
  g963
  (
    n994,
    n803,
    n885,
    n837,
    n866
  );


  xor
  g964
  (
    n984,
    n851,
    n807,
    n838,
    n868
  );


  and
  g965
  (
    n999,
    n852,
    n835,
    n861,
    n879
  );


  nand
  g966
  (
    n996,
    n864,
    n882,
    n860,
    n875
  );


  and
  g967
  (
    n997,
    n898,
    n844,
    n800,
    n901
  );


  or
  g968
  (
    n981,
    n903,
    n857,
    n862,
    n874
  );


  nand
  g969
  (
    n975,
    n873,
    n856,
    n843,
    n848
  );


  and
  g970
  (
    n977,
    n863,
    n846,
    n818,
    n804
  );


  nor
  g971
  (
    n985,
    n886,
    n828,
    n900,
    n805
  );


  nor
  g972
  (
    n993,
    n812,
    n881,
    n865,
    n815
  );


  xnor
  g973
  (
    n982,
    n890,
    n892,
    n817,
    n895
  );


  xnor
  g974
  (
    n1002,
    n919,
    n921,
    n977,
    n920
  );


  xnor
  g975
  (
    n1003,
    n914,
    n918,
    n911,
    n912
  );


  nand
  g976
  (
    n1004,
    n908,
    n976,
    n915,
    n975
  );


  and
  g977
  (
    n1001,
    n909,
    n917,
    n913,
    n916
  );


  nand
  g978
  (
    n1000,
    n910,
    n974,
    n973,
    n922
  );


  buf
  g979
  (
    n1010,
    n1004
  );


  not
  g980
  (
    n1013,
    n1004
  );


  buf
  g981
  (
    n1011,
    n1002
  );


  not
  g982
  (
    n1008,
    n1003
  );


  buf
  g983
  (
    n1006,
    n1001
  );


  buf
  g984
  (
    n1007,
    n923
  );


  not
  g985
  (
    n1012,
    n1003
  );


  not
  g986
  (
    n1009,
    n1000
  );


  buf
  g987
  (
    n1005,
    n1004
  );


  xor
  g988
  (
    n1018,
    n622,
    n622,
    n1012,
    n927
  );


  xor
  g989
  (
    n1017,
    n930,
    n925,
    n621
  );


  and
  g990
  (
    n1015,
    n620,
    n928,
    n929,
    n1008
  );


  or
  g991
  (
    n1021,
    n421,
    n1013,
    n924
  );


  or
  g992
  (
    n1019,
    n1010,
    n621,
    n1013
  );


  xnor
  g993
  (
    n1014,
    n931,
    n621,
    n1005,
    n932
  );


  xor
  g994
  (
    n1020,
    n620,
    n622,
    n926,
    n1006
  );


  nand
  g995
  (
    n1016,
    n1011,
    n1009,
    n620,
    n1007
  );


  xnor
  g996
  (
    n1022,
    n1019,
    n933,
    n1021,
    n1020
  );


  or
  g997
  (
    n1023,
    n939,
    n935,
    n938,
    n1022
  );


  and
  g998
  (
    n1024,
    n934,
    n1022,
    n937,
    n936
  );


  not
  g999
  (
    n1028,
    n1023
  );


  not
  g1000
  (
    n1030,
    n1024
  );


  xor
  g1001
  (
    n1029,
    n942,
    n941
  );


  or
  g1002
  (
    n1026,
    n943,
    n947,
    n1023
  );


  nand
  g1003
  (
    n1025,
    n1023,
    n1024
  );


  and
  g1004
  (
    n1031,
    n946,
    n945,
    n940
  );


  xnor
  g1005
  (
    n1027,
    n1023,
    n948,
    n944
  );


  and
  g1006
  (
    n1040,
    n123,
    n623,
    n1027,
    n1029
  );


  xnor
  g1007
  (
    n1052,
    n799,
    n950,
    n987,
    n997
  );


  xnor
  g1008
  (
    n1033,
    n1031,
    n797,
    n798,
    n1025
  );


  xor
  g1009
  (
    n1042,
    n121,
    n122,
    n1024,
    n996
  );


  xor
  g1010
  (
    n1047,
    n951,
    n796,
    n980,
    n1026
  );


  or
  g1011
  (
    n1044,
    n993,
    n1031,
    n1030,
    n798
  );


  or
  g1012
  (
    n1043,
    n1027,
    n623,
    n421
  );


  nor
  g1013
  (
    n1053,
    n122,
    n622,
    n796,
    n1031
  );


  and
  g1014
  (
    n1054,
    n1028,
    n421,
    n123,
    n1027
  );


  and
  g1015
  (
    n1035,
    n998,
    n1029,
    n1031,
    n991
  );


  or
  g1016
  (
    n1049,
    n960,
    n797,
    n956,
    n949
  );


  nor
  g1017
  (
    n1036,
    n1026,
    n988,
    n961,
    n986
  );


  nand
  g1018
  (
    n1032,
    n999,
    n1030,
    n982,
    n1028
  );


  nor
  g1019
  (
    n1050,
    n1026,
    n797,
    n981,
    n992
  );


  nand
  g1020
  (
    n1046,
    n798,
    n122,
    n958,
    n957
  );


  and
  g1021
  (
    n1037,
    n421,
    n798,
    n796,
    n979
  );


  nand
  g1022
  (
    n1034,
    n984,
    n122,
    n1030,
    n994
  );


  nand
  g1023
  (
    n1045,
    n1029,
    n623,
    n1028,
    n797
  );


  xor
  g1024
  (
    n1048,
    n978,
    n1026,
    n983,
    n959
  );


  nor
  g1025
  (
    n1039,
    n1030,
    n121,
    n1025,
    n954
  );


  nand
  g1026
  (
    n1051,
    n953,
    n955,
    n952,
    n123
  );


  nor
  g1027
  (
    n1041,
    n985,
    n989,
    n1027,
    n990
  );


  nand
  g1028
  (
    n1038,
    n1029,
    n1028,
    n123,
    n995
  );


  not
  g1029
  (
    n1055,
    n1048
  );


  or
  g1030
  (
    n1056,
    n1049,
    n1050,
    n1047
  );


  xor
  g1031
  (
    n1057,
    n422,
    n422,
    n1055,
    n1052
  );


  nor
  g1032
  (
    n1058,
    n962,
    n963,
    n1056
  );


  nand
  g1033
  (
    n1061,
    n1053,
    n965,
    n422
  );


  or
  g1034
  (
    n1059,
    n1051,
    n423,
    n966
  );


  or
  g1035
  (
    n1060,
    n964,
    n1056,
    n1054
  );


  nand
  g1036
  (
    n1065,
    n1060,
    n1057
  );


  or
  g1037
  (
    n1063,
    n1059,
    n124,
    n125
  );


  nor
  g1038
  (
    n1062,
    n124,
    n125,
    n967,
    n1058
  );


  or
  g1039
  (
    n1064,
    n125,
    n125,
    n124,
    n1061
  );


  nor
  g1040
  (
    n1066,
    n1064,
    n1065,
    n423
  );


  and
  g1041
  (
    n1067,
    n1062,
    n423,
    n1063
  );


  xnor
  g1042
  (
    n1068,
    n1066,
    n968,
    n969,
    n970
  );


  nand
  g1043
  (
    n1070,
    n1068,
    n799
  );


  and
  g1044
  (
    n1069,
    n1067,
    n1068,
    n799
  );


  nand
  g1045
  (
    n1071,
    n972,
    n1070,
    n971,
    n1069
  );


  xor
  KeyGate_0_0
  (
    n699,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n345,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n121,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n797,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n327,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n502,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n151,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n314,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n990,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n386,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n763,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n583,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n475,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n852,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n897,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n695,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n274,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n217,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n579,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n552,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n383,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n407,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n590,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n839,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n566,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n179,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n754,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n530,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n721,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n375,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n944,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n955,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

