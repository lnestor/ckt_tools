

module Stat_147_624
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n141,
  n149,
  n157,
  n162,
  n160,
  n165,
  n154,
  n151,
  n163,
  n158,
  n164,
  n150,
  n156,
  n161,
  n152,
  n153,
  n159,
  n155,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;
  output n141;output n149;output n157;output n162;output n160;output n165;output n154;output n151;output n163;output n158;output n164;output n150;output n156;output n161;output n152;output n153;output n159;output n155;
  wire n19;wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n51,
    n2
  );


  buf
  g1
  (
    n44,
    n6
  );


  not
  g2
  (
    n59,
    n10
  );


  not
  g3
  (
    n46,
    n12
  );


  buf
  g4
  (
    n38,
    n1
  );


  not
  g5
  (
    n39,
    n9
  );


  buf
  g6
  (
    n32,
    n10
  );


  buf
  g7
  (
    n58,
    n9
  );


  not
  g8
  (
    n55,
    n7
  );


  not
  g9
  (
    n31,
    n5
  );


  not
  g10
  (
    n35,
    n8
  );


  buf
  g11
  (
    n63,
    n8
  );


  buf
  g12
  (
    n20,
    n11
  );


  buf
  g13
  (
    n52,
    n6
  );


  not
  g14
  (
    n56,
    n11
  );


  not
  g15
  (
    n24,
    n7
  );


  not
  g16
  (
    n50,
    n2
  );


  not
  g17
  (
    n21,
    n12
  );


  buf
  g18
  (
    n53,
    n3
  );


  not
  g19
  (
    n49,
    n4
  );


  not
  g20
  (
    n26,
    n5
  );


  buf
  g21
  (
    n47,
    n5
  );


  not
  g22
  (
    n28,
    n3
  );


  buf
  g23
  (
    n43,
    n10
  );


  buf
  g24
  (
    n64,
    n2
  );


  buf
  g25
  (
    n19,
    n7
  );


  buf
  g26
  (
    n34,
    n1
  );


  not
  g27
  (
    n57,
    n5
  );


  not
  g28
  (
    n62,
    n3
  );


  buf
  g29
  (
    n29,
    n1
  );


  not
  g30
  (
    n30,
    n2
  );


  not
  g31
  (
    n33,
    n10
  );


  buf
  g32
  (
    n22,
    n4
  );


  not
  g33
  (
    n23,
    n8
  );


  not
  g34
  (
    n40,
    n4
  );


  not
  g35
  (
    n37,
    n6
  );


  buf
  g36
  (
    n25,
    n9
  );


  buf
  g37
  (
    n60,
    n9
  );


  not
  g38
  (
    n45,
    n6
  );


  not
  g39
  (
    n27,
    n3
  );


  buf
  g40
  (
    n54,
    n11
  );


  not
  g41
  (
    n48,
    n1
  );


  not
  g42
  (
    n41,
    n8
  );


  not
  g43
  (
    n42,
    n11
  );


  not
  g44
  (
    n36,
    n4
  );


  buf
  g45
  (
    n61,
    n7
  );


  xor
  g46
  (
    n65,
    n19,
    n20
  );


  xnor
  g47
  (
    n66,
    n20,
    n19
  );


  buf
  g48
  (
    n68,
    n66
  );


  buf
  g49
  (
    n69,
    n66
  );


  not
  g50
  (
    n67,
    n66
  );


  not
  g51
  (
    n70,
    n66
  );


  or
  g52
  (
    n83,
    n13,
    n17
  );


  xnor
  g53
  (
    n77,
    n15,
    n67
  );


  xor
  g54
  (
    n84,
    n69,
    n15
  );


  xor
  g55
  (
    n78,
    n70,
    n68
  );


  nand
  g56
  (
    n82,
    n70,
    n67
  );


  xnor
  g57
  (
    n71,
    n12,
    n17
  );


  buf
  g58
  (
    n73,
    n18
  );


  not
  g59
  (
    n85,
    n70
  );


  xor
  g60
  (
    n74,
    n14,
    n69
  );


  xnor
  g61
  (
    n81,
    n16,
    n14
  );


  buf
  g62
  (
    n76,
    n16
  );


  nor
  g63
  (
    n72,
    n68,
    n13,
    n67
  );


  and
  g64
  (
    n75,
    n16,
    n15,
    n69,
    n12
  );


  or
  g65
  (
    n80,
    n68,
    n17,
    n69
  );


  xor
  g66
  (
    n86,
    n18,
    n67,
    n68,
    n14
  );


  nor
  g67
  (
    n79,
    n14,
    n13,
    n18,
    n15
  );


  nand
  g68
  (
    n147,
    n62,
    n22,
    n82
  );


  xnor
  g69
  (
    n109,
    n29,
    n76,
    n75
  );


  nand
  g70
  (
    n148,
    n21,
    n28,
    n55
  );


  and
  g71
  (
    n125,
    n86,
    n30,
    n36
  );


  xor
  g72
  (
    n126,
    n42,
    n72,
    n27
  );


  and
  g73
  (
    n138,
    n42,
    n74,
    n40
  );


  and
  g74
  (
    n95,
    n58,
    n86,
    n33
  );


  and
  g75
  (
    n117,
    n22,
    n45,
    n30
  );


  nand
  g76
  (
    n141,
    n43,
    n76,
    n55,
    n72
  );


  and
  g77
  (
    n142,
    n60,
    n77,
    n27,
    n85
  );


  and
  g78
  (
    n100,
    n51,
    n86,
    n24,
    n71
  );


  xor
  g79
  (
    n89,
    n82,
    n32,
    n37,
    n57
  );


  and
  g80
  (
    n130,
    n51,
    n43,
    n40,
    n78
  );


  nor
  g81
  (
    n110,
    n42,
    n46,
    n78,
    n44
  );


  xor
  g82
  (
    n116,
    n40,
    n79,
    n53,
    n64
  );


  or
  g83
  (
    n122,
    n82,
    n42,
    n83,
    n64
  );


  xnor
  g84
  (
    n129,
    n27,
    n39,
    n76,
    n37
  );


  xnor
  g85
  (
    n137,
    n35,
    n61,
    n62,
    n32
  );


  and
  g86
  (
    n96,
    n34,
    n82,
    n25,
    n23
  );


  and
  g87
  (
    n90,
    n72,
    n73,
    n21,
    n58
  );


  nor
  g88
  (
    n91,
    n59,
    n21,
    n52,
    n74
  );


  nand
  g89
  (
    n88,
    n23,
    n60,
    n74,
    n56
  );


  or
  g90
  (
    n120,
    n77,
    n33,
    n47,
    n61
  );


  xor
  g91
  (
    n102,
    n79,
    n35,
    n45,
    n22
  );


  xor
  g92
  (
    n139,
    n58,
    n56,
    n71,
    n85
  );


  nor
  g93
  (
    n121,
    n38,
    n43,
    n75,
    n31
  );


  or
  g94
  (
    n105,
    n60,
    n25,
    n52,
    n40
  );


  xnor
  g95
  (
    n104,
    n36,
    n44,
    n51,
    n85
  );


  nand
  g96
  (
    n144,
    n80,
    n52,
    n32,
    n61
  );


  and
  g97
  (
    n101,
    n46,
    n83,
    n61,
    n76
  );


  xor
  g98
  (
    n113,
    n28,
    n80,
    n72,
    n71
  );


  nor
  g99
  (
    n115,
    n33,
    n74,
    n77,
    n50
  );


  xor
  g100
  (
    n143,
    n63,
    n83,
    n28
  );


  or
  g101
  (
    n106,
    n84,
    n36,
    n75,
    n30
  );


  xor
  g102
  (
    n112,
    n73,
    n53,
    n41,
    n80
  );


  nor
  g103
  (
    n107,
    n37,
    n59,
    n47,
    n45
  );


  and
  g104
  (
    n99,
    n54,
    n85,
    n34,
    n59
  );


  or
  g105
  (
    n140,
    n62,
    n59,
    n26,
    n57
  );


  or
  g106
  (
    n93,
    n48,
    n39,
    n23,
    n45
  );


  nor
  g107
  (
    n123,
    n47,
    n24,
    n64,
    n39
  );


  nand
  g108
  (
    n134,
    n63,
    n33,
    n56,
    n47
  );


  xor
  g109
  (
    n128,
    n62,
    n30,
    n48,
    n37
  );


  or
  g110
  (
    n124,
    n39,
    n26,
    n48
  );


  xnor
  g111
  (
    n132,
    n29,
    n31,
    n77,
    n35
  );


  and
  g112
  (
    n111,
    n84,
    n79,
    n54,
    n28
  );


  nand
  g113
  (
    n87,
    n86,
    n48,
    n23,
    n29
  );


  xnor
  g114
  (
    n133,
    n53,
    n22,
    n51,
    n43
  );


  or
  g115
  (
    n103,
    n53,
    n55,
    n56,
    n84
  );


  nor
  g116
  (
    n94,
    n41,
    n50,
    n44,
    n46
  );


  nand
  g117
  (
    n127,
    n75,
    n49,
    n25,
    n81
  );


  nor
  g118
  (
    n92,
    n29,
    n57,
    n21,
    n38
  );


  or
  g119
  (
    n118,
    n81,
    n35,
    n80,
    n36
  );


  and
  g120
  (
    n136,
    n54,
    n27,
    n73,
    n46
  );


  nor
  g121
  (
    n145,
    n73,
    n38,
    n24
  );


  nor
  g122
  (
    n146,
    n81,
    n50,
    n60,
    n79
  );


  xnor
  g123
  (
    n114,
    n34,
    n34,
    n50,
    n71
  );


  or
  g124
  (
    n135,
    n49,
    n31,
    n38,
    n25
  );


  xor
  g125
  (
    n131,
    n78,
    n49,
    n55
  );


  xnor
  g126
  (
    n97,
    n52,
    n81,
    n44,
    n54
  );


  and
  g127
  (
    n98,
    n57,
    n31,
    n41,
    n63
  );


  xor
  g128
  (
    n119,
    n78,
    n32,
    n84,
    n41
  );


  nor
  g129
  (
    n108,
    n26,
    n64,
    n58,
    n63
  );


  nand
  g130
  (
    n152,
    n98,
    n131,
    n147,
    n113
  );


  nor
  g131
  (
    n160,
    n90,
    n128,
    n144,
    n93
  );


  xnor
  g132
  (
    n163,
    n148,
    n147,
    n94,
    n140
  );


  nand
  g133
  (
    n158,
    n135,
    n147,
    n101,
    n141
  );


  xnor
  g134
  (
    n156,
    n121,
    n114,
    n89,
    n99
  );


  nand
  g135
  (
    n149,
    n136,
    n105,
    n110,
    n109
  );


  nand
  g136
  (
    n165,
    n104,
    n120,
    n118,
    n132
  );


  nor
  g137
  (
    n162,
    n112,
    n87,
    n88,
    n108
  );


  or
  g138
  (
    n161,
    n97,
    n129,
    n127,
    n96
  );


  nand
  g139
  (
    n155,
    n102,
    n148,
    n126,
    n125
  );


  or
  g140
  (
    n159,
    n148,
    n146,
    n103,
    n119
  );


  and
  g141
  (
    n164,
    n130,
    n91,
    n123,
    n106
  );


  and
  g142
  (
    AntiSAT_key_wire,
    n116,
    n107,
    n111,
    n95
  );


  nand
  g143
  (
    n151,
    n137,
    n100,
    n124,
    n122
  );


  nor
  g144
  (
    n154,
    n117,
    n147,
    n92,
    n145
  );


  xor
  g145
  (
    n153,
    n115,
    n138,
    n139,
    n134
  );


  or
  g146
  (
    n157,
    n143,
    n148,
    n133,
    n142
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_18
  (
    gbar_input_0_0,
    keyIn_0_18,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_19
  (
    gbar_input_0_1,
    keyIn_0_19,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_20
  (
    gbar_input_0_2,
    keyIn_0_20,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_21
  (
    gbar_input_0_3,
    keyIn_0_21,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_22
  (
    gbar_input_0_4,
    keyIn_0_22,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_23
  (
    gbar_input_0_5,
    keyIn_0_23,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_24
  (
    gbar_input_0_6,
    keyIn_0_24,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_25
  (
    gbar_input_0_7,
    keyIn_0_25,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_8,
    keyIn_0_26,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_9,
    keyIn_0_27,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_10,
    keyIn_0_28,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_11,
    keyIn_0_29,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_12,
    keyIn_0_30,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_13,
    keyIn_0_31,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_14,
    keyIn_0_32,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_15,
    keyIn_0_33,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_16,
    keyIn_0_34,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_17,
    keyIn_0_35,
    n18
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n150,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

