

module c1355
(
  G1,
  G10,
  G11,
  G12,
  G13,
  G1324,
  G1325,
  G1326,
  G1327,
  G1328,
  G1329,
  G1330,
  G1331,
  G1332,
  G1333,
  G1334,
  G1335,
  G1336,
  G1337,
  G1338,
  G1339,
  G1340,
  G1341,
  G1342,
  G1343,
  G1344,
  G1345,
  G1346,
  G1347,
  G1348,
  G1349,
  G1350,
  G1351,
  G1352,
  G1353,
  G1354,
  G1355,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G2,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G3,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G4,
  G40,
  G41,
  G5,
  G6,
  G7,
  G8,
  G9,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;
  output G1324;output G1325;output G1326;output G1327;output G1328;output G1329;output G1330;output G1331;output G1332;output G1333;output G1334;output G1335;output G1336;output G1337;output G1338;output G1339;output G1340;output G1341;output G1342;output G1343;output G1344;output G1345;output G1346;output G1347;output G1348;output G1349;output G1350;output G1351;output G1352;output G1353;output G1354;output G1355;
  wire G242;wire G245;wire G248;wire G251;wire G254;wire G257;wire G260;wire G263;wire G266;wire G269;wire G272;wire G275;wire G278;wire G281;wire G284;wire G287;wire G290;wire G293;wire G296;wire G299;wire G302;wire G305;wire G308;wire G311;wire G314;wire G317;wire G320;wire G323;wire G326;wire G329;wire G332;wire G335;wire G338;wire G341;wire G344;wire G347;wire G350;wire G353;wire G356;wire G359;wire G362;wire G363;wire G364;wire G365;wire G366;wire G367;wire G368;wire G369;wire G370;wire G371;wire G372;wire G373;wire G374;wire G375;wire G376;wire G377;wire G378;wire G379;wire G380;wire G381;wire G382;wire G383;wire G384;wire G385;wire G386;wire G387;wire G388;wire G389;wire G390;wire G391;wire G392;wire G393;wire G394;wire G395;wire G396;wire G397;wire G398;wire G399;wire G400;wire G401;wire G402;wire G403;wire G404;wire G405;wire G406;wire G407;wire G408;wire G409;wire G410;wire G411;wire G412;wire G413;wire G414;wire G415;wire G416;wire G417;wire G418;wire G419;wire G420;wire G421;wire G422;wire G423;wire G424;wire G425;wire G426;wire G429;wire G432;wire G435;wire G438;wire G441;wire G444;wire G447;wire G450;wire G453;wire G456;wire G459;wire G462;wire G465;wire G468;wire G471;wire G474;wire G477;wire G480;wire G483;wire G486;wire G489;wire G492;wire G495;wire G498;wire G501;wire G504;wire G507;wire G510;wire G513;wire G516;wire G519;wire G522;wire G525;wire G528;wire G531;wire G534;wire G537;wire G540;wire G543;wire G546;wire G549;wire G552;wire G555;wire G558;wire G561;wire G564;wire G567;wire G570;wire G571;wire G572;wire G573;wire G574;wire G575;wire G576;wire G577;wire G578;wire G579;wire G580;wire G581;wire G582;wire G583;wire G584;wire G585;wire G586;wire G587;wire G588;wire G589;wire G590;wire G591;wire G592;wire G593;wire G594;wire G595;wire G596;wire G597;wire G598;wire G599;wire G600;wire G601;wire G602;wire G607;wire G612;wire G617;wire G622;wire G627;wire G632;wire G637;wire G642;wire G645;wire G648;wire G651;wire G654;wire G657;wire G660;wire G663;wire G666;wire G669;wire G672;wire G675;wire G678;wire G681;wire G684;wire G687;wire G690;wire G691;wire G692;wire G693;wire G694;wire G695;wire G696;wire G697;wire G698;wire G699;wire G700;wire G701;wire G702;wire G703;wire G704;wire G705;wire G706;wire G709;wire G712;wire G715;wire G718;wire G721;wire G724;wire G727;wire G730;wire G733;wire G736;wire G739;wire G742;wire G745;wire G748;wire G751;wire G754;wire G755;wire G756;wire G757;wire G758;wire G759;wire G760;wire G761;wire G762;wire G763;wire G764;wire G765;wire G766;wire G767;wire G768;wire G769;wire G770;wire G773;wire G776;wire G779;wire G782;wire G785;wire G788;wire G791;wire G794;wire G797;wire G800;wire G803;wire G806;wire G809;wire G812;wire G815;wire G818;wire G819;wire G820;wire G821;wire G822;wire G823;wire G824;wire G825;wire G826;wire G827;wire G828;wire G829;wire G830;wire G831;wire G832;wire G833;wire G834;wire G847;wire G860;wire G873;wire G886;wire G899;wire G912;wire G925;wire G938;wire G939;wire G940;wire G941;wire G942;wire G943;wire G944;wire G945;wire G946;wire G947;wire G948;wire G949;wire G950;wire G951;wire G952;wire G953;wire G954;wire G955;wire G956;wire G957;wire G958;wire G959;wire G960;wire G961;wire G962;wire G963;wire G964;wire G965;wire G966;wire G967;wire G968;wire G969;wire G970;wire G971;wire G972;wire G973;wire G974;wire G975;wire G976;wire G977;wire G978;wire G979;wire G980;wire G981;wire G982;wire G983;wire G984;wire G985;wire G986;wire G991;wire G996;wire G1001;wire G1006;wire G1011;wire G1016;wire G1021;wire G1026;wire G1031;wire G1036;wire G1039;wire G1042;wire G1045;wire G1048;wire G1051;wire G1054;wire G1057;wire G1060;wire G1063;wire G1066;wire G1069;wire G1072;wire G1075;wire G1078;wire G1081;wire G1084;wire G1087;wire G1090;wire G1093;wire G1096;wire G1099;wire G1102;wire G1105;wire G1108;wire G1111;wire G1114;wire G1117;wire G1120;wire G1123;wire G1126;wire G1129;wire G1132;wire G1135;wire G1138;wire G1141;wire G1144;wire G1147;wire G1150;wire G1153;wire G1156;wire G1159;wire G1162;wire G1165;wire G1168;wire G1171;wire G1174;wire G1177;wire G1180;wire G1183;wire G1186;wire G1189;wire G1192;wire G1195;wire G1198;wire G1201;wire G1204;wire G1207;wire G1210;wire G1213;wire G1216;wire G1219;wire G1222;wire G1225;wire G1228;wire G1229;wire G1230;wire G1231;wire G1232;wire G1233;wire G1234;wire G1235;wire G1236;wire G1237;wire G1238;wire G1239;wire G1240;wire G1241;wire G1242;wire G1243;wire G1244;wire G1245;wire G1246;wire G1247;wire G1248;wire G1249;wire G1250;wire G1251;wire G1252;wire G1253;wire G1254;wire G1255;wire G1256;wire G1257;wire G1258;wire G1259;wire G1260;wire G1261;wire G1262;wire G1263;wire G1264;wire G1265;wire G1266;wire G1267;wire G1268;wire G1269;wire G1270;wire G1271;wire G1272;wire G1273;wire G1274;wire G1275;wire G1276;wire G1277;wire G1278;wire G1279;wire G1280;wire G1281;wire G1282;wire G1283;wire G1284;wire G1285;wire G1286;wire G1287;wire G1288;wire G1289;wire G1290;wire G1291;wire G1292;wire G1293;wire G1294;wire G1295;wire G1296;wire G1297;wire G1298;wire G1299;wire G1300;wire G1301;wire G1302;wire G1303;wire G1304;wire G1305;wire G1306;wire G1307;wire G1308;wire G1309;wire G1310;wire G1311;wire G1312;wire G1313;wire G1314;wire G1315;wire G1316;wire G1317;wire G1318;wire G1319;wire G1320;wire G1321;wire G1322;wire G1323;wire zip_xor_output_0;wire zip_xor_output_1;wire zip_xor_output_2;wire zip_xor_output_3;wire zip_xor_output_4;wire ha_0_0_sum;wire ha_0_0_carry;wire ha_1_0_sum;wire ha_1_0_carry;wire ha_1_1_sum;wire ha_1_1_carry;wire ha_2_0_sum;wire ha_2_0_carry;wire ha_2_1_sum;wire ha_2_1_carry;wire ha_2_2_sum;wire ha_2_2_carry;wire ha_3_0_sum;wire ha_3_0_carry;wire ha_3_1_sum;wire ha_3_1_carry;wire ha_3_2_sum;wire ha_3_2_carry;wire ha_3_3_sum;wire ha_3_3_carry;wire comparator_0_0;wire comparator_0_1;wire comparator_0_2;wire comparator_output;wire mask_xnor1_0;wire mask_xnor1_1;wire mask_xnor1_2;wire mask_xnor0_3;wire mask_xnor0_4;wire mask_and_0;wire mask_xnor0_0;wire mask_xnor1_4;wire mask_and_1;wire mask_xnor0_1;wire mask_xnor1_3;wire mask_and_2;wire mask_xnor0_2;wire mask_and_3;wire mask_and_4;wire mask_and_5;wire mask_and_6;wire mask_output;wire key_block_output;wire unmodified_output;

  and
  AND2_0
  (
    G242,
    G33,
    G41
  );


  and
  AND2_1
  (
    G245,
    G34,
    G41
  );


  and
  AND2_2
  (
    G248,
    G35,
    G41
  );


  and
  AND2_3
  (
    G251,
    G36,
    G41
  );


  and
  AND2_4
  (
    G254,
    G37,
    G41
  );


  and
  AND2_5
  (
    G257,
    G38,
    G41
  );


  and
  AND2_6
  (
    G260,
    G39,
    G41
  );


  and
  AND2_7
  (
    G263,
    G40,
    G41
  );


  nand
  NAND2_0
  (
    G266,
    G1,
    G2
  );


  nand
  NAND2_1
  (
    G269,
    G3,
    G4
  );


  nand
  NAND2_2
  (
    G272,
    G5,
    G6
  );


  nand
  NAND2_3
  (
    G275,
    G7,
    G8
  );


  nand
  NAND2_4
  (
    G278,
    G9,
    G10
  );


  nand
  NAND2_5
  (
    G281,
    G11,
    G12
  );


  nand
  NAND2_6
  (
    G284,
    G13,
    G14
  );


  nand
  NAND2_7
  (
    G287,
    G15,
    G16
  );


  nand
  NAND2_8
  (
    G290,
    G17,
    G18
  );


  nand
  NAND2_9
  (
    G293,
    G19,
    G20
  );


  nand
  NAND2_10
  (
    G296,
    G21,
    G22
  );


  nand
  NAND2_11
  (
    G299,
    G23,
    G24
  );


  nand
  NAND2_12
  (
    G302,
    G25,
    G26
  );


  nand
  NAND2_13
  (
    G305,
    G27,
    G28
  );


  nand
  NAND2_14
  (
    G308,
    G29,
    G30
  );


  nand
  NAND2_15
  (
    G311,
    G31,
    G32
  );


  nand
  NAND2_16
  (
    G314,
    G1,
    G5
  );


  nand
  NAND2_17
  (
    G317,
    G9,
    G13
  );


  nand
  NAND2_18
  (
    G320,
    G2,
    G6
  );


  nand
  NAND2_19
  (
    G323,
    G10,
    G14
  );


  nand
  NAND2_20
  (
    G326,
    G3,
    G7
  );


  nand
  NAND2_21
  (
    G329,
    G11,
    G15
  );


  nand
  NAND2_22
  (
    G332,
    G4,
    G8
  );


  nand
  NAND2_23
  (
    G335,
    G12,
    G16
  );


  nand
  NAND2_24
  (
    G338,
    G17,
    G21
  );


  nand
  NAND2_25
  (
    G341,
    G25,
    G29
  );


  nand
  NAND2_26
  (
    G344,
    G18,
    G22
  );


  nand
  NAND2_27
  (
    G347,
    G26,
    G30
  );


  nand
  NAND2_28
  (
    G350,
    G19,
    G23
  );


  nand
  NAND2_29
  (
    G353,
    G27,
    G31
  );


  nand
  NAND2_30
  (
    G356,
    G20,
    G24
  );


  nand
  NAND2_31
  (
    G359,
    G28,
    G32
  );


  nand
  NAND2_32
  (
    G362,
    G1,
    G266
  );


  nand
  NAND2_33
  (
    G363,
    G2,
    G266
  );


  nand
  NAND2_34
  (
    G364,
    G3,
    G269
  );


  nand
  NAND2_35
  (
    G365,
    G4,
    G269
  );


  nand
  NAND2_36
  (
    G366,
    G5,
    G272
  );


  nand
  NAND2_37
  (
    G367,
    G6,
    G272
  );


  nand
  NAND2_38
  (
    G368,
    G7,
    G275
  );


  nand
  NAND2_39
  (
    G369,
    G8,
    G275
  );


  nand
  NAND2_40
  (
    G370,
    G9,
    G278
  );


  nand
  NAND2_41
  (
    G371,
    G10,
    G278
  );


  nand
  NAND2_42
  (
    G372,
    G11,
    G281
  );


  nand
  NAND2_43
  (
    G373,
    G12,
    G281
  );


  nand
  NAND2_44
  (
    G374,
    G13,
    G284
  );


  nand
  NAND2_45
  (
    G375,
    G14,
    G284
  );


  nand
  NAND2_46
  (
    G376,
    G15,
    G287
  );


  nand
  NAND2_47
  (
    G377,
    G16,
    G287
  );


  nand
  NAND2_48
  (
    G378,
    G17,
    G290
  );


  nand
  NAND2_49
  (
    G379,
    G18,
    G290
  );


  nand
  NAND2_50
  (
    G380,
    G19,
    G293
  );


  nand
  NAND2_51
  (
    G381,
    G20,
    G293
  );


  nand
  NAND2_52
  (
    G382,
    G21,
    G296
  );


  nand
  NAND2_53
  (
    G383,
    G22,
    G296
  );


  nand
  NAND2_54
  (
    G384,
    G23,
    G299
  );


  nand
  NAND2_55
  (
    G385,
    G24,
    G299
  );


  nand
  NAND2_56
  (
    G386,
    G25,
    G302
  );


  nand
  NAND2_57
  (
    G387,
    G26,
    G302
  );


  nand
  NAND2_58
  (
    G388,
    G27,
    G305
  );


  nand
  NAND2_59
  (
    G389,
    G28,
    G305
  );


  nand
  NAND2_60
  (
    G390,
    G29,
    G308
  );


  nand
  NAND2_61
  (
    G391,
    G30,
    G308
  );


  nand
  NAND2_62
  (
    G392,
    G31,
    G311
  );


  nand
  NAND2_63
  (
    G393,
    G32,
    G311
  );


  nand
  NAND2_64
  (
    G394,
    G1,
    G314
  );


  nand
  NAND2_65
  (
    G395,
    G5,
    G314
  );


  nand
  NAND2_66
  (
    G396,
    G9,
    G317
  );


  nand
  NAND2_67
  (
    G397,
    G13,
    G317
  );


  nand
  NAND2_68
  (
    G398,
    G2,
    G320
  );


  nand
  NAND2_69
  (
    G399,
    G6,
    G320
  );


  nand
  NAND2_70
  (
    G400,
    G10,
    G323
  );


  nand
  NAND2_71
  (
    G401,
    G14,
    G323
  );


  nand
  NAND2_72
  (
    G402,
    G3,
    G326
  );


  nand
  NAND2_73
  (
    G403,
    G7,
    G326
  );


  nand
  NAND2_74
  (
    G404,
    G11,
    G329
  );


  nand
  NAND2_75
  (
    G405,
    G15,
    G329
  );


  nand
  NAND2_76
  (
    G406,
    G4,
    G332
  );


  nand
  NAND2_77
  (
    G407,
    G8,
    G332
  );


  nand
  NAND2_78
  (
    G408,
    G12,
    G335
  );


  nand
  NAND2_79
  (
    G409,
    G16,
    G335
  );


  nand
  NAND2_80
  (
    G410,
    G17,
    G338
  );


  nand
  NAND2_81
  (
    G411,
    G21,
    G338
  );


  nand
  NAND2_82
  (
    G412,
    G25,
    G341
  );


  nand
  NAND2_83
  (
    G413,
    G29,
    G341
  );


  nand
  NAND2_84
  (
    G414,
    G18,
    G344
  );


  nand
  NAND2_85
  (
    G415,
    G22,
    G344
  );


  nand
  NAND2_86
  (
    G416,
    G26,
    G347
  );


  nand
  NAND2_87
  (
    G417,
    G30,
    G347
  );


  nand
  NAND2_88
  (
    G418,
    G19,
    G350
  );


  nand
  NAND2_89
  (
    G419,
    G23,
    G350
  );


  nand
  NAND2_90
  (
    G420,
    G27,
    G353
  );


  nand
  NAND2_91
  (
    G421,
    G31,
    G353
  );


  nand
  NAND2_92
  (
    G422,
    G20,
    G356
  );


  nand
  NAND2_93
  (
    G423,
    G24,
    G356
  );


  nand
  NAND2_94
  (
    G424,
    G28,
    G359
  );


  nand
  NAND2_95
  (
    G425,
    G32,
    G359
  );


  nand
  NAND2_96
  (
    G426,
    G362,
    G363
  );


  nand
  NAND2_97
  (
    G429,
    G364,
    G365
  );


  nand
  NAND2_98
  (
    G432,
    G366,
    G367
  );


  nand
  NAND2_99
  (
    G435,
    G368,
    G369
  );


  nand
  NAND2_100
  (
    G438,
    G370,
    G371
  );


  nand
  NAND2_101
  (
    G441,
    G372,
    G373
  );


  nand
  NAND2_102
  (
    G444,
    G374,
    G375
  );


  nand
  NAND2_103
  (
    G447,
    G376,
    G377
  );


  nand
  NAND2_104
  (
    G450,
    G378,
    G379
  );


  nand
  NAND2_105
  (
    G453,
    G380,
    G381
  );


  nand
  NAND2_106
  (
    G456,
    G382,
    G383
  );


  nand
  NAND2_107
  (
    G459,
    G384,
    G385
  );


  nand
  NAND2_108
  (
    G462,
    G386,
    G387
  );


  nand
  NAND2_109
  (
    G465,
    G388,
    G389
  );


  nand
  NAND2_110
  (
    G468,
    G390,
    G391
  );


  nand
  NAND2_111
  (
    G471,
    G392,
    G393
  );


  nand
  NAND2_112
  (
    G474,
    G394,
    G395
  );


  nand
  NAND2_113
  (
    G477,
    G396,
    G397
  );


  nand
  NAND2_114
  (
    G480,
    G398,
    G399
  );


  nand
  NAND2_115
  (
    G483,
    G400,
    G401
  );


  nand
  NAND2_116
  (
    G486,
    G402,
    G403
  );


  nand
  NAND2_117
  (
    G489,
    G404,
    G405
  );


  nand
  NAND2_118
  (
    G492,
    G406,
    G407
  );


  nand
  NAND2_119
  (
    G495,
    G408,
    G409
  );


  nand
  NAND2_120
  (
    G498,
    G410,
    G411
  );


  nand
  NAND2_121
  (
    G501,
    G412,
    G413
  );


  nand
  NAND2_122
  (
    G504,
    G414,
    G415
  );


  nand
  NAND2_123
  (
    G507,
    G416,
    G417
  );


  nand
  NAND2_124
  (
    G510,
    G418,
    G419
  );


  nand
  NAND2_125
  (
    G513,
    G420,
    G421
  );


  nand
  NAND2_126
  (
    G516,
    G422,
    G423
  );


  nand
  NAND2_127
  (
    G519,
    G424,
    G425
  );


  nand
  NAND2_128
  (
    G522,
    G426,
    G429
  );


  nand
  NAND2_129
  (
    G525,
    G432,
    G435
  );


  nand
  NAND2_130
  (
    G528,
    G438,
    G441
  );


  nand
  NAND2_131
  (
    G531,
    G444,
    G447
  );


  nand
  NAND2_132
  (
    G534,
    G450,
    G453
  );


  nand
  NAND2_133
  (
    G537,
    G456,
    G459
  );


  nand
  NAND2_134
  (
    G540,
    G462,
    G465
  );


  nand
  NAND2_135
  (
    G543,
    G468,
    G471
  );


  nand
  NAND2_136
  (
    G546,
    G474,
    G477
  );


  nand
  NAND2_137
  (
    G549,
    G480,
    G483
  );


  nand
  NAND2_138
  (
    G552,
    G486,
    G489
  );


  nand
  NAND2_139
  (
    G555,
    G492,
    G495
  );


  nand
  NAND2_140
  (
    G558,
    G498,
    G501
  );


  nand
  NAND2_141
  (
    G561,
    G504,
    G507
  );


  nand
  NAND2_142
  (
    G564,
    G510,
    G513
  );


  nand
  NAND2_143
  (
    G567,
    G516,
    G519
  );


  nand
  NAND2_144
  (
    G570,
    G426,
    G522
  );


  nand
  NAND2_145
  (
    G571,
    G429,
    G522
  );


  nand
  NAND2_146
  (
    G572,
    G432,
    G525
  );


  nand
  NAND2_147
  (
    G573,
    G435,
    G525
  );


  nand
  NAND2_148
  (
    G574,
    G438,
    G528
  );


  nand
  NAND2_149
  (
    G575,
    G441,
    G528
  );


  nand
  NAND2_150
  (
    G576,
    G444,
    G531
  );


  nand
  NAND2_151
  (
    G577,
    G447,
    G531
  );


  nand
  NAND2_152
  (
    G578,
    G450,
    G534
  );


  nand
  NAND2_153
  (
    G579,
    G453,
    G534
  );


  nand
  NAND2_154
  (
    G580,
    G456,
    G537
  );


  nand
  NAND2_155
  (
    G581,
    G459,
    G537
  );


  nand
  NAND2_156
  (
    G582,
    G462,
    G540
  );


  nand
  NAND2_157
  (
    G583,
    G465,
    G540
  );


  nand
  NAND2_158
  (
    G584,
    G468,
    G543
  );


  nand
  NAND2_159
  (
    G585,
    G471,
    G543
  );


  nand
  NAND2_160
  (
    G586,
    G474,
    G546
  );


  nand
  NAND2_161
  (
    G587,
    G477,
    G546
  );


  nand
  NAND2_162
  (
    G588,
    G480,
    G549
  );


  nand
  NAND2_163
  (
    G589,
    G483,
    G549
  );


  nand
  NAND2_164
  (
    G590,
    G486,
    G552
  );


  nand
  NAND2_165
  (
    G591,
    G489,
    G552
  );


  nand
  NAND2_166
  (
    G592,
    G492,
    G555
  );


  nand
  NAND2_167
  (
    G593,
    G495,
    G555
  );


  nand
  NAND2_168
  (
    G594,
    G498,
    G558
  );


  nand
  NAND2_169
  (
    G595,
    G501,
    G558
  );


  nand
  NAND2_170
  (
    G596,
    G504,
    G561
  );


  nand
  NAND2_171
  (
    G597,
    G507,
    G561
  );


  nand
  NAND2_172
  (
    G598,
    G510,
    G564
  );


  nand
  NAND2_173
  (
    G599,
    G513,
    G564
  );


  nand
  NAND2_174
  (
    G600,
    G516,
    G567
  );


  nand
  NAND2_175
  (
    G601,
    G519,
    G567
  );


  nand
  NAND2_176
  (
    G602,
    G570,
    G571
  );


  nand
  NAND2_177
  (
    G607,
    G572,
    G573
  );


  nand
  NAND2_178
  (
    G612,
    G574,
    G575
  );


  nand
  NAND2_179
  (
    G617,
    G576,
    G577
  );


  nand
  NAND2_180
  (
    G622,
    G578,
    G579
  );


  nand
  NAND2_181
  (
    G627,
    G580,
    G581
  );


  nand
  NAND2_182
  (
    G632,
    G582,
    G583
  );


  nand
  NAND2_183
  (
    G637,
    G584,
    G585
  );


  nand
  NAND2_184
  (
    G642,
    G586,
    G587
  );


  nand
  NAND2_185
  (
    G645,
    G588,
    G589
  );


  nand
  NAND2_186
  (
    G648,
    G590,
    G591
  );


  nand
  NAND2_187
  (
    G651,
    G592,
    G593
  );


  nand
  NAND2_188
  (
    G654,
    G594,
    G595
  );


  nand
  NAND2_189
  (
    G657,
    G596,
    G597
  );


  nand
  NAND2_190
  (
    G660,
    G598,
    G599
  );


  nand
  NAND2_191
  (
    G663,
    G600,
    G601
  );


  nand
  NAND2_192
  (
    G666,
    G602,
    G607
  );


  nand
  NAND2_193
  (
    G669,
    G612,
    G617
  );


  nand
  NAND2_194
  (
    G672,
    G602,
    G612
  );


  nand
  NAND2_195
  (
    G675,
    G607,
    G617
  );


  nand
  NAND2_196
  (
    G678,
    G622,
    G627
  );


  nand
  NAND2_197
  (
    G681,
    G632,
    G637
  );


  nand
  NAND2_198
  (
    G684,
    G622,
    G632
  );


  nand
  NAND2_199
  (
    G687,
    G627,
    G637
  );


  nand
  NAND2_200
  (
    G690,
    G602,
    G666
  );


  nand
  NAND2_201
  (
    G691,
    G607,
    G666
  );


  nand
  NAND2_202
  (
    G692,
    G612,
    G669
  );


  nand
  NAND2_203
  (
    G693,
    G617,
    G669
  );


  nand
  NAND2_204
  (
    G694,
    G602,
    G672
  );


  nand
  NAND2_205
  (
    G695,
    G612,
    G672
  );


  nand
  NAND2_206
  (
    G696,
    G607,
    G675
  );


  nand
  NAND2_207
  (
    G697,
    G617,
    G675
  );


  nand
  NAND2_208
  (
    G698,
    G622,
    G678
  );


  nand
  NAND2_209
  (
    G699,
    G627,
    G678
  );


  nand
  NAND2_210
  (
    G700,
    G632,
    G681
  );


  nand
  NAND2_211
  (
    G701,
    G637,
    G681
  );


  nand
  NAND2_212
  (
    G702,
    G622,
    G684
  );


  nand
  NAND2_213
  (
    G703,
    G632,
    G684
  );


  nand
  NAND2_214
  (
    G704,
    G627,
    G687
  );


  nand
  NAND2_215
  (
    G705,
    G637,
    G687
  );


  nand
  NAND2_216
  (
    G706,
    G690,
    G691
  );


  nand
  NAND2_217
  (
    G709,
    G692,
    G693
  );


  nand
  NAND2_218
  (
    G712,
    G694,
    G695
  );


  nand
  NAND2_219
  (
    G715,
    G696,
    G697
  );


  nand
  NAND2_220
  (
    G718,
    G698,
    G699
  );


  nand
  NAND2_221
  (
    G721,
    G700,
    G701
  );


  nand
  NAND2_222
  (
    G724,
    G702,
    G703
  );


  nand
  NAND2_223
  (
    G727,
    G704,
    G705
  );


  nand
  NAND2_224
  (
    G730,
    G242,
    G718
  );


  nand
  NAND2_225
  (
    G733,
    G245,
    G721
  );


  nand
  NAND2_226
  (
    G736,
    G248,
    G724
  );


  nand
  NAND2_227
  (
    G739,
    G251,
    G727
  );


  nand
  NAND2_228
  (
    G742,
    G254,
    G706
  );


  nand
  NAND2_229
  (
    G745,
    G257,
    G709
  );


  nand
  NAND2_230
  (
    G748,
    G260,
    G712
  );


  nand
  NAND2_231
  (
    G751,
    G263,
    G715
  );


  nand
  NAND2_232
  (
    G754,
    G242,
    G730
  );


  nand
  NAND2_233
  (
    G755,
    G718,
    G730
  );


  nand
  NAND2_234
  (
    G756,
    G245,
    G733
  );


  nand
  NAND2_235
  (
    G757,
    G721,
    G733
  );


  nand
  NAND2_236
  (
    G758,
    G248,
    G736
  );


  nand
  NAND2_237
  (
    G759,
    G724,
    G736
  );


  nand
  NAND2_238
  (
    G760,
    G251,
    G739
  );


  nand
  NAND2_239
  (
    G761,
    G727,
    G739
  );


  nand
  NAND2_240
  (
    G762,
    G254,
    G742
  );


  nand
  NAND2_241
  (
    G763,
    G706,
    G742
  );


  nand
  NAND2_242
  (
    G764,
    G257,
    G745
  );


  nand
  NAND2_243
  (
    G765,
    G709,
    G745
  );


  nand
  NAND2_244
  (
    G766,
    G260,
    G748
  );


  nand
  NAND2_245
  (
    G767,
    G712,
    G748
  );


  nand
  NAND2_246
  (
    G768,
    G263,
    G751
  );


  nand
  NAND2_247
  (
    G769,
    G715,
    G751
  );


  nand
  NAND2_248
  (
    G770,
    G754,
    G755
  );


  nand
  NAND2_249
  (
    G773,
    G756,
    G757
  );


  nand
  NAND2_250
  (
    G776,
    G758,
    G759
  );


  nand
  NAND2_251
  (
    G779,
    G760,
    G761
  );


  nand
  NAND2_252
  (
    G782,
    G762,
    G763
  );


  nand
  NAND2_253
  (
    G785,
    G764,
    G765
  );


  nand
  NAND2_254
  (
    G788,
    G766,
    G767
  );


  nand
  NAND2_255
  (
    G791,
    G768,
    G769
  );


  nand
  NAND2_256
  (
    G794,
    G642,
    G770
  );


  nand
  NAND2_257
  (
    G797,
    G645,
    G773
  );


  nand
  NAND2_258
  (
    G800,
    G648,
    G776
  );


  nand
  NAND2_259
  (
    G803,
    G651,
    G779
  );


  nand
  NAND2_260
  (
    G806,
    G654,
    G782
  );


  nand
  NAND2_261
  (
    G809,
    G657,
    G785
  );


  nand
  NAND2_262
  (
    G812,
    G660,
    G788
  );


  nand
  NAND2_263
  (
    G815,
    G663,
    G791
  );


  nand
  NAND2_264
  (
    G818,
    G642,
    G794
  );


  nand
  NAND2_265
  (
    G819,
    G770,
    G794
  );


  nand
  NAND2_266
  (
    G820,
    G645,
    G797
  );


  nand
  NAND2_267
  (
    G821,
    G773,
    G797
  );


  nand
  NAND2_268
  (
    G822,
    G648,
    G800
  );


  nand
  NAND2_269
  (
    G823,
    G776,
    G800
  );


  nand
  NAND2_270
  (
    G824,
    G651,
    G803
  );


  nand
  NAND2_271
  (
    G825,
    G779,
    G803
  );


  nand
  NAND2_272
  (
    G826,
    G654,
    G806
  );


  nand
  NAND2_273
  (
    G827,
    G782,
    G806
  );


  nand
  NAND2_274
  (
    G828,
    G657,
    G809
  );


  nand
  NAND2_275
  (
    G829,
    G785,
    G809
  );


  nand
  NAND2_276
  (
    G830,
    G660,
    G812
  );


  nand
  NAND2_277
  (
    G831,
    G788,
    G812
  );


  nand
  NAND2_278
  (
    G832,
    G663,
    G815
  );


  nand
  NAND2_279
  (
    G833,
    G791,
    G815
  );


  nand
  NAND2_280
  (
    G834,
    G818,
    G819
  );


  nand
  NAND2_281
  (
    G847,
    G820,
    G821
  );


  nand
  NAND2_282
  (
    G860,
    G822,
    G823
  );


  nand
  NAND2_283
  (
    G873,
    G824,
    G825
  );


  nand
  NAND2_284
  (
    G886,
    G828,
    G829
  );


  nand
  NAND2_285
  (
    G899,
    G832,
    G833
  );


  nand
  NAND2_286
  (
    G912,
    G830,
    G831
  );


  nand
  NAND2_287
  (
    G925,
    G826,
    G827
  );


  not
  NOT_0
  (
    G938,
    G834
  );


  not
  NOT_1
  (
    G939,
    G847
  );


  not
  NOT_2
  (
    G940,
    G860
  );


  not
  NOT_3
  (
    G941,
    G834
  );


  not
  NOT_4
  (
    G942,
    G847
  );


  not
  NOT_5
  (
    G943,
    G873
  );


  not
  NOT_6
  (
    G944,
    G834
  );


  not
  NOT_7
  (
    G945,
    G860
  );


  not
  NOT_8
  (
    G946,
    G873
  );


  not
  NOT_9
  (
    G947,
    G847
  );


  not
  NOT_10
  (
    G948,
    G860
  );


  not
  NOT_11
  (
    G949,
    G873
  );


  not
  NOT_12
  (
    G950,
    G886
  );


  not
  NOT_13
  (
    G951,
    G899
  );


  not
  NOT_14
  (
    G952,
    G886
  );


  not
  NOT_15
  (
    G953,
    G912
  );


  not
  NOT_16
  (
    G954,
    G925
  );


  not
  NOT_17
  (
    G955,
    G899
  );


  not
  NOT_18
  (
    G956,
    G925
  );


  not
  NOT_19
  (
    G957,
    G912
  );


  not
  NOT_20
  (
    G958,
    G925
  );


  not
  NOT_21
  (
    G959,
    G886
  );


  not
  NOT_22
  (
    G960,
    G912
  );


  not
  NOT_23
  (
    G961,
    G925
  );


  not
  NOT_24
  (
    G962,
    G886
  );


  not
  NOT_25
  (
    G963,
    G899
  );


  not
  NOT_26
  (
    G964,
    G925
  );


  not
  NOT_27
  (
    G965,
    G912
  );


  not
  NOT_28
  (
    G966,
    G899
  );


  not
  NOT_29
  (
    G967,
    G886
  );


  not
  NOT_30
  (
    G968,
    G912
  );


  not
  NOT_31
  (
    G969,
    G899
  );


  not
  NOT_32
  (
    G970,
    G847
  );


  not
  NOT_33
  (
    G971,
    G873
  );


  not
  NOT_34
  (
    G972,
    G847
  );


  not
  NOT_35
  (
    G973,
    G860
  );


  not
  NOT_36
  (
    G974,
    G834
  );


  not
  NOT_37
  (
    G975,
    G873
  );


  not
  NOT_38
  (
    G976,
    G834
  );


  not
  NOT_39
  (
    G977,
    G860
  );


  and
  AND4_0
  (
    G978,
    G938,
    G939,
    G940,
    G873
  );


  and
  AND4_1
  (
    G979,
    G941,
    G942,
    G860,
    G943
  );


  and
  AND4_2
  (
    G980,
    G944,
    G847,
    G945,
    G946
  );


  and
  AND4_3
  (
    G981,
    G834,
    G947,
    G948,
    G949
  );


  and
  AND4_4
  (
    G982,
    G958,
    G959,
    G960,
    G899
  );


  and
  AND4_5
  (
    G983,
    G961,
    G962,
    G912,
    G963
  );


  and
  AND4_6
  (
    G984,
    G964,
    G886,
    G965,
    G966
  );


  and
  AND4_7
  (
    G985,
    G925,
    G967,
    G968,
    G969
  );


  or
  OR4_0
  (
    G986,
    G978,
    G979,
    G980,
    G981
  );


  or
  OR4_1
  (
    G991,
    G982,
    G983,
    G984,
    G985
  );


  and
  AND5_0
  (
    G996,
    G925,
    G950,
    G912,
    G951,
    G986
  );


  and
  AND5_1
  (
    G1001,
    G925,
    G952,
    G953,
    G899,
    G986
  );


  and
  AND5_2
  (
    G1006,
    G954,
    G886,
    G912,
    G955,
    G986
  );


  and
  AND5_3
  (
    G1011,
    G956,
    G886,
    G957,
    G899,
    G986
  );


  and
  AND5_4
  (
    G1016,
    G834,
    G970,
    G860,
    G971,
    G991
  );


  and
  AND5_5
  (
    G1021,
    G834,
    G972,
    G973,
    G873,
    G991
  );


  and
  AND5_6
  (
    G1026,
    G974,
    G847,
    G860,
    G975,
    G991
  );


  and
  AND5_7
  (
    G1031,
    G976,
    G847,
    G977,
    G873,
    G991
  );


  and
  AND2_8
  (
    G1036,
    G834,
    G996
  );


  and
  AND2_9
  (
    G1039,
    G847,
    G996
  );


  and
  AND2_10
  (
    G1042,
    G860,
    G996
  );


  and
  AND2_11
  (
    G1045,
    G873,
    G996
  );


  and
  AND2_12
  (
    G1048,
    G834,
    G1001
  );


  and
  AND2_13
  (
    G1051,
    G847,
    G1001
  );


  and
  AND2_14
  (
    G1054,
    G860,
    G1001
  );


  and
  AND2_15
  (
    G1057,
    G873,
    G1001
  );


  and
  AND2_16
  (
    G1060,
    G834,
    G1006
  );


  and
  AND2_17
  (
    G1063,
    G847,
    G1006
  );


  and
  AND2_18
  (
    G1066,
    G860,
    G1006
  );


  and
  AND2_19
  (
    G1069,
    G873,
    G1006
  );


  and
  AND2_20
  (
    G1072,
    G834,
    G1011
  );


  and
  AND2_21
  (
    G1075,
    G847,
    G1011
  );


  and
  AND2_22
  (
    G1078,
    G860,
    G1011
  );


  and
  AND2_23
  (
    G1081,
    G873,
    G1011
  );


  and
  AND2_24
  (
    G1084,
    G925,
    G1016
  );


  and
  AND2_25
  (
    G1087,
    G886,
    G1016
  );


  and
  AND2_26
  (
    G1090,
    G912,
    G1016
  );


  and
  AND2_27
  (
    G1093,
    G899,
    G1016
  );


  and
  AND2_28
  (
    G1096,
    G925,
    G1021
  );


  and
  AND2_29
  (
    G1099,
    G886,
    G1021
  );


  and
  AND2_30
  (
    G1102,
    G912,
    G1021
  );


  and
  AND2_31
  (
    G1105,
    G899,
    G1021
  );


  and
  AND2_32
  (
    G1108,
    G925,
    G1026
  );


  and
  AND2_33
  (
    G1111,
    G886,
    G1026
  );


  and
  AND2_34
  (
    G1114,
    G912,
    G1026
  );


  and
  AND2_35
  (
    G1117,
    G899,
    G1026
  );


  and
  AND2_36
  (
    G1120,
    G925,
    G1031
  );


  and
  AND2_37
  (
    G1123,
    G886,
    G1031
  );


  and
  AND2_38
  (
    G1126,
    G912,
    G1031
  );


  and
  AND2_39
  (
    G1129,
    G899,
    G1031
  );


  nand
  NAND2_288
  (
    G1132,
    G1,
    G1036
  );


  nand
  NAND2_289
  (
    G1135,
    G2,
    G1039
  );


  nand
  NAND2_290
  (
    G1138,
    G3,
    G1042
  );


  nand
  NAND2_291
  (
    G1141,
    G4,
    G1045
  );


  nand
  NAND2_292
  (
    G1144,
    G5,
    G1048
  );


  nand
  NAND2_293
  (
    G1147,
    G6,
    G1051
  );


  nand
  NAND2_294
  (
    G1150,
    G7,
    G1054
  );


  nand
  NAND2_295
  (
    G1153,
    G8,
    G1057
  );


  nand
  NAND2_296
  (
    G1156,
    G9,
    G1060
  );


  nand
  NAND2_297
  (
    G1159,
    G10,
    G1063
  );


  nand
  NAND2_298
  (
    G1162,
    G11,
    G1066
  );


  nand
  NAND2_299
  (
    G1165,
    G12,
    G1069
  );


  nand
  NAND2_300
  (
    G1168,
    G13,
    G1072
  );


  nand
  NAND2_301
  (
    G1171,
    G14,
    G1075
  );


  nand
  NAND2_302
  (
    G1174,
    G15,
    G1078
  );


  nand
  NAND2_303
  (
    G1177,
    G16,
    G1081
  );


  nand
  NAND2_304
  (
    G1180,
    G17,
    G1084
  );


  nand
  NAND2_305
  (
    G1183,
    G18,
    G1087
  );


  nand
  NAND2_306
  (
    G1186,
    G19,
    G1090
  );


  nand
  NAND2_307
  (
    G1189,
    G20,
    G1093
  );


  nand
  NAND2_308
  (
    G1192,
    G21,
    G1096
  );


  nand
  NAND2_309
  (
    G1195,
    G22,
    G1099
  );


  nand
  NAND2_310
  (
    G1198,
    G23,
    G1102
  );


  nand
  NAND2_311
  (
    G1201,
    G24,
    G1105
  );


  nand
  NAND2_312
  (
    G1204,
    G25,
    G1108
  );


  nand
  NAND2_313
  (
    G1207,
    G26,
    G1111
  );


  nand
  NAND2_314
  (
    G1210,
    G27,
    G1114
  );


  nand
  NAND2_315
  (
    G1213,
    G28,
    G1117
  );


  nand
  NAND2_316
  (
    G1216,
    G29,
    G1120
  );


  nand
  NAND2_317
  (
    G1219,
    G30,
    G1123
  );


  nand
  NAND2_318
  (
    G1222,
    G31,
    G1126
  );


  nand
  NAND2_319
  (
    G1225,
    G32,
    G1129
  );


  nand
  NAND2_320
  (
    G1228,
    G1,
    G1132
  );


  nand
  NAND2_321
  (
    G1229,
    G1036,
    G1132
  );


  nand
  NAND2_322
  (
    G1230,
    G2,
    G1135
  );


  nand
  NAND2_323
  (
    G1231,
    G1039,
    G1135
  );


  nand
  NAND2_324
  (
    G1232,
    G3,
    G1138
  );


  nand
  NAND2_325
  (
    G1233,
    G1042,
    G1138
  );


  nand
  NAND2_326
  (
    G1234,
    G4,
    G1141
  );


  nand
  NAND2_327
  (
    G1235,
    G1045,
    G1141
  );


  nand
  NAND2_328
  (
    G1236,
    G5,
    G1144
  );


  nand
  NAND2_329
  (
    G1237,
    G1048,
    G1144
  );


  nand
  NAND2_330
  (
    G1238,
    G6,
    G1147
  );


  nand
  NAND2_331
  (
    G1239,
    G1051,
    G1147
  );


  nand
  NAND2_332
  (
    G1240,
    G7,
    G1150
  );


  nand
  NAND2_333
  (
    G1241,
    G1054,
    G1150
  );


  nand
  NAND2_334
  (
    G1242,
    G8,
    G1153
  );


  nand
  NAND2_335
  (
    G1243,
    G1057,
    G1153
  );


  nand
  NAND2_336
  (
    G1244,
    G9,
    G1156
  );


  nand
  NAND2_337
  (
    G1245,
    G1060,
    G1156
  );


  nand
  NAND2_338
  (
    G1246,
    G10,
    G1159
  );


  nand
  NAND2_339
  (
    G1247,
    G1063,
    G1159
  );


  nand
  NAND2_340
  (
    G1248,
    G11,
    G1162
  );


  nand
  NAND2_341
  (
    G1249,
    G1066,
    G1162
  );


  nand
  NAND2_342
  (
    G1250,
    G12,
    G1165
  );


  nand
  NAND2_343
  (
    G1251,
    G1069,
    G1165
  );


  nand
  NAND2_344
  (
    G1252,
    G13,
    G1168
  );


  nand
  NAND2_345
  (
    G1253,
    G1072,
    G1168
  );


  nand
  NAND2_346
  (
    G1254,
    G14,
    G1171
  );


  nand
  NAND2_347
  (
    G1255,
    G1075,
    G1171
  );


  nand
  NAND2_348
  (
    G1256,
    G15,
    G1174
  );


  nand
  NAND2_349
  (
    G1257,
    G1078,
    G1174
  );


  nand
  NAND2_350
  (
    G1258,
    G16,
    G1177
  );


  nand
  NAND2_351
  (
    G1259,
    G1081,
    G1177
  );


  nand
  NAND2_352
  (
    G1260,
    G17,
    G1180
  );


  nand
  NAND2_353
  (
    G1261,
    G1084,
    G1180
  );


  nand
  NAND2_354
  (
    G1262,
    G18,
    G1183
  );


  nand
  NAND2_355
  (
    G1263,
    G1087,
    G1183
  );


  nand
  NAND2_356
  (
    G1264,
    G19,
    G1186
  );


  nand
  NAND2_357
  (
    G1265,
    G1090,
    G1186
  );


  nand
  NAND2_358
  (
    G1266,
    G20,
    G1189
  );


  nand
  NAND2_359
  (
    G1267,
    G1093,
    G1189
  );


  nand
  NAND2_360
  (
    G1268,
    G21,
    G1192
  );


  nand
  NAND2_361
  (
    G1269,
    G1096,
    G1192
  );


  nand
  NAND2_362
  (
    G1270,
    G22,
    G1195
  );


  nand
  NAND2_363
  (
    G1271,
    G1099,
    G1195
  );


  nand
  NAND2_364
  (
    G1272,
    G23,
    G1198
  );


  nand
  NAND2_365
  (
    G1273,
    G1102,
    G1198
  );


  nand
  NAND2_366
  (
    G1274,
    G24,
    G1201
  );


  nand
  NAND2_367
  (
    G1275,
    G1105,
    G1201
  );


  nand
  NAND2_368
  (
    G1276,
    G25,
    G1204
  );


  nand
  NAND2_369
  (
    G1277,
    G1108,
    G1204
  );


  nand
  NAND2_370
  (
    G1278,
    G26,
    G1207
  );


  nand
  NAND2_371
  (
    G1279,
    G1111,
    G1207
  );


  nand
  NAND2_372
  (
    G1280,
    G27,
    G1210
  );


  nand
  NAND2_373
  (
    G1281,
    G1114,
    G1210
  );


  nand
  NAND2_374
  (
    G1282,
    G28,
    G1213
  );


  nand
  NAND2_375
  (
    G1283,
    G1117,
    G1213
  );


  nand
  NAND2_376
  (
    G1284,
    G29,
    G1216
  );


  nand
  NAND2_377
  (
    G1285,
    G1120,
    G1216
  );


  nand
  NAND2_378
  (
    G1286,
    G30,
    G1219
  );


  nand
  NAND2_379
  (
    G1287,
    G1123,
    G1219
  );


  nand
  NAND2_380
  (
    G1288,
    G31,
    G1222
  );


  nand
  NAND2_381
  (
    G1289,
    G1126,
    G1222
  );


  nand
  NAND2_382
  (
    G1290,
    G32,
    G1225
  );


  nand
  NAND2_383
  (
    G1291,
    G1129,
    G1225
  );


  nand
  NAND2_384
  (
    G1292,
    G1228,
    G1229
  );


  nand
  NAND2_385
  (
    G1293,
    G1230,
    G1231
  );


  nand
  NAND2_386
  (
    G1294,
    G1232,
    G1233
  );


  nand
  NAND2_387
  (
    G1295,
    G1234,
    G1235
  );


  nand
  NAND2_388
  (
    G1296,
    G1236,
    G1237
  );


  nand
  NAND2_389
  (
    G1297,
    G1238,
    G1239
  );


  nand
  NAND2_390
  (
    G1298,
    G1240,
    G1241
  );


  nand
  NAND2_391
  (
    G1299,
    G1242,
    G1243
  );


  nand
  NAND2_392
  (
    G1300,
    G1244,
    G1245
  );


  nand
  NAND2_393
  (
    G1301,
    G1246,
    G1247
  );


  nand
  NAND2_394
  (
    G1302,
    G1248,
    G1249
  );


  nand
  NAND2_395
  (
    G1303,
    G1250,
    G1251
  );


  nand
  NAND2_396
  (
    G1304,
    G1252,
    G1253
  );


  nand
  NAND2_397
  (
    G1305,
    G1254,
    G1255
  );


  nand
  NAND2_398
  (
    G1306,
    G1256,
    G1257
  );


  nand
  NAND2_399
  (
    G1307,
    G1258,
    G1259
  );


  nand
  NAND2_400
  (
    G1308,
    G1260,
    G1261
  );


  nand
  NAND2_401
  (
    G1309,
    G1262,
    G1263
  );


  nand
  NAND2_402
  (
    G1310,
    G1264,
    G1265
  );


  nand
  NAND2_403
  (
    G1311,
    G1266,
    G1267
  );


  nand
  NAND2_404
  (
    G1312,
    G1268,
    G1269
  );


  nand
  NAND2_405
  (
    G1313,
    G1270,
    G1271
  );


  nand
  NAND2_406
  (
    G1314,
    G1272,
    G1273
  );


  nand
  NAND2_407
  (
    G1315,
    G1274,
    G1275
  );


  nand
  NAND2_408
  (
    G1316,
    G1276,
    G1277
  );


  nand
  NAND2_409
  (
    G1317,
    G1278,
    G1279
  );


  nand
  NAND2_410
  (
    G1318,
    G1280,
    G1281
  );


  nand
  NAND2_411
  (
    G1319,
    G1282,
    G1283
  );


  nand
  NAND2_412
  (
    G1320,
    G1284,
    G1285
  );


  nand
  NAND2_413
  (
    G1321,
    G1286,
    G1287
  );


  nand
  NAND2_414
  (
    G1322,
    G1288,
    G1289
  );


  nand
  NAND2_415
  (
    G1323,
    G1290,
    G1291
  );


  not
  NOT_40
  (
    G1324,
    G1292
  );


  not
  NOT_41
  (
    G1325,
    G1293
  );


  not
  NOT_42
  (
    G1326,
    G1294
  );


  not
  NOT_43
  (
    G1327,
    G1295
  );


  not
  NOT_44
  (
    G1328,
    G1296
  );


  not
  NOT_45
  (
    G1329,
    G1297
  );


  not
  NOT_46
  (
    G1330,
    G1298
  );


  not
  NOT_47
  (
    G1331,
    G1299
  );


  not
  NOT_48
  (
    G1332,
    G1300
  );


  not
  NOT_49
  (
    G1333,
    G1301
  );


  not
  NOT_50
  (
    G1334,
    G1302
  );


  not
  NOT_51
  (
    unmodified_output,
    G1303
  );


  not
  NOT_52
  (
    G1336,
    G1304
  );


  not
  NOT_53
  (
    G1337,
    G1305
  );


  not
  NOT_54
  (
    G1338,
    G1306
  );


  not
  NOT_55
  (
    G1339,
    G1307
  );


  not
  NOT_56
  (
    G1340,
    G1308
  );


  not
  NOT_57
  (
    G1341,
    G1309
  );


  not
  NOT_58
  (
    G1342,
    G1310
  );


  not
  NOT_59
  (
    G1343,
    G1311
  );


  not
  NOT_60
  (
    G1344,
    G1312
  );


  not
  NOT_61
  (
    G1345,
    G1313
  );


  not
  NOT_62
  (
    G1346,
    G1314
  );


  not
  NOT_63
  (
    G1347,
    G1315
  );


  not
  NOT_64
  (
    G1348,
    G1316
  );


  not
  NOT_65
  (
    G1349,
    G1317
  );


  not
  NOT_66
  (
    G1350,
    G1318
  );


  not
  NOT_67
  (
    G1351,
    G1319
  );


  not
  NOT_68
  (
    G1352,
    G1320
  );


  not
  NOT_69
  (
    G1353,
    G1321
  );


  not
  NOT_70
  (
    G1354,
    G1322
  );


  not
  NOT_71
  (
    G1355,
    G1323
  );


  xor
  zip_xor_0
  (
    zip_xor_output_0,
    keyIn_0_0,
    G1
  );


  xor
  zip_xor_1
  (
    zip_xor_output_1,
    keyIn_0_1,
    G2
  );


  xor
  zip_xor_2
  (
    zip_xor_output_2,
    keyIn_0_2,
    G3
  );


  xor
  zip_xor_3
  (
    zip_xor_output_3,
    keyIn_0_3,
    G4
  );


  xor
  zip_xor_4
  (
    zip_xor_output_4,
    keyIn_0_4,
    G5
  );


  xor
  ha_0_0_sum
  (
    ha_0_0_sum,
    zip_xor_output_0,
    zip_xor_output_1
  );


  and
  ha_0_0_carry
  (
    ha_0_0_carry,
    zip_xor_output_0,
    zip_xor_output_1
  );


  xor
  ha_1_0_sum
  (
    ha_1_0_sum,
    zip_xor_output_2,
    ha_0_0_sum
  );


  and
  ha_1_0_carry
  (
    ha_1_0_carry,
    zip_xor_output_2,
    ha_0_0_sum
  );


  xor
  ha_1_1_sum
  (
    ha_1_1_sum,
    ha_1_0_carry,
    ha_0_0_carry
  );


  and
  ha_1_1_carry
  (
    ha_1_1_carry,
    ha_1_0_carry,
    ha_0_0_carry
  );


  xor
  ha_2_0_sum
  (
    ha_2_0_sum,
    zip_xor_output_3,
    ha_1_0_sum
  );


  and
  ha_2_0_carry
  (
    ha_2_0_carry,
    zip_xor_output_3,
    ha_1_0_sum
  );


  xor
  ha_2_1_sum
  (
    ha_2_1_sum,
    ha_2_0_carry,
    ha_1_1_sum
  );


  and
  ha_2_1_carry
  (
    ha_2_1_carry,
    ha_2_0_carry,
    ha_1_1_sum
  );


  xor
  ha_2_2_sum
  (
    ha_2_2_sum,
    ha_2_1_carry,
    ha_1_1_carry
  );


  and
  ha_2_2_carry
  (
    ha_2_2_carry,
    ha_2_1_carry,
    ha_1_1_carry
  );


  xor
  ha_3_0_sum
  (
    ha_3_0_sum,
    zip_xor_output_4,
    ha_2_0_sum
  );


  and
  ha_3_0_carry
  (
    ha_3_0_carry,
    zip_xor_output_4,
    ha_2_0_sum
  );


  xor
  ha_3_1_sum
  (
    ha_3_1_sum,
    ha_3_0_carry,
    ha_2_1_sum
  );


  and
  ha_3_1_carry
  (
    ha_3_1_carry,
    ha_3_0_carry,
    ha_2_1_sum
  );


  xor
  ha_3_2_sum
  (
    ha_3_2_sum,
    ha_3_1_carry,
    ha_2_2_sum
  );


  and
  ha_3_2_carry
  (
    ha_3_2_carry,
    ha_3_1_carry,
    ha_2_2_sum
  );


  xor
  ha_3_3_sum
  (
    ha_3_3_sum,
    ha_3_2_carry,
    ha_2_2_carry
  );


  and
  ha_3_3_carry
  (
    ha_3_3_carry,
    ha_3_2_carry,
    ha_2_2_carry
  );


  xnor
  comparator_0_0
  (
    comparator_0_0,
    ha_3_0_sum,
    0
  );


  xnor
  comparator_0_1
  (
    comparator_0_1,
    ha_3_1_sum,
    0
  );


  xnor
  comparator_0_2
  (
    comparator_0_2,
    ha_3_2_sum,
    0
  );


  and
  comparator_and
  (
    comparator_output,
    comparator_0_0,
    comparator_0_1,
    comparator_0_2
  );


  xnor
  mask_xnor1_0
  (
    mask_xnor1_0,
    keyIn_0_0,
    1
  );


  xnor
  mask_xnor1_1
  (
    mask_xnor1_1,
    keyIn_0_1,
    1
  );


  xnor
  mask_xnor1_2
  (
    mask_xnor1_2,
    keyIn_0_2,
    1
  );


  xnor
  mask_xnor0_3
  (
    mask_xnor0_3,
    keyIn_0_3,
    0
  );


  xnor
  mask_xnor0_4
  (
    mask_xnor0_4,
    keyIn_0_4,
    0
  );


  and
  mask_and_0
  (
    mask_and_0,
    mask_xnor1_0,
    mask_xnor1_1,
    mask_xnor1_2,
    mask_xnor0_3,
    mask_xnor0_4
  );


  xnor
  mask_xnor0_0
  (
    mask_xnor0_0,
    keyIn_0_0,
    0
  );


  xnor
  mask_xnor1_4
  (
    mask_xnor1_4,
    keyIn_0_4,
    1
  );


  and
  mask_and_1
  (
    mask_and_1,
    mask_xnor0_0,
    mask_xnor1_1,
    mask_xnor1_2,
    mask_xnor0_3,
    mask_xnor1_4
  );


  xnor
  mask_xnor0_1
  (
    mask_xnor0_1,
    keyIn_0_1,
    0
  );


  xnor
  mask_xnor1_3
  (
    mask_xnor1_3,
    keyIn_0_3,
    1
  );


  and
  mask_and_2
  (
    mask_and_2,
    mask_xnor1_0,
    mask_xnor0_1,
    mask_xnor1_2,
    mask_xnor1_3,
    mask_xnor1_4
  );


  xnor
  mask_xnor0_2
  (
    mask_xnor0_2,
    keyIn_0_2,
    0
  );


  and
  mask_and_3
  (
    mask_and_3,
    mask_xnor0_0,
    mask_xnor1_1,
    mask_xnor0_2,
    mask_xnor0_3,
    mask_xnor1_4
  );


  and
  mask_and_4
  (
    mask_and_4,
    mask_xnor1_0,
    mask_xnor0_1,
    mask_xnor0_2,
    mask_xnor0_3,
    mask_xnor1_4
  );


  and
  mask_and_5
  (
    mask_and_5,
    mask_xnor1_0,
    mask_xnor0_1,
    mask_xnor1_2,
    mask_xnor1_3,
    mask_xnor0_4
  );


  and
  mask_and_6
  (
    mask_and_6,
    mask_xnor0_0,
    mask_xnor0_1,
    mask_xnor1_2,
    mask_xnor1_3,
    mask_xnor0_4
  );


  nor
  mask_output
  (
    mask_output,
    mask_and_0,
    mask_and_1,
    mask_and_2,
    mask_and_3,
    mask_and_4,
    mask_and_5,
    mask_and_6
  );


  and
  key_block_output
  (
    key_block_output,
    comparator_output,
    mask_output
  );


  xor
  flip_it
  (
    G1335,
    key_block_output,
    unmodified_output
  );


endmodule

