

module Stat_4000_361
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2762,
  n2753,
  n2764,
  n2768,
  n2761,
  n2759,
  n2754,
  n2760,
  n2758,
  n2763,
  n2755,
  n2756,
  n2766,
  n4032,
  n4025,
  n4022,
  n4026,
  n4014,
  n4031,
  n4021,
  n4015,
  n4019,
  n4023,
  n4027,
  n4020,
  n4024,
  n4018,
  n4030,
  n4028,
  n4016,
  n4029,
  n4017,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n2762;output n2753;output n2764;output n2768;output n2761;output n2759;output n2754;output n2760;output n2758;output n2763;output n2755;output n2756;output n2766;output n4032;output n4025;output n4022;output n4026;output n4014;output n4031;output n4021;output n4015;output n4019;output n4023;output n4027;output n4020;output n4024;output n4018;output n4030;output n4028;output n4016;output n4029;output n4017;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2757;wire n2765;wire n2767;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire n3011;wire n3012;wire n3013;wire n3014;wire n3015;wire n3016;wire n3017;wire n3018;wire n3019;wire n3020;wire n3021;wire n3022;wire n3023;wire n3024;wire n3025;wire n3026;wire n3027;wire n3028;wire n3029;wire n3030;wire n3031;wire n3032;wire n3033;wire n3034;wire n3035;wire n3036;wire n3037;wire n3038;wire n3039;wire n3040;wire n3041;wire n3042;wire n3043;wire n3044;wire n3045;wire n3046;wire n3047;wire n3048;wire n3049;wire n3050;wire n3051;wire n3052;wire n3053;wire n3054;wire n3055;wire n3056;wire n3057;wire n3058;wire n3059;wire n3060;wire n3061;wire n3062;wire n3063;wire n3064;wire n3065;wire n3066;wire n3067;wire n3068;wire n3069;wire n3070;wire n3071;wire n3072;wire n3073;wire n3074;wire n3075;wire n3076;wire n3077;wire n3078;wire n3079;wire n3080;wire n3081;wire n3082;wire n3083;wire n3084;wire n3085;wire n3086;wire n3087;wire n3088;wire n3089;wire n3090;wire n3091;wire n3092;wire n3093;wire n3094;wire n3095;wire n3096;wire n3097;wire n3098;wire n3099;wire n3100;wire n3101;wire n3102;wire n3103;wire n3104;wire n3105;wire n3106;wire n3107;wire n3108;wire n3109;wire n3110;wire n3111;wire n3112;wire n3113;wire n3114;wire n3115;wire n3116;wire n3117;wire n3118;wire n3119;wire n3120;wire n3121;wire n3122;wire n3123;wire n3124;wire n3125;wire n3126;wire n3127;wire n3128;wire n3129;wire n3130;wire n3131;wire n3132;wire n3133;wire n3134;wire n3135;wire n3136;wire n3137;wire n3138;wire n3139;wire n3140;wire n3141;wire n3142;wire n3143;wire n3144;wire n3145;wire n3146;wire n3147;wire n3148;wire n3149;wire n3150;wire n3151;wire n3152;wire n3153;wire n3154;wire n3155;wire n3156;wire n3157;wire n3158;wire n3159;wire n3160;wire n3161;wire n3162;wire n3163;wire n3164;wire n3165;wire n3166;wire n3167;wire n3168;wire n3169;wire n3170;wire n3171;wire n3172;wire n3173;wire n3174;wire n3175;wire n3176;wire n3177;wire n3178;wire n3179;wire n3180;wire n3181;wire n3182;wire n3183;wire n3184;wire n3185;wire n3186;wire n3187;wire n3188;wire n3189;wire n3190;wire n3191;wire n3192;wire n3193;wire n3194;wire n3195;wire n3196;wire n3197;wire n3198;wire n3199;wire n3200;wire n3201;wire n3202;wire n3203;wire n3204;wire n3205;wire n3206;wire n3207;wire n3208;wire n3209;wire n3210;wire n3211;wire n3212;wire n3213;wire n3214;wire n3215;wire n3216;wire n3217;wire n3218;wire n3219;wire n3220;wire n3221;wire n3222;wire n3223;wire n3224;wire n3225;wire n3226;wire n3227;wire n3228;wire n3229;wire n3230;wire n3231;wire n3232;wire n3233;wire n3234;wire n3235;wire n3236;wire n3237;wire n3238;wire n3239;wire n3240;wire n3241;wire n3242;wire n3243;wire n3244;wire n3245;wire n3246;wire n3247;wire n3248;wire n3249;wire n3250;wire n3251;wire n3252;wire n3253;wire n3254;wire n3255;wire n3256;wire n3257;wire n3258;wire n3259;wire n3260;wire n3261;wire n3262;wire n3263;wire n3264;wire n3265;wire n3266;wire n3267;wire n3268;wire n3269;wire n3270;wire n3271;wire n3272;wire n3273;wire n3274;wire n3275;wire n3276;wire n3277;wire n3278;wire n3279;wire n3280;wire n3281;wire n3282;wire n3283;wire n3284;wire n3285;wire n3286;wire n3287;wire n3288;wire n3289;wire n3290;wire n3291;wire n3292;wire n3293;wire n3294;wire n3295;wire n3296;wire n3297;wire n3298;wire n3299;wire n3300;wire n3301;wire n3302;wire n3303;wire n3304;wire n3305;wire n3306;wire n3307;wire n3308;wire n3309;wire n3310;wire n3311;wire n3312;wire n3313;wire n3314;wire n3315;wire n3316;wire n3317;wire n3318;wire n3319;wire n3320;wire n3321;wire n3322;wire n3323;wire n3324;wire n3325;wire n3326;wire n3327;wire n3328;wire n3329;wire n3330;wire n3331;wire n3332;wire n3333;wire n3334;wire n3335;wire n3336;wire n3337;wire n3338;wire n3339;wire n3340;wire n3341;wire n3342;wire n3343;wire n3344;wire n3345;wire n3346;wire n3347;wire n3348;wire n3349;wire n3350;wire n3351;wire n3352;wire n3353;wire n3354;wire n3355;wire n3356;wire n3357;wire n3358;wire n3359;wire n3360;wire n3361;wire n3362;wire n3363;wire n3364;wire n3365;wire n3366;wire n3367;wire n3368;wire n3369;wire n3370;wire n3371;wire n3372;wire n3373;wire n3374;wire n3375;wire n3376;wire n3377;wire n3378;wire n3379;wire n3380;wire n3381;wire n3382;wire n3383;wire n3384;wire n3385;wire n3386;wire n3387;wire n3388;wire n3389;wire n3390;wire n3391;wire n3392;wire n3393;wire n3394;wire n3395;wire n3396;wire n3397;wire n3398;wire n3399;wire n3400;wire n3401;wire n3402;wire n3403;wire n3404;wire n3405;wire n3406;wire n3407;wire n3408;wire n3409;wire n3410;wire n3411;wire n3412;wire n3413;wire n3414;wire n3415;wire n3416;wire n3417;wire n3418;wire n3419;wire n3420;wire n3421;wire n3422;wire n3423;wire n3424;wire n3425;wire n3426;wire n3427;wire n3428;wire n3429;wire n3430;wire n3431;wire n3432;wire n3433;wire n3434;wire n3435;wire n3436;wire n3437;wire n3438;wire n3439;wire n3440;wire n3441;wire n3442;wire n3443;wire n3444;wire n3445;wire n3446;wire n3447;wire n3448;wire n3449;wire n3450;wire n3451;wire n3452;wire n3453;wire n3454;wire n3455;wire n3456;wire n3457;wire n3458;wire n3459;wire n3460;wire n3461;wire n3462;wire n3463;wire n3464;wire n3465;wire n3466;wire n3467;wire n3468;wire n3469;wire n3470;wire n3471;wire n3472;wire n3473;wire n3474;wire n3475;wire n3476;wire n3477;wire n3478;wire n3479;wire n3480;wire n3481;wire n3482;wire n3483;wire n3484;wire n3485;wire n3486;wire n3487;wire n3488;wire n3489;wire n3490;wire n3491;wire n3492;wire n3493;wire n3494;wire n3495;wire n3496;wire n3497;wire n3498;wire n3499;wire n3500;wire n3501;wire n3502;wire n3503;wire n3504;wire n3505;wire n3506;wire n3507;wire n3508;wire n3509;wire n3510;wire n3511;wire n3512;wire n3513;wire n3514;wire n3515;wire n3516;wire n3517;wire n3518;wire n3519;wire n3520;wire n3521;wire n3522;wire n3523;wire n3524;wire n3525;wire n3526;wire n3527;wire n3528;wire n3529;wire n3530;wire n3531;wire n3532;wire n3533;wire n3534;wire n3535;wire n3536;wire n3537;wire n3538;wire n3539;wire n3540;wire n3541;wire n3542;wire n3543;wire n3544;wire n3545;wire n3546;wire n3547;wire n3548;wire n3549;wire n3550;wire n3551;wire n3552;wire n3553;wire n3554;wire n3555;wire n3556;wire n3557;wire n3558;wire n3559;wire n3560;wire n3561;wire n3562;wire n3563;wire n3564;wire n3565;wire n3566;wire n3567;wire n3568;wire n3569;wire n3570;wire n3571;wire n3572;wire n3573;wire n3574;wire n3575;wire n3576;wire n3577;wire n3578;wire n3579;wire n3580;wire n3581;wire n3582;wire n3583;wire n3584;wire n3585;wire n3586;wire n3587;wire n3588;wire n3589;wire n3590;wire n3591;wire n3592;wire n3593;wire n3594;wire n3595;wire n3596;wire n3597;wire n3598;wire n3599;wire n3600;wire n3601;wire n3602;wire n3603;wire n3604;wire n3605;wire n3606;wire n3607;wire n3608;wire n3609;wire n3610;wire n3611;wire n3612;wire n3613;wire n3614;wire n3615;wire n3616;wire n3617;wire n3618;wire n3619;wire n3620;wire n3621;wire n3622;wire n3623;wire n3624;wire n3625;wire n3626;wire n3627;wire n3628;wire n3629;wire n3630;wire n3631;wire n3632;wire n3633;wire n3634;wire n3635;wire n3636;wire n3637;wire n3638;wire n3639;wire n3640;wire n3641;wire n3642;wire n3643;wire n3644;wire n3645;wire n3646;wire n3647;wire n3648;wire n3649;wire n3650;wire n3651;wire n3652;wire n3653;wire n3654;wire n3655;wire n3656;wire n3657;wire n3658;wire n3659;wire n3660;wire n3661;wire n3662;wire n3663;wire n3664;wire n3665;wire n3666;wire n3667;wire n3668;wire n3669;wire n3670;wire n3671;wire n3672;wire n3673;wire n3674;wire n3675;wire n3676;wire n3677;wire n3678;wire n3679;wire n3680;wire n3681;wire n3682;wire n3683;wire n3684;wire n3685;wire n3686;wire n3687;wire n3688;wire n3689;wire n3690;wire n3691;wire n3692;wire n3693;wire n3694;wire n3695;wire n3696;wire n3697;wire n3698;wire n3699;wire n3700;wire n3701;wire n3702;wire n3703;wire n3704;wire n3705;wire n3706;wire n3707;wire n3708;wire n3709;wire n3710;wire n3711;wire n3712;wire n3713;wire n3714;wire n3715;wire n3716;wire n3717;wire n3718;wire n3719;wire n3720;wire n3721;wire n3722;wire n3723;wire n3724;wire n3725;wire n3726;wire n3727;wire n3728;wire n3729;wire n3730;wire n3731;wire n3732;wire n3733;wire n3734;wire n3735;wire n3736;wire n3737;wire n3738;wire n3739;wire n3740;wire n3741;wire n3742;wire n3743;wire n3744;wire n3745;wire n3746;wire n3747;wire n3748;wire n3749;wire n3750;wire n3751;wire n3752;wire n3753;wire n3754;wire n3755;wire n3756;wire n3757;wire n3758;wire n3759;wire n3760;wire n3761;wire n3762;wire n3763;wire n3764;wire n3765;wire n3766;wire n3767;wire n3768;wire n3769;wire n3770;wire n3771;wire n3772;wire n3773;wire n3774;wire n3775;wire n3776;wire n3777;wire n3778;wire n3779;wire n3780;wire n3781;wire n3782;wire n3783;wire n3784;wire n3785;wire n3786;wire n3787;wire n3788;wire n3789;wire n3790;wire n3791;wire n3792;wire n3793;wire n3794;wire n3795;wire n3796;wire n3797;wire n3798;wire n3799;wire n3800;wire n3801;wire n3802;wire n3803;wire n3804;wire n3805;wire n3806;wire n3807;wire n3808;wire n3809;wire n3810;wire n3811;wire n3812;wire n3813;wire n3814;wire n3815;wire n3816;wire n3817;wire n3818;wire n3819;wire n3820;wire n3821;wire n3822;wire n3823;wire n3824;wire n3825;wire n3826;wire n3827;wire n3828;wire n3829;wire n3830;wire n3831;wire n3832;wire n3833;wire n3834;wire n3835;wire n3836;wire n3837;wire n3838;wire n3839;wire n3840;wire n3841;wire n3842;wire n3843;wire n3844;wire n3845;wire n3846;wire n3847;wire n3848;wire n3849;wire n3850;wire n3851;wire n3852;wire n3853;wire n3854;wire n3855;wire n3856;wire n3857;wire n3858;wire n3859;wire n3860;wire n3861;wire n3862;wire n3863;wire n3864;wire n3865;wire n3866;wire n3867;wire n3868;wire n3869;wire n3870;wire n3871;wire n3872;wire n3873;wire n3874;wire n3875;wire n3876;wire n3877;wire n3878;wire n3879;wire n3880;wire n3881;wire n3882;wire n3883;wire n3884;wire n3885;wire n3886;wire n3887;wire n3888;wire n3889;wire n3890;wire n3891;wire n3892;wire n3893;wire n3894;wire n3895;wire n3896;wire n3897;wire n3898;wire n3899;wire n3900;wire n3901;wire n3902;wire n3903;wire n3904;wire n3905;wire n3906;wire n3907;wire n3908;wire n3909;wire n3910;wire n3911;wire n3912;wire n3913;wire n3914;wire n3915;wire n3916;wire n3917;wire n3918;wire n3919;wire n3920;wire n3921;wire n3922;wire n3923;wire n3924;wire n3925;wire n3926;wire n3927;wire n3928;wire n3929;wire n3930;wire n3931;wire n3932;wire n3933;wire n3934;wire n3935;wire n3936;wire n3937;wire n3938;wire n3939;wire n3940;wire n3941;wire n3942;wire n3943;wire n3944;wire n3945;wire n3946;wire n3947;wire n3948;wire n3949;wire n3950;wire n3951;wire n3952;wire n3953;wire n3954;wire n3955;wire n3956;wire n3957;wire n3958;wire n3959;wire n3960;wire n3961;wire n3962;wire n3963;wire n3964;wire n3965;wire n3966;wire n3967;wire n3968;wire n3969;wire n3970;wire n3971;wire n3972;wire n3973;wire n3974;wire n3975;wire n3976;wire n3977;wire n3978;wire n3979;wire n3980;wire n3981;wire n3982;wire n3983;wire n3984;wire n3985;wire n3986;wire n3987;wire n3988;wire n3989;wire n3990;wire n3991;wire n3992;wire n3993;wire n3994;wire n3995;wire n3996;wire n3997;wire n3998;wire n3999;wire n4000;wire n4001;wire n4002;wire n4003;wire n4004;wire n4005;wire n4006;wire n4007;wire n4008;wire n4009;wire n4010;wire n4011;wire n4012;wire n4013;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n133,
    n23
  );


  not
  g1
  (
    n104,
    n27
  );


  not
  g2
  (
    n82,
    n11
  );


  buf
  g3
  (
    n100,
    n12
  );


  buf
  g4
  (
    n40,
    n1
  );


  not
  g5
  (
    n66,
    n13
  );


  buf
  g6
  (
    n38,
    n10
  );


  buf
  g7
  (
    n111,
    n8
  );


  buf
  g8
  (
    n34,
    n21
  );


  buf
  g9
  (
    n139,
    n26
  );


  buf
  g10
  (
    n36,
    n5
  );


  not
  g11
  (
    n84,
    n3
  );


  buf
  g12
  (
    n49,
    n20
  );


  buf
  g13
  (
    n65,
    n4
  );


  not
  g14
  (
    n144,
    n25
  );


  not
  g15
  (
    n59,
    n14
  );


  not
  g16
  (
    n113,
    n7
  );


  buf
  g17
  (
    n126,
    n8
  );


  buf
  g18
  (
    n138,
    n2
  );


  not
  g19
  (
    n122,
    n23
  );


  buf
  g20
  (
    n117,
    n21
  );


  not
  g21
  (
    n78,
    n27
  );


  buf
  g22
  (
    n55,
    n24
  );


  not
  g23
  (
    n119,
    n7
  );


  buf
  g24
  (
    n115,
    n1
  );


  not
  g25
  (
    n60,
    n24
  );


  buf
  g26
  (
    n44,
    n1
  );


  buf
  g27
  (
    n64,
    n2
  );


  not
  g28
  (
    n103,
    n18
  );


  not
  g29
  (
    n128,
    n6
  );


  buf
  g30
  (
    n109,
    n28
  );


  buf
  g31
  (
    n54,
    n4
  );


  buf
  g32
  (
    n63,
    n23
  );


  not
  g33
  (
    n43,
    n28
  );


  not
  g34
  (
    n123,
    n28
  );


  buf
  g35
  (
    n107,
    n19
  );


  buf
  g36
  (
    n85,
    n6
  );


  buf
  g37
  (
    n106,
    n10
  );


  buf
  g38
  (
    n86,
    n17
  );


  not
  g39
  (
    n71,
    n16
  );


  not
  g40
  (
    n70,
    n17
  );


  not
  g41
  (
    n50,
    n9
  );


  buf
  g42
  (
    n80,
    n7
  );


  not
  g43
  (
    n95,
    n14
  );


  buf
  g44
  (
    n125,
    n12
  );


  not
  g45
  (
    n62,
    n29
  );


  buf
  g46
  (
    n94,
    n25
  );


  not
  g47
  (
    n68,
    n3
  );


  not
  g48
  (
    n33,
    n23
  );


  not
  g49
  (
    n48,
    n11
  );


  not
  g50
  (
    n47,
    n16
  );


  not
  g51
  (
    n130,
    n21
  );


  buf
  g52
  (
    n92,
    n9
  );


  not
  g53
  (
    n136,
    n24
  );


  buf
  g54
  (
    n46,
    n11
  );


  buf
  g55
  (
    n114,
    n20
  );


  not
  g56
  (
    n69,
    n14
  );


  buf
  g57
  (
    n77,
    n10
  );


  not
  g58
  (
    n98,
    n17
  );


  not
  g59
  (
    n35,
    n2
  );


  not
  g60
  (
    n140,
    n19
  );


  not
  g61
  (
    n121,
    n5
  );


  buf
  g62
  (
    n116,
    n5
  );


  buf
  g63
  (
    n89,
    n8
  );


  buf
  g64
  (
    n90,
    n22
  );


  buf
  g65
  (
    n131,
    n15
  );


  not
  g66
  (
    n53,
    n12
  );


  not
  g67
  (
    n52,
    n26
  );


  not
  g68
  (
    n112,
    n18
  );


  buf
  g69
  (
    n37,
    n1
  );


  buf
  g70
  (
    n45,
    n9
  );


  buf
  g71
  (
    n135,
    n15
  );


  buf
  g72
  (
    n58,
    n6
  );


  not
  g73
  (
    n51,
    n17
  );


  buf
  g74
  (
    n97,
    n28
  );


  not
  g75
  (
    n132,
    n16
  );


  not
  g76
  (
    n137,
    n4
  );


  buf
  g77
  (
    n141,
    n12
  );


  buf
  g78
  (
    n105,
    n29
  );


  buf
  g79
  (
    n75,
    n9
  );


  buf
  g80
  (
    n129,
    n6
  );


  buf
  g81
  (
    n143,
    n27
  );


  buf
  g82
  (
    n61,
    n18
  );


  not
  g83
  (
    n41,
    n10
  );


  buf
  g84
  (
    n146,
    n3
  );


  buf
  g85
  (
    n118,
    n22
  );


  not
  g86
  (
    n81,
    n20
  );


  buf
  g87
  (
    n96,
    n11
  );


  not
  g88
  (
    n87,
    n18
  );


  buf
  g89
  (
    n101,
    n14
  );


  buf
  g90
  (
    n83,
    n27
  );


  buf
  g91
  (
    n67,
    n15
  );


  not
  g92
  (
    n57,
    n24
  );


  buf
  g93
  (
    n93,
    n8
  );


  buf
  g94
  (
    n73,
    n19
  );


  buf
  g95
  (
    n76,
    n20
  );


  buf
  g96
  (
    n91,
    n22
  );


  buf
  g97
  (
    n79,
    n16
  );


  buf
  g98
  (
    n102,
    n13
  );


  not
  g99
  (
    n42,
    n19
  );


  buf
  g100
  (
    n134,
    n3
  );


  not
  g101
  (
    n88,
    n26
  );


  not
  g102
  (
    n99,
    n25
  );


  buf
  g103
  (
    n127,
    n2
  );


  buf
  g104
  (
    n142,
    n22
  );


  not
  g105
  (
    n120,
    n26
  );


  not
  g106
  (
    n124,
    n13
  );


  not
  g107
  (
    n108,
    n5
  );


  buf
  g108
  (
    n74,
    n15
  );


  not
  g109
  (
    n72,
    n25
  );


  buf
  g110
  (
    n56,
    n13
  );


  not
  g111
  (
    n110,
    n21
  );


  buf
  g112
  (
    n145,
    n7
  );


  buf
  g113
  (
    n39,
    n4
  );


  buf
  g114
  (
    n425,
    n115
  );


  not
  g115
  (
    n489,
    n48
  );


  not
  g116
  (
    n152,
    n98
  );


  not
  g117
  (
    n276,
    n133
  );


  not
  g118
  (
    n217,
    n33
  );


  buf
  g119
  (
    n340,
    n107
  );


  buf
  g120
  (
    n428,
    n39
  );


  buf
  g121
  (
    n474,
    n41
  );


  not
  g122
  (
    n297,
    n131
  );


  not
  g123
  (
    n374,
    n92
  );


  not
  g124
  (
    n324,
    n104
  );


  not
  g125
  (
    n499,
    n38
  );


  buf
  g126
  (
    n481,
    n109
  );


  buf
  g127
  (
    n422,
    n134
  );


  buf
  g128
  (
    n375,
    n63
  );


  not
  g129
  (
    n345,
    n70
  );


  not
  g130
  (
    n326,
    n77
  );


  buf
  g131
  (
    n407,
    n63
  );


  not
  g132
  (
    n284,
    n53
  );


  not
  g133
  (
    n336,
    n86
  );


  buf
  g134
  (
    n164,
    n110
  );


  buf
  g135
  (
    n175,
    n137
  );


  not
  g136
  (
    n271,
    n125
  );


  buf
  g137
  (
    n313,
    n109
  );


  buf
  g138
  (
    n494,
    n69
  );


  buf
  g139
  (
    n317,
    n127
  );


  buf
  g140
  (
    n495,
    n40
  );


  buf
  g141
  (
    n200,
    n141
  );


  buf
  g142
  (
    n176,
    n111
  );


  buf
  g143
  (
    n258,
    n100
  );


  buf
  g144
  (
    n199,
    n136
  );


  not
  g145
  (
    n268,
    n41
  );


  not
  g146
  (
    n372,
    n39
  );


  buf
  g147
  (
    n437,
    n128
  );


  not
  g148
  (
    n201,
    n77
  );


  buf
  g149
  (
    n150,
    n131
  );


  not
  g150
  (
    n177,
    n37
  );


  not
  g151
  (
    n490,
    n145
  );


  buf
  g152
  (
    n212,
    n100
  );


  not
  g153
  (
    n189,
    n103
  );


  buf
  g154
  (
    n487,
    n114
  );


  buf
  g155
  (
    n230,
    n117
  );


  buf
  g156
  (
    n445,
    n59
  );


  not
  g157
  (
    n251,
    n58
  );


  not
  g158
  (
    n391,
    n146
  );


  not
  g159
  (
    n226,
    n120
  );


  not
  g160
  (
    n392,
    n89
  );


  buf
  g161
  (
    n298,
    n81
  );


  buf
  g162
  (
    n309,
    n119
  );


  buf
  g163
  (
    n304,
    n61
  );


  not
  g164
  (
    n224,
    n136
  );


  not
  g165
  (
    n486,
    n137
  );


  buf
  g166
  (
    n332,
    n102
  );


  buf
  g167
  (
    n368,
    n78
  );


  not
  g168
  (
    n412,
    n85
  );


  not
  g169
  (
    n341,
    n53
  );


  not
  g170
  (
    n496,
    n37
  );


  buf
  g171
  (
    n397,
    n97
  );


  not
  g172
  (
    n352,
    n50
  );


  not
  g173
  (
    n254,
    n40
  );


  not
  g174
  (
    n315,
    n136
  );


  not
  g175
  (
    n156,
    n92
  );


  not
  g176
  (
    n167,
    n130
  );


  not
  g177
  (
    n381,
    n45
  );


  not
  g178
  (
    n196,
    n45
  );


  not
  g179
  (
    n311,
    n52
  );


  buf
  g180
  (
    n447,
    n127
  );


  buf
  g181
  (
    n228,
    n114
  );


  not
  g182
  (
    n274,
    n133
  );


  buf
  g183
  (
    n163,
    n94
  );


  buf
  g184
  (
    n371,
    n54
  );


  buf
  g185
  (
    n299,
    n74
  );


  not
  g186
  (
    n373,
    n39
  );


  not
  g187
  (
    n263,
    n103
  );


  not
  g188
  (
    n294,
    n64
  );


  not
  g189
  (
    n367,
    n60
  );


  buf
  g190
  (
    n168,
    n135
  );


  not
  g191
  (
    n355,
    n135
  );


  not
  g192
  (
    n227,
    n113
  );


  buf
  g193
  (
    n148,
    n49
  );


  not
  g194
  (
    n248,
    n47
  );


  not
  g195
  (
    n151,
    n29
  );


  buf
  g196
  (
    n153,
    n76
  );


  not
  g197
  (
    n165,
    n142
  );


  buf
  g198
  (
    n443,
    n107
  );


  not
  g199
  (
    n436,
    n38
  );


  buf
  g200
  (
    n300,
    n44
  );


  buf
  g201
  (
    n270,
    n45
  );


  buf
  g202
  (
    n488,
    n139
  );


  not
  g203
  (
    n213,
    n54
  );


  not
  g204
  (
    n416,
    n121
  );


  buf
  g205
  (
    n361,
    n129
  );


  buf
  g206
  (
    n190,
    n135
  );


  buf
  g207
  (
    n158,
    n49
  );


  not
  g208
  (
    n203,
    n96
  );


  not
  g209
  (
    n380,
    n70
  );


  buf
  g210
  (
    n257,
    n84
  );


  not
  g211
  (
    n262,
    n97
  );


  not
  g212
  (
    n386,
    n94
  );


  buf
  g213
  (
    n245,
    n79
  );


  buf
  g214
  (
    n387,
    n132
  );


  buf
  g215
  (
    n344,
    n139
  );


  buf
  g216
  (
    n218,
    n77
  );


  not
  g217
  (
    n384,
    n93
  );


  buf
  g218
  (
    n316,
    n46
  );


  buf
  g219
  (
    n382,
    n124
  );


  not
  g220
  (
    n467,
    n141
  );


  not
  g221
  (
    n348,
    n42
  );


  buf
  g222
  (
    n255,
    n63
  );


  buf
  g223
  (
    n149,
    n112
  );


  not
  g224
  (
    n339,
    n66
  );


  not
  g225
  (
    n264,
    n53
  );


  not
  g226
  (
    n337,
    n78
  );


  buf
  g227
  (
    n184,
    n84
  );


  not
  g228
  (
    n356,
    n50
  );


  buf
  g229
  (
    n259,
    n143
  );


  not
  g230
  (
    n272,
    n55
  );


  not
  g231
  (
    n232,
    n141
  );


  not
  g232
  (
    n308,
    n46
  );


  not
  g233
  (
    n191,
    n112
  );


  buf
  g234
  (
    n266,
    n40
  );


  not
  g235
  (
    n281,
    n90
  );


  buf
  g236
  (
    n415,
    n84
  );


  buf
  g237
  (
    n208,
    n58
  );


  buf
  g238
  (
    n484,
    n142
  );


  buf
  g239
  (
    n478,
    n126
  );


  not
  g240
  (
    n362,
    n115
  );


  not
  g241
  (
    n430,
    n115
  );


  not
  g242
  (
    n358,
    n74
  );


  not
  g243
  (
    n314,
    n71
  );


  not
  g244
  (
    n366,
    n93
  );


  not
  g245
  (
    n461,
    n64
  );


  not
  g246
  (
    n243,
    n103
  );


  not
  g247
  (
    n222,
    n56
  );


  not
  g248
  (
    n347,
    n82
  );


  buf
  g249
  (
    n493,
    n114
  );


  not
  g250
  (
    n231,
    n92
  );


  not
  g251
  (
    n290,
    n118
  );


  buf
  g252
  (
    n498,
    n112
  );


  buf
  g253
  (
    n477,
    n125
  );


  not
  g254
  (
    n179,
    n93
  );


  buf
  g255
  (
    n390,
    n33
  );


  buf
  g256
  (
    n157,
    n123
  );


  not
  g257
  (
    n269,
    n78
  );


  buf
  g258
  (
    n301,
    n67
  );


  buf
  g259
  (
    n174,
    n51
  );


  not
  g260
  (
    n320,
    n115
  );


  not
  g261
  (
    n160,
    n128
  );


  not
  g262
  (
    n240,
    n113
  );


  buf
  g263
  (
    n460,
    n73
  );


  not
  g264
  (
    n349,
    n57
  );


  not
  g265
  (
    n406,
    n124
  );


  buf
  g266
  (
    n473,
    n95
  );


  buf
  g267
  (
    n480,
    n61
  );


  buf
  g268
  (
    n210,
    n46
  );


  not
  g269
  (
    n220,
    n121
  );


  buf
  g270
  (
    n318,
    n66
  );


  buf
  g271
  (
    n171,
    n145
  );


  buf
  g272
  (
    n395,
    n123
  );


  buf
  g273
  (
    n396,
    n41
  );


  not
  g274
  (
    n181,
    n71
  );


  buf
  g275
  (
    n260,
    n139
  );


  buf
  g276
  (
    n154,
    n125
  );


  not
  g277
  (
    n379,
    n123
  );


  not
  g278
  (
    n328,
    n46
  );


  not
  g279
  (
    n286,
    n138
  );


  not
  g280
  (
    n334,
    n66
  );


  buf
  g281
  (
    n434,
    n54
  );


  buf
  g282
  (
    n305,
    n66
  );


  not
  g283
  (
    n369,
    n83
  );


  not
  g284
  (
    n161,
    n91
  );


  buf
  g285
  (
    n435,
    n129
  );


  buf
  g286
  (
    n453,
    n107
  );


  not
  g287
  (
    n408,
    n87
  );


  not
  g288
  (
    n424,
    n42
  );


  buf
  g289
  (
    n197,
    n59
  );


  not
  g290
  (
    n330,
    n78
  );


  not
  g291
  (
    n198,
    n101
  );


  buf
  g292
  (
    n492,
    n34
  );


  not
  g293
  (
    n187,
    n140
  );


  buf
  g294
  (
    n239,
    n47
  );


  buf
  g295
  (
    n289,
    n89
  );


  not
  g296
  (
    n433,
    n98
  );


  not
  g297
  (
    n456,
    n43
  );


  buf
  g298
  (
    n469,
    n83
  );


  buf
  g299
  (
    n223,
    n44
  );


  buf
  g300
  (
    n458,
    n136
  );


  not
  g301
  (
    n354,
    n43
  );


  buf
  g302
  (
    n182,
    n85
  );


  not
  g303
  (
    n173,
    n110
  );


  not
  g304
  (
    n439,
    n81
  );


  not
  g305
  (
    n421,
    n55
  );


  not
  g306
  (
    n296,
    n44
  );


  not
  g307
  (
    n327,
    n58
  );


  not
  g308
  (
    n357,
    n102
  );


  buf
  g309
  (
    n265,
    n121
  );


  not
  g310
  (
    n398,
    n144
  );


  not
  g311
  (
    n429,
    n93
  );


  buf
  g312
  (
    n470,
    n81
  );


  not
  g313
  (
    n393,
    n128
  );


  not
  g314
  (
    n147,
    n35
  );


  not
  g315
  (
    n476,
    n81
  );


  not
  g316
  (
    n359,
    n108
  );


  not
  g317
  (
    n244,
    n51
  );


  not
  g318
  (
    n394,
    n108
  );


  buf
  g319
  (
    n225,
    n102
  );


  not
  g320
  (
    n186,
    n72
  );


  not
  g321
  (
    n440,
    n123
  );


  not
  g322
  (
    n388,
    n36
  );


  not
  g323
  (
    n293,
    n131
  );


  not
  g324
  (
    n295,
    n139
  );


  buf
  g325
  (
    n465,
    n77
  );


  not
  g326
  (
    n485,
    n87
  );


  buf
  g327
  (
    n275,
    n60
  );


  buf
  g328
  (
    n180,
    n88
  );


  buf
  g329
  (
    n249,
    n99
  );


  not
  g330
  (
    n472,
    n48
  );


  not
  g331
  (
    n221,
    n119
  );


  buf
  g332
  (
    n491,
    n36
  );


  not
  g333
  (
    n235,
    n59
  );


  buf
  g334
  (
    n162,
    n130
  );


  buf
  g335
  (
    n463,
    n140
  );


  not
  g336
  (
    n242,
    n135
  );


  buf
  g337
  (
    n444,
    n72
  );


  not
  g338
  (
    n455,
    n42
  );


  not
  g339
  (
    n418,
    n68
  );


  not
  g340
  (
    n457,
    n60
  );


  not
  g341
  (
    n400,
    n88
  );


  not
  g342
  (
    n307,
    n122
  );


  buf
  g343
  (
    n404,
    n51
  );


  not
  g344
  (
    n172,
    n144
  );


  not
  g345
  (
    n338,
    n83
  );


  not
  g346
  (
    n178,
    n88
  );


  buf
  g347
  (
    n449,
    n49
  );


  not
  g348
  (
    n287,
    n76
  );


  not
  g349
  (
    n383,
    n36
  );


  buf
  g350
  (
    n282,
    n34
  );


  not
  g351
  (
    n432,
    n65
  );


  not
  g352
  (
    n376,
    n117
  );


  buf
  g353
  (
    n363,
    n120
  );


  buf
  g354
  (
    n331,
    n100
  );


  buf
  g355
  (
    n323,
    n35
  );


  buf
  g356
  (
    n419,
    n126
  );


  buf
  g357
  (
    n319,
    n90
  );


  buf
  g358
  (
    n216,
    n69
  );


  not
  g359
  (
    n325,
    n39
  );


  buf
  g360
  (
    n303,
    n52
  );


  not
  g361
  (
    n399,
    n98
  );


  buf
  g362
  (
    n378,
    n100
  );


  not
  g363
  (
    n291,
    n104
  );


  not
  g364
  (
    n497,
    n137
  );


  not
  g365
  (
    n267,
    n143
  );


  not
  g366
  (
    n464,
    n128
  );


  not
  g367
  (
    n310,
    n85
  );


  not
  g368
  (
    n285,
    n57
  );


  buf
  g369
  (
    n402,
    n41
  );


  not
  g370
  (
    n219,
    n64
  );


  not
  g371
  (
    n483,
    n47
  );


  not
  g372
  (
    n401,
    n140
  );


  buf
  g373
  (
    n370,
    n64
  );


  not
  g374
  (
    n280,
    n109
  );


  not
  g375
  (
    n389,
    n106
  );


  not
  g376
  (
    n364,
    n145
  );


  buf
  g377
  (
    n322,
    n122
  );


  not
  g378
  (
    n482,
    n65
  );


  buf
  g379
  (
    n170,
    n105
  );


  buf
  g380
  (
    n195,
    n143
  );


  buf
  g381
  (
    n417,
    n102
  );


  not
  g382
  (
    n194,
    n103
  );


  buf
  g383
  (
    n377,
    n49
  );


  buf
  g384
  (
    n204,
    n55
  );


  buf
  g385
  (
    n188,
    n91
  );


  buf
  g386
  (
    n350,
    n99
  );


  buf
  g387
  (
    n253,
    n108
  );


  not
  g388
  (
    n214,
    n86
  );


  buf
  g389
  (
    n343,
    n62
  );


  not
  g390
  (
    n209,
    n43
  );


  buf
  g391
  (
    n360,
    n84
  );


  buf
  g392
  (
    n306,
    n73
  );


  not
  g393
  (
    n252,
    n101
  );


  buf
  g394
  (
    n312,
    n80
  );


  buf
  g395
  (
    n420,
    n96
  );


  buf
  g396
  (
    n169,
    n56
  );


  not
  g397
  (
    n475,
    n76
  );


  buf
  g398
  (
    n468,
    n109
  );


  not
  g399
  (
    n205,
    n70
  );


  buf
  g400
  (
    n385,
    n33
  );


  buf
  g401
  (
    n450,
    n111
  );


  not
  g402
  (
    n155,
    n70
  );


  buf
  g403
  (
    n166,
    n131
  );


  not
  g404
  (
    n441,
    n134
  );


  not
  g405
  (
    n193,
    n107
  );


  buf
  g406
  (
    n448,
    n76
  );


  buf
  g407
  (
    n283,
    n47
  );


  buf
  g408
  (
    n241,
    n111
  );


  not
  g409
  (
    n466,
    n130
  );


  not
  g410
  (
    n335,
    n90
  );


  not
  g411
  (
    n454,
    n99
  );


  not
  g412
  (
    n438,
    n132
  );


  buf
  g413
  (
    n159,
    n105
  );


  buf
  g414
  (
    n446,
    n44
  );


  not
  g415
  (
    n215,
    n67
  );


  buf
  g416
  (
    n403,
    n105
  );


  buf
  g417
  (
    n471,
    n120
  );


  buf
  g418
  (
    n273,
    n62
  );


  buf
  g419
  (
    n353,
    n120
  );


  not
  g420
  (
    n250,
    n94
  );


  buf
  g421
  (
    n321,
    n112
  );


  not
  g422
  (
    n414,
    n59
  );


  not
  g423
  (
    n452,
    n117
  );


  not
  g424
  (
    n236,
    n34
  );


  not
  g425
  (
    n292,
    n113
  );


  buf
  g426
  (
    n426,
    n116
  );


  buf
  g427
  (
    n423,
    n35
  );


  buf
  g428
  (
    n183,
    n40
  );


  buf
  g429
  (
    n238,
    n116
  );


  not
  g430
  (
    n211,
    n113
  );


  buf
  g431
  (
    n479,
    n129
  );


  buf
  g432
  (
    n410,
    n67
  );


  nor
  g433
  (
    n234,
    n116,
    n119,
    n54,
    n133
  );


  nor
  g434
  (
    n427,
    n72,
    n96,
    n138,
    n122
  );


  and
  g435
  (
    n185,
    n56,
    n129,
    n36,
    n34
  );


  and
  g436
  (
    n462,
    n57,
    n43,
    n61,
    n138
  );


  and
  g437
  (
    n261,
    n55,
    n63,
    n82,
    n62
  );


  or
  g438
  (
    n431,
    n74,
    n48,
    n134,
    n79
  );


  or
  g439
  (
    n278,
    n106,
    n80,
    n137,
    n119
  );


  nand
  g440
  (
    n288,
    n37,
    n50,
    n79,
    n65
  );


  or
  g441
  (
    n413,
    n88,
    n132,
    n52,
    n122
  );


  or
  g442
  (
    n247,
    n69,
    n50,
    n71,
    n29
  );


  and
  g443
  (
    n229,
    n98,
    n118,
    n130,
    n45
  );


  or
  g444
  (
    n333,
    n68,
    n96,
    n141,
    n62
  );


  and
  g445
  (
    n351,
    n110,
    n86,
    n95,
    n80
  );


  xnor
  g446
  (
    n451,
    n138,
    n53,
    n33,
    n97
  );


  or
  g447
  (
    n206,
    n48,
    n73,
    n91,
    n75
  );


  nand
  g448
  (
    n442,
    n121,
    n124,
    n72,
    n142
  );


  or
  g449
  (
    n237,
    n126,
    n124,
    n105,
    n82
  );


  or
  g450
  (
    n233,
    n106,
    n133,
    n74,
    n132
  );


  xor
  g451
  (
    n202,
    n75,
    n127,
    n68,
    n140
  );


  and
  g452
  (
    n277,
    n106,
    n101,
    n116,
    n111
  );


  and
  g453
  (
    n192,
    n73,
    n95,
    n90,
    n57
  );


  xor
  g454
  (
    n411,
    n117,
    n51,
    n143,
    n87
  );


  or
  g455
  (
    n329,
    n61,
    n125,
    n145,
    n82
  );


  or
  g456
  (
    n207,
    n58,
    n83,
    n56,
    n142
  );


  nor
  g457
  (
    n302,
    n38,
    n79,
    n60,
    n99
  );


  xnor
  g458
  (
    n346,
    n91,
    n38,
    n75,
    n71
  );


  nor
  g459
  (
    n365,
    n104,
    n101,
    n127,
    n144
  );


  and
  g460
  (
    n459,
    n86,
    n52,
    n65,
    n134
  );


  or
  g461
  (
    n256,
    n89,
    n114,
    n67,
    n35
  );


  xor
  g462
  (
    n405,
    n108,
    n89,
    n85,
    n75
  );


  and
  g463
  (
    n409,
    n97,
    n118,
    n94,
    n104
  );


  nor
  g464
  (
    n342,
    n95,
    n37,
    n126,
    n118
  );


  and
  g465
  (
    n279,
    n69,
    n68,
    n80,
    n42
  );


  xnor
  g466
  (
    n246,
    n92,
    n110,
    n144,
    n87
  );


  and
  g467
  (
    n515,
    n156,
    n160,
    n163
  );


  or
  g468
  (
    n508,
    n152,
    n154,
    n158,
    n161
  );


  nand
  g469
  (
    n503,
    n151,
    n154,
    n161,
    n155
  );


  xnor
  g470
  (
    n505,
    n148,
    n155,
    n159,
    n162
  );


  xor
  g471
  (
    n511,
    n156,
    n153,
    n149,
    n155
  );


  nand
  g472
  (
    n513,
    n151,
    n154,
    n163,
    n153
  );


  or
  g473
  (
    n504,
    n157,
    n158,
    n147
  );


  and
  g474
  (
    n501,
    n149,
    n147,
    n150,
    n158
  );


  xor
  g475
  (
    n506,
    n162,
    n152,
    n149,
    n159
  );


  and
  g476
  (
    n509,
    n148,
    n157,
    n153,
    n156
  );


  nand
  g477
  (
    n500,
    n159,
    n162,
    n160,
    n151
  );


  or
  g478
  (
    n514,
    n148,
    n162,
    n161,
    n150
  );


  and
  g479
  (
    n507,
    n157,
    n150,
    n154,
    n153
  );


  nand
  g480
  (
    n502,
    n159,
    n160,
    n150,
    n149
  );


  xor
  g481
  (
    n510,
    n151,
    n157,
    n152,
    n158
  );


  nor
  g482
  (
    n512,
    n152,
    n156,
    n155,
    n161
  );


  buf
  g483
  (
    n516,
    n500
  );


  buf
  g484
  (
    n517,
    n516
  );


  buf
  g485
  (
    n518,
    n517
  );


  not
  g486
  (
    n519,
    n518
  );


  buf
  g487
  (
    n522,
    n519
  );


  not
  g488
  (
    n520,
    n519
  );


  not
  g489
  (
    n521,
    n519
  );


  not
  g490
  (
    n523,
    n519
  );


  and
  g491
  (
    n525,
    n522,
    n522,
    n520,
    n521
  );


  or
  g492
  (
    n529,
    n522,
    n520,
    n517,
    n165
  );


  and
  g493
  (
    n526,
    n163,
    n163,
    n164,
    n520
  );


  and
  g494
  (
    n524,
    n521,
    n522,
    n165,
    n164
  );


  xnor
  g495
  (
    n528,
    n523,
    n165,
    n521,
    n164
  );


  xor
  g496
  (
    n527,
    n517,
    n164,
    n521,
    n520
  );


  nor
  g497
  (
    n534,
    n527,
    n516,
    n166,
    n529
  );


  nor
  g498
  (
    n532,
    n168,
    n168,
    n525,
    n167
  );


  nand
  g499
  (
    n533,
    n167,
    n524,
    n528,
    n527
  );


  xor
  g500
  (
    n531,
    n523,
    n167,
    n168,
    n527
  );


  and
  g501
  (
    n538,
    n516,
    n166,
    n523
  );


  nor
  g502
  (
    n536,
    n165,
    n525,
    n526,
    n528
  );


  nand
  g503
  (
    n537,
    n30,
    n167,
    n526,
    n529
  );


  or
  g504
  (
    n535,
    n168,
    n517,
    n525,
    n529
  );


  or
  g505
  (
    n530,
    n528,
    n523,
    n166,
    n526
  );


  not
  g506
  (
    n540,
    n530
  );


  and
  g507
  (
    n539,
    n531,
    n530
  );


  not
  g508
  (
    n542,
    n540
  );


  buf
  g509
  (
    n543,
    n539
  );


  not
  g510
  (
    n541,
    n539
  );


  not
  g511
  (
    n545,
    n539
  );


  not
  g512
  (
    n544,
    n539
  );


  nor
  g513
  (
    n549,
    n541,
    n544,
    n543
  );


  nand
  g514
  (
    n548,
    n30,
    n542,
    n544
  );


  nand
  g515
  (
    n547,
    n542,
    n541
  );


  nand
  g516
  (
    n546,
    n543,
    n543,
    n542,
    n544
  );


  buf
  g517
  (
    n553,
    n548
  );


  buf
  g518
  (
    n552,
    n546
  );


  buf
  g519
  (
    n550,
    n546
  );


  buf
  g520
  (
    n557,
    n549
  );


  not
  g521
  (
    n554,
    n547
  );


  buf
  g522
  (
    n555,
    n546
  );


  not
  g523
  (
    n560,
    n549
  );


  not
  g524
  (
    n558,
    n548
  );


  not
  g525
  (
    n556,
    n549
  );


  buf
  g526
  (
    n559,
    n547
  );


  buf
  g527
  (
    n561,
    n547
  );


  buf
  g528
  (
    n551,
    n548
  );


  and
  g529
  (
    n586,
    n192,
    n554,
    n188,
    n178
  );


  xor
  g530
  (
    n599,
    n175,
    n553,
    n183,
    n171
  );


  nand
  g531
  (
    n583,
    n202,
    n203,
    n188,
    n190
  );


  nor
  g532
  (
    n609,
    n169,
    n202,
    n177,
    n199
  );


  nand
  g533
  (
    n594,
    n183,
    n179,
    n187,
    n181
  );


  xor
  g534
  (
    n598,
    n201,
    n195,
    n172,
    n174
  );


  or
  g535
  (
    n605,
    n558,
    n172,
    n190,
    n175
  );


  nand
  g536
  (
    n568,
    n182,
    n551,
    n196,
    n552
  );


  and
  g537
  (
    n597,
    n171,
    n185,
    n201,
    n172
  );


  xnor
  g538
  (
    n590,
    n561,
    n169,
    n559,
    n170
  );


  nor
  g539
  (
    n578,
    n169,
    n204,
    n184,
    n186
  );


  and
  g540
  (
    n607,
    n558,
    n180,
    n200,
    n181
  );


  xnor
  g541
  (
    n565,
    n186,
    n554,
    n561,
    n556
  );


  and
  g542
  (
    n592,
    n176,
    n176,
    n558,
    n191
  );


  nand
  g543
  (
    n601,
    n181,
    n192,
    n173,
    n189
  );


  and
  g544
  (
    n582,
    n204,
    n550,
    n195,
    n177
  );


  xnor
  g545
  (
    n570,
    n176,
    n560,
    n561,
    n559
  );


  xnor
  g546
  (
    n585,
    n553,
    n550,
    n173,
    n202
  );


  and
  g547
  (
    n572,
    n194,
    n191,
    n555,
    n553
  );


  nor
  g548
  (
    n593,
    n560,
    n187,
    n178,
    n179
  );


  and
  g549
  (
    n584,
    n183,
    n180,
    n194,
    n175
  );


  xnor
  g550
  (
    n563,
    n177,
    n170,
    n557,
    n203
  );


  xnor
  g551
  (
    n589,
    n197,
    n178,
    n198,
    n554
  );


  nand
  g552
  (
    n566,
    n551,
    n174,
    n175,
    n189
  );


  xnor
  g553
  (
    n580,
    n557,
    n193,
    n169,
    n190
  );


  nand
  g554
  (
    n569,
    n188,
    n200,
    n182,
    n186
  );


  or
  g555
  (
    n577,
    n558,
    n189,
    n557,
    n201
  );


  xor
  g556
  (
    n591,
    n196,
    n194,
    n197,
    n204
  );


  nor
  g557
  (
    n574,
    n559,
    n196,
    n555,
    n185
  );


  nor
  g558
  (
    n604,
    n198,
    n195,
    n550
  );


  xor
  g559
  (
    n562,
    n198,
    n197,
    n200,
    n552
  );


  xor
  g560
  (
    n581,
    n179,
    n172,
    n184,
    n183
  );


  xor
  g561
  (
    n575,
    n184,
    n190,
    n192,
    n199
  );


  or
  g562
  (
    n603,
    n184,
    n185,
    n196,
    n180
  );


  and
  g563
  (
    n573,
    n191,
    n203,
    n556,
    n174
  );


  nand
  g564
  (
    n571,
    n195,
    n559,
    n552,
    n553
  );


  and
  g565
  (
    n600,
    n198,
    n187,
    n202,
    n185
  );


  nor
  g566
  (
    n567,
    n177,
    n180,
    n174,
    n201
  );


  nand
  g567
  (
    n579,
    n551,
    n555,
    n193,
    n556
  );


  and
  g568
  (
    n596,
    n203,
    n178,
    n176,
    n556
  );


  nand
  g569
  (
    n587,
    n173,
    n193,
    n187,
    n200
  );


  and
  g570
  (
    n602,
    n186,
    n179,
    n192,
    n181
  );


  or
  g571
  (
    n595,
    n194,
    n560,
    n552
  );


  nand
  g572
  (
    n606,
    n554,
    n189,
    n170,
    n171
  );


  nor
  g573
  (
    n608,
    n555,
    n188,
    n193,
    n182
  );


  nand
  g574
  (
    n588,
    n173,
    n199,
    n557,
    n561
  );


  xor
  g575
  (
    n576,
    n551,
    n191,
    n171,
    n199
  );


  and
  g576
  (
    n564,
    n182,
    n197,
    n204,
    n170
  );


  buf
  g577
  (
    n664,
    n595
  );


  not
  g578
  (
    n616,
    n586
  );


  not
  g579
  (
    n699,
    n588
  );


  buf
  g580
  (
    n720,
    n565
  );


  buf
  g581
  (
    n621,
    n583
  );


  not
  g582
  (
    n690,
    n562
  );


  not
  g583
  (
    n721,
    n568
  );


  not
  g584
  (
    n704,
    n601
  );


  buf
  g585
  (
    n733,
    n597
  );


  not
  g586
  (
    n652,
    n580
  );


  not
  g587
  (
    n674,
    n571
  );


  buf
  g588
  (
    n680,
    n580
  );


  buf
  g589
  (
    n613,
    n513
  );


  not
  g590
  (
    n626,
    n509
  );


  not
  g591
  (
    n705,
    n586
  );


  buf
  g592
  (
    n666,
    n567
  );


  buf
  g593
  (
    n646,
    n506
  );


  not
  g594
  (
    n713,
    n577
  );


  buf
  g595
  (
    n678,
    n577
  );


  not
  g596
  (
    n641,
    n577
  );


  not
  g597
  (
    n676,
    n582
  );


  buf
  g598
  (
    n660,
    n605
  );


  not
  g599
  (
    n686,
    n601
  );


  buf
  g600
  (
    n696,
    n586
  );


  not
  g601
  (
    n681,
    n571
  );


  not
  g602
  (
    n724,
    n590
  );


  buf
  g603
  (
    n628,
    n584
  );


  not
  g604
  (
    n706,
    n594
  );


  not
  g605
  (
    n632,
    n606
  );


  not
  g606
  (
    n730,
    n593
  );


  not
  g607
  (
    n619,
    n594
  );


  not
  g608
  (
    n715,
    n585
  );


  buf
  g609
  (
    n645,
    n599
  );


  not
  g610
  (
    n630,
    n602
  );


  not
  g611
  (
    n659,
    n569
  );


  buf
  g612
  (
    n668,
    n583
  );


  not
  g613
  (
    n639,
    n566
  );


  buf
  g614
  (
    n656,
    n569
  );


  buf
  g615
  (
    n643,
    n565
  );


  not
  g616
  (
    n635,
    n576
  );


  buf
  g617
  (
    n732,
    n570
  );


  not
  g618
  (
    n722,
    n587
  );


  buf
  g619
  (
    n672,
    n589
  );


  buf
  g620
  (
    n693,
    n586
  );


  not
  g621
  (
    n687,
    n604
  );


  not
  g622
  (
    n711,
    n601
  );


  not
  g623
  (
    n634,
    n564
  );


  not
  g624
  (
    n633,
    n584
  );


  buf
  g625
  (
    n663,
    n570
  );


  not
  g626
  (
    n682,
    n579
  );


  not
  g627
  (
    n725,
    n591
  );


  not
  g628
  (
    n649,
    n593
  );


  buf
  g629
  (
    n661,
    n580
  );


  buf
  g630
  (
    n677,
    n597
  );


  buf
  g631
  (
    n654,
    n607
  );


  not
  g632
  (
    n618,
    n576
  );


  buf
  g633
  (
    n617,
    n572
  );


  not
  g634
  (
    n665,
    n514
  );


  buf
  g635
  (
    n614,
    n591
  );


  buf
  g636
  (
    n650,
    n503
  );


  not
  g637
  (
    n729,
    n562
  );


  not
  g638
  (
    n636,
    n563
  );


  not
  g639
  (
    n638,
    n563
  );


  buf
  g640
  (
    n651,
    n576
  );


  not
  g641
  (
    n723,
    n564
  );


  buf
  g642
  (
    n710,
    n600
  );


  not
  g643
  (
    n670,
    n578
  );


  not
  g644
  (
    n731,
    n595
  );


  not
  g645
  (
    n727,
    n593
  );


  buf
  g646
  (
    n689,
    n595
  );


  buf
  g647
  (
    n655,
    n574
  );


  buf
  g648
  (
    n648,
    n599
  );


  not
  g649
  (
    n640,
    n596
  );


  not
  g650
  (
    n698,
    n603
  );


  buf
  g651
  (
    n703,
    n531
  );


  buf
  g652
  (
    n673,
    n581
  );


  not
  g653
  (
    n615,
    n591
  );


  buf
  g654
  (
    n700,
    n607
  );


  buf
  g655
  (
    n714,
    n592
  );


  buf
  g656
  (
    n669,
    n585
  );


  not
  g657
  (
    n702,
    n578
  );


  not
  g658
  (
    n712,
    n573
  );


  buf
  g659
  (
    n709,
    n570
  );


  not
  g660
  (
    n691,
    n602
  );


  buf
  g661
  (
    n627,
    n590
  );


  not
  g662
  (
    n695,
    n588
  );


  buf
  g663
  (
    n622,
    n510
  );


  buf
  g664
  (
    n629,
    n567
  );


  buf
  g665
  (
    n620,
    n507
  );


  buf
  g666
  (
    n692,
    n512
  );


  buf
  g667
  (
    n701,
    n597
  );


  not
  g668
  (
    n625,
    n575
  );


  not
  g669
  (
    n657,
    n592
  );


  buf
  g670
  (
    n662,
    n595
  );


  buf
  g671
  (
    n647,
    n501
  );


  not
  g672
  (
    n726,
    n568
  );


  nor
  g673
  (
    n624,
    n598,
    n596,
    n585,
    n566
  );


  and
  g674
  (
    n684,
    n563,
    n504,
    n571,
    n594
  );


  and
  g675
  (
    n667,
    n584,
    n609,
    n565
  );


  xnor
  g676
  (
    n718,
    n598,
    n568,
    n600,
    n572
  );


  nor
  g677
  (
    n623,
    n591,
    n587,
    n575,
    n608
  );


  xor
  g678
  (
    n728,
    n562,
    n587,
    n605,
    n585
  );


  nor
  g679
  (
    n658,
    n605,
    n579,
    n563,
    n578
  );


  or
  g680
  (
    n716,
    n606,
    n568,
    n605,
    n581
  );


  xnor
  g681
  (
    n612,
    n594,
    n590,
    n573,
    n571
  );


  and
  g682
  (
    n685,
    n565,
    n505,
    n502,
    n581
  );


  nand
  g683
  (
    n611,
    n603,
    n572,
    n604,
    n599
  );


  nand
  g684
  (
    n717,
    n608,
    n600,
    n575,
    n602
  );


  xor
  g685
  (
    n679,
    n593,
    n603,
    n592,
    n596
  );


  xor
  g686
  (
    n653,
    n607,
    n607,
    n601,
    n600
  );


  nor
  g687
  (
    n631,
    n597,
    n598,
    n604,
    n582
  );


  nor
  g688
  (
    n697,
    n581,
    n564,
    n570,
    n569
  );


  or
  g689
  (
    n694,
    n562,
    n579,
    n566,
    n602
  );


  xor
  g690
  (
    n675,
    n598,
    n589,
    n604,
    n587
  );


  xnor
  g691
  (
    n688,
    n589,
    n575,
    n574,
    n582
  );


  nand
  g692
  (
    n610,
    n582,
    n567,
    n589,
    n564
  );


  and
  g693
  (
    n708,
    n588,
    n590,
    n508,
    n603
  );


  xnor
  g694
  (
    n644,
    n588,
    n531,
    n583,
    n592
  );


  nor
  g695
  (
    n707,
    n596,
    n569,
    n608
  );


  nor
  g696
  (
    n719,
    n566,
    n578,
    n576,
    n573
  );


  nor
  g697
  (
    n637,
    n609,
    n606,
    n599
  );


  and
  g698
  (
    n642,
    n584,
    n583,
    n580,
    n574
  );


  xor
  g699
  (
    n683,
    n567,
    n609,
    n572,
    n574
  );


  xor
  g700
  (
    n671,
    n573,
    n577,
    n579,
    n511
  );


  buf
  g701
  (
    n775,
    n624
  );


  buf
  g702
  (
    n737,
    n624
  );


  buf
  g703
  (
    n752,
    n622
  );


  buf
  g704
  (
    n791,
    n614
  );


  not
  g705
  (
    n788,
    n620
  );


  buf
  g706
  (
    n773,
    n618
  );


  buf
  g707
  (
    n756,
    n613
  );


  buf
  g708
  (
    n750,
    n619
  );


  buf
  g709
  (
    n792,
    n616
  );


  not
  g710
  (
    n751,
    n612
  );


  not
  g711
  (
    n754,
    n614
  );


  not
  g712
  (
    n741,
    n621
  );


  not
  g713
  (
    n745,
    n615
  );


  buf
  g714
  (
    n736,
    n610
  );


  not
  g715
  (
    n738,
    n611
  );


  not
  g716
  (
    n783,
    n611
  );


  buf
  g717
  (
    n740,
    n617
  );


  buf
  g718
  (
    n744,
    n619
  );


  not
  g719
  (
    n748,
    n617
  );


  buf
  g720
  (
    n774,
    n623
  );


  buf
  g721
  (
    n780,
    n612
  );


  not
  g722
  (
    n766,
    n613
  );


  not
  g723
  (
    n759,
    n620
  );


  not
  g724
  (
    n776,
    n617
  );


  not
  g725
  (
    n755,
    n611
  );


  not
  g726
  (
    n743,
    n623
  );


  not
  g727
  (
    n765,
    n622
  );


  not
  g728
  (
    n735,
    n622
  );


  buf
  g729
  (
    n757,
    n621
  );


  not
  g730
  (
    n781,
    n610
  );


  not
  g731
  (
    n764,
    n610
  );


  buf
  g732
  (
    n763,
    n613
  );


  not
  g733
  (
    n784,
    n612
  );


  not
  g734
  (
    n778,
    n618
  );


  buf
  g735
  (
    n771,
    n622
  );


  not
  g736
  (
    n749,
    n624
  );


  not
  g737
  (
    n785,
    n614
  );


  not
  g738
  (
    n768,
    n615
  );


  buf
  g739
  (
    n762,
    n616
  );


  buf
  g740
  (
    n777,
    n620
  );


  buf
  g741
  (
    n739,
    n615
  );


  buf
  g742
  (
    n753,
    n613
  );


  not
  g743
  (
    n772,
    n623
  );


  buf
  g744
  (
    n746,
    n611
  );


  buf
  g745
  (
    n734,
    n614
  );


  buf
  g746
  (
    n787,
    n616
  );


  buf
  g747
  (
    n769,
    n621
  );


  buf
  g748
  (
    n793,
    n615
  );


  buf
  g749
  (
    n747,
    n621
  );


  not
  g750
  (
    n767,
    n624
  );


  buf
  g751
  (
    n761,
    n619
  );


  buf
  g752
  (
    n758,
    n616
  );


  buf
  g753
  (
    n742,
    n618
  );


  buf
  g754
  (
    n760,
    n617
  );


  buf
  g755
  (
    n789,
    n620
  );


  buf
  g756
  (
    n779,
    n619
  );


  not
  g757
  (
    n790,
    n618
  );


  buf
  g758
  (
    n786,
    n610
  );


  not
  g759
  (
    n782,
    n612
  );


  not
  g760
  (
    n770,
    n623
  );


  buf
  g761
  (
    n918,
    n765
  );


  not
  g762
  (
    n988,
    n705
  );


  buf
  g763
  (
    n902,
    n695
  );


  buf
  g764
  (
    n992,
    n650
  );


  buf
  g765
  (
    n874,
    n745
  );


  buf
  g766
  (
    n834,
    n719
  );


  buf
  g767
  (
    n1006,
    n626
  );


  not
  g768
  (
    n937,
    n747
  );


  buf
  g769
  (
    n839,
    n788
  );


  not
  g770
  (
    n1007,
    n734
  );


  not
  g771
  (
    n982,
    n773
  );


  buf
  g772
  (
    n861,
    n785
  );


  buf
  g773
  (
    n961,
    n626
  );


  buf
  g774
  (
    n821,
    n660
  );


  buf
  g775
  (
    n997,
    n736
  );


  buf
  g776
  (
    n947,
    n689
  );


  not
  g777
  (
    n846,
    n651
  );


  not
  g778
  (
    n919,
    n628
  );


  not
  g779
  (
    n1011,
    n662
  );


  buf
  g780
  (
    n842,
    n787
  );


  not
  g781
  (
    n893,
    n679
  );


  not
  g782
  (
    n930,
    n747
  );


  not
  g783
  (
    n969,
    n745
  );


  not
  g784
  (
    n841,
    n678
  );


  buf
  g785
  (
    n803,
    n772
  );


  buf
  g786
  (
    n940,
    n695
  );


  not
  g787
  (
    n941,
    n750
  );


  not
  g788
  (
    n858,
    n776
  );


  not
  g789
  (
    n876,
    n736
  );


  not
  g790
  (
    n825,
    n637
  );


  not
  g791
  (
    n901,
    n642
  );


  not
  g792
  (
    n807,
    n634
  );


  buf
  g793
  (
    n847,
    n674
  );


  buf
  g794
  (
    n907,
    n727
  );


  not
  g795
  (
    n855,
    n713
  );


  not
  g796
  (
    n826,
    n703
  );


  not
  g797
  (
    n996,
    n713
  );


  buf
  g798
  (
    n1009,
    n750
  );


  buf
  g799
  (
    n921,
    n771
  );


  buf
  g800
  (
    n913,
    n756
  );


  buf
  g801
  (
    n799,
    n704
  );


  buf
  g802
  (
    n1000,
    n715
  );


  not
  g803
  (
    n884,
    n671
  );


  buf
  g804
  (
    n891,
    n741
  );


  buf
  g805
  (
    n990,
    n720
  );


  buf
  g806
  (
    n849,
    n749
  );


  not
  g807
  (
    n833,
    n752
  );


  not
  g808
  (
    n968,
    n668
  );


  not
  g809
  (
    n822,
    n672
  );


  not
  g810
  (
    n868,
    n768
  );


  not
  g811
  (
    n945,
    n685
  );


  not
  g812
  (
    n844,
    n753
  );


  not
  g813
  (
    n1018,
    n725
  );


  buf
  g814
  (
    n854,
    n730
  );


  buf
  g815
  (
    n932,
    n675
  );


  buf
  g816
  (
    n900,
    n700
  );


  not
  g817
  (
    n999,
    n645
  );


  not
  g818
  (
    n828,
    n724
  );


  buf
  g819
  (
    n1026,
    n755
  );


  buf
  g820
  (
    n956,
    n726
  );


  buf
  g821
  (
    n994,
    n694
  );


  buf
  g822
  (
    n811,
    n783
  );


  not
  g823
  (
    n818,
    n670
  );


  buf
  g824
  (
    n963,
    n721
  );


  buf
  g825
  (
    n971,
    n701
  );


  buf
  g826
  (
    n910,
    n694
  );


  not
  g827
  (
    n860,
    n789
  );


  not
  g828
  (
    n960,
    n676
  );


  buf
  g829
  (
    n889,
    n672
  );


  buf
  g830
  (
    n843,
    n773
  );


  not
  g831
  (
    n806,
    n625
  );


  buf
  g832
  (
    n878,
    n713
  );


  buf
  g833
  (
    n829,
    n743
  );


  not
  g834
  (
    n865,
    n637
  );


  not
  g835
  (
    n899,
    n744
  );


  buf
  g836
  (
    n1031,
    n770
  );


  not
  g837
  (
    n863,
    n708
  );


  buf
  g838
  (
    n836,
    n658
  );


  buf
  g839
  (
    n815,
    n747
  );


  not
  g840
  (
    n974,
    n725
  );


  not
  g841
  (
    n816,
    n690
  );


  not
  g842
  (
    n904,
    n766
  );


  not
  g843
  (
    n898,
    n660
  );


  buf
  g844
  (
    n949,
    n760
  );


  buf
  g845
  (
    n911,
    n744
  );


  not
  g846
  (
    n1020,
    n756
  );


  buf
  g847
  (
    n1023,
    n684
  );


  not
  g848
  (
    n859,
    n740
  );


  buf
  g849
  (
    n897,
    n682
  );


  buf
  g850
  (
    n948,
    n642
  );


  not
  g851
  (
    n795,
    n667
  );


  not
  g852
  (
    n905,
    n754
  );


  buf
  g853
  (
    n944,
    n761
  );


  not
  g854
  (
    n951,
    n645
  );


  not
  g855
  (
    n942,
    n732
  );


  or
  g856
  (
    n838,
    n764,
    n766,
    n793
  );


  xor
  g857
  (
    n810,
    n729,
    n751,
    n748,
    n681
  );


  or
  g858
  (
    n877,
    n739,
    n763,
    n793,
    n790
  );


  or
  g859
  (
    n1005,
    n731,
    n670,
    n711,
    n730
  );


  and
  g860
  (
    n853,
    n791,
    n630,
    n740,
    n745
  );


  nor
  g861
  (
    n1013,
    n681,
    n740,
    n721,
    n655
  );


  xnor
  g862
  (
    n857,
    n712,
    n754,
    n667,
    n631
  );


  nand
  g863
  (
    n1012,
    n632,
    n722,
    n786,
    n742
  );


  xnor
  g864
  (
    n1001,
    n711,
    n680,
    n663,
    n638
  );


  and
  g865
  (
    n1025,
    n667,
    n689,
    n752,
    n755
  );


  nand
  g866
  (
    n946,
    n692,
    n639,
    n698,
    n743
  );


  nand
  g867
  (
    n896,
    n649,
    n641,
    n718,
    n626
  );


  or
  g868
  (
    n991,
    n708,
    n774,
    n685,
    n757
  );


  or
  g869
  (
    n979,
    n731,
    n663,
    n686,
    n775
  );


  or
  g870
  (
    n882,
    n655,
    n632,
    n669,
    n658
  );


  or
  g871
  (
    n985,
    n776,
    n710,
    n769,
    n761
  );


  and
  g872
  (
    n809,
    n635,
    n668,
    n633,
    n714
  );


  nor
  g873
  (
    n903,
    n733,
    n728,
    n688,
    n775
  );


  xor
  g874
  (
    n819,
    n702,
    n770,
    n647,
    n691
  );


  nor
  g875
  (
    n831,
    n715,
    n644,
    n730,
    n726
  );


  nor
  g876
  (
    n962,
    n778,
    n656,
    n639,
    n647
  );


  xnor
  g877
  (
    n915,
    n687,
    n714,
    n740,
    n644
  );


  xnor
  g878
  (
    n796,
    n640,
    n771,
    n788,
    n680
  );


  nor
  g879
  (
    n808,
    n715,
    n628,
    n711,
    n741
  );


  xor
  g880
  (
    n804,
    n716,
    n702,
    n707,
    n665
  );


  nor
  g881
  (
    n812,
    n648,
    n634,
    n726,
    n636
  );


  xor
  g882
  (
    n801,
    n791,
    n679,
    n779,
    n657
  );


  and
  g883
  (
    n794,
    n655,
    n676,
    n767,
    n640
  );


  nor
  g884
  (
    n805,
    n748,
    n672,
    n741,
    n771
  );


  nand
  g885
  (
    n802,
    n786,
    n652,
    n772,
    n700
  );


  or
  g886
  (
    n923,
    n675,
    n651,
    n686,
    n669
  );


  xnor
  g887
  (
    n845,
    n700,
    n735,
    n710,
    n773
  );


  nand
  g888
  (
    n953,
    n723,
    n677,
    n777,
    n691
  );


  nand
  g889
  (
    n824,
    n675,
    n704,
    n700,
    n787
  );


  xor
  g890
  (
    n970,
    n779,
    n713,
    n648,
    n674
  );


  or
  g891
  (
    n866,
    n783,
    n699,
    n697,
    n715
  );


  and
  g892
  (
    n935,
    n703,
    n779,
    n695,
    n759
  );


  or
  g893
  (
    n936,
    n785,
    n789,
    n788,
    n631
  );


  and
  g894
  (
    n952,
    n664,
    n748,
    n708,
    n765
  );


  xor
  g895
  (
    n883,
    n736,
    n690,
    n671,
    n729
  );


  nor
  g896
  (
    n1032,
    n656,
    n658,
    n652,
    n678
  );


  xor
  g897
  (
    n797,
    n755,
    n659,
    n639,
    n703
  );


  and
  g898
  (
    n1033,
    n791,
    n629,
    n785,
    n681
  );


  xnor
  g899
  (
    n1017,
    n650,
    n688,
    n792,
    n728
  );


  xor
  g900
  (
    n840,
    n673,
    n742,
    n635,
    n637
  );


  and
  g901
  (
    n1028,
    n721,
    n711,
    n784,
    n695
  );


  nand
  g902
  (
    n1014,
    n646,
    n640,
    n678,
    n772
  );


  xor
  g903
  (
    n958,
    n656,
    n636,
    n634,
    n780
  );


  nand
  g904
  (
    n931,
    n742,
    n789,
    n696,
    n764
  );


  xnor
  g905
  (
    n798,
    n643,
    n727,
    n757,
    n627
  );


  or
  g906
  (
    n995,
    n723,
    n774,
    n722
  );


  xor
  g907
  (
    n1022,
    n646,
    n756,
    n749,
    n657
  );


  xnor
  g908
  (
    n954,
    n629,
    n647,
    n652,
    n786
  );


  xnor
  g909
  (
    n870,
    n709,
    n752,
    n732,
    n627
  );


  or
  g910
  (
    n966,
    n754,
    n774,
    n677,
    n672
  );


  or
  g911
  (
    n976,
    n662,
    n746,
    n632,
    n739
  );


  xnor
  g912
  (
    n892,
    n753,
    n630,
    n710
  );


  nor
  g913
  (
    n875,
    n678,
    n653,
    n768,
    n771
  );


  nand
  g914
  (
    n1003,
    n661,
    n699,
    n660,
    n653
  );


  xnor
  g915
  (
    n1027,
    n707,
    n669,
    n666,
    n728
  );


  nor
  g916
  (
    n943,
    n665,
    n757,
    n784,
    n651
  );


  xnor
  g917
  (
    n1015,
    n758,
    n707,
    n738,
    n639
  );


  xnor
  g918
  (
    n983,
    n694,
    n705,
    n655,
    n686
  );


  nor
  g919
  (
    n820,
    n760,
    n634,
    n630,
    n790
  );


  and
  g920
  (
    n869,
    n765,
    n707,
    n706,
    n730
  );


  or
  g921
  (
    n873,
    n642,
    n724,
    n738,
    n752
  );


  nor
  g922
  (
    n978,
    n699,
    n687,
    n646,
    n793
  );


  nor
  g923
  (
    n1008,
    n671,
    n781,
    n654,
    n744
  );


  or
  g924
  (
    n817,
    n632,
    n782,
    n743,
    n641
  );


  xor
  g925
  (
    n973,
    n661,
    n675,
    n729,
    n702
  );


  xor
  g926
  (
    n964,
    n629,
    n732,
    n763,
    n755
  );


  nand
  g927
  (
    n981,
    n709,
    n769,
    n725,
    n684
  );


  nor
  g928
  (
    n823,
    n779,
    n758,
    n763,
    n629
  );


  nand
  g929
  (
    n926,
    n719,
    n654,
    n705,
    n734
  );


  and
  g930
  (
    n885,
    n714,
    n735,
    n762,
    n751
  );


  nand
  g931
  (
    n975,
    n633,
    n656,
    n691,
    n653
  );


  or
  g932
  (
    n827,
    n788,
    n665,
    n676,
    n768
  );


  xnor
  g933
  (
    n895,
    n652,
    n724,
    n782,
    n739
  );


  nand
  g934
  (
    n906,
    n728,
    n743,
    n705,
    n737
  );


  xnor
  g935
  (
    n1004,
    n793,
    n647,
    n777,
    n698
  );


  xnor
  g936
  (
    n950,
    n669,
    n716,
    n770,
    n649
  );


  xnor
  g937
  (
    n888,
    n709,
    n770,
    n626,
    n682
  );


  xor
  g938
  (
    n1024,
    n654,
    n691,
    n648,
    n667
  );


  or
  g939
  (
    n881,
    n763,
    n680,
    n760,
    n759
  );


  xnor
  g940
  (
    n852,
    n638,
    n693,
    n631,
    n737
  );


  nor
  g941
  (
    n917,
    n659,
    n720,
    n736,
    n641
  );


  xor
  g942
  (
    n924,
    n633,
    n718,
    n712,
    n664
  );


  or
  g943
  (
    n939,
    n758,
    n701,
    n750,
    n727
  );


  and
  g944
  (
    n984,
    n663,
    n687,
    n659,
    n719
  );


  and
  g945
  (
    n894,
    n745,
    n685,
    n635,
    n653
  );


  nand
  g946
  (
    n925,
    n679,
    n682,
    n686,
    n670
  );


  xor
  g947
  (
    n862,
    n780,
    n769,
    n751,
    n692
  );


  and
  g948
  (
    n933,
    n688,
    n778,
    n733,
    n723
  );


  xnor
  g949
  (
    n1029,
    n792,
    n764,
    n697,
    n744
  );


  nand
  g950
  (
    n887,
    n712,
    n670,
    n640,
    n625
  );


  and
  g951
  (
    n938,
    n768,
    n762,
    n777,
    n765
  );


  or
  g952
  (
    n922,
    n792,
    n679,
    n631,
    n646
  );


  or
  g953
  (
    n959,
    n689,
    n657,
    n690,
    n716
  );


  xor
  g954
  (
    n1002,
    n699,
    n790,
    n703,
    n706
  );


  and
  g955
  (
    n851,
    n685,
    n701,
    n693,
    n683
  );


  and
  g956
  (
    n998,
    n766,
    n697,
    n791,
    n739
  );


  and
  g957
  (
    n1019,
    n658,
    n753,
    n761,
    n775
  );


  nand
  g958
  (
    n800,
    n729,
    n698,
    n688,
    n751
  );


  and
  g959
  (
    n1010,
    n749,
    n746,
    n776,
    n754
  );


  or
  g960
  (
    n871,
    n781,
    n782,
    n674,
    n666
  );


  nand
  g961
  (
    n880,
    n790,
    n627,
    n636,
    n787
  );


  xor
  g962
  (
    n872,
    n761,
    n648,
    n708,
    n717
  );


  nor
  g963
  (
    n986,
    n760,
    n757,
    n666,
    n684
  );


  xor
  g964
  (
    n916,
    n778,
    n738,
    n784,
    n668
  );


  nor
  g965
  (
    n856,
    n726,
    n683,
    n662,
    n702
  );


  xor
  g966
  (
    n1021,
    n735,
    n644,
    n732,
    n780
  );


  nor
  g967
  (
    n908,
    n734,
    n735,
    n764,
    n643
  );


  or
  g968
  (
    n814,
    n698,
    n709,
    n696,
    n676
  );


  xor
  g969
  (
    n957,
    n681,
    n767,
    n692,
    n759
  );


  or
  g970
  (
    n890,
    n665,
    n682,
    n717,
    n792
  );


  nand
  g971
  (
    n867,
    n787,
    n786,
    n780,
    n668
  );


  xor
  g972
  (
    n848,
    n674,
    n762,
    n649,
    n673
  );


  or
  g973
  (
    n832,
    n654,
    n714,
    n633,
    n748
  );


  and
  g974
  (
    n987,
    n673,
    n784,
    n696,
    n785
  );


  nor
  g975
  (
    n928,
    n737,
    n717,
    n789,
    n663
  );


  nor
  g976
  (
    n879,
    n638,
    n719,
    n683,
    n783
  );


  nand
  g977
  (
    n929,
    n645,
    n661,
    n718,
    n766
  );


  xor
  g978
  (
    n909,
    n716,
    n649,
    n758,
    n693
  );


  and
  g979
  (
    n965,
    n693,
    n753,
    n625,
    n731
  );


  and
  g980
  (
    n980,
    n772,
    n644,
    n637,
    n643
  );


  and
  g981
  (
    n912,
    n664,
    n697,
    n625,
    n778
  );


  nand
  g982
  (
    n977,
    n659,
    n692,
    n721,
    n727
  );


  nand
  g983
  (
    n993,
    n704,
    n774,
    n635,
    n642
  );


  nand
  g984
  (
    n927,
    n767,
    n775,
    n741,
    n650
  );


  nor
  g985
  (
    n934,
    n641,
    n746,
    n756,
    n677
  );


  xnor
  g986
  (
    n955,
    n737,
    n684,
    n722,
    n636
  );


  xnor
  g987
  (
    n1030,
    n738,
    n696,
    n776,
    n628
  );


  nand
  g988
  (
    n967,
    n731,
    n734,
    n627,
    n762
  );


  xor
  g989
  (
    n835,
    n720,
    n720,
    n717,
    n759
  );


  xor
  g990
  (
    n972,
    n650,
    n694,
    n769,
    n706
  );


  nand
  g991
  (
    n920,
    n773,
    n643,
    n749,
    n651
  );


  and
  g992
  (
    n864,
    n660,
    n746,
    n689,
    n645
  );


  and
  g993
  (
    n830,
    n664,
    n704,
    n683,
    n782
  );


  xor
  g994
  (
    n813,
    n628,
    n677,
    n638,
    n661
  );


  xnor
  g995
  (
    n989,
    n781,
    n671,
    n690,
    n712
  );


  xnor
  g996
  (
    n1016,
    n718,
    n680,
    n725,
    n630
  );


  or
  g997
  (
    n837,
    n701,
    n657,
    n742,
    n767
  );


  and
  g998
  (
    n914,
    n673,
    n783,
    n666,
    n724
  );


  xnor
  g999
  (
    n886,
    n687,
    n747,
    n723,
    n781
  );


  nor
  g1000
  (
    n850,
    n750,
    n706,
    n777,
    n662
  );


  buf
  g1001
  (
    n1805,
    n956
  );


  buf
  g1002
  (
    n1488,
    n974
  );


  not
  g1003
  (
    n1412,
    n845
  );


  buf
  g1004
  (
    n1608,
    n893
  );


  not
  g1005
  (
    n1565,
    n896
  );


  buf
  g1006
  (
    n1388,
    n965
  );


  buf
  g1007
  (
    n1788,
    n968
  );


  buf
  g1008
  (
    n1784,
    n961
  );


  buf
  g1009
  (
    n1764,
    n899
  );


  not
  g1010
  (
    n1660,
    n909
  );


  not
  g1011
  (
    n1334,
    n901
  );


  buf
  g1012
  (
    n1760,
    n1009
  );


  buf
  g1013
  (
    n1898,
    n930
  );


  not
  g1014
  (
    n1065,
    n834
  );


  buf
  g1015
  (
    n1228,
    n1014
  );


  not
  g1016
  (
    n1540,
    n945
  );


  not
  g1017
  (
    n1441,
    n967
  );


  not
  g1018
  (
    n1477,
    n1025
  );


  buf
  g1019
  (
    n1593,
    n866
  );


  buf
  g1020
  (
    n1309,
    n855
  );


  not
  g1021
  (
    n1380,
    n996
  );


  not
  g1022
  (
    n1212,
    n888
  );


  buf
  g1023
  (
    n1532,
    n907
  );


  buf
  g1024
  (
    n1816,
    n934
  );


  buf
  g1025
  (
    n1268,
    n936
  );


  not
  g1026
  (
    n1740,
    n880
  );


  buf
  g1027
  (
    n1545,
    n868
  );


  not
  g1028
  (
    n1774,
    n829
  );


  not
  g1029
  (
    n1790,
    n1007
  );


  not
  g1030
  (
    n1156,
    n996
  );


  not
  g1031
  (
    n1499,
    n799
  );


  not
  g1032
  (
    n1042,
    n948
  );


  not
  g1033
  (
    n1289,
    n1018
  );


  not
  g1034
  (
    n1688,
    n796
  );


  not
  g1035
  (
    n1104,
    n841
  );


  buf
  g1036
  (
    n1553,
    n1017
  );


  buf
  g1037
  (
    n1038,
    n944
  );


  buf
  g1038
  (
    n1452,
    n902
  );


  not
  g1039
  (
    n1480,
    n903
  );


  buf
  g1040
  (
    n1373,
    n801
  );


  buf
  g1041
  (
    n1625,
    n946
  );


  buf
  g1042
  (
    n1709,
    n949
  );


  not
  g1043
  (
    n1219,
    n925
  );


  buf
  g1044
  (
    n1485,
    n848
  );


  buf
  g1045
  (
    n1066,
    n863
  );


  buf
  g1046
  (
    n1721,
    n892
  );


  not
  g1047
  (
    n1749,
    n814
  );


  not
  g1048
  (
    n1283,
    n972
  );


  not
  g1049
  (
    n1511,
    n865
  );


  not
  g1050
  (
    n1270,
    n969
  );


  buf
  g1051
  (
    n1391,
    n946
  );


  not
  g1052
  (
    n1750,
    n800
  );


  buf
  g1053
  (
    n1433,
    n976
  );


  not
  g1054
  (
    n1569,
    n908
  );


  not
  g1055
  (
    n1514,
    n997
  );


  not
  g1056
  (
    n1258,
    n991
  );


  buf
  g1057
  (
    n1801,
    n986
  );


  buf
  g1058
  (
    n1686,
    n1005
  );


  buf
  g1059
  (
    n1910,
    n985
  );


  buf
  g1060
  (
    n1053,
    n1021
  );


  not
  g1061
  (
    n1503,
    n1012
  );


  not
  g1062
  (
    n1827,
    n962
  );


  not
  g1063
  (
    n1554,
    n941
  );


  not
  g1064
  (
    n1186,
    n906
  );


  not
  g1065
  (
    n1497,
    n1008
  );


  buf
  g1066
  (
    n1176,
    n1025
  );


  buf
  g1067
  (
    n1142,
    n799
  );


  buf
  g1068
  (
    n1658,
    n912
  );


  not
  g1069
  (
    n1639,
    n889
  );


  buf
  g1070
  (
    n1466,
    n807
  );


  buf
  g1071
  (
    n1573,
    n997
  );


  buf
  g1072
  (
    n1733,
    n813
  );


  buf
  g1073
  (
    n1317,
    n963
  );


  buf
  g1074
  (
    n1201,
    n206
  );


  not
  g1075
  (
    n1071,
    n829
  );


  not
  g1076
  (
    n1439,
    n927
  );


  buf
  g1077
  (
    n1077,
    n805
  );


  buf
  g1078
  (
    n1567,
    n797
  );


  not
  g1079
  (
    n1339,
    n823
  );


  buf
  g1080
  (
    n1505,
    n821
  );


  buf
  g1081
  (
    n1035,
    n812
  );


  buf
  g1082
  (
    n1907,
    n839
  );


  not
  g1083
  (
    n1891,
    n869
  );


  not
  g1084
  (
    n1881,
    n1016
  );


  not
  g1085
  (
    n1534,
    n966
  );


  buf
  g1086
  (
    n1550,
    n1020
  );


  not
  g1087
  (
    n1926,
    n922
  );


  buf
  g1088
  (
    n1860,
    n1006
  );


  not
  g1089
  (
    n1671,
    n988
  );


  not
  g1090
  (
    n1747,
    n821
  );


  not
  g1091
  (
    n1251,
    n846
  );


  buf
  g1092
  (
    n1135,
    n1007
  );


  not
  g1093
  (
    n1397,
    n850
  );


  not
  g1094
  (
    n1803,
    n835
  );


  not
  g1095
  (
    n1654,
    n837
  );


  not
  g1096
  (
    n1130,
    n1022
  );


  buf
  g1097
  (
    n1861,
    n861
  );


  not
  g1098
  (
    n1606,
    n827
  );


  not
  g1099
  (
    n1165,
    n1002
  );


  buf
  g1100
  (
    n1196,
    n999
  );


  buf
  g1101
  (
    n1664,
    n857
  );


  not
  g1102
  (
    n1325,
    n926
  );


  buf
  g1103
  (
    n1638,
    n994
  );


  buf
  g1104
  (
    n1349,
    n945
  );


  buf
  g1105
  (
    n1779,
    n985
  );


  not
  g1106
  (
    n1442,
    n848
  );


  buf
  g1107
  (
    n1248,
    n848
  );


  buf
  g1108
  (
    n1762,
    n1008
  );


  not
  g1109
  (
    n1166,
    n836
  );


  buf
  g1110
  (
    n1387,
    n930
  );


  not
  g1111
  (
    n1657,
    n816
  );


  not
  g1112
  (
    n1546,
    n917
  );


  not
  g1113
  (
    n1647,
    n846
  );


  buf
  g1114
  (
    n1605,
    n827
  );


  not
  g1115
  (
    n1555,
    n966
  );


  buf
  g1116
  (
    n1456,
    n878
  );


  buf
  g1117
  (
    n1102,
    n886
  );


  buf
  g1118
  (
    n1913,
    n1013
  );


  buf
  g1119
  (
    n1644,
    n943
  );


  not
  g1120
  (
    n1359,
    n978
  );


  buf
  g1121
  (
    n1524,
    n939
  );


  not
  g1122
  (
    n1254,
    n896
  );


  not
  g1123
  (
    n1875,
    n951
  );


  not
  g1124
  (
    n1318,
    n1020
  );


  buf
  g1125
  (
    n1735,
    n982
  );


  buf
  g1126
  (
    n1160,
    n1021
  );


  not
  g1127
  (
    n1703,
    n820
  );


  buf
  g1128
  (
    n1210,
    n885
  );


  not
  g1129
  (
    n1474,
    n808
  );


  not
  g1130
  (
    n1313,
    n846
  );


  not
  g1131
  (
    n1675,
    n993
  );


  not
  g1132
  (
    n1879,
    n205
  );


  buf
  g1133
  (
    n1095,
    n1015
  );


  buf
  g1134
  (
    n1134,
    n865
  );


  not
  g1135
  (
    n1842,
    n916
  );


  buf
  g1136
  (
    n1247,
    n841
  );


  buf
  g1137
  (
    n1106,
    n1008
  );


  buf
  g1138
  (
    n1508,
    n861
  );


  buf
  g1139
  (
    n1336,
    n926
  );


  not
  g1140
  (
    n1314,
    n884
  );


  buf
  g1141
  (
    n1737,
    n825
  );


  buf
  g1142
  (
    n1817,
    n835
  );


  buf
  g1143
  (
    n1195,
    n950
  );


  not
  g1144
  (
    n1140,
    n887
  );


  buf
  g1145
  (
    n1406,
    n1019
  );


  buf
  g1146
  (
    n1108,
    n966
  );


  not
  g1147
  (
    n1164,
    n840
  );


  buf
  g1148
  (
    n1171,
    n890
  );


  not
  g1149
  (
    n1202,
    n951
  );


  buf
  g1150
  (
    n1579,
    n882
  );


  not
  g1151
  (
    n1386,
    n953
  );


  not
  g1152
  (
    n1791,
    n1004
  );


  not
  g1153
  (
    n1263,
    n845
  );


  not
  g1154
  (
    n1487,
    n795
  );


  buf
  g1155
  (
    n1304,
    n819
  );


  buf
  g1156
  (
    n1620,
    n1007
  );


  buf
  g1157
  (
    n1244,
    n925
  );


  buf
  g1158
  (
    n1473,
    n999
  );


  not
  g1159
  (
    n1830,
    n842
  );


  not
  g1160
  (
    n1138,
    n823
  );


  not
  g1161
  (
    n1179,
    n1010
  );


  buf
  g1162
  (
    n1547,
    n872
  );


  buf
  g1163
  (
    n1281,
    n1016
  );


  buf
  g1164
  (
    n1401,
    n862
  );


  not
  g1165
  (
    n1865,
    n921
  );


  buf
  g1166
  (
    n1706,
    n956
  );


  buf
  g1167
  (
    n1836,
    n854
  );


  buf
  g1168
  (
    n1746,
    n1012
  );


  buf
  g1169
  (
    n1670,
    n819
  );


  buf
  g1170
  (
    n1720,
    n963
  );


  not
  g1171
  (
    n1435,
    n1013
  );


  buf
  g1172
  (
    n1416,
    n988
  );


  not
  g1173
  (
    n1049,
    n802
  );


  not
  g1174
  (
    n1343,
    n997
  );


  buf
  g1175
  (
    n1848,
    n857
  );


  not
  g1176
  (
    n1856,
    n911
  );


  buf
  g1177
  (
    n1502,
    n881
  );


  not
  g1178
  (
    n1455,
    n856
  );


  buf
  g1179
  (
    n1612,
    n862
  );


  buf
  g1180
  (
    n1837,
    n876
  );


  not
  g1181
  (
    n1105,
    n950
  );


  not
  g1182
  (
    n1903,
    n812
  );


  buf
  g1183
  (
    n1125,
    n834
  );


  buf
  g1184
  (
    n1815,
    n206
  );


  not
  g1185
  (
    n1252,
    n951
  );


  buf
  g1186
  (
    n1577,
    n818
  );


  not
  g1187
  (
    n1440,
    n924
  );


  buf
  g1188
  (
    n1491,
    n967
  );


  buf
  g1189
  (
    n1494,
    n815
  );


  buf
  g1190
  (
    n1080,
    n794
  );


  buf
  g1191
  (
    n1460,
    n900
  );


  buf
  g1192
  (
    n1797,
    n1028
  );


  not
  g1193
  (
    n1124,
    n990
  );


  not
  g1194
  (
    n1759,
    n998
  );


  not
  g1195
  (
    n1927,
    n1024
  );


  not
  g1196
  (
    n1451,
    n868
  );


  buf
  g1197
  (
    n1233,
    n998
  );


  buf
  g1198
  (
    n1128,
    n916
  );


  buf
  g1199
  (
    n1398,
    n987
  );


  buf
  g1200
  (
    n1344,
    n1022
  );


  buf
  g1201
  (
    n1590,
    n930
  );


  not
  g1202
  (
    n1697,
    n1001
  );


  buf
  g1203
  (
    n1752,
    n829
  );


  buf
  g1204
  (
    n1168,
    n892
  );


  not
  g1205
  (
    n1831,
    n997
  );


  not
  g1206
  (
    n1857,
    n986
  );


  buf
  g1207
  (
    n1624,
    n979
  );


  buf
  g1208
  (
    n1197,
    n911
  );


  not
  g1209
  (
    n1372,
    n986
  );


  buf
  g1210
  (
    n1381,
    n874
  );


  not
  g1211
  (
    n1234,
    n879
  );


  buf
  g1212
  (
    n1613,
    n947
  );


  not
  g1213
  (
    n1450,
    n983
  );


  buf
  g1214
  (
    n1086,
    n947
  );


  buf
  g1215
  (
    n1526,
    n998
  );


  buf
  g1216
  (
    n1161,
    n971
  );


  not
  g1217
  (
    n1810,
    n928
  );


  not
  g1218
  (
    n1900,
    n830
  );


  not
  g1219
  (
    n1719,
    n879
  );


  not
  g1220
  (
    n1043,
    n801
  );


  not
  g1221
  (
    n1932,
    n968
  );


  buf
  g1222
  (
    n1562,
    n1005
  );


  not
  g1223
  (
    n1117,
    n918
  );


  not
  g1224
  (
    n1859,
    n920
  );


  not
  g1225
  (
    n1256,
    n904
  );


  not
  g1226
  (
    n1649,
    n877
  );


  buf
  g1227
  (
    n1522,
    n876
  );


  buf
  g1228
  (
    n1635,
    n795
  );


  buf
  g1229
  (
    n1286,
    n1011
  );


  not
  g1230
  (
    n1328,
    n831
  );


  buf
  g1231
  (
    n1715,
    n1000
  );


  not
  g1232
  (
    n1229,
    n878
  );


  buf
  g1233
  (
    n1418,
    n938
  );


  not
  g1234
  (
    n1659,
    n1030
  );


  buf
  g1235
  (
    n1911,
    n946
  );


  not
  g1236
  (
    n1482,
    n840
  );


  not
  g1237
  (
    n1915,
    n992
  );


  not
  g1238
  (
    n1097,
    n952
  );


  not
  g1239
  (
    n1299,
    n900
  );


  not
  g1240
  (
    n1366,
    n842
  );


  not
  g1241
  (
    n1871,
    n839
  );


  buf
  g1242
  (
    n1517,
    n942
  );


  not
  g1243
  (
    n1887,
    n1000
  );


  buf
  g1244
  (
    n1350,
    n847
  );


  buf
  g1245
  (
    n1240,
    n884
  );


  not
  g1246
  (
    n1463,
    n1026
  );


  buf
  g1247
  (
    n1708,
    n849
  );


  not
  g1248
  (
    n1157,
    n863
  );


  buf
  g1249
  (
    n1807,
    n974
  );


  not
  g1250
  (
    n1408,
    n861
  );


  not
  g1251
  (
    n1754,
    n835
  );


  buf
  g1252
  (
    n1518,
    n864
  );


  buf
  g1253
  (
    n1434,
    n923
  );


  buf
  g1254
  (
    n1712,
    n1030
  );


  buf
  g1255
  (
    n1217,
    n980
  );


  not
  g1256
  (
    n1870,
    n918
  );


  buf
  g1257
  (
    n1409,
    n983
  );


  not
  g1258
  (
    n1100,
    n808
  );


  not
  g1259
  (
    n1149,
    n812
  );


  not
  g1260
  (
    n1415,
    n205
  );


  buf
  g1261
  (
    n1483,
    n938
  );


  not
  g1262
  (
    n1855,
    n1024
  );


  buf
  g1263
  (
    n1211,
    n1004
  );


  not
  g1264
  (
    n1583,
    n976
  );


  buf
  g1265
  (
    n1589,
    n864
  );


  buf
  g1266
  (
    n1162,
    n1027
  );


  buf
  g1267
  (
    n1262,
    n925
  );


  buf
  g1268
  (
    n1702,
    n957
  );


  not
  g1269
  (
    n1853,
    n828
  );


  buf
  g1270
  (
    n1255,
    n877
  );


  buf
  g1271
  (
    n1832,
    n850
  );


  not
  g1272
  (
    n1330,
    n873
  );


  not
  g1273
  (
    n1191,
    n820
  );


  not
  g1274
  (
    n1884,
    n961
  );


  not
  g1275
  (
    n1716,
    n916
  );


  buf
  g1276
  (
    n1352,
    n844
  );


  not
  g1277
  (
    n1669,
    n816
  );


  not
  g1278
  (
    n1713,
    n889
  );


  not
  g1279
  (
    n1402,
    n905
  );


  not
  g1280
  (
    n1449,
    n884
  );


  buf
  g1281
  (
    n1552,
    n919
  );


  buf
  g1282
  (
    n1661,
    n804
  );


  not
  g1283
  (
    n1814,
    n823
  );


  buf
  g1284
  (
    n1689,
    n1013
  );


  not
  g1285
  (
    n1148,
    n955
  );


  not
  g1286
  (
    n1465,
    n981
  );


  not
  g1287
  (
    n1253,
    n881
  );


  buf
  g1288
  (
    n1642,
    n875
  );


  buf
  g1289
  (
    n1489,
    n901
  );


  buf
  g1290
  (
    n1628,
    n1010
  );


  not
  g1291
  (
    n1429,
    n853
  );


  not
  g1292
  (
    n1290,
    n907
  );


  not
  g1293
  (
    n1621,
    n1004
  );


  buf
  g1294
  (
    n1428,
    n994
  );


  not
  g1295
  (
    n1698,
    n1006
  );


  not
  g1296
  (
    n1458,
    n845
  );


  buf
  g1297
  (
    n1756,
    n1008
  );


  buf
  g1298
  (
    n1591,
    n920
  );


  not
  g1299
  (
    n1650,
    n1022
  );


  buf
  g1300
  (
    n1885,
    n806
  );


  buf
  g1301
  (
    n1793,
    n921
  );


  not
  g1302
  (
    n1530,
    n970
  );


  not
  g1303
  (
    n1092,
    n993
  );


  not
  g1304
  (
    n1395,
    n1014
  );


  buf
  g1305
  (
    n1150,
    n961
  );


  buf
  g1306
  (
    n1223,
    n928
  );


  buf
  g1307
  (
    n1531,
    n924
  );


  not
  g1308
  (
    n1348,
    n892
  );


  not
  g1309
  (
    n1777,
    n815
  );


  buf
  g1310
  (
    n1193,
    n968
  );


  not
  g1311
  (
    n1772,
    n1023
  );


  buf
  g1312
  (
    n1582,
    n837
  );


  not
  g1313
  (
    n1789,
    n989
  );


  buf
  g1314
  (
    n1250,
    n866
  );


  not
  g1315
  (
    n1781,
    n1002
  );


  buf
  g1316
  (
    n1739,
    n883
  );


  not
  g1317
  (
    n1420,
    n899
  );


  not
  g1318
  (
    n1766,
    n870
  );


  not
  g1319
  (
    n1923,
    n1030
  );


  not
  g1320
  (
    n1340,
    n835
  );


  not
  g1321
  (
    n1404,
    n1020
  );


  not
  g1322
  (
    n1652,
    n911
  );


  buf
  g1323
  (
    n1082,
    n836
  );


  not
  g1324
  (
    n1634,
    n854
  );


  not
  g1325
  (
    n1167,
    n881
  );


  not
  g1326
  (
    n1111,
    n966
  );


  buf
  g1327
  (
    n1385,
    n814
  );


  buf
  g1328
  (
    n1691,
    n971
  );


  buf
  g1329
  (
    n1367,
    n840
  );


  buf
  g1330
  (
    n1151,
    n890
  );


  not
  g1331
  (
    n1414,
    n914
  );


  not
  g1332
  (
    n1265,
    n1017
  );


  not
  g1333
  (
    n1901,
    n849
  );


  not
  g1334
  (
    n1575,
    n844
  );


  buf
  g1335
  (
    n1034,
    n816
  );


  not
  g1336
  (
    n1558,
    n1021
  );


  buf
  g1337
  (
    n1630,
    n1023
  );


  not
  g1338
  (
    n1479,
    n943
  );


  buf
  g1339
  (
    n1360,
    n885
  );


  not
  g1340
  (
    n1776,
    n942
  );


  buf
  g1341
  (
    n1858,
    n1018
  );


  not
  g1342
  (
    n1492,
    n893
  );


  not
  g1343
  (
    n1623,
    n804
  );


  not
  g1344
  (
    n1852,
    n914
  );


  buf
  g1345
  (
    n1431,
    n811
  );


  buf
  g1346
  (
    n1734,
    n1012
  );


  not
  g1347
  (
    n1184,
    n830
  );


  not
  g1348
  (
    n1237,
    n811
  );


  buf
  g1349
  (
    n1358,
    n1003
  );


  not
  g1350
  (
    n1561,
    n1001
  );


  not
  g1351
  (
    n1353,
    n951
  );


  not
  g1352
  (
    n1795,
    n908
  );


  buf
  g1353
  (
    n1653,
    n953
  );


  not
  g1354
  (
    n1292,
    n897
  );


  buf
  g1355
  (
    n1332,
    n960
  );


  buf
  g1356
  (
    n1666,
    n798
  );


  not
  g1357
  (
    n1556,
    n907
  );


  not
  g1358
  (
    n1103,
    n919
  );


  buf
  g1359
  (
    n1321,
    n936
  );


  buf
  g1360
  (
    n1758,
    n832
  );


  not
  g1361
  (
    n1773,
    n964
  );


  buf
  g1362
  (
    n1778,
    n826
  );


  buf
  g1363
  (
    n1761,
    n843
  );


  not
  g1364
  (
    n1368,
    n795
  );


  not
  g1365
  (
    n1728,
    n944
  );


  not
  g1366
  (
    n1717,
    n870
  );


  buf
  g1367
  (
    n1896,
    n886
  );


  buf
  g1368
  (
    n1341,
    n968
  );


  buf
  g1369
  (
    n1120,
    n995
  );


  not
  g1370
  (
    n1403,
    n939
  );


  not
  g1371
  (
    n1207,
    n919
  );


  buf
  g1372
  (
    n1445,
    n803
  );


  buf
  g1373
  (
    n1806,
    n879
  );


  buf
  g1374
  (
    n1496,
    n920
  );


  buf
  g1375
  (
    n1394,
    n948
  );


  buf
  g1376
  (
    n1690,
    n1029
  );


  buf
  g1377
  (
    n1113,
    n935
  );


  not
  g1378
  (
    n1521,
    n921
  );


  buf
  g1379
  (
    n1298,
    n940
  );


  buf
  g1380
  (
    n1059,
    n823
  );


  not
  g1381
  (
    n1566,
    n850
  );


  buf
  g1382
  (
    n1844,
    n1028
  );


  buf
  g1383
  (
    n1763,
    n821
  );


  not
  g1384
  (
    n1227,
    n1003
  );


  not
  g1385
  (
    n1061,
    n955
  );


  not
  g1386
  (
    n1301,
    n932
  );


  buf
  g1387
  (
    n1087,
    n903
  );


  not
  g1388
  (
    n1796,
    n833
  );


  buf
  g1389
  (
    n1743,
    n882
  );


  not
  g1390
  (
    n1279,
    n826
  );


  not
  g1391
  (
    n1099,
    n926
  );


  not
  g1392
  (
    n1916,
    n979
  );


  buf
  g1393
  (
    n1529,
    n838
  );


  buf
  g1394
  (
    n1745,
    n898
  );


  not
  g1395
  (
    n1570,
    n872
  );


  not
  g1396
  (
    n1182,
    n941
  );


  not
  g1397
  (
    n1622,
    n924
  );


  not
  g1398
  (
    n1362,
    n928
  );


  not
  g1399
  (
    n1088,
    n802
  );


  not
  g1400
  (
    n1147,
    n916
  );


  buf
  g1401
  (
    n1109,
    n849
  );


  buf
  g1402
  (
    n1096,
    n852
  );


  buf
  g1403
  (
    n1090,
    n812
  );


  not
  g1404
  (
    n1192,
    n937
  );


  not
  g1405
  (
    n1158,
    n989
  );


  buf
  g1406
  (
    n1269,
    n891
  );


  buf
  g1407
  (
    n1051,
    n1026
  );


  buf
  g1408
  (
    n1854,
    n809
  );


  not
  g1409
  (
    n1930,
    n1032
  );


  not
  g1410
  (
    n1375,
    n980
  );


  buf
  g1411
  (
    n1116,
    n995
  );


  buf
  g1412
  (
    n1890,
    n800
  );


  not
  g1413
  (
    n1285,
    n806
  );


  not
  g1414
  (
    n1742,
    n1028
  );


  buf
  g1415
  (
    n1925,
    n895
  );


  not
  g1416
  (
    n1469,
    n1000
  );


  buf
  g1417
  (
    n1094,
    n943
  );


  not
  g1418
  (
    n1548,
    n1010
  );


  not
  g1419
  (
    n1346,
    n990
  );


  buf
  g1420
  (
    n1040,
    n902
  );


  not
  g1421
  (
    n1235,
    n1028
  );


  not
  g1422
  (
    n1039,
    n1010
  );


  not
  g1423
  (
    n1272,
    n969
  );


  buf
  g1424
  (
    n1711,
    n841
  );


  not
  g1425
  (
    n1417,
    n987
  );


  not
  g1426
  (
    n1519,
    n936
  );


  not
  g1427
  (
    n1423,
    n889
  );


  buf
  g1428
  (
    n1324,
    n990
  );


  buf
  g1429
  (
    n1284,
    n930
  );


  buf
  g1430
  (
    n1845,
    n870
  );


  not
  g1431
  (
    n1347,
    n1011
  );


  buf
  g1432
  (
    n1867,
    n1015
  );


  buf
  g1433
  (
    n1457,
    n796
  );


  not
  g1434
  (
    n1327,
    n818
  );


  buf
  g1435
  (
    n1663,
    n1001
  );


  not
  g1436
  (
    n1533,
    n992
  );


  not
  g1437
  (
    n1126,
    n887
  );


  buf
  g1438
  (
    n1137,
    n842
  );


  buf
  g1439
  (
    n1770,
    n1014
  );


  buf
  g1440
  (
    n1243,
    n910
  );


  not
  g1441
  (
    n1563,
    n924
  );


  not
  g1442
  (
    n1453,
    n949
  );


  buf
  g1443
  (
    n1895,
    n933
  );


  buf
  g1444
  (
    n1800,
    n945
  );


  not
  g1445
  (
    n1390,
    n957
  );


  not
  g1446
  (
    n1581,
    n858
  );


  buf
  g1447
  (
    n1536,
    n960
  );


  not
  g1448
  (
    n1363,
    n854
  );


  not
  g1449
  (
    n1655,
    n796
  );


  not
  g1450
  (
    n1645,
    n1003
  );


  buf
  g1451
  (
    n1677,
    n847
  );


  buf
  g1452
  (
    n1114,
    n929
  );


  buf
  g1453
  (
    n1592,
    n901
  );


  buf
  g1454
  (
    n1924,
    n827
  );


  not
  g1455
  (
    n1089,
    n899
  );


  not
  g1456
  (
    n1904,
    n819
  );


  not
  g1457
  (
    n1241,
    n1006
  );


  buf
  g1458
  (
    n1424,
    n817
  );


  not
  g1459
  (
    n1851,
    n844
  );


  not
  g1460
  (
    n1929,
    n824
  );


  buf
  g1461
  (
    n1393,
    n922
  );


  not
  g1462
  (
    n1389,
    n822
  );


  buf
  g1463
  (
    n1303,
    n833
  );


  not
  g1464
  (
    n1769,
    n852
  );


  not
  g1465
  (
    n1041,
    n828
  );


  not
  g1466
  (
    n1432,
    n949
  );


  not
  g1467
  (
    n1308,
    n830
  );


  not
  g1468
  (
    n1154,
    n862
  );


  not
  g1469
  (
    n1280,
    n984
  );


  buf
  g1470
  (
    n1484,
    n1031
  );


  buf
  g1471
  (
    n1906,
    n798
  );


  buf
  g1472
  (
    n1539,
    n813
  );


  buf
  g1473
  (
    n1732,
    n834
  );


  buf
  g1474
  (
    n1369,
    n988
  );


  buf
  g1475
  (
    n1786,
    n898
  );


  buf
  g1476
  (
    n1356,
    n867
  );


  buf
  g1477
  (
    n1333,
    n861
  );


  not
  g1478
  (
    n1062,
    n804
  );


  not
  g1479
  (
    n1446,
    n805
  );


  not
  g1480
  (
    n1679,
    n868
  );


  buf
  g1481
  (
    n1276,
    n914
  );


  buf
  g1482
  (
    n1199,
    n984
  );


  buf
  g1483
  (
    n1611,
    n985
  );


  not
  g1484
  (
    n1467,
    n959
  );


  not
  g1485
  (
    n1685,
    n910
  );


  not
  g1486
  (
    n1873,
    n940
  );


  not
  g1487
  (
    n1825,
    n839
  );


  buf
  g1488
  (
    n1568,
    n1000
  );


  not
  g1489
  (
    n1205,
    n958
  );


  not
  g1490
  (
    n1821,
    n863
  );


  not
  g1491
  (
    n1464,
    n1009
  );


  not
  g1492
  (
    n1232,
    n902
  );


  not
  g1493
  (
    n1218,
    n931
  );


  not
  g1494
  (
    n1872,
    n978
  );


  buf
  g1495
  (
    n1354,
    n971
  );


  not
  g1496
  (
    n1601,
    n983
  );


  not
  g1497
  (
    n1928,
    n915
  );


  not
  g1498
  (
    n1101,
    n953
  );


  buf
  g1499
  (
    n1081,
    n859
  );


  buf
  g1500
  (
    n1180,
    n885
  );


  buf
  g1501
  (
    n1886,
    n874
  );


  not
  g1502
  (
    n1425,
    n851
  );


  buf
  g1503
  (
    n1617,
    n940
  );


  not
  g1504
  (
    n1785,
    n848
  );


  buf
  g1505
  (
    n1183,
    n976
  );


  buf
  g1506
  (
    n1172,
    n847
  );


  buf
  g1507
  (
    n1905,
    n939
  );


  not
  g1508
  (
    n1525,
    n836
  );


  buf
  g1509
  (
    n1122,
    n896
  );


  buf
  g1510
  (
    n1616,
    n814
  );


  not
  g1511
  (
    n1880,
    n843
  );


  not
  g1512
  (
    n1323,
    n982
  );


  buf
  g1513
  (
    n1278,
    n952
  );


  buf
  g1514
  (
    n1036,
    n859
  );


  buf
  g1515
  (
    n1692,
    n955
  );


  buf
  g1516
  (
    n1091,
    n929
  );


  buf
  g1517
  (
    n1874,
    n869
  );


  not
  g1518
  (
    n1107,
    n963
  );


  not
  g1519
  (
    n1242,
    n947
  );


  not
  g1520
  (
    n1069,
    n866
  );


  buf
  g1521
  (
    n1236,
    n965
  );


  not
  g1522
  (
    n1922,
    n1003
  );


  buf
  g1523
  (
    n1046,
    n998
  );


  not
  g1524
  (
    n1787,
    n895
  );


  buf
  g1525
  (
    n1054,
    n826
  );


  buf
  g1526
  (
    n1588,
    n945
  );


  not
  g1527
  (
    n1571,
    n940
  );


  buf
  g1528
  (
    n1294,
    n901
  );


  not
  g1529
  (
    n1603,
    n831
  );


  not
  g1530
  (
    n1152,
    n909
  );


  buf
  g1531
  (
    n1259,
    n876
  );


  buf
  g1532
  (
    n1731,
    n933
  );


  not
  g1533
  (
    n1510,
    n825
  );


  buf
  g1534
  (
    n1214,
    n958
  );


  not
  g1535
  (
    n1410,
    n991
  );


  buf
  g1536
  (
    n1123,
    n205
  );


  not
  g1537
  (
    n1288,
    n1019
  );


  buf
  g1538
  (
    n1730,
    n841
  );


  not
  g1539
  (
    n1405,
    n860
  );


  buf
  g1540
  (
    n1310,
    n898
  );


  buf
  g1541
  (
    n1413,
    n912
  );


  buf
  g1542
  (
    n1899,
    n844
  );


  buf
  g1543
  (
    n1818,
    n805
  );


  buf
  g1544
  (
    n1687,
    n1014
  );


  buf
  g1545
  (
    n1799,
    n867
  );


  buf
  g1546
  (
    n1118,
    n851
  );


  not
  g1547
  (
    n1572,
    n818
  );


  not
  g1548
  (
    n1277,
    n904
  );


  not
  g1549
  (
    n1908,
    n956
  );


  not
  g1550
  (
    n1382,
    n979
  );


  buf
  g1551
  (
    n1824,
    n960
  );


  not
  g1552
  (
    n1057,
    n1002
  );


  buf
  g1553
  (
    n1238,
    n833
  );


  buf
  g1554
  (
    n1864,
    n890
  );


  not
  g1555
  (
    n1834,
    n915
  );


  not
  g1556
  (
    n1364,
    n813
  );


  buf
  g1557
  (
    n1882,
    n946
  );


  buf
  g1558
  (
    n1765,
    n884
  );


  not
  g1559
  (
    n1501,
    n965
  );


  not
  g1560
  (
    n1329,
    n959
  );


  not
  g1561
  (
    n1194,
    n954
  );


  not
  g1562
  (
    n1921,
    n937
  );


  buf
  g1563
  (
    n1724,
    n897
  );


  not
  g1564
  (
    n1631,
    n975
  );


  buf
  g1565
  (
    n1037,
    n855
  );


  buf
  g1566
  (
    n1163,
    n991
  );


  buf
  g1567
  (
    n1468,
    n808
  );


  buf
  g1568
  (
    n1609,
    n887
  );


  not
  g1569
  (
    n1643,
    n818
  );


  not
  g1570
  (
    n1131,
    n919
  );


  buf
  g1571
  (
    n1678,
    n972
  );


  not
  g1572
  (
    n1542,
    n984
  );


  not
  g1573
  (
    n1129,
    n978
  );


  not
  g1574
  (
    n1121,
    n853
  );


  buf
  g1575
  (
    n1931,
    n1006
  );


  not
  g1576
  (
    n1868,
    n964
  );


  buf
  g1577
  (
    n1798,
    n798
  );


  buf
  g1578
  (
    n1295,
    n871
  );


  not
  g1579
  (
    n1181,
    n891
  );


  not
  g1580
  (
    n1917,
    n994
  );


  buf
  g1581
  (
    n1153,
    n963
  );


  not
  g1582
  (
    n1437,
    n965
  );


  buf
  g1583
  (
    n1374,
    n912
  );


  not
  g1584
  (
    n1209,
    n803
  );


  buf
  g1585
  (
    n1768,
    n880
  );


  not
  g1586
  (
    n1804,
    n978
  );


  buf
  g1587
  (
    n1681,
    n977
  );


  not
  g1588
  (
    n1188,
    n868
  );


  buf
  g1589
  (
    n1271,
    n914
  );


  buf
  g1590
  (
    n1538,
    n954
  );


  buf
  g1591
  (
    n1718,
    n863
  );


  not
  g1592
  (
    n1063,
    n913
  );


  buf
  g1593
  (
    n1377,
    n855
  );


  not
  g1594
  (
    n1741,
    n1031
  );


  buf
  g1595
  (
    n1411,
    n941
  );


  not
  g1596
  (
    n1672,
    n909
  );


  not
  g1597
  (
    n1312,
    n953
  );


  buf
  g1598
  (
    n1897,
    n958
  );


  not
  g1599
  (
    n1863,
    n871
  );


  not
  g1600
  (
    n1444,
    n866
  );


  not
  g1601
  (
    n1627,
    n969
  );


  buf
  g1602
  (
    n1755,
    n967
  );


  buf
  g1603
  (
    n1537,
    n860
  );


  not
  g1604
  (
    n1607,
    n794
  );


  not
  g1605
  (
    n1888,
    n1033
  );


  not
  g1606
  (
    n1355,
    n852
  );


  not
  g1607
  (
    n1792,
    n820
  );


  not
  g1608
  (
    n1478,
    n796
  );


  not
  g1609
  (
    n1127,
    n895
  );


  not
  g1610
  (
    n1093,
    n999
  );


  buf
  g1611
  (
    n1682,
    n880
  );


  buf
  g1612
  (
    n1811,
    n971
  );


  not
  g1613
  (
    n1378,
    n964
  );


  buf
  g1614
  (
    n1472,
    n949
  );


  not
  g1615
  (
    n1300,
    n872
  );


  not
  g1616
  (
    n1751,
    n903
  );


  buf
  g1617
  (
    n1632,
    n900
  );


  buf
  g1618
  (
    n1676,
    n898
  );


  buf
  g1619
  (
    n1461,
    n932
  );


  buf
  g1620
  (
    n1808,
    n843
  );


  not
  g1621
  (
    n1215,
    n904
  );


  buf
  g1622
  (
    n1748,
    n921
  );


  buf
  g1623
  (
    n1351,
    n939
  );


  buf
  g1624
  (
    n1169,
    n935
  );


  not
  g1625
  (
    n1399,
    n1033
  );


  not
  g1626
  (
    n1665,
    n804
  );


  not
  g1627
  (
    n1574,
    n874
  );


  not
  g1628
  (
    n1224,
    n815
  );


  buf
  g1629
  (
    n1342,
    n905
  );


  not
  g1630
  (
    n1838,
    n824
  );


  not
  g1631
  (
    n1841,
    n955
  );


  not
  g1632
  (
    n1597,
    n960
  );


  not
  g1633
  (
    n1757,
    n1032
  );


  buf
  g1634
  (
    n1714,
    n913
  );


  buf
  g1635
  (
    n1058,
    n1021
  );


  not
  g1636
  (
    n1584,
    n1002
  );


  not
  g1637
  (
    n1523,
    n803
  );


  not
  g1638
  (
    n1208,
    n881
  );


  buf
  g1639
  (
    n1878,
    n925
  );


  not
  g1640
  (
    n1723,
    n869
  );


  not
  g1641
  (
    n1119,
    n934
  );


  buf
  g1642
  (
    n1544,
    n895
  );


  buf
  g1643
  (
    n1115,
    n878
  );


  not
  g1644
  (
    n1287,
    n908
  );


  buf
  g1645
  (
    n1315,
    n992
  );


  not
  g1646
  (
    n1471,
    n917
  );


  not
  g1647
  (
    n1370,
    n954
  );


  not
  g1648
  (
    n1869,
    n1013
  );


  not
  g1649
  (
    n1430,
    n837
  );


  buf
  g1650
  (
    n1504,
    n800
  );


  buf
  g1651
  (
    n1662,
    n808
  );


  not
  g1652
  (
    n1267,
    n976
  );


  not
  g1653
  (
    n1699,
    n980
  );


  buf
  g1654
  (
    n1599,
    n1015
  );


  not
  g1655
  (
    n1133,
    n903
  );


  not
  g1656
  (
    n1337,
    n950
  );


  buf
  g1657
  (
    n1710,
    n937
  );


  not
  g1658
  (
    n1700,
    n944
  );


  not
  g1659
  (
    n1459,
    n893
  );


  buf
  g1660
  (
    n1527,
    n816
  );


  buf
  g1661
  (
    n1070,
    n917
  );


  buf
  g1662
  (
    n1909,
    n827
  );


  buf
  g1663
  (
    n1707,
    n972
  );


  not
  g1664
  (
    n1443,
    n1015
  );


  buf
  g1665
  (
    n1206,
    n894
  );


  buf
  g1666
  (
    n1422,
    n806
  );


  buf
  g1667
  (
    n1306,
    n988
  );


  buf
  g1668
  (
    n1174,
    n869
  );


  not
  g1669
  (
    n1683,
    n875
  );


  buf
  g1670
  (
    n1307,
    n894
  );


  not
  g1671
  (
    n1705,
    n909
  );


  not
  g1672
  (
    n1146,
    n967
  );


  not
  g1673
  (
    n1668,
    n832
  );


  not
  g1674
  (
    n1222,
    n800
  );


  buf
  g1675
  (
    n1516,
    n952
  );


  not
  g1676
  (
    n1319,
    n883
  );


  buf
  g1677
  (
    n1225,
    n957
  );


  buf
  g1678
  (
    n1083,
    n834
  );


  buf
  g1679
  (
    n1667,
    n819
  );


  not
  g1680
  (
    n1684,
    n973
  );


  buf
  g1681
  (
    n1595,
    n995
  );


  not
  g1682
  (
    n1419,
    n941
  );


  buf
  g1683
  (
    n1361,
    n932
  );


  buf
  g1684
  (
    n1078,
    n891
  );


  not
  g1685
  (
    n1475,
    n989
  );


  not
  g1686
  (
    n1780,
    n908
  );


  buf
  g1687
  (
    n1226,
    n836
  );


  not
  g1688
  (
    n1919,
    n850
  );


  buf
  g1689
  (
    n1220,
    n912
  );


  buf
  g1690
  (
    n1738,
    n803
  );


  buf
  g1691
  (
    n1767,
    n851
  );


  buf
  g1692
  (
    n1213,
    n794
  );


  buf
  g1693
  (
    n1819,
    n913
  );


  not
  g1694
  (
    n1641,
    n975
  );


  not
  g1695
  (
    n1143,
    n934
  );


  not
  g1696
  (
    n1454,
    n814
  );


  buf
  g1697
  (
    n1618,
    n845
  );


  buf
  g1698
  (
    n1331,
    n832
  );


  not
  g1699
  (
    n1136,
    n882
  );


  buf
  g1700
  (
    n1187,
    n897
  );


  not
  g1701
  (
    n1701,
    n906
  );


  not
  g1702
  (
    n1203,
    n996
  );


  not
  g1703
  (
    n1231,
    n831
  );


  not
  g1704
  (
    n1839,
    n829
  );


  buf
  g1705
  (
    n1829,
    n905
  );


  buf
  g1706
  (
    n1541,
    n858
  );


  buf
  g1707
  (
    n1520,
    n913
  );


  not
  g1708
  (
    n1894,
    n956
  );


  not
  g1709
  (
    n1470,
    n927
  );


  buf
  g1710
  (
    n1615,
    n838
  );


  not
  g1711
  (
    n1828,
    n959
  );


  not
  g1712
  (
    n1802,
    n981
  );


  not
  g1713
  (
    n1889,
    n867
  );


  not
  g1714
  (
    n1175,
    n900
  );


  buf
  g1715
  (
    n1076,
    n852
  );


  not
  g1716
  (
    n1216,
    n947
  );


  buf
  g1717
  (
    n1629,
    n797
  );


  not
  g1718
  (
    n1651,
    n889
  );


  buf
  g1719
  (
    n1067,
    n853
  );


  not
  g1720
  (
    n1840,
    n907
  );


  buf
  g1721
  (
    n1426,
    n809
  );


  not
  g1722
  (
    n1221,
    n917
  );


  not
  g1723
  (
    n1052,
    n985
  );


  not
  g1724
  (
    n1291,
    n846
  );


  buf
  g1725
  (
    n1693,
    n857
  );


  not
  g1726
  (
    n1112,
    n923
  );


  not
  g1727
  (
    n1230,
    n888
  );


  buf
  g1728
  (
    n1736,
    n872
  );


  buf
  g1729
  (
    n1585,
    n974
  );


  not
  g1730
  (
    n1535,
    n799
  );


  buf
  g1731
  (
    n1835,
    n942
  );


  not
  g1732
  (
    n1297,
    n920
  );


  buf
  g1733
  (
    n1155,
    n931
  );


  not
  g1734
  (
    n1075,
    n935
  );


  buf
  g1735
  (
    n1602,
    n1022
  );


  buf
  g1736
  (
    n1178,
    n885
  );


  not
  g1737
  (
    n1648,
    n1029
  );


  not
  g1738
  (
    n1189,
    n995
  );


  not
  g1739
  (
    n1775,
    n1005
  );


  not
  g1740
  (
    n1177,
    n839
  );


  buf
  g1741
  (
    n1823,
    n822
  );


  not
  g1742
  (
    n1902,
    n973
  );


  not
  g1743
  (
    n1098,
    n1031
  );


  not
  g1744
  (
    n1877,
    n932
  );


  not
  g1745
  (
    n1822,
    n1032
  );


  not
  g1746
  (
    n1316,
    n856
  );


  not
  g1747
  (
    n1170,
    n1024
  );


  buf
  g1748
  (
    n1072,
    n888
  );


  not
  g1749
  (
    n1345,
    n886
  );


  buf
  g1750
  (
    n1085,
    n1027
  );


  buf
  g1751
  (
    n1260,
    n831
  );


  buf
  g1752
  (
    n1379,
    n958
  );


  not
  g1753
  (
    n1132,
    n897
  );


  buf
  g1754
  (
    n1833,
    n1020
  );


  buf
  g1755
  (
    n1302,
    n893
  );


  not
  g1756
  (
    n1481,
    n798
  );


  buf
  g1757
  (
    n1141,
    n938
  );


  not
  g1758
  (
    n1576,
    n840
  );


  buf
  g1759
  (
    n1726,
    n825
  );


  not
  g1760
  (
    n1246,
    n1032
  );


  buf
  g1761
  (
    n1050,
    n981
  );


  not
  g1762
  (
    n1674,
    n918
  );


  buf
  g1763
  (
    n1594,
    n959
  );


  buf
  g1764
  (
    n1551,
    n891
  );


  not
  g1765
  (
    n1598,
    n822
  );


  not
  g1766
  (
    n1190,
    n994
  );


  buf
  g1767
  (
    n1296,
    n843
  );


  buf
  g1768
  (
    n1311,
    n817
  );


  not
  g1769
  (
    n1557,
    n797
  );


  buf
  g1770
  (
    n1498,
    n1018
  );


  buf
  g1771
  (
    n1704,
    n929
  );


  not
  g1772
  (
    n1392,
    n894
  );


  buf
  g1773
  (
    n1421,
    n922
  );


  buf
  g1774
  (
    n1320,
    n1026
  );


  buf
  g1775
  (
    n1274,
    n822
  );


  buf
  g1776
  (
    n1600,
    n877
  );


  buf
  g1777
  (
    n1809,
    n824
  );


  not
  g1778
  (
    n1812,
    n887
  );


  buf
  g1779
  (
    n1145,
    n964
  );


  not
  g1780
  (
    n1139,
    n892
  );


  buf
  g1781
  (
    n1578,
    n993
  );


  not
  g1782
  (
    n1384,
    n910
  );


  buf
  g1783
  (
    n1204,
    n981
  );


  buf
  g1784
  (
    n1729,
    n973
  );


  buf
  g1785
  (
    n1694,
    n873
  );


  not
  g1786
  (
    n1656,
    n847
  );


  not
  g1787
  (
    n1543,
    n824
  );


  buf
  g1788
  (
    n1055,
    n896
  );


  buf
  g1789
  (
    n1846,
    n802
  );


  not
  g1790
  (
    n1326,
    n980
  );


  buf
  g1791
  (
    n1866,
    n931
  );


  buf
  g1792
  (
    n1794,
    n986
  );


  buf
  g1793
  (
    n1673,
    n943
  );


  not
  g1794
  (
    n1862,
    n1001
  );


  not
  g1795
  (
    n1448,
    n826
  );


  buf
  g1796
  (
    n1322,
    n973
  );


  buf
  g1797
  (
    n1245,
    n828
  );


  buf
  g1798
  (
    n1293,
    n874
  );


  buf
  g1799
  (
    n1564,
    n1027
  );


  buf
  g1800
  (
    n1239,
    n811
  );


  not
  g1801
  (
    n1640,
    n1012
  );


  not
  g1802
  (
    n1365,
    n933
  );


  not
  g1803
  (
    n1376,
    n810
  );


  buf
  g1804
  (
    n1056,
    n928
  );


  not
  g1805
  (
    n1068,
    n983
  );


  not
  g1806
  (
    n1725,
    n996
  );


  not
  g1807
  (
    n1438,
    n815
  );


  buf
  g1808
  (
    n1893,
    n1019
  );


  buf
  g1809
  (
    n1826,
    n972
  );


  buf
  g1810
  (
    n1074,
    n857
  );


  not
  g1811
  (
    n1513,
    n991
  );


  not
  g1812
  (
    n1876,
    n927
  );


  not
  g1813
  (
    n1783,
    n952
  );


  buf
  g1814
  (
    n1680,
    n950
  );


  buf
  g1815
  (
    n1587,
    n833
  );


  not
  g1816
  (
    n1273,
    n961
  );


  not
  g1817
  (
    n1305,
    n838
  );


  not
  g1818
  (
    n1462,
    n982
  );


  not
  g1819
  (
    n1264,
    n948
  );


  buf
  g1820
  (
    n1849,
    n873
  );


  buf
  g1821
  (
    n1727,
    n1026
  );


  buf
  g1822
  (
    n1695,
    n865
  );


  not
  g1823
  (
    n1486,
    n1031
  );


  buf
  g1824
  (
    n1753,
    n855
  );


  not
  g1825
  (
    n1257,
    n797
  );


  buf
  g1826
  (
    n1782,
    n856
  );


  not
  g1827
  (
    n1490,
    n989
  );


  buf
  g1828
  (
    n1580,
    n878
  );


  buf
  g1829
  (
    n1559,
    n206
  );


  buf
  g1830
  (
    n1500,
    n1009
  );


  not
  g1831
  (
    n1507,
    n876
  );


  buf
  g1832
  (
    n1528,
    n969
  );


  not
  g1833
  (
    n1614,
    n888
  );


  not
  g1834
  (
    n1509,
    n923
  );


  buf
  g1835
  (
    n1610,
    n856
  );


  buf
  g1836
  (
    n1447,
    n871
  );


  not
  g1837
  (
    n1820,
    n864
  );


  buf
  g1838
  (
    n1144,
    n825
  );


  buf
  g1839
  (
    n1198,
    n858
  );


  buf
  g1840
  (
    n1357,
    n1027
  );


  buf
  g1841
  (
    n1047,
    n970
  );


  buf
  g1842
  (
    n1060,
    n894
  );


  not
  g1843
  (
    n1512,
    n809
  );


  buf
  g1844
  (
    n1396,
    n886
  );


  buf
  g1845
  (
    n1586,
    n934
  );


  not
  g1846
  (
    n1436,
    n832
  );


  buf
  g1847
  (
    n1912,
    n1017
  );


  buf
  g1848
  (
    n1560,
    n1004
  );


  not
  g1849
  (
    n1084,
    n987
  );


  not
  g1850
  (
    n1079,
    n990
  );


  buf
  g1851
  (
    n1159,
    n1023
  );


  not
  g1852
  (
    n1847,
    n820
  );


  buf
  g1853
  (
    n1335,
    n1011
  );


  buf
  g1854
  (
    n1771,
    n1017
  );


  buf
  g1855
  (
    n1843,
    n883
  );


  buf
  g1856
  (
    n1596,
    n801
  );


  buf
  g1857
  (
    n1626,
    n938
  );


  not
  g1858
  (
    n1249,
    n1011
  );


  not
  g1859
  (
    n1371,
    n911
  );


  buf
  g1860
  (
    n1636,
    n799
  );


  not
  g1861
  (
    n1646,
    n877
  );


  not
  g1862
  (
    n1637,
    n865
  );


  not
  g1863
  (
    n1619,
    n807
  );


  not
  g1864
  (
    n1282,
    n927
  );


  buf
  g1865
  (
    n1185,
    n975
  );


  not
  g1866
  (
    n1515,
    n880
  );


  nor
  g1867
  (
    n1493,
    n970,
    n854,
    n922
  );


  and
  g1868
  (
    n1549,
    n882,
    n902,
    n851
  );


  nand
  g1869
  (
    n1427,
    n984,
    n975,
    n905
  );


  nand
  g1870
  (
    n1200,
    n1018,
    n795,
    n871
  );


  nand
  g1871
  (
    n1920,
    n1007,
    n873,
    n1016
  );


  or
  g1872
  (
    n1048,
    n853,
    n817,
    n948
  );


  nor
  g1873
  (
    n1266,
    n875,
    n809,
    n830
  );


  xor
  g1874
  (
    n1110,
    n992,
    n879,
    n918
  );


  nor
  g1875
  (
    n1338,
    n1023,
    n860,
    n979
  );


  or
  g1876
  (
    n1850,
    n929,
    n205,
    n935
  );


  or
  g1877
  (
    n1064,
    n860,
    n1029,
    n904
  );


  nor
  g1878
  (
    n1506,
    n915,
    n899,
    n1030
  );


  xnor
  g1879
  (
    n1918,
    n1019,
    n805,
    n974
  );


  and
  g1880
  (
    n1400,
    n883,
    n864,
    n794
  );


  xnor
  g1881
  (
    n1914,
    n944,
    n915,
    n890
  );


  xnor
  g1882
  (
    n1383,
    n859,
    n206,
    n1025
  );


  and
  g1883
  (
    n1892,
    n1025,
    n862,
    n875
  );


  xor
  g1884
  (
    n1604,
    n999,
    n813,
    n962
  );


  or
  g1885
  (
    n1275,
    n1005,
    n828,
    n910
  );


  and
  g1886
  (
    n1476,
    n867,
    n937,
    n970
  );


  xor
  g1887
  (
    n1633,
    n810,
    n838,
    n977
  );


  xnor
  g1888
  (
    n1696,
    n802,
    n1009,
    n811
  );


  nor
  g1889
  (
    n1261,
    n859,
    n936,
    n977
  );


  or
  g1890
  (
    n1045,
    n801,
    n962,
    n957
  );


  xnor
  g1891
  (
    n1407,
    n807,
    n817,
    n1016
  );


  or
  g1892
  (
    n1744,
    n923,
    n962,
    n906
  );


  nand
  g1893
  (
    n1073,
    n842,
    n810
  );


  and
  g1894
  (
    n1722,
    n931,
    n977,
    n858
  );


  nand
  g1895
  (
    n1813,
    n837,
    n982,
    n954
  );


  nand
  g1896
  (
    n1044,
    n993,
    n906,
    n849
  );


  nor
  g1897
  (
    n1883,
    n987,
    n821,
    n942
  );


  xnor
  g1898
  (
    n1173,
    n807,
    n1029,
    n933
  );


  xnor
  g1899
  (
    n1495,
    n870,
    n926,
    n1024,
    n806
  );


  xor
  g1900
  (
    n2084,
    n1082,
    n1186,
    n1735
  );


  xor
  g1901
  (
    n2244,
    n1659,
    n1156,
    n1437,
    n1417
  );


  nand
  g1902
  (
    n2697,
    n1146,
    n1399,
    n1220,
    n1585
  );


  xor
  g1903
  (
    n2397,
    n1346,
    n1281,
    n1656,
    n1185
  );


  or
  g1904
  (
    n2711,
    n1103,
    n1732,
    n1120,
    n1076
  );


  xnor
  g1905
  (
    n2615,
    n1807,
    n1358,
    n1336,
    n1266
  );


  xnor
  g1906
  (
    n2309,
    n1178,
    n1188,
    n1176,
    n1706
  );


  or
  g1907
  (
    n2398,
    n1324,
    n1783,
    n1795,
    n1694
  );


  or
  g1908
  (
    n2435,
    n1230,
    n1742,
    n1763,
    n1535
  );


  or
  g1909
  (
    n1938,
    n1166,
    n1125,
    n1423,
    n1208
  );


  nor
  g1910
  (
    n2195,
    n1067,
    n1677,
    n1571,
    n1311
  );


  xor
  g1911
  (
    n2692,
    n1062,
    n1739,
    n1795,
    n1451
  );


  nand
  g1912
  (
    n2015,
    n1661,
    n1455,
    n1382,
    n1192
  );


  or
  g1913
  (
    n2274,
    n1169,
    n1534,
    n1712,
    n1422
  );


  xnor
  g1914
  (
    n2667,
    n1075,
    n1179,
    n1771,
    n1346
  );


  nand
  g1915
  (
    n2461,
    n1352,
    n1545,
    n1195,
    n1085
  );


  xnor
  g1916
  (
    n1992,
    n1080,
    n1734,
    n1751,
    n1321
  );


  xor
  g1917
  (
    n2108,
    n1247,
    n1410,
    n1427,
    n1531
  );


  or
  g1918
  (
    n2634,
    n1777,
    n1598,
    n1190,
    n1352
  );


  and
  g1919
  (
    n2395,
    n1604,
    n1220,
    n1675,
    n1124
  );


  xor
  g1920
  (
    n2064,
    n1038,
    n1422,
    n1465,
    n1775
  );


  and
  g1921
  (
    n2591,
    n1513,
    n1250,
    n1563,
    n1369
  );


  nor
  g1922
  (
    n1956,
    n1314,
    n1760,
    n1761,
    n1521
  );


  or
  g1923
  (
    n2059,
    n1774,
    n1188,
    n1418,
    n1757
  );


  nand
  g1924
  (
    n1975,
    n1625,
    n1169,
    n1395,
    n1663
  );


  and
  g1925
  (
    n2500,
    n1601,
    n1734,
    n1496,
    n1568
  );


  nand
  g1926
  (
    n2463,
    n1345,
    n1063,
    n1387,
    n1343
  );


  xnor
  g1927
  (
    n2297,
    n1302,
    n1574,
    n1060,
    n1350
  );


  or
  g1928
  (
    n2004,
    n1493,
    n1064,
    n1375,
    n1357
  );


  xor
  g1929
  (
    n2608,
    n1583,
    n1653,
    n1678,
    n1652
  );


  nor
  g1930
  (
    n2504,
    n1184,
    n1402,
    n1610,
    n1651
  );


  or
  g1931
  (
    n2536,
    n1722,
    n1042,
    n1263,
    n1100
  );


  xor
  g1932
  (
    n2329,
    n1713,
    n1339,
    n1401,
    n1649
  );


  or
  g1933
  (
    n2558,
    n1802,
    n1136,
    n1037,
    n1631
  );


  xor
  g1934
  (
    n2382,
    n1615,
    n1390,
    n1593,
    n1808
  );


  xor
  g1935
  (
    n2164,
    n1264,
    n1260,
    n1764,
    n1378
  );


  and
  g1936
  (
    n2386,
    n1265,
    n1454,
    n1198,
    n1039
  );


  nor
  g1937
  (
    n2285,
    n1479,
    n1473,
    n1302,
    n1203
  );


  nand
  g1938
  (
    n2264,
    n1380,
    n1574,
    n1576,
    n1351
  );


  xor
  g1939
  (
    n2013,
    n1391,
    n1787,
    n1256,
    n1561
  );


  xor
  g1940
  (
    n2054,
    n1652,
    n1773,
    n1072,
    n1551
  );


  and
  g1941
  (
    n2073,
    n1334,
    n1495,
    n1534,
    n1369
  );


  or
  g1942
  (
    n2121,
    n1109,
    n1519,
    n1779,
    n1811
  );


  xnor
  g1943
  (
    n2646,
    n1555,
    n1676,
    n1049,
    n1587
  );


  or
  g1944
  (
    n2304,
    n1799,
    n1543,
    n1444,
    n1148
  );


  xor
  g1945
  (
    n2036,
    n1558,
    n1773,
    n1578,
    n1241
  );


  xor
  g1946
  (
    n2700,
    n1104,
    n1575,
    n1442,
    n1165
  );


  nor
  g1947
  (
    n2277,
    n1072,
    n1558,
    n1272,
    n1532
  );


  or
  g1948
  (
    n2431,
    n1703,
    n1488,
    n1424,
    n1101
  );


  xor
  g1949
  (
    n2506,
    n1759,
    n1358,
    n1168,
    n1098
  );


  nor
  g1950
  (
    n2550,
    n1112,
    n1433,
    n1051,
    n1742
  );


  xor
  g1951
  (
    n2189,
    n1484,
    n1274,
    n1053,
    n1648
  );


  nand
  g1952
  (
    n2203,
    n1132,
    n1233,
    n1609,
    n1653
  );


  xor
  g1953
  (
    n2284,
    n1151,
    n1544,
    n1228,
    n1066
  );


  or
  g1954
  (
    n2582,
    n1277,
    n1465,
    n1720,
    n1252
  );


  nand
  g1955
  (
    n2460,
    n1702,
    n1660,
    n1177,
    n1300
  );


  nor
  g1956
  (
    n2633,
    n1528,
    n1406,
    n1525,
    n1124
  );


  nand
  g1957
  (
    n2508,
    n1528,
    n1294,
    n1290,
    n1092
  );


  xor
  g1958
  (
    n2464,
    n1420,
    n1171,
    n1224,
    n1239
  );


  xnor
  g1959
  (
    n2282,
    n1562,
    n1584,
    n1489,
    n1154
  );


  and
  g1960
  (
    n2450,
    n1749,
    n1274,
    n1679,
    n1547
  );


  and
  g1961
  (
    n2167,
    n1636,
    n1448,
    n1769,
    n1625
  );


  nor
  g1962
  (
    n2596,
    n1074,
    n1787,
    n1442,
    n1622
  );


  xnor
  g1963
  (
    n2628,
    n1350,
    n1473,
    n1323,
    n1393
  );


  xor
  g1964
  (
    n2131,
    n1511,
    n1689,
    n1272,
    n1095
  );


  nor
  g1965
  (
    n2622,
    n1740,
    n1626,
    n1596,
    n1756
  );


  or
  g1966
  (
    n2410,
    n1556,
    n1097,
    n1748,
    n1034
  );


  nor
  g1967
  (
    n1987,
    n1683,
    n1532,
    n1563,
    n1799
  );


  nor
  g1968
  (
    n2241,
    n1642,
    n1335,
    n1595,
    n1500
  );


  and
  g1969
  (
    n2002,
    n1809,
    n1198,
    n1329,
    n1776
  );


  nor
  g1970
  (
    n2128,
    n1097,
    n1524,
    n1348,
    n1446
  );


  or
  g1971
  (
    n2540,
    n1754,
    n1499,
    n1758,
    n1716
  );


  or
  g1972
  (
    n2296,
    n1048,
    n1428,
    n1274,
    n1493
  );


  nor
  g1973
  (
    n2000,
    n1476,
    n1267,
    n1123,
    n1303
  );


  or
  g1974
  (
    n2513,
    n1543,
    n1260,
    n1212,
    n1470
  );


  nor
  g1975
  (
    n2173,
    n1401,
    n1405,
    n1625,
    n1301
  );


  and
  g1976
  (
    n2486,
    n1781,
    n1608,
    n1584,
    n1783
  );


  xnor
  g1977
  (
    n1937,
    n1110,
    n1452,
    n1475,
    n1180
  );


  and
  g1978
  (
    n2141,
    n1441,
    n1785,
    n1774,
    n1810
  );


  or
  g1979
  (
    n2246,
    n1318,
    n1586,
    n1441,
    n1699
  );


  nor
  g1980
  (
    n2401,
    n1651,
    n1306,
    n1072,
    n1333
  );


  xnor
  g1981
  (
    n2368,
    n1328,
    n1379,
    n1275,
    n1711
  );


  xor
  g1982
  (
    n2010,
    n1500,
    n1328,
    n1333,
    n1107
  );


  nor
  g1983
  (
    n2514,
    n1338,
    n1224,
    n1214,
    n1755
  );


  or
  g1984
  (
    n2299,
    n1753,
    n1132,
    n1529,
    n1645
  );


  nand
  g1985
  (
    n2685,
    n1608,
    n1287,
    n1659,
    n1719
  );


  xor
  g1986
  (
    n2288,
    n1514,
    n1668,
    n1508
  );


  and
  g1987
  (
    n2447,
    n1436,
    n1414,
    n1622,
    n1555
  );


  or
  g1988
  (
    n2367,
    n1768,
    n1046,
    n1609,
    n1623
  );


  nor
  g1989
  (
    n2592,
    n1232,
    n1541,
    n1315,
    n1106
  );


  nand
  g1990
  (
    n2116,
    n1067,
    n1232,
    n1327,
    n1757
  );


  xnor
  g1991
  (
    n2194,
    n1197,
    n1763,
    n1693,
    n1092
  );


  nand
  g1992
  (
    n2370,
    n1607,
    n1603,
    n1399,
    n1778
  );


  and
  g1993
  (
    n2267,
    n1572,
    n1811,
    n1059,
    n1470
  );


  and
  g1994
  (
    n1952,
    n1035,
    n1092,
    n1405,
    n1649
  );


  and
  g1995
  (
    n2130,
    n1749,
    n1679,
    n1776,
    n1638
  );


  nand
  g1996
  (
    n2125,
    n1691,
    n1622,
    n1069,
    n1088
  );


  xnor
  g1997
  (
    n1953,
    n1692,
    n1797,
    n1071,
    n1058
  );


  or
  g1998
  (
    n1978,
    n1666,
    n1808,
    n1597,
    n1081
  );


  nand
  g1999
  (
    n2146,
    n1188,
    n1498,
    n1283,
    n1211
  );


  xnor
  g2000
  (
    n2122,
    n1335,
    n1380,
    n1141,
    n1392
  );


  xnor
  g2001
  (
    n2415,
    n1223,
    n1668,
    n1542,
    n1132
  );


  and
  g2002
  (
    n2567,
    n1525,
    n1313,
    n1720,
    n1674
  );


  or
  g2003
  (
    n1970,
    n1554,
    n1644,
    n1076,
    n1738
  );


  xnor
  g2004
  (
    n2623,
    n1633,
    n1783,
    n1577,
    n1699
  );


  or
  g2005
  (
    n2377,
    n1323,
    n1185,
    n1251,
    n1504
  );


  and
  g2006
  (
    n2494,
    n1223,
    n1312,
    n1447,
    n1416
  );


  or
  g2007
  (
    n2616,
    n1173,
    n1172,
    n1094,
    n1405
  );


  nand
  g2008
  (
    n2578,
    n1049,
    n1188,
    n1166,
    n1327
  );


  nor
  g2009
  (
    n2559,
    n1299,
    n1643,
    n1616,
    n1763
  );


  nand
  g2010
  (
    n2156,
    n1111,
    n1759,
    n1151,
    n1413
  );


  or
  g2011
  (
    n2318,
    n1662,
    n1562,
    n1714,
    n1812
  );


  and
  g2012
  (
    n2373,
    n1406,
    n1371,
    n1209,
    n1540
  );


  nand
  g2013
  (
    n2477,
    n1549,
    n1372,
    n1531,
    n1581
  );


  nor
  g2014
  (
    n2242,
    n1345,
    n1687,
    n1083,
    n1144
  );


  nor
  g2015
  (
    n2154,
    n1156,
    n1294,
    n1431,
    n1552
  );


  xnor
  g2016
  (
    n1982,
    n1467,
    n1304,
    n1317,
    n1348
  );


  nand
  g2017
  (
    n1983,
    n1586,
    n1094,
    n1637,
    n1269
  );


  or
  g2018
  (
    n1996,
    n1358,
    n1284,
    n1502,
    n1483
  );


  xor
  g2019
  (
    n2570,
    n1733,
    n1137,
    n1627,
    n1322
  );


  xnor
  g2020
  (
    n2606,
    n1702,
    n1326,
    n1655,
    n1090
  );


  nand
  g2021
  (
    n2511,
    n1527,
    n1798,
    n1170,
    n1066
  );


  or
  g2022
  (
    n2519,
    n1526,
    n1801,
    n1265,
    n207
  );


  xnor
  g2023
  (
    n2038,
    n1489,
    n1628,
    n1313,
    n1302
  );


  nand
  g2024
  (
    n2594,
    n1393,
    n1181,
    n1349,
    n1670
  );


  xor
  g2025
  (
    n2200,
    n1047,
    n1571,
    n1428,
    n1359
  );


  nand
  g2026
  (
    n2201,
    n1497,
    n1548,
    n1696,
    n1754
  );


  xnor
  g2027
  (
    n2308,
    n1043,
    n1080,
    n1787,
    n1636
  );


  nor
  g2028
  (
    n2351,
    n1114,
    n1400,
    n1781,
    n1534
  );


  and
  g2029
  (
    n2483,
    n1535,
    n1716,
    n1428,
    n1644
  );


  xor
  g2030
  (
    n2019,
    n1241,
    n1096,
    n1572,
    n1417
  );


  and
  g2031
  (
    n2380,
    n1340,
    n1042,
    n1136,
    n1270
  );


  xnor
  g2032
  (
    n2071,
    n1146,
    n1129,
    n1087,
    n1235
  );


  or
  g2033
  (
    n2181,
    n1582,
    n1320,
    n1161,
    n1581
  );


  xor
  g2034
  (
    n2509,
    n1561,
    n1054,
    n1207,
    n1648
  );


  and
  g2035
  (
    n2683,
    n1206,
    n1162,
    n1139,
    n1343
  );


  or
  g2036
  (
    n2432,
    n1123,
    n1485,
    n1448,
    n1529
  );


  xnor
  g2037
  (
    n2003,
    n1453,
    n1727,
    n1170,
    n1382
  );


  and
  g2038
  (
    n2466,
    n1193,
    n1201,
    n1115,
    n1399
  );


  and
  g2039
  (
    n2429,
    n1622,
    n1039,
    n1720,
    n1271
  );


  nand
  g2040
  (
    n2114,
    n1790,
    n1532,
    n1788,
    n1231
  );


  and
  g2041
  (
    n2406,
    n1397,
    n1464,
    n1388,
    n1443
  );


  nor
  g2042
  (
    n2037,
    n1505,
    n1284,
    n1048,
    n1740
  );


  nand
  g2043
  (
    n2340,
    n1583,
    n1665,
    n1139,
    n1035
  );


  or
  g2044
  (
    n2497,
    n1458,
    n1225,
    n1758,
    n1436
  );


  and
  g2045
  (
    n2222,
    n1593,
    n1557,
    n1349,
    n1548
  );


  or
  g2046
  (
    n2074,
    n1615,
    n1635,
    n1769,
    n1459
  );


  nor
  g2047
  (
    n2310,
    n1214,
    n1580,
    n1745,
    n1194
  );


  xnor
  g2048
  (
    n2279,
    n1719,
    n1507,
    n1376,
    n1313
  );


  xnor
  g2049
  (
    n2488,
    n1064,
    n1662,
    n1271,
    n1377
  );


  xor
  g2050
  (
    n2350,
    n1672,
    n1367,
    n1756,
    n1093
  );


  or
  g2051
  (
    n2110,
    n1399,
    n1419,
    n1598,
    n1062
  );


  xnor
  g2052
  (
    n2694,
    n1318,
    n1468,
    n1400,
    n1577
  );


  and
  g2053
  (
    n2672,
    n1461,
    n1189,
    n1069,
    n1467
  );


  and
  g2054
  (
    n1990,
    n1568,
    n1796,
    n1243,
    n1540
  );


  nor
  g2055
  (
    n1967,
    n1409,
    n1531,
    n1173,
    n1190
  );


  nand
  g2056
  (
    n2365,
    n1626,
    n1698,
    n1630,
    n1497
  );


  nor
  g2057
  (
    n2276,
    n1395,
    n1071,
    n1630,
    n1761
  );


  nand
  g2058
  (
    n2040,
    n1354,
    n1062,
    n1111,
    n1640
  );


  xor
  g2059
  (
    n2046,
    n1454,
    n1707,
    n1342,
    n1482
  );


  nand
  g2060
  (
    n2053,
    n1363,
    n1303,
    n1357,
    n1569
  );


  or
  g2061
  (
    n1965,
    n1375,
    n1283,
    n1455,
    n1110
  );


  xnor
  g2062
  (
    n2171,
    n1721,
    n1138,
    n1656,
    n1248
  );


  xor
  g2063
  (
    n1991,
    n1495,
    n1639,
    n1263,
    n1529
  );


  or
  g2064
  (
    n2357,
    n1145,
    n1328,
    n1370,
    n1122
  );


  xnor
  g2065
  (
    n2078,
    n1465,
    n1088,
    n1716,
    n1404
  );


  xnor
  g2066
  (
    n2187,
    n1213,
    n1619,
    n1217,
    n1485
  );


  or
  g2067
  (
    n2058,
    n1492,
    n1121,
    n1076,
    n1212
  );


  nor
  g2068
  (
    n2233,
    n1793,
    n1181,
    n1654,
    n1202
  );


  and
  g2069
  (
    n2144,
    n1481,
    n1106,
    n1259,
    n1053
  );


  nor
  g2070
  (
    n2600,
    n1114,
    n1353,
    n1129,
    n1766
  );


  and
  g2071
  (
    n2521,
    n1700,
    n1550,
    n1088,
    n1295
  );


  or
  g2072
  (
    n2707,
    n1731,
    n1699,
    n1714,
    n1055
  );


  xnor
  g2073
  (
    n2556,
    n1759,
    n1527,
    n1273,
    n1376
  );


  and
  g2074
  (
    n2027,
    n1486,
    n1566,
    n1180,
    n1084
  );


  xnor
  g2075
  (
    n2321,
    n1448,
    n1548,
    n1582,
    n1517
  );


  nand
  g2076
  (
    n2314,
    n1639,
    n1533,
    n1715,
    n1695
  );


  nor
  g2077
  (
    n2315,
    n1431,
    n1116,
    n1404,
    n1080
  );


  or
  g2078
  (
    n2664,
    n1713,
    n1330,
    n1681,
    n1496
  );


  nand
  g2079
  (
    n2192,
    n1724,
    n1729,
    n1230,
    n1163
  );


  and
  g2080
  (
    n2434,
    n1711,
    n1340,
    n1723,
    n1232
  );


  xnor
  g2081
  (
    n1933,
    n1794,
    n1619,
    n1070,
    n1307
  );


  nor
  g2082
  (
    n2176,
    n1592,
    n1785,
    n1209,
    n1649
  );


  or
  g2083
  (
    n2327,
    n1553,
    n1118,
    n1121,
    n1152
  );


  or
  g2084
  (
    n2455,
    n1202,
    n1653,
    n1425,
    n1694
  );


  xor
  g2085
  (
    n2115,
    n1392,
    n1726,
    n1383,
    n1524
  );


  xor
  g2086
  (
    n2501,
    n1466,
    n1771,
    n1046,
    n1698
  );


  nor
  g2087
  (
    n2618,
    n1752,
    n1045,
    n1200,
    n1124
  );


  xnor
  g2088
  (
    n2089,
    n1471,
    n1526,
    n1595,
    n1470
  );


  xor
  g2089
  (
    n2405,
    n1199,
    n1585,
    n1486,
    n1398
  );


  and
  g2090
  (
    n2095,
    n1749,
    n1486,
    n1772,
    n1100
  );


  nand
  g2091
  (
    n2641,
    n1252,
    n1598,
    n1370,
    n207
  );


  xor
  g2092
  (
    n2021,
    n1180,
    n1275,
    n1704,
    n207
  );


  or
  g2093
  (
    n2030,
    n1337,
    n1567,
    n1252,
    n1181
  );


  xor
  g2094
  (
    n2665,
    n1278,
    n1266,
    n1364,
    n1708
  );


  xor
  g2095
  (
    n2290,
    n1035,
    n1682,
    n1095,
    n1124
  );


  and
  g2096
  (
    n2417,
    n1314,
    n1353,
    n1292,
    n1182
  );


  or
  g2097
  (
    n2298,
    n1127,
    n1246,
    n1638,
    n1089
  );


  or
  g2098
  (
    n2348,
    n1728,
    n1097,
    n1311,
    n1058
  );


  nor
  g2099
  (
    n1943,
    n1688,
    n1384,
    n1202,
    n1061
  );


  nor
  g2100
  (
    n2048,
    n1730,
    n1418,
    n1375,
    n1276
  );


  nand
  g2101
  (
    n2364,
    n1162,
    n1221,
    n1798,
    n1588
  );


  nor
  g2102
  (
    n2198,
    n1247,
    n1165,
    n1386,
    n1146
  );


  and
  g2103
  (
    n2081,
    n1435,
    n1775,
    n1385,
    n1737
  );


  nand
  g2104
  (
    n2250,
    n1796,
    n1403,
    n1371,
    n1730
  );


  xnor
  g2105
  (
    n2485,
    n1195,
    n1750,
    n1341,
    n1166
  );


  or
  g2106
  (
    n2433,
    n1189,
    n1426,
    n1163,
    n1128
  );


  xor
  g2107
  (
    n2462,
    n1600,
    n1704,
    n1616,
    n1772
  );


  and
  g2108
  (
    n2561,
    n1260,
    n1175,
    n1469,
    n1233
  );


  and
  g2109
  (
    n2269,
    n1500,
    n1289,
    n1547,
    n1747
  );


  xnor
  g2110
  (
    n2693,
    n1491,
    n1279,
    n1705,
    n1103
  );


  nor
  g2111
  (
    n1966,
    n1510,
    n1464,
    n1410,
    n1648
  );


  or
  g2112
  (
    n2517,
    n1248,
    n1565,
    n1200,
    n1686
  );


  and
  g2113
  (
    n2292,
    n1733,
    n1538,
    n1421,
    n1245
  );


  xnor
  g2114
  (
    n2470,
    n1604,
    n1609,
    n1658,
    n1541
  );


  nor
  g2115
  (
    n2468,
    n1257,
    n1514,
    n1606,
    n1559
  );


  and
  g2116
  (
    n2422,
    n1116,
    n1352,
    n1633,
    n1139
  );


  xnor
  g2117
  (
    n2619,
    n1158,
    n1312,
    n1620,
    n1424
  );


  and
  g2118
  (
    n2230,
    n1095,
    n1794,
    n1410,
    n1222
  );


  xnor
  g2119
  (
    n1981,
    n1147,
    n1035,
    n1766,
    n1708
  );


  nand
  g2120
  (
    n2597,
    n1255,
    n1136,
    n1283,
    n1522
  );


  or
  g2121
  (
    n2403,
    n1618,
    n1074,
    n1034,
    n1145
  );


  nand
  g2122
  (
    n2023,
    n1371,
    n1348,
    n1294,
    n1544
  );


  nand
  g2123
  (
    n2480,
    n1559,
    n1119,
    n1542,
    n1624
  );


  and
  g2124
  (
    n2101,
    n1402,
    n1789,
    n1090,
    n1728
  );


  and
  g2125
  (
    n2043,
    n1312,
    n1498,
    n1618,
    n1134
  );


  xnor
  g2126
  (
    n2695,
    n1770,
    n1242,
    n1494,
    n1244
  );


  or
  g2127
  (
    n2137,
    n1125,
    n1671,
    n1299,
    n1113
  );


  nor
  g2128
  (
    n2252,
    n1746,
    n1295,
    n1431,
    n1791
  );


  xor
  g2129
  (
    n2082,
    n1490,
    n1350,
    n1447,
    n1627
  );


  or
  g2130
  (
    n2247,
    n1434,
    n1099,
    n1417,
    n1320
  );


  and
  g2131
  (
    n2243,
    n1791,
    n1785,
    n1152,
    n1381
  );


  or
  g2132
  (
    n1936,
    n1133,
    n1080,
    n1114,
    n1258
  );


  xor
  g2133
  (
    n1957,
    n1334,
    n1475,
    n1057,
    n1114
  );


  xnor
  g2134
  (
    n2305,
    n1616,
    n1594,
    n1237,
    n30
  );


  xnor
  g2135
  (
    n2153,
    n1108,
    n1722,
    n1590,
    n1600
  );


  or
  g2136
  (
    n2272,
    n1157,
    n1324,
    n1109,
    n1050
  );


  nor
  g2137
  (
    n2202,
    n1699,
    n1782,
    n1486,
    n1503
  );


  or
  g2138
  (
    n2366,
    n1236,
    n1106,
    n1490,
    n1376
  );


  and
  g2139
  (
    n2307,
    n1246,
    n1226,
    n1108,
    n1384
  );


  nand
  g2140
  (
    n1958,
    n1740,
    n1520,
    n1499,
    n1047
  );


  nand
  g2141
  (
    n2520,
    n1667,
    n1146,
    n1050,
    n1807
  );


  nand
  g2142
  (
    n2343,
    n1045,
    n1151,
    n1512,
    n1631
  );


  or
  g2143
  (
    n2065,
    n1393,
    n1562,
    n1701,
    n1082
  );


  nor
  g2144
  (
    n2278,
    n1646,
    n1556,
    n1404,
    n1767
  );


  xnor
  g2145
  (
    n2636,
    n1531,
    n1744,
    n1073,
    n1403
  );


  or
  g2146
  (
    n2313,
    n1306,
    n1356,
    n1767,
    n1200
  );


  xor
  g2147
  (
    n2286,
    n1527,
    n1440,
    n1354,
    n1171
  );


  xnor
  g2148
  (
    n2527,
    n1102,
    n1552,
    n1279,
    n1178
  );


  nor
  g2149
  (
    n2656,
    n1420,
    n1639,
    n1319,
    n1281
  );


  xor
  g2150
  (
    n1947,
    n1253,
    n1086,
    n1204,
    n1712
  );


  xnor
  g2151
  (
    n2639,
    n1413,
    n1083,
    n30,
    n1455
  );


  xor
  g2152
  (
    n2449,
    n1650,
    n1518,
    n1780,
    n1117
  );


  nor
  g2153
  (
    n2174,
    n1330,
    n1784,
    n1329,
    n1462
  );


  xnor
  g2154
  (
    n2621,
    n1409,
    n1735,
    n1786,
    n1610
  );


  or
  g2155
  (
    n2086,
    n1750,
    n1361,
    n1656,
    n1642
  );


  xor
  g2156
  (
    n2251,
    n1580,
    n1520,
    n1794,
    n1767
  );


  or
  g2157
  (
    n2576,
    n1731,
    n1351,
    n1460,
    n1396
  );


  nor
  g2158
  (
    n2452,
    n1645,
    n1808,
    n1287,
    n1437
  );


  and
  g2159
  (
    n2360,
    n1284,
    n1276,
    n1390,
    n1508
  );


  nor
  g2160
  (
    n2706,
    n1739,
    n1074,
    n1147,
    n1496
  );


  or
  g2161
  (
    n2407,
    n1440,
    n1803,
    n1046,
    n1480
  );


  xor
  g2162
  (
    n2391,
    n1322,
    n1621,
    n1637,
    n1785
  );


  xnor
  g2163
  (
    n2162,
    n1587,
    n1446,
    n1203,
    n1065
  );


  nand
  g2164
  (
    n2522,
    n1643,
    n1700,
    n1739,
    n1483
  );


  nor
  g2165
  (
    n2443,
    n1601,
    n1712,
    n1367,
    n1130
  );


  xor
  g2166
  (
    n2336,
    n1249,
    n1613,
    n1372,
    n1652
  );


  and
  g2167
  (
    n2487,
    n1091,
    n1354,
    n1734,
    n1253
  );


  nor
  g2168
  (
    n2206,
    n1471,
    n1669,
    n1515,
    n1723
  );


  and
  g2169
  (
    n2651,
    n1178,
    n1378,
    n1245,
    n1388
  );


  nor
  g2170
  (
    n2354,
    n1333,
    n1401,
    n1509,
    n1606
  );


  xor
  g2171
  (
    n2001,
    n1496,
    n1044,
    n1355,
    n1733
  );


  xnor
  g2172
  (
    n2642,
    n1154,
    n1670,
    n1647,
    n1554
  );


  xnor
  g2173
  (
    n2635,
    n1433,
    n1569,
    n1059,
    n1636
  );


  or
  g2174
  (
    n1955,
    n1284,
    n1160,
    n1212,
    n1755
  );


  and
  g2175
  (
    n2150,
    n1752,
    n1477,
    n1220,
    n1191
  );


  and
  g2176
  (
    n2438,
    n1690,
    n1511,
    n1457,
    n1252
  );


  and
  g2177
  (
    n2547,
    n1615,
    n1384,
    n1765,
    n1149
  );


  and
  g2178
  (
    n2042,
    n1104,
    n1297,
    n1754,
    n1782
  );


  xnor
  g2179
  (
    n2177,
    n1254,
    n1323,
    n1130,
    n1729
  );


  or
  g2180
  (
    n2640,
    n1492,
    n1089,
    n1348,
    n1043
  );


  xnor
  g2181
  (
    n1940,
    n1445,
    n1203,
    n1347,
    n1308
  );


  nor
  g2182
  (
    n2257,
    n1328,
    n1161,
    n1727,
    n1478
  );


  and
  g2183
  (
    n2648,
    n1469,
    n1148,
    n1282,
    n1568
  );


  nand
  g2184
  (
    n2258,
    n1266,
    n1458,
    n1421,
    n1585
  );


  nor
  g2185
  (
    n2142,
    n1571,
    n1741,
    n1374,
    n1629
  );


  nand
  g2186
  (
    n2515,
    n1774,
    n1747,
    n1310,
    n1130
  );


  or
  g2187
  (
    n2151,
    n1754,
    n1264,
    n1630,
    n1733
  );


  xnor
  g2188
  (
    n2542,
    n1481,
    n1477,
    n1517,
    n1456
  );


  or
  g2189
  (
    n2049,
    n1594,
    n1672,
    n1810,
    n1507
  );


  xor
  g2190
  (
    n2311,
    n1153,
    n1330,
    n1617,
    n1307
  );


  or
  g2191
  (
    n2476,
    n1261,
    n1205,
    n1487,
    n1565
  );


  or
  g2192
  (
    n1968,
    n1064,
    n1131,
    n1570,
    n1492
  );


  xor
  g2193
  (
    n2317,
    n1276,
    n1233,
    n1499,
    n1682
  );


  and
  g2194
  (
    n2262,
    n1671,
    n1709,
    n1098,
    n1770
  );


  xnor
  g2195
  (
    n2524,
    n1107,
    n1193,
    n1331,
    n1387
  );


  xor
  g2196
  (
    n2041,
    n1429,
    n1349,
    n1341,
    n1418
  );


  xnor
  g2197
  (
    n2611,
    n1256,
    n1753,
    n1089,
    n1309
  );


  nand
  g2198
  (
    n2280,
    n1174,
    n1478,
    n1623,
    n1514
  );


  nor
  g2199
  (
    n2676,
    n1079,
    n1504,
    n1506,
    n1788
  );


  nor
  g2200
  (
    n1959,
    n1711,
    n1265,
    n1421,
    n1459
  );


  and
  g2201
  (
    n2179,
    n1503,
    n1613,
    n1614,
    n1408
  );


  xnor
  g2202
  (
    n2214,
    n1644,
    n1757,
    n1407,
    n1415
  );


  and
  g2203
  (
    n2421,
    n1771,
    n1708,
    n1603,
    n1129
  );


  or
  g2204
  (
    n2035,
    n1738,
    n1578,
    n1147,
    n1536
  );


  nand
  g2205
  (
    n2363,
    n1700,
    n1663,
    n1651,
    n1290
  );


  or
  g2206
  (
    n2390,
    n1383,
    n1669,
    n1762,
    n1277
  );


  xnor
  g2207
  (
    n2458,
    n1094,
    n1185,
    n1245,
    n1286
  );


  xnor
  g2208
  (
    n2579,
    n1159,
    n1489,
    n1793,
    n1336
  );


  xnor
  g2209
  (
    n2178,
    n1176,
    n1539,
    n1374,
    n1761
  );


  or
  g2210
  (
    n2068,
    n1373,
    n1108,
    n1670,
    n1047
  );


  or
  g2211
  (
    n2165,
    n1100,
    n1298,
    n1056,
    n1179
  );


  xnor
  g2212
  (
    n2045,
    n1221,
    n1451,
    n1254,
    n1466
  );


  xor
  g2213
  (
    n2669,
    n1301,
    n1153,
    n1404,
    n1257
  );


  xor
  g2214
  (
    n2496,
    n1150,
    n1512,
    n1237,
    n1362
  );


  xnor
  g2215
  (
    n2448,
    n1145,
    n1473,
    n1034,
    n1142
  );


  xor
  g2216
  (
    n2698,
    n1791,
    n1407,
    n1057,
    n1579
  );


  xor
  g2217
  (
    n2630,
    n1691,
    n1435,
    n1427,
    n1300
  );


  and
  g2218
  (
    n2238,
    n1809,
    n1261,
    n1479,
    n1459
  );


  xnor
  g2219
  (
    n2427,
    n1406,
    n1779,
    n1258,
    n1103
  );


  and
  g2220
  (
    n2529,
    n1105,
    n1084,
    n1692,
    n1627
  );


  and
  g2221
  (
    n2103,
    n1262,
    n1319,
    n1050,
    n1589
  );


  and
  g2222
  (
    n2612,
    n1034,
    n1582,
    n1610,
    n1665
  );


  nand
  g2223
  (
    n1935,
    n1784,
    n1732,
    n1331,
    n1641
  );


  nor
  g2224
  (
    n2323,
    n1250,
    n1536,
    n1322,
    n1667
  );


  nor
  g2225
  (
    n2209,
    n1183,
    n1192,
    n1676,
    n1056
  );


  nand
  g2226
  (
    n2020,
    n1577,
    n1641,
    n1683,
    n1712
  );


  nor
  g2227
  (
    n2017,
    n1636,
    n1424,
    n1392,
    n1504
  );


  nand
  g2228
  (
    n2557,
    n1044,
    n1665,
    n1140,
    n1674
  );


  xnor
  g2229
  (
    n2374,
    n1211,
    n1253,
    n1234,
    n1591
  );


  nand
  g2230
  (
    n2361,
    n1275,
    n1308,
    n1160,
    n1755
  );


  xnor
  g2231
  (
    n2356,
    n1429,
    n1465,
    n1194,
    n1593
  );


  nand
  g2232
  (
    n2007,
    n1335,
    n1808,
    n1387,
    n1128
  );


  nand
  g2233
  (
    n2538,
    n1319,
    n1060,
    n1681,
    n1508
  );


  and
  g2234
  (
    n2129,
    n1172,
    n1552,
    n1261,
    n1336
  );


  nand
  g2235
  (
    n2120,
    n1540,
    n1390,
    n1691,
    n1385
  );


  or
  g2236
  (
    n2590,
    n1722,
    n1723,
    n1807,
    n1676
  );


  nand
  g2237
  (
    n2024,
    n1301,
    n1262,
    n1099,
    n1800
  );


  nand
  g2238
  (
    n2281,
    n1674,
    n1614,
    n1546,
    n1077
  );


  or
  g2239
  (
    n2553,
    n1067,
    n1100,
    n1331,
    n1172
  );


  nor
  g2240
  (
    n2259,
    n1507,
    n1049,
    n1066,
    n1725
  );


  or
  g2241
  (
    n2076,
    n1432,
    n1250,
    n1279,
    n1276
  );


  xor
  g2242
  (
    n2338,
    n1305,
    n1189,
    n1196,
    n1579
  );


  nand
  g2243
  (
    n2631,
    n1505,
    n1575,
    n1213,
    n1632
  );


  xnor
  g2244
  (
    n2320,
    n1242,
    n1394,
    n1502,
    n1443
  );


  or
  g2245
  (
    n2545,
    n1236,
    n1073,
    n1690,
    n1389
  );


  xnor
  g2246
  (
    n2333,
    n1614,
    n1506,
    n1398,
    n1099
  );


  and
  g2247
  (
    n2493,
    n1718,
    n1494,
    n1201,
    n1576
  );


  or
  g2248
  (
    n2474,
    n1694,
    n1745,
    n1222,
    n1216
  );


  or
  g2249
  (
    n2117,
    n1371,
    n1036,
    n1717,
    n1145
  );


  nand
  g2250
  (
    n2335,
    n1219,
    n1775,
    n1207,
    n1112
  );


  and
  g2251
  (
    n2352,
    n1444,
    n1721,
    n1487,
    n1047
  );


  nand
  g2252
  (
    n2255,
    n1590,
    n1635,
    n1474,
    n1093
  );


  nor
  g2253
  (
    n2525,
    n1359,
    n1137,
    n1296,
    n1693
  );


  or
  g2254
  (
    n1997,
    n1790,
    n1254,
    n1525,
    n1581
  );


  xnor
  g2255
  (
    n2196,
    n1642,
    n1195,
    n1240,
    n1096
  );


  and
  g2256
  (
    n2118,
    n1053,
    n1628,
    n1143,
    n1166
  );


  or
  g2257
  (
    n2688,
    n1489,
    n1272,
    n1375,
    n1689
  );


  nor
  g2258
  (
    n2534,
    n1206,
    n1588,
    n1070,
    n1519
  );


  and
  g2259
  (
    n2489,
    n1705,
    n1344,
    n1129,
    n1090
  );


  nand
  g2260
  (
    n1945,
    n1559,
    n1718,
    n1792,
    n1293
  );


  nand
  g2261
  (
    n2625,
    n1084,
    n1302,
    n1184,
    n1201
  );


  nor
  g2262
  (
    n1946,
    n1196,
    n1640,
    n1359,
    n1563
  );


  nor
  g2263
  (
    n2109,
    n1234,
    n1460,
    n1238,
    n1551
  );


  or
  g2264
  (
    n2413,
    n1688,
    n1223,
    n1515,
    n1453
  );


  or
  g2265
  (
    n2119,
    n1571,
    n1368,
    n1476,
    n1657
  );


  xnor
  g2266
  (
    n2712,
    n1419,
    n1477,
    n1511,
    n1264
  );


  xor
  g2267
  (
    n2428,
    n1322,
    n1363,
    n1321,
    n1451
  );


  nand
  g2268
  (
    n2376,
    n1187,
    n1282,
    n1292,
    n1556
  );


  xor
  g2269
  (
    n2342,
    n1162,
    n1771,
    n1460,
    n1377
  );


  nor
  g2270
  (
    n2457,
    n1268,
    n1060,
    n1225,
    n1163
  );


  nand
  g2271
  (
    n2140,
    n1038,
    n1545,
    n1430,
    n1197
  );


  and
  g2272
  (
    n2093,
    n1228,
    n1447,
    n1123,
    n1068
  );


  or
  g2273
  (
    n2414,
    n1546,
    n1087,
    n1629,
    n1312
  );


  xor
  g2274
  (
    n2148,
    n1645,
    n1659,
    n1726,
    n1760
  );


  and
  g2275
  (
    n2126,
    n1739,
    n1347,
    n1373,
    n1307
  );


  xor
  g2276
  (
    n2523,
    n1728,
    n1137,
    n1437,
    n1062
  );


  or
  g2277
  (
    n2124,
    n1171,
    n1192,
    n1247,
    n1385
  );


  or
  g2278
  (
    n2102,
    n1481,
    n1528,
    n1275,
    n1240
  );


  xor
  g2279
  (
    n1964,
    n1741,
    n1612,
    n1117,
    n1633
  );


  xor
  g2280
  (
    n2554,
    n1579,
    n1599,
    n1742,
    n1181
  );


  nand
  g2281
  (
    n2349,
    n1196,
    n1458,
    n1197,
    n1420
  );


  nand
  g2282
  (
    n2632,
    n1721,
    n1565,
    n1804,
    n1426
  );


  xor
  g2283
  (
    n2339,
    n1635,
    n1148,
    n1230,
    n1554
  );


  nor
  g2284
  (
    n2453,
    n1456,
    n1093,
    n1592,
    n1133
  );


  xor
  g2285
  (
    n2647,
    n1516,
    n1782,
    n1498,
    n1341
  );


  or
  g2286
  (
    n2345,
    n1295,
    n1217,
    n1668,
    n1131
  );


  xnor
  g2287
  (
    n2445,
    n1161,
    n1809,
    n1501,
    n1681
  );


  xnor
  g2288
  (
    n1974,
    n1685,
    n1363,
    n1726,
    n1164
  );


  xor
  g2289
  (
    n2372,
    n1757,
    n1434,
    n1318,
    n1154
  );


  and
  g2290
  (
    n1948,
    n1494,
    n1037,
    n1355,
    n1523
  );


  nand
  g2291
  (
    n2237,
    n1337,
    n1411,
    n1214,
    n1325
  );


  nor
  g2292
  (
    n2139,
    n1340,
    n1039,
    n1600,
    n1173
  );


  nor
  g2293
  (
    n2145,
    n1117,
    n1101,
    n1408,
    n1609
  );


  nand
  g2294
  (
    n2604,
    n1714,
    n1247,
    n1557,
    n1353
  );


  or
  g2295
  (
    n2703,
    n1647,
    n1515,
    n1251,
    n1567
  );


  and
  g2296
  (
    n2186,
    n1311,
    n1416,
    n1411,
    n1664
  );


  xor
  g2297
  (
    n1942,
    n1199,
    n1397,
    n1091,
    n1655
  );


  or
  g2298
  (
    n2637,
    n1731,
    n1079,
    n1155,
    n1282
  );


  xnor
  g2299
  (
    n2510,
    n1521,
    n1464,
    n1105,
    n1792
  );


  xor
  g2300
  (
    n2265,
    n1162,
    n1081,
    n1251,
    n1318
  );


  or
  g2301
  (
    n2679,
    n1158,
    n1797,
    n1519,
    n1692
  );


  xnor
  g2302
  (
    n2507,
    n1411,
    n1438,
    n1172,
    n1780
  );


  nor
  g2303
  (
    n2072,
    n1122,
    n1667,
    n1365,
    n1285
  );


  or
  g2304
  (
    n1994,
    n1468,
    n1143,
    n1338,
    n1719
  );


  xnor
  g2305
  (
    n2666,
    n1484,
    n1096,
    n1799,
    n1155
  );


  and
  g2306
  (
    n2260,
    n1516,
    n1540,
    n1491,
    n1412
  );


  and
  g2307
  (
    n2454,
    n1075,
    n1634,
    n1119,
    n1569
  );


  nor
  g2308
  (
    n2107,
    n1150,
    n1420,
    n1533,
    n1602
  );


  xor
  g2309
  (
    n2302,
    n1642,
    n1332,
    n1267,
    n1463
  );


  nor
  g2310
  (
    n2499,
    n1353,
    n1766,
    n1612,
    n1213
  );


  xor
  g2311
  (
    n2400,
    n1573,
    n1576,
    n1314,
    n1396
  );


  nor
  g2312
  (
    n2353,
    n1745,
    n1143,
    n1703,
    n1594
  );


  xor
  g2313
  (
    n2465,
    n1475,
    n1293,
    n1061,
    n1142
  );


  xnor
  g2314
  (
    n2052,
    n1244,
    n1366,
    n1356,
    n1445
  );


  and
  g2315
  (
    n1984,
    n1439,
    n1370,
    n1582,
    n1794
  );


  nand
  g2316
  (
    n2369,
    n1789,
    n1446,
    n1775,
    n1135
  );


  xnor
  g2317
  (
    n2392,
    n1086,
    n1578,
    n1366,
    n1432
  );


  nand
  g2318
  (
    n2595,
    n1327,
    n1706,
    n1326,
    n1296
  );


  nor
  g2319
  (
    n2098,
    n1605,
    n1338,
    n1083,
    n1445
  );


  xnor
  g2320
  (
    n2166,
    n1463,
    n1265,
    n1649,
    n1291
  );


  and
  g2321
  (
    n2127,
    n1359,
    n1346,
    n1216,
    n1355
  );


  nor
  g2322
  (
    n2658,
    n1297,
    n1788,
    n1407,
    n1285
  );


  nand
  g2323
  (
    n2325,
    n1811,
    n1707,
    n1538,
    n1510
  );


  xnor
  g2324
  (
    n1993,
    n1628,
    n1042,
    n1365,
    n1654
  );


  nor
  g2325
  (
    n2426,
    n1305,
    n1159,
    n1076,
    n1229
  );


  or
  g2326
  (
    n2051,
    n1415,
    n1641,
    n1321,
    n1055
  );


  xnor
  g2327
  (
    n2191,
    n1654,
    n1155,
    n1127,
    n1520
  );


  or
  g2328
  (
    n2344,
    n1456,
    n1672,
    n1792,
    n1235
  );


  nand
  g2329
  (
    n2518,
    n1781,
    n1409,
    n1219,
    n1439
  );


  or
  g2330
  (
    n2652,
    n1408,
    n1418,
    n1697,
    n1227
  );


  and
  g2331
  (
    n2589,
    n1085,
    n1256,
    n1524,
    n1584
  );


  nor
  g2332
  (
    n2423,
    n1673,
    n1272,
    n1706,
    n1599
  );


  xnor
  g2333
  (
    n1954,
    n1117,
    n1403,
    n1232,
    n1068
  );


  xor
  g2334
  (
    n2541,
    n1780,
    n1426,
    n1281,
    n1725
  );


  or
  g2335
  (
    n2531,
    n1419,
    n1099,
    n1439,
    n1812
  );


  or
  g2336
  (
    n2549,
    n1595,
    n1676,
    n1416,
    n1593
  );


  nand
  g2337
  (
    n2094,
    n1337,
    n1714,
    n1177,
    n1360
  );


  xnor
  g2338
  (
    n2087,
    n1762,
    n1107,
    n1661,
    n1374
  );


  and
  g2339
  (
    n2270,
    n1539,
    n1368,
    n1180,
    n1432
  );


  nand
  g2340
  (
    n2055,
    n1559,
    n1227,
    n1475,
    n1539
  );


  nor
  g2341
  (
    n2439,
    n1752,
    n1068,
    n1560,
    n1550
  );


  and
  g2342
  (
    n2492,
    n1193,
    n1037,
    n1748,
    n1541
  );


  or
  g2343
  (
    n2212,
    n1576,
    n1211,
    n1268,
    n1377
  );


  nor
  g2344
  (
    n2029,
    n1210,
    n1317,
    n1536,
    n1243
  );


  xor
  g2345
  (
    n2404,
    n1494,
    n1138,
    n1516,
    n1215
  );


  nand
  g2346
  (
    n2228,
    n1046,
    n1542,
    n1620,
    n1204
  );


  nor
  g2347
  (
    n2505,
    n1158,
    n1619,
    n1655,
    n1456
  );


  xor
  g2348
  (
    n2396,
    n1717,
    n1633,
    n1347,
    n1167
  );


  xor
  g2349
  (
    n2436,
    n1581,
    n1201,
    n1389,
    n1537
  );


  or
  g2350
  (
    n2469,
    n1552,
    n1379,
    n1665,
    n1555
  );


  or
  g2351
  (
    n2528,
    n1055,
    n1213,
    n1705,
    n1590
  );


  or
  g2352
  (
    n2326,
    n1096,
    n1743,
    n1042,
    n1502
  );


  xor
  g2353
  (
    n1962,
    n1206,
    n1516,
    n1608,
    n1565
  );


  xnor
  g2354
  (
    n2418,
    n1072,
    n1805,
    n1454,
    n1430
  );


  or
  g2355
  (
    n2512,
    n1105,
    n1159,
    n1193,
    n1186
  );


  xor
  g2356
  (
    n2028,
    n1527,
    n1717,
    n1445,
    n1167
  );


  nand
  g2357
  (
    n2009,
    n1366,
    n1514,
    n1750,
    n1697
  );


  xnor
  g2358
  (
    n2713,
    n1223,
    n1538,
    n1729,
    n1646
  );


  or
  g2359
  (
    n2088,
    n1397,
    n1696,
    n1278,
    n1471
  );


  nor
  g2360
  (
    n2245,
    n1748,
    n1286,
    n1134,
    n1678
  );


  or
  g2361
  (
    n2586,
    n1764,
    n1680,
    n1512,
    n1078
  );


  xnor
  g2362
  (
    n2134,
    n1236,
    n1187,
    n1800,
    n1696
  );


  xnor
  g2363
  (
    n2551,
    n1382,
    n1325,
    n1746,
    n1227
  );


  and
  g2364
  (
    n2168,
    n1602,
    n1139,
    n1377,
    n1591
  );


  or
  g2365
  (
    n2099,
    n1118,
    n1488,
    n1671,
    n1468
  );


  and
  g2366
  (
    n1969,
    n1149,
    n1367,
    n1656,
    n1693
  );


  nor
  g2367
  (
    n2319,
    n1573,
    n1085,
    n1688,
    n1433
  );


  xnor
  g2368
  (
    n2018,
    n1809,
    n1618,
    n1191,
    n1684
  );


  or
  g2369
  (
    n2221,
    n1584,
    n1064,
    n1106,
    n1262
  );


  nand
  g2370
  (
    n2409,
    n1397,
    n1378,
    n1664,
    n1718
  );


  or
  g2371
  (
    n2562,
    n1640,
    n1255,
    n1141,
    n1177
  );


  nand
  g2372
  (
    n2620,
    n1677,
    n1791,
    n1470,
    n1452
  );


  xnor
  g2373
  (
    n2607,
    n1566,
    n1205,
    n1198,
    n1078
  );


  xnor
  g2374
  (
    n2657,
    n1607,
    n1415,
    n1184,
    n1115
  );


  or
  g2375
  (
    n2175,
    n1658,
    n1324,
    n1510,
    n1680
  );


  or
  g2376
  (
    n2456,
    n1310,
    n1703,
    n1157,
    n1250
  );


  nand
  g2377
  (
    n2384,
    n1270,
    n1570,
    n1280,
    n1563
  );


  xor
  g2378
  (
    n2603,
    n1332,
    n1812,
    n1036,
    n1457
  );


  xor
  g2379
  (
    n2502,
    n1550,
    n1183,
    n1786,
    n1675
  );


  nor
  g2380
  (
    n2475,
    n1753,
    n1273,
    n1658,
    n1725
  );


  and
  g2381
  (
    n2025,
    n1696,
    n1679,
    n1689,
    n1773
  );


  nor
  g2382
  (
    n2389,
    n1621,
    n1474,
    n1732,
    n1589
  );


  and
  g2383
  (
    n2580,
    n1317,
    n1522,
    n1136,
    n1768
  );


  nor
  g2384
  (
    n2673,
    n1189,
    n1111,
    n1639,
    n1789
  );


  nor
  g2385
  (
    n2273,
    n1481,
    n1427,
    n1115,
    n1480
  );


  xnor
  g2386
  (
    n2324,
    n1412,
    n1341,
    n1095,
    n1291
  );


  xnor
  g2387
  (
    n2008,
    n1077,
    n1362,
    n1546,
    n1632
  );


  nand
  g2388
  (
    n2213,
    n1566,
    n1506,
    n1380,
    n1668
  );


  xnor
  g2389
  (
    n2132,
    n1122,
    n1568,
    n1586,
    n1128
  );


  xnor
  g2390
  (
    n2012,
    n1112,
    n1521,
    n1555,
    n1661
  );


  nor
  g2391
  (
    n1950,
    n1126,
    n1580,
    n1048,
    n1283
  );


  and
  g2392
  (
    n2322,
    n1196,
    n1255,
    n1562,
    n1179
  );


  xnor
  g2393
  (
    n2106,
    n1560,
    n1798,
    n1233,
    n1218
  );


  xor
  g2394
  (
    n2624,
    n1345,
    n1184,
    n1303,
    n1141
  );


  xnor
  g2395
  (
    n2617,
    n1800,
    n1393,
    n1660,
    n1510
  );


  or
  g2396
  (
    n2565,
    n1294,
    n1372,
    n1395,
    n1502
  );


  xor
  g2397
  (
    n2332,
    n1056,
    n1164,
    n1340,
    n1174
  );


  xnor
  g2398
  (
    n2682,
    n1043,
    n1629,
    n1589,
    n1646
  );


  xor
  g2399
  (
    n2204,
    n1713,
    n1737,
    n1264,
    n1235
  );


  and
  g2400
  (
    n2601,
    n1434,
    n1432,
    n1708,
    n1547
  );


  or
  g2401
  (
    n2552,
    n1611,
    n1509,
    n1285,
    n1280
  );


  xnor
  g2402
  (
    n2047,
    n1177,
    n1518,
    n1616,
    n1772
  );


  or
  g2403
  (
    n2147,
    n1165,
    n1787,
    n1478,
    n1638
  );


  or
  g2404
  (
    n2484,
    n1142,
    n1650,
    n1805,
    n1543
  );


  and
  g2405
  (
    n2253,
    n1611,
    n1705,
    n1173,
    n1338
  );


  and
  g2406
  (
    n2705,
    n1635,
    n1374,
    n1227,
    n1756
  );


  xnor
  g2407
  (
    n2613,
    n1425,
    n1779,
    n1711,
    n1744
  );


  nor
  g2408
  (
    n2543,
    n1360,
    n1490,
    n1354,
    n1692
  );


  xnor
  g2409
  (
    n2143,
    n1732,
    n1690,
    n1493,
    n1517
  );


  or
  g2410
  (
    n1973,
    n1168,
    n1675,
    n1280,
    n1384
  );


  and
  g2411
  (
    n2033,
    n1597,
    n1422,
    n1661,
    n1724
  );


  xor
  g2412
  (
    n2234,
    n1098,
    n1701,
    n1263,
    n1747
  );


  nand
  g2413
  (
    n2063,
    n1681,
    n1673,
    n31,
    n1402
  );


  nand
  g2414
  (
    n2231,
    n1795,
    n1450,
    n1410,
    n1137
  );


  or
  g2415
  (
    n2684,
    n1672,
    n1241,
    n1505,
    n1239
  );


  xnor
  g2416
  (
    n2275,
    n1467,
    n1277,
    n1724,
    n1194
  );


  nand
  g2417
  (
    n2287,
    n1436,
    n1744,
    n1810,
    n1134
  );


  nor
  g2418
  (
    n2424,
    n1678,
    n1626,
    n1097,
    n1634
  );


  xnor
  g2419
  (
    n2208,
    n1619,
    n1730,
    n1606,
    n1645
  );


  xnor
  g2420
  (
    n2473,
    n1789,
    n1387,
    n1599,
    n1747
  );


  nor
  g2421
  (
    n2687,
    n1518,
    n1430,
    n1291,
    n1295
  );


  nand
  g2422
  (
    n2005,
    n1218,
    n1686,
    n1772,
    n1238
  );


  or
  g2423
  (
    n2585,
    n1449,
    n1237,
    n1783,
    n1564
  );


  and
  g2424
  (
    n2660,
    n1101,
    n1266,
    n1413,
    n1607
  );


  nor
  g2425
  (
    n2440,
    n1483,
    n1406,
    n1239,
    n1691
  );


  nor
  g2426
  (
    n2123,
    n1090,
    n1155,
    n1368,
    n1381
  );


  nor
  g2427
  (
    n2185,
    n1135,
    n1624,
    n1426,
    n1298
  );


  and
  g2428
  (
    n2219,
    n1051,
    n1071,
    n1140,
    n1174
  );


  and
  g2429
  (
    n2239,
    n1135,
    n1573,
    n1778,
    n1390
  );


  xnor
  g2430
  (
    n2539,
    n1702,
    n1546,
    n1052,
    n1596
  );


  and
  g2431
  (
    n2188,
    n1485,
    n1769,
    n1806,
    n1102
  );


  xor
  g2432
  (
    n2199,
    n1458,
    n1545,
    n1700,
    n1485
  );


  xor
  g2433
  (
    n2224,
    n1085,
    n1776,
    n1597,
    n1289
  );


  xnor
  g2434
  (
    n2482,
    n1329,
    n1351,
    n1055,
    n1509
  );


  nand
  g2435
  (
    n1998,
    n1472,
    n1727,
    n1438,
    n1495
  );


  or
  g2436
  (
    n2060,
    n1365,
    n1356,
    n1806,
    n1240
  );


  nor
  g2437
  (
    n2205,
    n1666,
    n1585,
    n1463,
    n1101
  );


  xor
  g2438
  (
    n1986,
    n1206,
    n1605,
    n1332,
    n1462
  );


  and
  g2439
  (
    n2643,
    n1442,
    n1156,
    n1394,
    n1290
  );


  nand
  g2440
  (
    n2419,
    n1463,
    n1330,
    n1104,
    n1036
  );


  xor
  g2441
  (
    n2587,
    n1103,
    n1075,
    n1479,
    n1534
  );


  nand
  g2442
  (
    n2626,
    n1560,
    n1623,
    n1081,
    n1127
  );


  xnor
  g2443
  (
    n2229,
    n1460,
    n1443,
    n1105,
    n1760
  );


  xor
  g2444
  (
    n2070,
    n1369,
    n1685,
    n1270,
    n1183
  );


  xnor
  g2445
  (
    n2371,
    n1720,
    n1663,
    n1040,
    n1685
  );


  or
  g2446
  (
    n2211,
    n1394,
    n1620,
    n1625,
    n1536
  );


  or
  g2447
  (
    n2574,
    n1063,
    n1200,
    n1073,
    n1530
  );


  xor
  g2448
  (
    n2183,
    n1203,
    n1104,
    n1244,
    n1300
  );


  and
  g2449
  (
    n2689,
    n1144,
    n1218,
    n1373,
    n1511
  );


  nand
  g2450
  (
    n1963,
    n1143,
    n1226,
    n1706,
    n1766
  );


  xor
  g2451
  (
    n2248,
    n1765,
    n1504,
    n1041,
    n1446
  );


  xor
  g2452
  (
    n2564,
    n1241,
    n1535,
    n1217,
    n1144
  );


  xor
  g2453
  (
    n2034,
    n1518,
    n1664,
    n1737,
    n1674
  );


  or
  g2454
  (
    n2702,
    n1715,
    n1777,
    n1476,
    n1602
  );


  and
  g2455
  (
    n2526,
    n1271,
    n1612,
    n1098,
    n1491
  );


  nor
  g2456
  (
    n2083,
    n1513,
    n1325,
    n1288,
    n1780
  );


  nor
  g2457
  (
    n2331,
    n1575,
    n1709,
    n1053,
    n1216
  );


  xor
  g2458
  (
    n2709,
    n1362,
    n1134,
    n1082,
    n1488
  );


  xor
  g2459
  (
    n2271,
    n1561,
    n1405,
    n1274,
    n1624
  );


  xor
  g2460
  (
    n2334,
    n1362,
    n1515,
    n1560,
    n1225
  );


  and
  g2461
  (
    n2416,
    n1803,
    n1744,
    n1326,
    n1778
  );


  and
  g2462
  (
    n2385,
    n1226,
    n1423,
    n1522,
    n1461
  );


  and
  g2463
  (
    n2681,
    n1159,
    n1419,
    n1273,
    n1613
  );


  and
  g2464
  (
    n2437,
    n1807,
    n1641,
    n1178,
    n1240
  );


  xnor
  g2465
  (
    n2533,
    n1480,
    n1423,
    n1229,
    n1689
  );


  nor
  g2466
  (
    n2548,
    n1503,
    n1723,
    n1066,
    n1054
  );


  xnor
  g2467
  (
    n2235,
    n1564,
    n1315,
    n1082,
    n1052
  );


  xor
  g2468
  (
    n2161,
    n1479,
    n1120,
    n1396,
    n1378
  );


  or
  g2469
  (
    n2560,
    n1415,
    n1798,
    n1430,
    n1236
  );


  and
  g2470
  (
    n2655,
    n1190,
    n1634,
    n1191,
    n1438
  );


  or
  g2471
  (
    n2481,
    n1683,
    n1110,
    n1102,
    n1158
  );


  nand
  g2472
  (
    n2472,
    n1411,
    n1667,
    n1690,
    n1709
  );


  nand
  g2473
  (
    n2358,
    n1071,
    n1684,
    n1441,
    n1677
  );


  xor
  g2474
  (
    n2471,
    n1395,
    n1569,
    n1288,
    n1537
  );


  and
  g2475
  (
    n2678,
    n1759,
    n1482,
    n1786,
    n1542
  );


  and
  g2476
  (
    n2256,
    n1321,
    n1287,
    n1208,
    n1586
  );


  nand
  g2477
  (
    n2441,
    n1601,
    n1126,
    n1734,
    n1210
  );


  xnor
  g2478
  (
    n2210,
    n1315,
    n1599,
    n1075,
    n1049
  );


  and
  g2479
  (
    n2563,
    n1501,
    n1658,
    n1601,
    n1278
  );


  xor
  g2480
  (
    n2157,
    n1500,
    n1631,
    n207,
    n1222
  );


  nand
  g2481
  (
    n2050,
    n1171,
    n1777,
    n1438,
    n1425
  );


  or
  g2482
  (
    n2680,
    n1614,
    n1385,
    n1306,
    n1660
  );


  xnor
  g2483
  (
    n2016,
    n1621,
    n1651,
    n1195,
    n1087
  );


  nor
  g2484
  (
    n2675,
    n1800,
    n1796,
    n1237,
    n1774
  );


  or
  g2485
  (
    n2223,
    n1309,
    n1267,
    n1767,
    n1402
  );


  nand
  g2486
  (
    n2495,
    n1300,
    n1564,
    n1592,
    n1311
  );


  and
  g2487
  (
    n2207,
    n1382,
    n1242,
    n1160,
    n1113
  );


  nor
  g2488
  (
    n2593,
    n1149,
    n1743,
    n1235,
    n1684
  );


  and
  g2489
  (
    n2627,
    n1561,
    n1663,
    n1804,
    n1444
  );


  and
  g2490
  (
    n2602,
    n1618,
    n1434,
    n1738,
    n1135
  );


  nand
  g2491
  (
    n2644,
    n1413,
    n1784,
    n1327,
    n1792
  );


  nand
  g2492
  (
    n2091,
    n1253,
    n1669,
    n1715,
    n1255
  );


  or
  g2493
  (
    n2249,
    n1424,
    n1357,
    n1535,
    n1611
  );


  or
  g2494
  (
    n2544,
    n1519,
    n1169,
    n1498,
    n1174
  );


  nor
  g2495
  (
    n2546,
    n1793,
    n1133,
    n1249,
    n1407
  );


  nor
  g2496
  (
    n2062,
    n1660,
    n1543,
    n1142,
    n1736
  );


  xnor
  g2497
  (
    n2346,
    n1414,
    n1127,
    n1745,
    n1530
  );


  xnor
  g2498
  (
    n2263,
    n1065,
    n1040,
    n1449,
    n1461
  );


  nor
  g2499
  (
    n2184,
    n1388,
    n1175,
    n1768,
    n1607
  );


  or
  g2500
  (
    n2677,
    n1482,
    n1449,
    n1238,
    n1521
  );


  and
  g2501
  (
    n1995,
    n1743,
    n1679,
    n1344,
    n1779
  );


  and
  g2502
  (
    n2588,
    n1163,
    n1296,
    n1453,
    n1811
  );


  or
  g2503
  (
    n2444,
    n1111,
    n1710,
    n1682,
    n1790
  );


  xnor
  g2504
  (
    n2172,
    n1762,
    n1186,
    n1215,
    n1693
  );


  xnor
  g2505
  (
    n2022,
    n1335,
    n1228,
    n1637,
    n1659
  );


  or
  g2506
  (
    n2571,
    n1260,
    n1238,
    n1389,
    n1455
  );


  xor
  g2507
  (
    n1979,
    n1452,
    n1799,
    n1538,
    n1617
  );


  or
  g2508
  (
    n2155,
    n1680,
    n1731,
    n1316,
    n1069
  );


  and
  g2509
  (
    n2069,
    n1539,
    n1466,
    n1067,
    n1234
  );


  nor
  g2510
  (
    n2566,
    n1487,
    n1164,
    n1657,
    n1773
  );


  or
  g2511
  (
    n2659,
    n1214,
    n1391,
    n1459,
    n1450
  );


  nand
  g2512
  (
    n2306,
    n1447,
    n1334,
    n1727,
    n1205
  );


  nand
  g2513
  (
    n2430,
    n1451,
    n1670,
    n1152,
    n1383
  );


  xnor
  g2514
  (
    n2080,
    n1695,
    n1719,
    n1632,
    n1215
  );


  or
  g2515
  (
    n2710,
    n1507,
    n1333,
    n1313,
    n1259
  );


  nand
  g2516
  (
    n1976,
    n1591,
    n1680,
    n1051,
    n1412
  );


  or
  g2517
  (
    n2328,
    n1468,
    n1038,
    n1323,
    n1638
  );


  xnor
  g2518
  (
    n2614,
    n1762,
    n1244,
    n1113,
    n1701
  );


  and
  g2519
  (
    n2216,
    n1128,
    n1182,
    n1373,
    n1503
  );


  xnor
  g2520
  (
    n2294,
    n1140,
    n1043,
    n1108,
    n1296
  );


  nand
  g2521
  (
    n1989,
    n1567,
    n1208,
    n1478,
    n1078
  );


  nand
  g2522
  (
    n2378,
    n1443,
    n1526,
    n1039,
    n1729
  );


  nand
  g2523
  (
    n2160,
    n1597,
    n1219,
    n1249,
    n1057
  );


  nor
  g2524
  (
    n2425,
    n1509,
    n1057,
    n1687,
    n1472
  );


  and
  g2525
  (
    n1944,
    n1758,
    n1697,
    n1304,
    n1273
  );


  xor
  g2526
  (
    n2663,
    n1605,
    n1627,
    n1740,
    n1544
  );


  xnor
  g2527
  (
    n1939,
    n1435,
    n1688,
    n1730,
    n1401
  );


  or
  g2528
  (
    n2699,
    n1755,
    n1782,
    n1441,
    n1626
  );


  nand
  g2529
  (
    n2381,
    n1588,
    n1702,
    n1396,
    n1556
  );


  and
  g2530
  (
    n2066,
    n1138,
    n1736,
    n1176,
    n1036
  );


  nor
  g2531
  (
    n2555,
    n1474,
    n1218,
    n1081,
    n1695
  );


  nor
  g2532
  (
    n2077,
    n1457,
    n1339,
    n1574,
    n1592
  );


  nor
  g2533
  (
    n1980,
    n1624,
    n1570,
    n1298,
    n1269
  );


  nor
  g2534
  (
    n2674,
    n1435,
    n1256,
    n1583,
    n1760
  );


  nand
  g2535
  (
    n2303,
    n1344,
    n1806,
    n1109,
    n1551
  );


  nor
  g2536
  (
    n2236,
    n1643,
    n1068,
    n1647,
    n1147
  );


  nand
  g2537
  (
    n2090,
    n1074,
    n1224,
    n1242,
    n1286
  );


  xnor
  g2538
  (
    n2696,
    n1343,
    n1381,
    n1490,
    n1183
  );


  nor
  g2539
  (
    n2569,
    n1186,
    n1617,
    n1462,
    n1640
  );


  nor
  g2540
  (
    n2362,
    n1116,
    n1041,
    n1793,
    n1226
  );


  or
  g2541
  (
    n2535,
    n1192,
    n1153,
    n1342,
    n1765
  );


  xnor
  g2542
  (
    n2096,
    n1425,
    n1753,
    n1224,
    n1336
  );


  xnor
  g2543
  (
    n2283,
    n1306,
    n1717,
    n1205,
    n1187
  );


  nand
  g2544
  (
    n2218,
    n1709,
    n1271,
    n1077,
    n1191
  );


  and
  g2545
  (
    n2530,
    n1041,
    n1148,
    n1677,
    n1157
  );


  xnor
  g2546
  (
    n2006,
    n1344,
    n1310,
    n1752,
    n1683
  );


  nand
  g2547
  (
    n2169,
    n1054,
    n1230,
    n1229,
    n1093
  );


  and
  g2548
  (
    n2411,
    n1533,
    n1077,
    n1170,
    n1777
  );


  nor
  g2549
  (
    n1988,
    n1528,
    n1220,
    n1450,
    n1694
  );


  nor
  g2550
  (
    n2097,
    n1360,
    n1505,
    n1125,
    n1400
  );


  nand
  g2551
  (
    n2408,
    n1497,
    n1288,
    n1648,
    n1805
  );


  xnor
  g2552
  (
    n2226,
    n1229,
    n1083,
    n1666,
    n1370
  );


  or
  g2553
  (
    n2387,
    n1750,
    n1742,
    n1386,
    n1564
  );


  or
  g2554
  (
    n2503,
    n1052,
    n1796,
    n1089,
    n1484
  );


  nor
  g2555
  (
    n2182,
    n1710,
    n1112,
    n1231,
    n1126
  );


  and
  g2556
  (
    n2394,
    n1572,
    n1728,
    n1292,
    n1741
  );


  or
  g2557
  (
    n2113,
    n1429,
    n1154,
    n1150,
    n1088
  );


  nand
  g2558
  (
    n2668,
    n1725,
    n1751,
    n1197,
    n1379
  );


  xnor
  g2559
  (
    n2459,
    n1286,
    n1684,
    n1204,
    n1389
  );


  xnor
  g2560
  (
    n2092,
    n1544,
    n1248,
    n1501,
    n1209
  );


  xnor
  g2561
  (
    n2584,
    n1632,
    n1381,
    n1249,
    n1257
  );


  nor
  g2562
  (
    n2225,
    n1351,
    n1073,
    n1182,
    n1263
  );


  xor
  g2563
  (
    n2159,
    n1471,
    n1603,
    n1185,
    n1453
  );


  nor
  g2564
  (
    n2316,
    n1480,
    n1449,
    n1770,
    n1169
  );


  xor
  g2565
  (
    n2490,
    n1219,
    n1259,
    n1363,
    n1450
  );


  and
  g2566
  (
    n2650,
    n1629,
    n1605,
    n1268,
    n1558
  );


  or
  g2567
  (
    n2379,
    n1331,
    n1469,
    n1710,
    n1259
  );


  and
  g2568
  (
    n2295,
    n1059,
    n1687,
    n1092,
    n1579
  );


  xor
  g2569
  (
    n2654,
    n1412,
    n1476,
    n1301,
    n1078
  );


  nand
  g2570
  (
    n2057,
    n1217,
    n1123,
    n1454,
    n1590
  );


  and
  g2571
  (
    n1934,
    n1715,
    n1292,
    n1653,
    n1602
  );


  or
  g2572
  (
    n2190,
    n1492,
    n1257,
    n1199,
    n1063
  );


  xnor
  g2573
  (
    n2330,
    n1686,
    n1675,
    n1364,
    n1671
  );


  and
  g2574
  (
    n1960,
    n1735,
    n1685,
    n1277,
    n1140
  );


  xnor
  g2575
  (
    n2577,
    n1644,
    n1604,
    n1710,
    n1210
  );


  xor
  g2576
  (
    n2479,
    n1059,
    n1231,
    n1687,
    n1778
  );


  and
  g2577
  (
    n2609,
    n1698,
    n1383,
    n1472,
    n1493
  );


  xnor
  g2578
  (
    n2704,
    n1513,
    n1058,
    n1795,
    n1654
  );


  nor
  g2579
  (
    n1951,
    n1246,
    n1669,
    n1349,
    n1804
  );


  nand
  g2580
  (
    n2446,
    n1572,
    n1251,
    n1491,
    n1061
  );


  nand
  g2581
  (
    n2691,
    n1797,
    n1126,
    n1678,
    n1339
  );


  nand
  g2582
  (
    n1985,
    n1594,
    n1666,
    n1118,
    n1423
  );


  xnor
  g2583
  (
    n2180,
    n1115,
    n1769,
    n1646,
    n1065
  );


  and
  g2584
  (
    n2044,
    n1802,
    n1628,
    n1361,
    n1537
  );


  nand
  g2585
  (
    n2383,
    n1523,
    n1347,
    n1216,
    n1319
  );


  xor
  g2586
  (
    n2661,
    n1231,
    n1379,
    n1282,
    n1574
  );


  and
  g2587
  (
    n2031,
    n1484,
    n1329,
    n1091,
    n1701
  );


  nor
  g2588
  (
    n2232,
    n1530,
    n1400,
    n1290,
    n1595
  );


  or
  g2589
  (
    n2573,
    n1523,
    n1788,
    n1721,
    n1801
  );


  xor
  g2590
  (
    n2388,
    n1611,
    n1086,
    n1621,
    n1304
  );


  xor
  g2591
  (
    n2670,
    n1768,
    n1291,
    n1604,
    n1187
  );


  nand
  g2592
  (
    n2293,
    n1596,
    n1190,
    n1234,
    n1452
  );


  or
  g2593
  (
    n2610,
    n1179,
    n1487,
    n1293,
    n1650
  );


  xnor
  g2594
  (
    n2032,
    n1613,
    n1320,
    n1269,
    n1297
  );


  xor
  g2595
  (
    n2629,
    n1051,
    n1526,
    n1810,
    n1297
  );


  xor
  g2596
  (
    n2163,
    n1603,
    n1427,
    n1610,
    n1802
  );


  xnor
  g2597
  (
    n2136,
    n1472,
    n1703,
    n1041,
    n1337
  );


  nand
  g2598
  (
    n1961,
    n1364,
    n1748,
    n1138,
    n1391
  );


  nor
  g2599
  (
    n2402,
    n1469,
    n1736,
    n1054,
    n1060
  );


  xor
  g2600
  (
    n2347,
    n1523,
    n1243,
    n1547,
    n1279
  );


  xor
  g2601
  (
    n2104,
    n1121,
    n1482,
    n1365,
    n1416
  );


  xor
  g2602
  (
    n2498,
    n1770,
    n1324,
    n1784,
    n1352
  );


  and
  g2603
  (
    n1949,
    n1361,
    n1686,
    n1596,
    n1160
  );


  nand
  g2604
  (
    n2220,
    n1141,
    n1278,
    n1506,
    n1107
  );


  or
  g2605
  (
    n2197,
    n1804,
    n1575,
    n1157,
    n1392
  );


  or
  g2606
  (
    n2268,
    n1303,
    n1167,
    n1513,
    n1551
  );


  xnor
  g2607
  (
    n2039,
    n1040,
    n1304,
    n1545,
    n1339
  );


  or
  g2608
  (
    n2575,
    n1467,
    n1367,
    n1761,
    n1287
  );


  xnor
  g2609
  (
    n2671,
    n1358,
    n1298,
    n1751,
    n1221
  );


  xor
  g2610
  (
    n2375,
    n1408,
    n1038,
    n1553,
    n1537
  );


  xnor
  g2611
  (
    n2266,
    n1580,
    n1697,
    n1464,
    n1461
  );


  or
  g2612
  (
    n2491,
    n1346,
    n1125,
    n1655,
    n1132
  );


  nand
  g2613
  (
    n2079,
    n1345,
    n1110,
    n1802,
    n1079
  );


  xnor
  g2614
  (
    n2653,
    n1606,
    n1598,
    n1525,
    n1431
  );


  xnor
  g2615
  (
    n2227,
    n1781,
    n1222,
    n1662,
    n1372
  );


  xor
  g2616
  (
    n2014,
    n1215,
    n1488,
    n1119,
    n1746
  );


  and
  g2617
  (
    n2568,
    n1102,
    n1207,
    n1394,
    n1749
  );


  xnor
  g2618
  (
    n2056,
    n1239,
    n1803,
    n1168,
    n1524
  );


  and
  g2619
  (
    n2061,
    n1386,
    n1091,
    n1317,
    n1790
  );


  or
  g2620
  (
    n2075,
    n1210,
    n1704,
    n1554,
    n1221
  );


  or
  g2621
  (
    n2291,
    n1288,
    n1440,
    n1070,
    n1501
  );


  and
  g2622
  (
    n2686,
    n1164,
    n1332,
    n1398,
    n1299
  );


  nor
  g2623
  (
    n2240,
    n1268,
    n1803,
    n1087,
    n1364
  );


  or
  g2624
  (
    n2026,
    n1388,
    n1751,
    n1558,
    n1726
  );


  nor
  g2625
  (
    n2105,
    n1657,
    n1199,
    n1617,
    n1550
  );


  nand
  g2626
  (
    n2261,
    n1293,
    n1522,
    n1786,
    n1368
  );


  nand
  g2627
  (
    n2649,
    n1258,
    n1600,
    n1167,
    n1360
  );


  or
  g2628
  (
    n2085,
    n1130,
    n1254,
    n1532,
    n1116
  );


  and
  g2629
  (
    n2701,
    n1549,
    n1724,
    n1119,
    n1361
  );


  xor
  g2630
  (
    n2583,
    n1207,
    n1308,
    n1805,
    n1591
  );


  and
  g2631
  (
    n1977,
    n1520,
    n1497,
    n1150,
    n1553
  );


  nand
  g2632
  (
    n2393,
    n1391,
    n1326,
    n1466,
    n1289
  );


  or
  g2633
  (
    n2215,
    n1289,
    n1156,
    n1120,
    n1588
  );


  xnor
  g2634
  (
    n2100,
    n1707,
    n1713,
    n1718,
    n1495
  );


  xor
  g2635
  (
    n1971,
    n1765,
    n1662,
    n1620,
    n1315
  );


  xor
  g2636
  (
    n2193,
    n1414,
    n1357,
    n1673,
    n1409
  );


  nor
  g2637
  (
    n2605,
    n1549,
    n1630,
    n1258,
    n1070
  );


  nor
  g2638
  (
    n2412,
    n1577,
    n1056,
    n1168,
    n1735
  );


  nand
  g2639
  (
    n2599,
    n1615,
    n1801,
    n1716,
    n1439
  );


  xor
  g2640
  (
    n2532,
    n1084,
    n1436,
    n1695,
    n1176
  );


  xnor
  g2641
  (
    n2149,
    n1131,
    n1299,
    n1448,
    n1320
  );


  nor
  g2642
  (
    n2300,
    n1566,
    n1170,
    n1270,
    n1109
  );


  xor
  g2643
  (
    n2451,
    n1417,
    n1211,
    n1801,
    n1305
  );


  and
  g2644
  (
    n2359,
    n1444,
    n1316,
    n1623,
    n1631
  );


  xor
  g2645
  (
    n2399,
    n1262,
    n1587,
    n1133,
    n1647
  );


  xor
  g2646
  (
    n2067,
    n1483,
    n1517,
    n1202,
    n1122
  );


  xor
  g2647
  (
    n2254,
    n1161,
    n1573,
    n1144,
    n1369
  );


  nand
  g2648
  (
    n2420,
    n1533,
    n1280,
    n1776,
    n1118
  );


  and
  g2649
  (
    n2662,
    n1429,
    n1756,
    n1309,
    n1583
  );


  xnor
  g2650
  (
    n2638,
    n1428,
    n1553,
    n1310,
    n1499
  );


  xnor
  g2651
  (
    n2572,
    n1052,
    n1153,
    n1746,
    n1040
  );


  xnor
  g2652
  (
    n1972,
    n1198,
    n1797,
    n1664,
    n1704
  );


  nor
  g2653
  (
    n2301,
    n1131,
    n1806,
    n1342,
    n1758
  );


  xnor
  g2654
  (
    n2170,
    n1529,
    n1037,
    n1044,
    n1589
  );


  xnor
  g2655
  (
    n2112,
    n1421,
    n1652,
    n1743,
    n1228
  );


  or
  g2656
  (
    n2645,
    n1086,
    n1608,
    n1763,
    n1212
  );


  xor
  g2657
  (
    n2011,
    n1682,
    n1812,
    n1587,
    n1637
  );


  nor
  g2658
  (
    n2138,
    n1334,
    n1398,
    n1737,
    n1194
  );


  nor
  g2659
  (
    n2133,
    n1567,
    n1243,
    n1442,
    n1325
  );


  xor
  g2660
  (
    n2158,
    n1376,
    n1182,
    n1650,
    n1121
  );


  or
  g2661
  (
    n2537,
    n1403,
    n1094,
    n1120,
    n1149
  );


  xor
  g2662
  (
    n2217,
    n1305,
    n1204,
    n1285,
    n1065
  );


  xnor
  g2663
  (
    n2111,
    n1549,
    n1414,
    n1079,
    n1175
  );


  xnor
  g2664
  (
    n2312,
    n1308,
    n1437,
    n1350,
    n1045
  );


  xnor
  g2665
  (
    n2708,
    n1045,
    n1741,
    n1356,
    n1474
  );


  nand
  g2666
  (
    n2478,
    n1281,
    n1261,
    n1061,
    n1433
  );


  nor
  g2667
  (
    n2442,
    n1316,
    n1248,
    n1225,
    n1044
  );


  nand
  g2668
  (
    n2598,
    n1050,
    n1355,
    n1764,
    n1152
  );


  nor
  g2669
  (
    n2289,
    n1657,
    n1245,
    n1578,
    n1165
  );


  or
  g2670
  (
    n2581,
    n1530,
    n1151,
    n1612,
    n1698
  );


  nor
  g2671
  (
    n2690,
    n1113,
    n1440,
    n1557,
    n1316
  );


  xor
  g2672
  (
    n2341,
    n1738,
    n1386,
    n1541,
    n1764
  );


  or
  g2673
  (
    n1999,
    n1457,
    n1058,
    n1557,
    n1462
  );


  and
  g2674
  (
    n2355,
    n1269,
    n1175,
    n1209,
    n1673
  );


  nor
  g2675
  (
    n2337,
    n1063,
    n1342,
    n1548,
    n1707
  );


  xor
  g2676
  (
    n2516,
    n1267,
    n1570,
    n1643,
    n1307
  );


  or
  g2677
  (
    n2467,
    n1309,
    n1736,
    n1208,
    n1512
  );


  xnor
  g2678
  (
    n2135,
    n1477,
    n1473,
    n1069,
    n1048
  );


  and
  g2679
  (
    n1941,
    n1246,
    n1314,
    n1422,
    n1634
  );


  nand
  g2680
  (
    n2152,
    n1722,
    n1343,
    n1366,
    n1380
  );


  nor
  g2681
  (
    n2719,
    n1942,
    n1952,
    n1960,
    n1982
  );


  xnor
  g2682
  (
    n2718,
    n1934,
    n1988,
    n1963,
    n1935
  );


  and
  g2683
  (
    n2714,
    n1989,
    n1945,
    n1951,
    n1953
  );


  nand
  g2684
  (
    n2728,
    n1973,
    n1961,
    n1940,
    n1970
  );


  xnor
  g2685
  (
    n2717,
    n1978,
    n1977,
    n1991,
    n1958
  );


  and
  g2686
  (
    n2715,
    n1938,
    n1947,
    n1986,
    n1992
  );


  nand
  g2687
  (
    n2726,
    n1974,
    n1948,
    n1981,
    n1962
  );


  xor
  g2688
  (
    n2725,
    n1967,
    n1957,
    n1969,
    n1966
  );


  and
  g2689
  (
    n2720,
    n1949,
    n1936,
    n1984,
    n1975
  );


  or
  g2690
  (
    n2722,
    n1976,
    n1968,
    n1956,
    n1985
  );


  xor
  g2691
  (
    n2716,
    n1954,
    n1950,
    n1971,
    n1937
  );


  nor
  g2692
  (
    n2723,
    n1959,
    n1943,
    n1990,
    n1939
  );


  nand
  g2693
  (
    n2721,
    n1987,
    n1983,
    n1941,
    n1955
  );


  or
  g2694
  (
    n2724,
    n1965,
    n1979,
    n1980,
    n1946
  );


  xnor
  g2695
  (
    n2727,
    n1933,
    n1964,
    n1944,
    n1972
  );


  not
  g2696
  (
    n2731,
    n208
  );


  buf
  g2697
  (
    n2730,
    n2714
  );


  nor
  g2698
  (
    n2729,
    n2716,
    n208,
    n2715
  );


  xnor
  g2699
  (
    n2738,
    n534,
    n2730,
    n536
  );


  or
  g2700
  (
    n2737,
    n532,
    n537,
    n2731
  );


  nor
  g2701
  (
    n2733,
    n2729,
    n535,
    n532
  );


  xnor
  g2702
  (
    n2734,
    n2730,
    n534,
    n536
  );


  nor
  g2703
  (
    n2740,
    n2731,
    n536,
    n2730,
    n537
  );


  or
  g2704
  (
    n2735,
    n532,
    n533,
    n531
  );


  and
  g2705
  (
    n2736,
    n533,
    n535,
    n532,
    n2731
  );


  or
  g2706
  (
    n2739,
    n534,
    n2731,
    n533,
    n535
  );


  or
  g2707
  (
    n2732,
    n2730,
    n2729
  );


  buf
  g2708
  (
    n2743,
    n2732
  );


  buf
  g2709
  (
    n2750,
    n2733
  );


  not
  g2710
  (
    n2745,
    n2734
  );


  not
  g2711
  (
    n2746,
    n2733
  );


  not
  g2712
  (
    n2749,
    n2736
  );


  buf
  g2713
  (
    n2747,
    n2735
  );


  buf
  g2714
  (
    n2752,
    n2736
  );


  not
  g2715
  (
    n2748,
    n2733
  );


  not
  g2716
  (
    n2741,
    n208
  );


  not
  g2717
  (
    n2751,
    n2734
  );


  nor
  g2718
  (
    n2742,
    n2733,
    n2735
  );


  xor
  g2719
  (
    n2744,
    n2734,
    n2735
  );


  nand
  g2720
  (
    n2766,
    n2742,
    n2752,
    n2736
  );


  xor
  g2721
  (
    n2765,
    n2746,
    n2739,
    n2752,
    n2747
  );


  xnor
  g2722
  (
    n2768,
    n2748,
    n2745,
    n2741
  );


  or
  g2723
  (
    n2758,
    n2737,
    n2747,
    n2749,
    n2739
  );


  nor
  g2724
  (
    n2767,
    n2738,
    n2743,
    n2749,
    n2747
  );


  and
  g2725
  (
    n2761,
    n2743,
    n2745,
    n2738,
    n2737
  );


  xnor
  g2726
  (
    n2753,
    n2750,
    n2750,
    n2739,
    n2752
  );


  nand
  g2727
  (
    n2754,
    n2746,
    n2744,
    n2749
  );


  xnor
  g2728
  (
    n2760,
    n2744,
    n2742,
    n2746,
    n2750
  );


  nand
  g2729
  (
    n2757,
    n2751,
    n2743,
    n2750,
    n2741
  );


  and
  g2730
  (
    n2764,
    n2746,
    n2738,
    n2751,
    n2748
  );


  nand
  g2731
  (
    n2762,
    n2737,
    n2745,
    n2736,
    n2744
  );


  and
  g2732
  (
    n2756,
    n2740,
    n2747,
    n2748
  );


  or
  g2733
  (
    n2755,
    n2744,
    n2751,
    n2738,
    n2739
  );


  xor
  g2734
  (
    n2763,
    n2737,
    n2751,
    n2742
  );


  xnor
  g2735
  (
    n2759,
    n2741,
    n2743,
    n2745,
    n2740
  );


  xnor
  g2736
  (
    n2769,
    n2766,
    n146
  );


  not
  g2737
  (
    n2771,
    n209
  );


  nand
  g2738
  (
    n2772,
    n208,
    n2769
  );


  xnor
  g2739
  (
    n2770,
    n2769,
    n209
  );


  not
  g2740
  (
    n2776,
    n2771
  );


  not
  g2741
  (
    n2780,
    n515
  );


  not
  g2742
  (
    n2781,
    n514
  );


  not
  g2743
  (
    n2778,
    n2770
  );


  buf
  g2744
  (
    n2775,
    n2771
  );


  not
  g2745
  (
    n2777,
    n515
  );


  or
  g2746
  (
    n2773,
    n2771,
    n514
  );


  xor
  g2747
  (
    n2774,
    n515,
    n2770,
    n2772
  );


  or
  g2748
  (
    n2779,
    n2772,
    n2740,
    n2770
  );


  or
  g2749
  (
    n2783,
    n2773,
    n2774,
    n2775
  );


  nand
  g2750
  (
    n2784,
    n2774,
    n2773,
    n2775
  );


  nand
  g2751
  (
    n2782,
    n2775,
    n2775,
    n2773,
    n2774
  );


  not
  g2752
  (
    n2792,
    n2783
  );


  buf
  g2753
  (
    n2791,
    n2784
  );


  not
  g2754
  (
    n2785,
    n2782
  );


  not
  g2755
  (
    n2794,
    n2784
  );


  not
  g2756
  (
    n2790,
    n2784
  );


  buf
  g2757
  (
    n2786,
    n2783
  );


  buf
  g2758
  (
    n2787,
    n2784
  );


  buf
  g2759
  (
    n2788,
    n2782
  );


  buf
  g2760
  (
    n2789,
    n2783
  );


  not
  g2761
  (
    n2793,
    n2783
  );


  buf
  g2762
  (
    n2826,
    n210
  );


  buf
  g2763
  (
    n2812,
    n2788
  );


  buf
  g2764
  (
    n2831,
    n2790
  );


  not
  g2765
  (
    n2825,
    n2780
  );


  buf
  g2766
  (
    n2820,
    n2789
  );


  buf
  g2767
  (
    n2809,
    n2777
  );


  xor
  g2768
  (
    n2810,
    n2779,
    n2786,
    n2776
  );


  and
  g2769
  (
    n2822,
    n2790,
    n2791,
    n2720
  );


  or
  g2770
  (
    n2821,
    n2778,
    n545,
    n31
  );


  and
  g2771
  (
    n2827,
    n213,
    n538,
    n545
  );


  or
  g2772
  (
    n2808,
    n2777,
    n32,
    n213
  );


  xor
  g2773
  (
    n2802,
    n2789,
    n2776,
    n540
  );


  xnor
  g2774
  (
    n2804,
    n2788,
    n2794,
    n2786
  );


  xnor
  g2775
  (
    n2798,
    n733,
    n2717,
    n2794
  );


  and
  g2776
  (
    n2834,
    n2793,
    n212,
    n518
  );


  xnor
  g2777
  (
    n2805,
    n540,
    n2719,
    n2791
  );


  nor
  g2778
  (
    n2803,
    n2718,
    n2792,
    n733
  );


  nor
  g2779
  (
    n2830,
    n211,
    n210,
    n2792
  );


  nor
  g2780
  (
    n2823,
    n32,
    n211,
    n2780
  );


  and
  g2781
  (
    n2817,
    n2779,
    n545,
    n2793
  );


  and
  g2782
  (
    n2811,
    n2789,
    n2790,
    n2768
  );


  or
  g2783
  (
    n2800,
    n2788,
    n2793,
    n2780
  );


  xnor
  g2784
  (
    n2799,
    n2786,
    n544,
    n1033
  );


  xor
  g2785
  (
    n2819,
    n2781,
    n2787,
    n2792
  );


  or
  g2786
  (
    n2828,
    n545,
    n516,
    n212
  );


  xor
  g2787
  (
    n2814,
    n2781,
    n2785,
    n2780
  );


  xnor
  g2788
  (
    n2796,
    n2787,
    n2776,
    n2781
  );


  xor
  g2789
  (
    n2832,
    n2794,
    n2790,
    n2776
  );


  nor
  g2790
  (
    n2801,
    n1033,
    n518,
    n211
  );


  nor
  g2791
  (
    n2807,
    n2791,
    n2789,
    n31
  );


  nor
  g2792
  (
    n2806,
    n2779,
    n2778,
    n32
  );


  or
  g2793
  (
    n2816,
    n2779,
    n32,
    n2777
  );


  xnor
  g2794
  (
    n2818,
    n210,
    n211,
    n2781
  );


  xnor
  g2795
  (
    n2813,
    n2721,
    n212,
    n2785
  );


  xnor
  g2796
  (
    n2829,
    n2767,
    n518,
    n2778
  );


  nand
  g2797
  (
    n2795,
    n2794,
    n2786,
    n538
  );


  xor
  g2798
  (
    n2815,
    n2787,
    n2793,
    n2788,
    n2791
  );


  xnor
  g2799
  (
    n2833,
    n2787,
    n538,
    n212,
    n2792
  );


  nor
  g2800
  (
    n2824,
    n2785,
    n2778,
    n540,
    n537
  );


  xnor
  g2801
  (
    n2797,
    n31,
    n210,
    n2785,
    n2777
  );


  xnor
  g2802
  (
    n2903,
    n1825,
    n2810,
    n1885,
    n1849
  );


  nor
  g2803
  (
    n2971,
    n1880,
    n1932,
    n1828,
    n1906
  );


  xnor
  g2804
  (
    n2992,
    n2826,
    n2809,
    n1870,
    n1882
  );


  and
  g2805
  (
    n2945,
    n1896,
    n2819,
    n1847,
    n2808
  );


  xor
  g2806
  (
    n2917,
    n1830,
    n1879,
    n2811,
    n1818
  );


  nor
  g2807
  (
    n2876,
    n1858,
    n2795,
    n1886,
    n1910
  );


  nor
  g2808
  (
    n2927,
    n1913,
    n2807,
    n1882,
    n1921
  );


  xor
  g2809
  (
    n2994,
    n1887,
    n1825,
    n2833,
    n2822
  );


  and
  g2810
  (
    n2862,
    n1919,
    n2797,
    n1820,
    n1877
  );


  xnor
  g2811
  (
    n2850,
    n1900,
    n1880,
    n1897,
    n1844
  );


  or
  g2812
  (
    n2861,
    n1918,
    n1881,
    n1889,
    n1878
  );


  and
  g2813
  (
    n2961,
    n2801,
    n1814,
    n1862,
    n1893
  );


  nand
  g2814
  (
    n2976,
    n1924,
    n2822,
    n2817,
    n1901
  );


  nand
  g2815
  (
    n2886,
    n1874,
    n1928,
    n1888,
    n1903
  );


  xor
  g2816
  (
    n2949,
    n1831,
    n1904,
    n1834,
    n2829
  );


  or
  g2817
  (
    n2879,
    n1919,
    n2825,
    n1892,
    n1836
  );


  nand
  g2818
  (
    n2912,
    n1871,
    n2829,
    n1923,
    n1901
  );


  xor
  g2819
  (
    n2874,
    n1908,
    n2804,
    n1918,
    n1845
  );


  xor
  g2820
  (
    n2911,
    n1895,
    n1906,
    n1892,
    n2800
  );


  nor
  g2821
  (
    n2944,
    n1832,
    n2817,
    n1820,
    n1888
  );


  nand
  g2822
  (
    n2856,
    n1922,
    n1918,
    n2827,
    n1816
  );


  and
  g2823
  (
    n2887,
    n2813,
    n1883,
    n2805,
    n1823
  );


  xnor
  g2824
  (
    n2939,
    n1845,
    n1857,
    n2800,
    n1925
  );


  or
  g2825
  (
    n2851,
    n1840,
    n1865,
    n2804,
    n2806
  );


  xor
  g2826
  (
    n2923,
    n1890,
    n1828,
    n1918,
    n1823
  );


  nand
  g2827
  (
    n2891,
    n1829,
    n1850,
    n2830,
    n1855
  );


  nor
  g2828
  (
    n2942,
    n1814,
    n1816,
    n2823,
    n1881
  );


  xor
  g2829
  (
    n2979,
    n2834,
    n1913,
    n1925,
    n1852
  );


  and
  g2830
  (
    n2962,
    n1815,
    n1832,
    n2825,
    n1924
  );


  nand
  g2831
  (
    n2986,
    n1850,
    n1916,
    n1931,
    n1846
  );


  xor
  g2832
  (
    n2924,
    n1883,
    n1817,
    n1900,
    n1875
  );


  nor
  g2833
  (
    n2852,
    n1841,
    n1840,
    n1865,
    n1858
  );


  or
  g2834
  (
    n2985,
    n1864,
    n1895,
    n1877,
    n1817
  );


  or
  g2835
  (
    n2837,
    n2834,
    n1815,
    n1907,
    n1912
  );


  xor
  g2836
  (
    n2920,
    n1813,
    n1817,
    n2817,
    n2820
  );


  nand
  g2837
  (
    n2877,
    n1897,
    n1869,
    n1822,
    n1889
  );


  nor
  g2838
  (
    n2965,
    n2801,
    n2809,
    n1826,
    n2797
  );


  or
  g2839
  (
    n2964,
    n1853,
    n1829,
    n1849,
    n1913
  );


  nor
  g2840
  (
    n2846,
    n1822,
    n1830,
    n2822,
    n1927
  );


  nor
  g2841
  (
    n2875,
    n2810,
    n1825,
    n1917,
    n1862
  );


  xnor
  g2842
  (
    n2901,
    n1909,
    n2830,
    n2831,
    n1814
  );


  and
  g2843
  (
    n2931,
    n2814,
    n2834,
    n1927,
    n1903
  );


  and
  g2844
  (
    n2839,
    n1838,
    n2824,
    n1846,
    n1867
  );


  xnor
  g2845
  (
    n2935,
    n1915,
    n1888,
    n1862,
    n1838
  );


  nor
  g2846
  (
    n2922,
    n1894,
    n2815,
    n1866,
    n2809
  );


  nor
  g2847
  (
    n2878,
    n2811,
    n2834,
    n1865,
    n2831
  );


  nor
  g2848
  (
    n2840,
    n1901,
    n1863,
    n1931,
    n1860
  );


  xnor
  g2849
  (
    n2937,
    n1875,
    n1891,
    n1833,
    n1894
  );


  nand
  g2850
  (
    n2854,
    n1922,
    n1879,
    n1932,
    n1844
  );


  and
  g2851
  (
    n2870,
    n1846,
    n1914,
    n1921,
    n1821
  );


  xor
  g2852
  (
    n2848,
    n1842,
    n2812,
    n1883,
    n1904
  );


  xnor
  g2853
  (
    n2904,
    n1824,
    n1887,
    n2798,
    n2809
  );


  nor
  g2854
  (
    n2892,
    n1823,
    n1867,
    n1837,
    n1929
  );


  or
  g2855
  (
    n2882,
    n1885,
    n1895,
    n1821,
    n1909
  );


  xor
  g2856
  (
    n2914,
    n2795,
    n1908,
    n1913,
    n1863
  );


  xor
  g2857
  (
    n2950,
    n1911,
    n1871,
    n2810,
    n2812
  );


  nand
  g2858
  (
    n2990,
    n1834,
    n1826,
    n2812,
    n1860
  );


  or
  g2859
  (
    n2955,
    n1880,
    n1869,
    n2823,
    n1877
  );


  and
  g2860
  (
    n2981,
    n1903,
    n1836,
    n1849,
    n1855
  );


  xnor
  g2861
  (
    n2858,
    n2796,
    n2821,
    n1860,
    n1837
  );


  nand
  g2862
  (
    n2889,
    n1853,
    n2828,
    n1932,
    n1899
  );


  or
  g2863
  (
    n2863,
    n2798,
    n1857,
    n2818,
    n1884
  );


  and
  g2864
  (
    n2940,
    n1883,
    n1886,
    n2806,
    n1854
  );


  or
  g2865
  (
    n2991,
    n1857,
    n1905,
    n1861,
    n1821
  );


  and
  g2866
  (
    n2957,
    n1827,
    n1843,
    n1901,
    n1825
  );


  nand
  g2867
  (
    n2841,
    n2818,
    n1837,
    n2821,
    n1872
  );


  xor
  g2868
  (
    n2982,
    n1886,
    n1894,
    n1899,
    n1926
  );


  or
  g2869
  (
    n2910,
    n1854,
    n1835,
    n2797,
    n2799
  );


  or
  g2870
  (
    n2993,
    n2799,
    n1841,
    n2797,
    n2795
  );


  or
  g2871
  (
    n2946,
    n1893,
    n1831,
    n1929,
    n1824
  );


  nand
  g2872
  (
    n2954,
    n1921,
    n1925,
    n2814,
    n1890
  );


  or
  g2873
  (
    n2835,
    n1838,
    n1890,
    n1859,
    n1826
  );


  and
  g2874
  (
    n2936,
    n1818,
    n1930,
    n1856,
    n1904
  );


  nor
  g2875
  (
    n2968,
    n1856,
    n1885,
    n1822,
    n2816
  );


  nor
  g2876
  (
    n2934,
    n2802,
    n2803,
    n2823,
    n1914
  );


  and
  g2877
  (
    n2867,
    n1912,
    n1912,
    n2796,
    n2818
  );


  and
  g2878
  (
    n2869,
    n1823,
    n2802,
    n1888,
    n1931
  );


  nand
  g2879
  (
    n2943,
    n1842,
    n2804,
    n1844,
    n2825
  );


  or
  g2880
  (
    n2972,
    n1881,
    n2819,
    n2827,
    n1900
  );


  and
  g2881
  (
    n2970,
    n1873,
    n1924,
    n1868,
    n1836
  );


  and
  g2882
  (
    n2983,
    n1919,
    n1878,
    n1907,
    n2801
  );


  xor
  g2883
  (
    n2894,
    n1872,
    n2828,
    n2796,
    n1866
  );


  or
  g2884
  (
    n2906,
    n1861,
    n1851,
    n2819,
    n1844
  );


  or
  g2885
  (
    n2909,
    n2833,
    n1892,
    n1819,
    n1840
  );


  or
  g2886
  (
    n2843,
    n1873,
    n2803,
    n2825,
    n1835
  );


  nor
  g2887
  (
    n2872,
    n1893,
    n1911,
    n2826,
    n1896
  );


  nand
  g2888
  (
    n2919,
    n1829,
    n1843,
    n2833,
    n1905
  );


  xor
  g2889
  (
    n2926,
    n1868,
    n1889,
    n1850,
    n1824
  );


  and
  g2890
  (
    n2947,
    n2800,
    n1876,
    n1890,
    n1879
  );


  or
  g2891
  (
    n2888,
    n1902,
    n1900,
    n1911,
    n1873
  );


  and
  g2892
  (
    n2907,
    n1852,
    n2824,
    n1829,
    n1838
  );


  nand
  g2893
  (
    n2905,
    n2821,
    n1827,
    n1875,
    n2807
  );


  nand
  g2894
  (
    n2916,
    n1895,
    n1902,
    n1899,
    n1820
  );


  nand
  g2895
  (
    n2897,
    n1851,
    n1926,
    n1845,
    n1847
  );


  and
  g2896
  (
    n2842,
    n1827,
    n1836,
    n1859,
    n1874
  );


  or
  g2897
  (
    n2938,
    n2811,
    n1862,
    n1819,
    n1835
  );


  or
  g2898
  (
    n2951,
    n1909,
    n1928,
    n1917,
    n1908
  );


  nor
  g2899
  (
    n2975,
    n2826,
    n1866,
    n1867,
    n1842
  );


  or
  g2900
  (
    n2953,
    n1817,
    n1924,
    n2832,
    n1884
  );


  xnor
  g2901
  (
    n2978,
    n1833,
    n1898,
    n1912,
    n2816
  );


  nand
  g2902
  (
    n2928,
    n1930,
    n1914,
    n1858,
    n1926
  );


  xnor
  g2903
  (
    n2845,
    n1848,
    n1818,
    n1893,
    n1821
  );


  or
  g2904
  (
    n2896,
    n1902,
    n1869,
    n2810,
    n2815
  );


  xor
  g2905
  (
    n2974,
    n2832,
    n1870,
    n1906,
    n2820
  );


  and
  g2906
  (
    n2956,
    n1898,
    n1864,
    n1847,
    n1875
  );


  xor
  g2907
  (
    n2925,
    n1872,
    n1813,
    n1925,
    n2833
  );


  or
  g2908
  (
    n2849,
    n1815,
    n1834,
    n1920,
    n1915
  );


  nand
  g2909
  (
    n2963,
    n2830,
    n2800,
    n2821,
    n1840
  );


  or
  g2910
  (
    n2880,
    n1921,
    n1832,
    n2805,
    n1885
  );


  and
  g2911
  (
    n2853,
    n2811,
    n1841,
    n2832,
    n1905
  );


  xnor
  g2912
  (
    n2960,
    n1927,
    n1882,
    n1894,
    n2830
  );


  xor
  g2913
  (
    n2895,
    n1891,
    n2822,
    n1926,
    n1869
  );


  and
  g2914
  (
    n2948,
    n1928,
    n1820,
    n1863,
    n1824
  );


  nor
  g2915
  (
    n2918,
    n1864,
    n1850,
    n2799,
    n2813
  );


  xnor
  g2916
  (
    n2989,
    n2832,
    n1907,
    n2824,
    n1867
  );


  xnor
  g2917
  (
    n2973,
    n1928,
    n1851,
    n1864,
    n1922
  );


  nand
  g2918
  (
    n2988,
    n1911,
    n1833,
    n2819,
    n2820
  );


  xor
  g2919
  (
    n2987,
    n1874,
    n1871,
    n1816,
    n1863
  );


  or
  g2920
  (
    n2921,
    n2799,
    n1866,
    n1814,
    n1932
  );


  xnor
  g2921
  (
    n2857,
    n1855,
    n2828,
    n2805,
    n1846
  );


  xnor
  g2922
  (
    n2860,
    n2815,
    n1828,
    n2814,
    n1910
  );


  xor
  g2923
  (
    n2847,
    n1930,
    n1923,
    n1839
  );


  xnor
  g2924
  (
    n2885,
    n1892,
    n1930,
    n2803,
    n1871
  );


  xnor
  g2925
  (
    n2967,
    n1915,
    n1903,
    n1891,
    n1819
  );


  nand
  g2926
  (
    n2966,
    n2827,
    n1891,
    n1906,
    n1822
  );


  nand
  g2927
  (
    n2952,
    n2826,
    n1855,
    n1914,
    n2795
  );


  xor
  g2928
  (
    n2871,
    n2798,
    n1856,
    n2806,
    n2824
  );


  nor
  g2929
  (
    n2958,
    n1857,
    n1832,
    n1905,
    n1860
  );


  nand
  g2930
  (
    n2929,
    n1909,
    n1816,
    n1876,
    n1815
  );


  and
  g2931
  (
    n2844,
    n2802,
    n1910,
    n1897,
    n1853
  );


  or
  g2932
  (
    n2884,
    n2831,
    n1898,
    n1878,
    n1916
  );


  nand
  g2933
  (
    n2933,
    n1861,
    n2808,
    n2807,
    n2814
  );


  xor
  g2934
  (
    n2890,
    n1870,
    n1842,
    n1898,
    n1813
  );


  nor
  g2935
  (
    n2859,
    n1849,
    n2803,
    n1931,
    n1830
  );


  xor
  g2936
  (
    n2941,
    n1843,
    n1878,
    n1910,
    n1856
  );


  nor
  g2937
  (
    n2866,
    n1848,
    n1922,
    n1841,
    n1884
  );


  xor
  g2938
  (
    n2898,
    n2823,
    n1920,
    n1896
  );


  xnor
  g2939
  (
    n2980,
    n1873,
    n1851,
    n2829,
    n2808
  );


  xnor
  g2940
  (
    n2977,
    n1872,
    n1916,
    n1876
  );


  xnor
  g2941
  (
    n2900,
    n1877,
    n1834,
    n1853,
    n1848
  );


  and
  g2942
  (
    n2899,
    n1868,
    n1826,
    n1813,
    n1847
  );


  xnor
  g2943
  (
    n2873,
    n2804,
    n1828,
    n2813,
    n1819
  );


  xnor
  g2944
  (
    n2959,
    n2827,
    n1904,
    n1868,
    n1831
  );


  xnor
  g2945
  (
    n2913,
    n2796,
    n1848,
    n1839,
    n1870
  );


  xor
  g2946
  (
    n2908,
    n2812,
    n1839,
    n1929,
    n1859
  );


  nor
  g2947
  (
    n2984,
    n2817,
    n1884,
    n1831,
    n1876
  );


  nand
  g2948
  (
    n2915,
    n1859,
    n1852,
    n1854,
    n2802
  );


  nand
  g2949
  (
    n2838,
    n2816,
    n1854,
    n1889,
    n2815
  );


  xor
  g2950
  (
    n2836,
    n1865,
    n1818,
    n1917,
    n2807
  );


  nand
  g2951
  (
    n2930,
    n2801,
    n1915,
    n1917,
    n1887
  );


  nand
  g2952
  (
    n2893,
    n2818,
    n1843,
    n1830,
    n1929
  );


  or
  g2953
  (
    n2969,
    n1852,
    n1874,
    n2808,
    n1919
  );


  nand
  g2954
  (
    n2865,
    n1927,
    n1835,
    n1880,
    n2829
  );


  xor
  g2955
  (
    n2883,
    n1899,
    n2805,
    n2798,
    n1923
  );


  nor
  g2956
  (
    n2902,
    n1907,
    n1882,
    n1920,
    n1827
  );


  xor
  g2957
  (
    n2864,
    n1897,
    n1839,
    n1902,
    n2831
  );


  xor
  g2958
  (
    n2932,
    n1837,
    n1833,
    n1845,
    n1879
  );


  xor
  g2959
  (
    n2855,
    n1896,
    n1861,
    n1886,
    n1881
  );


  and
  g2960
  (
    n2881,
    n2820,
    n2806,
    n1887,
    n1908
  );


  nand
  g2961
  (
    n2868,
    n2828,
    n2813,
    n2816,
    n1858
  );


  xor
  g2962
  (
    n3370,
    n325,
    n248,
    n308,
    n419
  );


  and
  g2963
  (
    n3068,
    n2911,
    n420,
    n2948,
    n2946
  );


  nor
  g2964
  (
    n3138,
    n463,
    n2978,
    n2994,
    n417
  );


  or
  g2965
  (
    n3162,
    n2884,
    n2942,
    n289,
    n2854
  );


  xnor
  g2966
  (
    n3232,
    n477,
    n2965,
    n2849,
    n246
  );


  nand
  g2967
  (
    n3381,
    n462,
    n2306,
    n423,
    n332
  );


  or
  g2968
  (
    n3085,
    n421,
    n319,
    n308,
    n2923
  );


  and
  g2969
  (
    n3482,
    n2976,
    n488,
    n2149,
    n2448
  );


  nor
  g2970
  (
    n3112,
    n286,
    n250,
    n2950,
    n236
  );


  xor
  g2971
  (
    n3366,
    n440,
    n390,
    n2952,
    n418
  );


  xnor
  g2972
  (
    n3211,
    n415,
    n473,
    n2883,
    n2240
  );


  xor
  g2973
  (
    n3461,
    n2676,
    n370,
    n232,
    n292
  );


  xnor
  g2974
  (
    n3516,
    n2712,
    n267,
    n2983,
    n313
  );


  or
  g2975
  (
    n3186,
    n368,
    n2414,
    n2883,
    n2486
  );


  xnor
  g2976
  (
    n3227,
    n441,
    n364,
    n215,
    n381
  );


  and
  g2977
  (
    n3149,
    n2247,
    n2711,
    n2261,
    n280
  );


  and
  g2978
  (
    n3304,
    n2275,
    n275,
    n2972,
    n2940
  );


  xor
  g2979
  (
    n3428,
    n538,
    n2957,
    n382,
    n465
  );


  and
  g2980
  (
    n3209,
    n266,
    n2098,
    n2987,
    n452
  );


  xor
  g2981
  (
    n3564,
    n378,
    n2856,
    n2071,
    n420
  );


  or
  g2982
  (
    n3494,
    n2858,
    n2699,
    n2170,
    n330
  );


  xor
  g2983
  (
    n3574,
    n223,
    n328,
    n2287,
    n2076
  );


  or
  g2984
  (
    n3390,
    n2061,
    n2485,
    n261,
    n464
  );


  nand
  g2985
  (
    n3414,
    n2498,
    n2915,
    n454,
    n2701
  );


  or
  g2986
  (
    n3386,
    n2955,
    n2914,
    n2106,
    n326
  );


  nor
  g2987
  (
    n3114,
    n222,
    n407,
    n2954,
    n216
  );


  or
  g2988
  (
    n3441,
    n2908,
    n2129,
    n474,
    n277
  );


  and
  g2989
  (
    n3631,
    n406,
    n278,
    n398,
    n2537
  );


  or
  g2990
  (
    n3193,
    n2520,
    n2175,
    n2544,
    n2911
  );


  xnor
  g2991
  (
    n3405,
    n2627,
    n2662,
    n491,
    n2346
  );


  xor
  g2992
  (
    n3244,
    n2942,
    n225,
    n2257,
    n437
  );


  and
  g2993
  (
    n3240,
    n2991,
    n2471,
    n2702,
    n2423
  );


  nor
  g2994
  (
    n3460,
    n2194,
    n2236,
    n2880,
    n2200
  );


  xor
  g2995
  (
    n3127,
    n2379,
    n2920,
    n423,
    n359
  );


  xnor
  g2996
  (
    n3348,
    n468,
    n2959,
    n2019,
    n2855
  );


  and
  g2997
  (
    n3418,
    n330,
    n238,
    n2837,
    n310
  );


  or
  g2998
  (
    n3293,
    n2523,
    n432,
    n2474,
    n2921
  );


  nand
  g2999
  (
    n3140,
    n2940,
    n2836,
    n490,
    n2843
  );


  xor
  g3000
  (
    n3259,
    n254,
    n2111,
    n2427,
    n2031
  );


  xnor
  g3001
  (
    n3133,
    n478,
    n407,
    n2699,
    n451
  );


  xnor
  g3002
  (
    n3358,
    n2943,
    n2630,
    n323,
    n2981
  );


  xor
  g3003
  (
    n3159,
    n2140,
    n2499,
    n2036,
    n342
  );


  xnor
  g3004
  (
    n3538,
    n2624,
    n407,
    n227,
    n495
  );


  nor
  g3005
  (
    n3148,
    n2697,
    n232,
    n334,
    n338
  );


  nor
  g3006
  (
    n3335,
    n2851,
    n2913,
    n2228,
    n2225
  );


  xor
  g3007
  (
    n3246,
    n451,
    n2659,
    n2862,
    n488
  );


  xnor
  g3008
  (
    n3583,
    n493,
    n452,
    n496,
    n488
  );


  xnor
  g3009
  (
    n3580,
    n2302,
    n2027,
    n2133,
    n2906
  );


  nor
  g3010
  (
    n3302,
    n2948,
    n2041,
    n2931,
    n2250
  );


  xor
  g3011
  (
    n3618,
    n2875,
    n2169,
    n2512,
    n2367
  );


  xor
  g3012
  (
    n3255,
    n2937,
    n2005,
    n306,
    n2905
  );


  xnor
  g3013
  (
    n3345,
    n2220,
    n2975,
    n405,
    n2099
  );


  and
  g3014
  (
    n3187,
    n2983,
    n2868,
    n413,
    n460
  );


  nand
  g3015
  (
    n3426,
    n316,
    n2882,
    n2304,
    n2962
  );


  xnor
  g3016
  (
    n3478,
    n369,
    n314,
    n2028,
    n2010
  );


  nand
  g3017
  (
    n3152,
    n247,
    n2430,
    n2872,
    n2290
  );


  xnor
  g3018
  (
    n3463,
    n2179,
    n2846,
    n2959,
    n257
  );


  nand
  g3019
  (
    n3183,
    n386,
    n405,
    n312,
    n2888
  );


  nor
  g3020
  (
    n3435,
    n2605,
    n274,
    n2586,
    n2337
  );


  or
  g3021
  (
    n3197,
    n2249,
    n286,
    n2957,
    n2879
  );


  or
  g3022
  (
    n3528,
    n241,
    n2875,
    n2503,
    n2424
  );


  nand
  g3023
  (
    n3089,
    n345,
    n326,
    n428,
    n226
  );


  nand
  g3024
  (
    n3589,
    n342,
    n289,
    n2269,
    n306
  );


  or
  g3025
  (
    n3242,
    n2172,
    n2277,
    n2968,
    n282
  );


  xor
  g3026
  (
    n3515,
    n2035,
    n446,
    n2453,
    n264
  );


  nor
  g3027
  (
    n3230,
    n2990,
    n485,
    n380,
    n2631
  );


  or
  g3028
  (
    n3353,
    n2984,
    n2695,
    n2000,
    n388
  );


  nor
  g3029
  (
    n3373,
    n322,
    n348,
    n2905,
    n380
  );


  xnor
  g3030
  (
    n3363,
    n2899,
    n2494,
    n2946,
    n2316
  );


  or
  g3031
  (
    n3216,
    n354,
    n348,
    n480,
    n2890
  );


  xnor
  g3032
  (
    n3623,
    n402,
    n279,
    n2393,
    n2913
  );


  or
  g3033
  (
    n3079,
    n485,
    n301,
    n2221,
    n2921
  );


  nor
  g3034
  (
    n3207,
    n2159,
    n2243,
    n2296,
    n2708
  );


  nor
  g3035
  (
    n3121,
    n2866,
    n2933,
    n2889,
    n2952
  );


  xnor
  g3036
  (
    n3493,
    n338,
    n2961,
    n477,
    n2901
  );


  nand
  g3037
  (
    n3451,
    n2860,
    n221,
    n2696,
    n367
  );


  xor
  g3038
  (
    n3597,
    n2969,
    n270,
    n2329,
    n2694
  );


  nor
  g3039
  (
    n3104,
    n225,
    n350,
    n2533,
    n2604
  );


  or
  g3040
  (
    n3459,
    n214,
    n2406,
    n327,
    n2935
  );


  xor
  g3041
  (
    n3380,
    n2156,
    n2990,
    n268,
    n2564
  );


  nor
  g3042
  (
    n3178,
    n400,
    n2854,
    n370,
    n2397
  );


  nor
  g3043
  (
    n3020,
    n215,
    n2325,
    n2206,
    n2909
  );


  xor
  g3044
  (
    n3297,
    n2363,
    n268,
    n475,
    n2873
  );


  and
  g3045
  (
    n3412,
    n374,
    n321,
    n2889,
    n494
  );


  or
  g3046
  (
    n3359,
    n2842,
    n2864,
    n375,
    n2846
  );


  and
  g3047
  (
    n3611,
    n450,
    n2874,
    n232,
    n2139
  );


  nand
  g3048
  (
    n3433,
    n2984,
    n423,
    n2917,
    n371
  );


  xor
  g3049
  (
    n3600,
    n272,
    n2878,
    n2925,
    n2887
  );


  or
  g3050
  (
    n3382,
    n468,
    n439,
    n2647,
    n411
  );


  nor
  g3051
  (
    n3462,
    n239,
    n380,
    n381,
    n418
  );


  xnor
  g3052
  (
    n3082,
    n349,
    n237,
    n2283,
    n471
  );


  nor
  g3053
  (
    n3423,
    n291,
    n2924,
    n2903,
    n314
  );


  xor
  g3054
  (
    n3453,
    n2601,
    n2929,
    n2880,
    n2378
  );


  or
  g3055
  (
    n3378,
    n2915,
    n2298,
    n318,
    n228
  );


  nor
  g3056
  (
    n3280,
    n2092,
    n481,
    n343,
    n325
  );


  or
  g3057
  (
    n3629,
    n2054,
    n2579,
    n466,
    n401
  );


  and
  g3058
  (
    n3064,
    n234,
    n296,
    n2590,
    n239
  );


  or
  g3059
  (
    n3278,
    n2978,
    n367,
    n2177,
    n425
  );


  nor
  g3060
  (
    n3111,
    n243,
    n468,
    n242,
    n453
  );


  or
  g3061
  (
    n3000,
    n284,
    n2632,
    n2124,
    n2847
  );


  xnor
  g3062
  (
    n3258,
    n2654,
    n2974,
    n490,
    n2922
  );


  or
  g3063
  (
    n3223,
    n2868,
    n2049,
    n2213,
    n415
  );


  nor
  g3064
  (
    n3265,
    n2923,
    n2876,
    n394,
    n2157
  );


  nand
  g3065
  (
    n3375,
    n480,
    n470,
    n2274,
    n2853
  );


  xnor
  g3066
  (
    n3274,
    n2864,
    n472,
    n319,
    n377
  );


  xnor
  g3067
  (
    n3102,
    n363,
    n422,
    n2938,
    n2706
  );


  xnor
  g3068
  (
    n3062,
    n2881,
    n245,
    n365,
    n2372
  );


  nor
  g3069
  (
    n3055,
    n2202,
    n2073,
    n428,
    n367
  );


  and
  g3070
  (
    n3628,
    n2581,
    n2961,
    n2192,
    n472
  );


  xor
  g3071
  (
    n3058,
    n2930,
    n321,
    n461,
    n234
  );


  and
  g3072
  (
    n3379,
    n2493,
    n2850,
    n2297,
    n2845
  );


  and
  g3073
  (
    n3003,
    n309,
    n2519,
    n473,
    n2925
  );


  and
  g3074
  (
    n3533,
    n340,
    n2853,
    n433,
    n314
  );


  nor
  g3075
  (
    n3267,
    n2695,
    n2839,
    n2895,
    n2417
  );


  and
  g3076
  (
    n3179,
    n216,
    n453,
    n2465,
    n2487
  );


  xnor
  g3077
  (
    n3550,
    n2836,
    n2617,
    n2838,
    n2058
  );


  nand
  g3078
  (
    n3282,
    n2855,
    n2538,
    n278,
    n258
  );


  nor
  g3079
  (
    n3552,
    n2915,
    n393,
    n466,
    n461
  );


  nor
  g3080
  (
    n3481,
    n2842,
    n2950,
    n246,
    n2894
  );


  nand
  g3081
  (
    n3237,
    n2929,
    n2902,
    n2932,
    n389
  );


  xor
  g3082
  (
    n3181,
    n471,
    n2875,
    n259,
    n400
  );


  and
  g3083
  (
    n3499,
    n2207,
    n2560,
    n2841,
    n458
  );


  nor
  g3084
  (
    n3101,
    n2947,
    n2844,
    n385,
    n2890
  );


  nand
  g3085
  (
    n3092,
    n399,
    n2693,
    n2307,
    n2399
  );


  nand
  g3086
  (
    n3588,
    n326,
    n327,
    n484,
    n276
  );


  or
  g3087
  (
    n3344,
    n2899,
    n2033,
    n289,
    n2983
  );


  nor
  g3088
  (
    n3530,
    n214,
    n2237,
    n2929,
    n2892
  );


  and
  g3089
  (
    n3044,
    n357,
    n255,
    n228,
    n221
  );


  xor
  g3090
  (
    n3005,
    n320,
    n2936,
    n385,
    n399
  );


  nand
  g3091
  (
    n3442,
    n485,
    n2566,
    n226,
    n298
  );


  or
  g3092
  (
    n3351,
    n456,
    n2917,
    n2232,
    n2573
  );


  nand
  g3093
  (
    n3213,
    n2850,
    n2864,
    n303,
    n2597
  );


  and
  g3094
  (
    n3444,
    n2021,
    n333,
    n401,
    n2368
  );


  nand
  g3095
  (
    n3142,
    n2398,
    n436,
    n2451,
    n285
  );


  nand
  g3096
  (
    n3024,
    n2989,
    n2059,
    n219,
    n264
  );


  xor
  g3097
  (
    n3201,
    n2935,
    n392,
    n2876,
    n2332
  );


  nand
  g3098
  (
    n3141,
    n373,
    n2039,
    n2475,
    n292
  );


  xor
  g3099
  (
    n3226,
    n2985,
    n2968,
    n244,
    n303
  );


  or
  g3100
  (
    n3483,
    n2936,
    n2701,
    n2842,
    n2886
  );


  and
  g3101
  (
    n3139,
    n375,
    n2112,
    n2884,
    n229
  );


  xnor
  g3102
  (
    n3457,
    n256,
    n2917,
    n364,
    n2419
  );


  xnor
  g3103
  (
    n3314,
    n2911,
    n385,
    n2945,
    n2359
  );


  xor
  g3104
  (
    n3252,
    n2375,
    n2847,
    n2898,
    n2958
  );


  xnor
  g3105
  (
    n3436,
    n2954,
    n2489,
    n2288,
    n2928
  );


  xnor
  g3106
  (
    n3249,
    n307,
    n487,
    n265,
    n2352
  );


  xnor
  g3107
  (
    n3250,
    n298,
    n236,
    n373,
    n2893
  );


  nor
  g3108
  (
    n3383,
    n386,
    n222,
    n347,
    n2705
  );


  and
  g3109
  (
    n3455,
    n2138,
    n2878,
    n339,
    n2510
  );


  xnor
  g3110
  (
    n3050,
    n497,
    n2318,
    n242,
    n2713
  );


  and
  g3111
  (
    n3376,
    n2979,
    n2069,
    n2933,
    n481
  );


  nor
  g3112
  (
    n3416,
    n491,
    n2428,
    n2280,
    n2967
  );


  nand
  g3113
  (
    n3155,
    n237,
    n455,
    n2480,
    n267
  );


  nor
  g3114
  (
    n3231,
    n388,
    n2246,
    n2979,
    n309
  );


  xor
  g3115
  (
    n3194,
    n2515,
    n2916,
    n2946,
    n2964
  );


  xor
  g3116
  (
    n3225,
    n2900,
    n2707,
    n2167,
    n2990
  );


  and
  g3117
  (
    n3347,
    n2987,
    n2893,
    n315,
    n2994
  );


  or
  g3118
  (
    n3484,
    n2550,
    n2704,
    n434,
    n2184
  );


  nor
  g3119
  (
    n3042,
    n2939,
    n337,
    n296,
    n2941
  );


  and
  g3120
  (
    n3610,
    n2918,
    n2931,
    n2835,
    n2964
  );


  nor
  g3121
  (
    n3001,
    n257,
    n2900,
    n2371,
    n445
  );


  xor
  g3122
  (
    n3184,
    n2867,
    n270,
    n333,
    n433
  );


  xor
  g3123
  (
    n3458,
    n2859,
    n331,
    n2044,
    n2852
  );


  and
  g3124
  (
    n3073,
    n2840,
    n2311,
    n248,
    n2122
  );


  xor
  g3125
  (
    n3596,
    n359,
    n2292,
    n2835,
    n2994
  );


  xor
  g3126
  (
    n3571,
    n216,
    n363,
    n2907,
    n2892
  );


  or
  g3127
  (
    n3339,
    n214,
    n437,
    n2950,
    n2365
  );


  xor
  g3128
  (
    n3254,
    n2037,
    n2658,
    n300,
    n410
  );


  or
  g3129
  (
    n3132,
    n2847,
    n464,
    n317,
    n427
  );


  and
  g3130
  (
    n3269,
    n2936,
    n2901,
    n283,
    n2610
  );


  and
  g3131
  (
    n3377,
    n2251,
    n357,
    n307,
    n403
  );


  nand
  g3132
  (
    n3584,
    n2421,
    n329,
    n2248,
    n2646
  );


  nand
  g3133
  (
    n3535,
    n2145,
    n495,
    n282,
    n472
  );


  or
  g3134
  (
    n3498,
    n2902,
    n2945,
    n2340,
    n338
  );


  or
  g3135
  (
    n3321,
    n2939,
    n2016,
    n2443,
    n261
  );


  or
  g3136
  (
    n3521,
    n325,
    n2458,
    n2949,
    n2906
  );


  or
  g3137
  (
    n3248,
    n2983,
    n2420,
    n347,
    n486
  );


  and
  g3138
  (
    n3061,
    n2858,
    n391,
    n213,
    n456
  );


  xor
  g3139
  (
    n3115,
    n381,
    n277,
    n443,
    n2850
  );


  xnor
  g3140
  (
    n3561,
    n297,
    n2038,
    n2075,
    n2856
  );


  nor
  g3141
  (
    n3427,
    n2353,
    n2518,
    n372,
    n2216
  );


  xnor
  g3142
  (
    n3276,
    n2879,
    n443,
    n2850,
    n243
  );


  xor
  g3143
  (
    n3558,
    n349,
    n2120,
    n2907,
    n2935
  );


  or
  g3144
  (
    n3595,
    n295,
    n2910,
    n260,
    n409
  );


  nor
  g3145
  (
    n3497,
    n233,
    n2980,
    n2703,
    n2198
  );


  xor
  g3146
  (
    n3326,
    n2691,
    n2703,
    n458,
    n2190
  );


  xnor
  g3147
  (
    n3220,
    n2976,
    n232,
    n2927,
    n2707
  );


  xor
  g3148
  (
    n3091,
    n2259,
    n2931,
    n294,
    n2118
  );


  and
  g3149
  (
    n3298,
    n268,
    n492,
    n2963,
    n331
  );


  xor
  g3150
  (
    n3257,
    n2657,
    n2123,
    n435,
    n2845
  );


  or
  g3151
  (
    n3431,
    n2985,
    n2125,
    n2879,
    n2293
  );


  xnor
  g3152
  (
    n3099,
    n335,
    n2947,
    n2963,
    n2971
  );


  xor
  g3153
  (
    n3475,
    n429,
    n2574,
    n2951,
    n2973
  );


  xor
  g3154
  (
    n3430,
    n2867,
    n226,
    n278,
    n2326
  );


  nor
  g3155
  (
    n3292,
    n280,
    n2583,
    n2050,
    n2908
  );


  nand
  g3156
  (
    n3158,
    n2386,
    n296,
    n2849,
    n2260
  );


  or
  g3157
  (
    n3320,
    n282,
    n440,
    n371,
    n281
  );


  xor
  g3158
  (
    n3546,
    n273,
    n255,
    n366,
    n433
  );


  nand
  g3159
  (
    n3434,
    n459,
    n219,
    n378,
    n2954
  );


  xor
  g3160
  (
    n3038,
    n394,
    n240,
    n404,
    n2128
  );


  nand
  g3161
  (
    n3272,
    n2835,
    n312,
    n2253,
    n2299
  );


  xor
  g3162
  (
    n3266,
    n2965,
    n2887,
    n2452,
    n382
  );


  xor
  g3163
  (
    n3367,
    n249,
    n248,
    n2018,
    n2439
  );


  nand
  g3164
  (
    n3425,
    n2843,
    n430,
    n2934,
    n457
  );


  nor
  g3165
  (
    n3054,
    n427,
    n2415,
    n496,
    n310
  );


  or
  g3166
  (
    n3217,
    n2578,
    n2433,
    n244,
    n2330
  );


  xor
  g3167
  (
    n3072,
    n2934,
    n2319,
    n231,
    n417
  );


  xor
  g3168
  (
    n3330,
    n2700,
    n429,
    n2844,
    n2881
  );


  nand
  g3169
  (
    n3466,
    n253,
    n2079,
    n354,
    n438
  );


  xnor
  g3170
  (
    n3598,
    n318,
    n2705,
    n430,
    n240
  );


  nor
  g3171
  (
    n3076,
    n324,
    n2582,
    n2838,
    n2350
  );


  xor
  g3172
  (
    n3349,
    n378,
    n220,
    n257,
    n2057
  );


  and
  g3173
  (
    n3137,
    n383,
    n263,
    n248,
    n2315
  );


  nand
  g3174
  (
    n3519,
    n224,
    n2966,
    n2880,
    n2690
  );


  xor
  g3175
  (
    n3361,
    n2392,
    n2703,
    n2976,
    n426
  );


  nor
  g3176
  (
    n3198,
    n413,
    n2943,
    n2933,
    n2837
  );


  nand
  g3177
  (
    n3300,
    n436,
    n354,
    n233,
    n384
  );


  nand
  g3178
  (
    n3243,
    n2535,
    n2700,
    n2703,
    n2920
  );


  xnor
  g3179
  (
    n3395,
    n384,
    n2854,
    n2977,
    n2960
  );


  or
  g3180
  (
    n3019,
    n2173,
    n2986,
    n2991,
    n2215
  );


  xor
  g3181
  (
    n3454,
    n2904,
    n257,
    n2857,
    n408
  );


  xnor
  g3182
  (
    n3513,
    n2483,
    n2877,
    n224,
    n2464
  );


  nand
  g3183
  (
    n3575,
    n2871,
    n395,
    n374,
    n2837
  );


  xnor
  g3184
  (
    n3568,
    n2110,
    n321,
    n2121,
    n292
  );


  xnor
  g3185
  (
    n3191,
    n351,
    n340,
    n385,
    n2638
  );


  nand
  g3186
  (
    n3236,
    n273,
    n2096,
    n467,
    n2154
  );


  nor
  g3187
  (
    n3371,
    n475,
    n2109,
    n2866,
    n2838
  );


  xnor
  g3188
  (
    n3200,
    n379,
    n479,
    n462,
    n2881
  );


  xor
  g3189
  (
    n3066,
    n2876,
    n2020,
    n2870,
    n2095
  );


  xnor
  g3190
  (
    n3356,
    n307,
    n2904,
    n425,
    n263
  );


  or
  g3191
  (
    n3017,
    n393,
    n2301,
    n331,
    n404
  );


  nand
  g3192
  (
    n3409,
    n2007,
    n2546,
    n421,
    n2218
  );


  or
  g3193
  (
    n3124,
    n2234,
    n2956,
    n2896,
    n341
  );


  or
  g3194
  (
    n3310,
    n2835,
    n377,
    n309,
    n2967
  );


  nor
  g3195
  (
    n3438,
    n2162,
    n2960,
    n2193,
    n2990
  );


  or
  g3196
  (
    n3545,
    n2664,
    n241,
    n2107,
    n301
  );


  or
  g3197
  (
    n3009,
    n2591,
    n395,
    n337,
    n217
  );


  and
  g3198
  (
    n3060,
    n2565,
    n2002,
    n2970,
    n2896
  );


  nand
  g3199
  (
    n3608,
    n2712,
    n2979,
    n263,
    n2844
  );


  or
  g3200
  (
    n3422,
    n2295,
    n1995,
    n2988,
    n2077
  );


  nand
  g3201
  (
    n3399,
    n469,
    n2629,
    n478,
    n2620
  );


  and
  g3202
  (
    n3202,
    n409,
    n329,
    n252,
    n415
  );


  nand
  g3203
  (
    n3372,
    n294,
    n2900,
    n306,
    n2067
  );


  nor
  g3204
  (
    n3027,
    n2839,
    n2648,
    n2572,
    n251
  );


  xor
  g3205
  (
    n3578,
    n332,
    n454,
    n2344,
    n2912
  );


  xor
  g3206
  (
    n3270,
    n228,
    n396,
    n382,
    n2239
  );


  or
  g3207
  (
    n3234,
    n431,
    n465,
    n287,
    n2993
  );


  nor
  g3208
  (
    n3403,
    n2407,
    n459,
    n308,
    n2937
  );


  and
  g3209
  (
    n3168,
    n459,
    n2974,
    n415,
    n2459
  );


  xor
  g3210
  (
    n3522,
    n2045,
    n2323,
    n241,
    n286
  );


  and
  g3211
  (
    n3603,
    n305,
    n358,
    n2022,
    n2914
  );


  nand
  g3212
  (
    n3008,
    n390,
    n2074,
    n250,
    n252
  );


  xor
  g3213
  (
    n3107,
    n445,
    n2147,
    n2476,
    n2861
  );


  xor
  g3214
  (
    n3113,
    n2273,
    n424,
    n2376,
    n2940
  );


  xnor
  g3215
  (
    n3262,
    n2984,
    n372,
    n2849,
    n2988
  );


  xor
  g3216
  (
    n3607,
    n448,
    n327,
    n2637,
    n2956
  );


  xnor
  g3217
  (
    n3354,
    n2963,
    n478,
    n2083,
    n2698
  );


  xor
  g3218
  (
    n3065,
    n2909,
    n2222,
    n2491,
    n2980
  );


  or
  g3219
  (
    n3296,
    n419,
    n451,
    n482,
    n2314
  );


  nand
  g3220
  (
    n3592,
    n2962,
    n380,
    n2023,
    n2644
  );


  xnor
  g3221
  (
    n3165,
    n2126,
    n2357,
    n2151,
    n2671
  );


  xor
  g3222
  (
    n3273,
    n2116,
    n321,
    n2900,
    n449
  );


  nor
  g3223
  (
    n3057,
    n2672,
    n2973,
    n2977,
    n496
  );


  nand
  g3224
  (
    n3456,
    n2896,
    n355,
    n253,
    n2705
  );


  nand
  g3225
  (
    n3539,
    n318,
    n2256,
    n2974,
    n323
  );


  nand
  g3226
  (
    n3486,
    n2103,
    n2987,
    n476,
    n2242
  );


  and
  g3227
  (
    n3264,
    n274,
    n2599,
    n341,
    n2015
  );


  xor
  g3228
  (
    n3318,
    n218,
    n2444,
    n2343,
    n2279
  );


  and
  g3229
  (
    n3328,
    n336,
    n467,
    n2258,
    n2947
  );


  nand
  g3230
  (
    n3573,
    n274,
    n2105,
    n2972,
    n2856
  );


  nor
  g3231
  (
    n3524,
    n239,
    n2066,
    n2992,
    n2043
  );


  xor
  g3232
  (
    n3447,
    n412,
    n298,
    n278,
    n2596
  );


  or
  g3233
  (
    n3450,
    n2543,
    n299,
    n235,
    n401
  );


  or
  g3234
  (
    n3180,
    n1997,
    n397,
    n343,
    n315
  );


  nand
  g3235
  (
    n3224,
    n2839,
    n2369,
    n2972,
    n2843
  );


  nor
  g3236
  (
    n3253,
    n2100,
    n2626,
    n2956,
    n293
  );


  xnor
  g3237
  (
    n3160,
    n333,
    n2466,
    n354,
    n434
  );


  nand
  g3238
  (
    n3540,
    n226,
    n391,
    n2361,
    n2348
  );


  or
  g3239
  (
    n3620,
    n448,
    n360,
    n376,
    n2142
  );


  nor
  g3240
  (
    n3408,
    n2871,
    n2677,
    n260,
    n290
  );


  and
  g3241
  (
    n3565,
    n484,
    n426,
    n2354,
    n2924
  );


  nand
  g3242
  (
    n3077,
    n221,
    n322,
    n331,
    n490
  );


  and
  g3243
  (
    n3541,
    n473,
    n2922,
    n361,
    n2978
  );


  nor
  g3244
  (
    n3315,
    n419,
    n2964,
    n2003,
    n2866
  );


  xnor
  g3245
  (
    n3313,
    n2166,
    n350,
    n2004,
    n2707
  );


  and
  g3246
  (
    n3199,
    n408,
    n320,
    n2913,
    n431
  );


  xnor
  g3247
  (
    n3281,
    n295,
    n2085,
    n2891,
    n440
  );


  xor
  g3248
  (
    n3134,
    n2910,
    n292,
    n2887,
    n2463
  );


  and
  g3249
  (
    n3083,
    n2863,
    n2992,
    n2693,
    n2847
  );


  nand
  g3250
  (
    n3510,
    n420,
    n2704,
    n2945,
    n335
  );


  xnor
  g3251
  (
    n3306,
    n343,
    n490,
    n334,
    n413
  );


  nand
  g3252
  (
    n3387,
    n220,
    n2117,
    n2209,
    n239
  );


  xor
  g3253
  (
    n3593,
    n407,
    n277,
    n330,
    n2700
  );


  or
  g3254
  (
    n3245,
    n2944,
    n2653,
    n485,
    n2390
  );


  nand
  g3255
  (
    n3150,
    n438,
    n368,
    n2255,
    n2934
  );


  and
  g3256
  (
    n3123,
    n359,
    n2882,
    n2187,
    n312
  );


  nor
  g3257
  (
    n3256,
    n313,
    n285,
    n2916,
    n2938
  );


  or
  g3258
  (
    n3411,
    n2639,
    n2370,
    n339,
    n495
  );


  or
  g3259
  (
    n3415,
    n2457,
    n471,
    n300,
    n335
  );


  xnor
  g3260
  (
    n3268,
    n276,
    n441,
    n2683
  );


  nor
  g3261
  (
    n3290,
    n2431,
    n2204,
    n2470,
    n378
  );


  xor
  g3262
  (
    n3452,
    n376,
    n2708,
    n404,
    n235
  );


  nor
  g3263
  (
    n3239,
    n497,
    n2901,
    n335,
    n421
  );


  nor
  g3264
  (
    n3566,
    n259,
    n2969,
    n2091,
    n2941
  );


  nand
  g3265
  (
    n3404,
    n263,
    n2872,
    n288,
    n2899
  );


  or
  g3266
  (
    n3324,
    n2959,
    n399,
    n2053,
    n260
  );


  or
  g3267
  (
    n3176,
    n2970,
    n2951,
    n2685,
    n282
  );


  nand
  g3268
  (
    n3175,
    n364,
    n2939,
    n465,
    n2196
  );


  xnor
  g3269
  (
    n3214,
    n2508,
    n2689,
    n317,
    n2481
  );


  xor
  g3270
  (
    n3503,
    n2926,
    n2148,
    n455,
    n2953
  );


  or
  g3271
  (
    n3156,
    n460,
    n346,
    n352,
    n408
  );


  xnor
  g3272
  (
    n3075,
    n2101,
    n2922,
    n2890,
    n2235
  );


  or
  g3273
  (
    n3170,
    n2971,
    n2373,
    n2882,
    n273
  );


  or
  g3274
  (
    n3472,
    n2913,
    n338,
    n2645,
    n2446
  );


  nand
  g3275
  (
    n3145,
    n2408,
    n476,
    n2956,
    n253
  );


  xor
  g3276
  (
    n3308,
    n2040,
    n2609,
    n290,
    n295
  );


  nor
  g3277
  (
    n3577,
    n2556,
    n2867,
    n458,
    n2072
  );


  nor
  g3278
  (
    n3049,
    n410,
    n2898,
    n347,
    n480
  );


  xnor
  g3279
  (
    n3518,
    n487,
    n324,
    n358,
    n2993
  );


  nor
  g3280
  (
    n3074,
    n364,
    n2014,
    n474,
    n2704
  );


  nand
  g3281
  (
    n3120,
    n350,
    n319,
    n2936,
    n242
  );


  xnor
  g3282
  (
    n3025,
    n2943,
    n302,
    n494,
    n2479
  );


  or
  g3283
  (
    n3398,
    n2294,
    n387,
    n2532,
    n390
  );


  nand
  g3284
  (
    n3247,
    n345,
    n2263,
    n293,
    n2905
  );


  or
  g3285
  (
    n3277,
    n2919,
    n489,
    n2840,
    n486
  );


  nand
  g3286
  (
    n3594,
    n426,
    n2602,
    n2898,
    n484
  );


  nand
  g3287
  (
    n3471,
    n325,
    n2080,
    n398,
    n2978
  );


  nand
  g3288
  (
    n3606,
    n2495,
    n271,
    n470,
    n2888
  );


  and
  g3289
  (
    n3036,
    n320,
    n2855,
    n474,
    n307
  );


  and
  g3290
  (
    n3086,
    n293,
    n2885,
    n2709,
    n2584
  );


  xnor
  g3291
  (
    n3014,
    n2017,
    n2836,
    n459,
    n2852
  );


  xor
  g3292
  (
    n3161,
    n489,
    n2866,
    n2908,
    n369
  );


  xor
  g3293
  (
    n3144,
    n222,
    n434,
    n2513,
    n350
  );


  xnor
  g3294
  (
    n3617,
    n2580,
    n2872,
    n2405,
    n311
  );


  xor
  g3295
  (
    n3343,
    n2137,
    n2855,
    n371,
    n2402
  );


  or
  g3296
  (
    n3185,
    n444,
    n342,
    n2034,
    n339
  );


  nand
  g3297
  (
    n3143,
    n397,
    n487,
    n2966,
    n2937
  );


  nand
  g3298
  (
    n3601,
    n2545,
    n265,
    n2851,
    n2921
  );


  and
  g3299
  (
    n2998,
    n2548,
    n2945,
    n2908,
    n2656
  );


  nand
  g3300
  (
    n3307,
    n2843,
    n445,
    n323,
    n2863
  );


  and
  g3301
  (
    n3291,
    n479,
    n2230,
    n2916,
    n456
  );


  and
  g3302
  (
    n3196,
    n427,
    n2967,
    n2231,
    n2891
  );


  and
  g3303
  (
    n3045,
    n388,
    n2526,
    n2661,
    n2853
  );


  xnor
  g3304
  (
    n3334,
    n2944,
    n265,
    n353,
    n409
  );


  xnor
  g3305
  (
    n3177,
    n315,
    n2199,
    n2455,
    n255
  );


  xor
  g3306
  (
    n3039,
    n2941,
    n2853,
    n2467,
    n2933
  );


  and
  g3307
  (
    n3400,
    n2701,
    n2384,
    n289,
    n291
  );


  or
  g3308
  (
    n3401,
    n308,
    n246,
    n2881,
    n448
  );


  nand
  g3309
  (
    n2997,
    n2924,
    n2366,
    n288,
    n284
  );


  or
  g3310
  (
    n3473,
    n234,
    n2891,
    n360,
    n2585
  );


  or
  g3311
  (
    n3251,
    n2982,
    n353,
    n2178,
    n2870
  );


  nand
  g3312
  (
    n3369,
    n384,
    n2973,
    n2869,
    n2387
  );


  xnor
  g3313
  (
    n3619,
    n2563,
    n411,
    n2852,
    n2943
  );


  xnor
  g3314
  (
    n3591,
    n2102,
    n272,
    n341,
    n2932
  );


  nand
  g3315
  (
    n3195,
    n2906,
    n2926,
    n2383,
    n2885
  );


  nor
  g3316
  (
    n3294,
    n373,
    n2987,
    n217,
    n2603
  );


  and
  g3317
  (
    n3167,
    n422,
    n2935,
    n355,
    n2897
  );


  nor
  g3318
  (
    n3260,
    n2951,
    n345,
    n247,
    n434
  );


  xnor
  g3319
  (
    n3621,
    n2401,
    n328,
    n2404,
    n362
  );


  xnor
  g3320
  (
    n3051,
    n450,
    n2883,
    n2915,
    n430
  );


  and
  g3321
  (
    n3029,
    n2836,
    n2906,
    n2865,
    n2410
  );


  xnor
  g3322
  (
    n3235,
    n2272,
    n2974,
    n295,
    n233
  );


  and
  g3323
  (
    n3118,
    n285,
    n422,
    n455,
    n2201
  );


  xnor
  g3324
  (
    n3616,
    n2912,
    n2525,
    n2278,
    n281
  );


  nor
  g3325
  (
    n3437,
    n220,
    n2957,
    n247,
    n2621
  );


  or
  g3326
  (
    n3069,
    n314,
    n259,
    n255,
    n2949
  );


  nor
  g3327
  (
    n3626,
    n357,
    n324,
    n2973,
    n2898
  );


  nand
  g3328
  (
    n3553,
    n2953,
    n2561,
    n2636,
    n2944
  );


  and
  g3329
  (
    n3443,
    n394,
    n401,
    n2289,
    n2961
  );


  nand
  g3330
  (
    n3215,
    n2338,
    n2497,
    n360,
    n1999
  );


  nor
  g3331
  (
    n3295,
    n2270,
    n262,
    n2171,
    n1996
  );


  xnor
  g3332
  (
    n3288,
    n319,
    n400,
    n2113,
    n414
  );


  nor
  g3333
  (
    n3586,
    n483,
    n2135,
    n2893,
    n2511
  );


  and
  g3334
  (
    n3534,
    n2713,
    n2971,
    n2197,
    n2660
  );


  xnor
  g3335
  (
    n3125,
    n486,
    n2930,
    n483,
    n2223
  );


  and
  g3336
  (
    n3128,
    n475,
    n251,
    n2084,
    n2953
  );


  nor
  g3337
  (
    n3053,
    n406,
    n2155,
    n2955,
    n2358
  );


  and
  g3338
  (
    n3261,
    n397,
    n2029,
    n2233,
    n379
  );


  nand
  g3339
  (
    n3590,
    n304,
    n392,
    n2865,
    n240
  );


  and
  g3340
  (
    n3350,
    n2962,
    n425,
    n230,
    n303
  );


  xor
  g3341
  (
    n3559,
    n2980,
    n2334,
    n410,
    n395
  );


  xor
  g3342
  (
    n3203,
    n2705,
    n2902,
    n2712,
    n322
  );


  nand
  g3343
  (
    n3543,
    n2211,
    n2426,
    n2699,
    n447
  );


  nand
  g3344
  (
    n3095,
    n475,
    n437,
    n2349,
    n2693
  );


  xnor
  g3345
  (
    n3100,
    n377,
    n2130,
    n224,
    n2529
  );


  xor
  g3346
  (
    n3043,
    n2968,
    n2970,
    n256,
    n299
  );


  nand
  g3347
  (
    n3572,
    n249,
    n472,
    n383,
    n429
  );


  xor
  g3348
  (
    n3037,
    n497,
    n392,
    n330,
    n2934
  );


  and
  g3349
  (
    n3492,
    n2902,
    n352,
    n2894,
    n2858
  );


  xor
  g3350
  (
    n3153,
    n2244,
    n281,
    n2667,
    n2642
  );


  nand
  g3351
  (
    n3560,
    n271,
    n2849,
    n2857,
    n2611
  );


  xnor
  g3352
  (
    n3507,
    n231,
    n2063,
    n2869,
    n404
  );


  nor
  g3353
  (
    n3479,
    n2612,
    n2445,
    n376,
    n2958
  );


  xor
  g3354
  (
    n3228,
    n480,
    n469,
    n231,
    n2473
  );


  nor
  g3355
  (
    n3011,
    n2174,
    n493,
    n2227,
    n474
  );


  and
  g3356
  (
    n3500,
    n2975,
    n276,
    n2669,
    n2869
  );


  nand
  g3357
  (
    n3322,
    n468,
    n2088,
    n242,
    n2895
  );


  nand
  g3358
  (
    n3346,
    n218,
    n288,
    n400,
    n2655
  );


  and
  g3359
  (
    n3013,
    n317,
    n274,
    n2394,
    n2490
  );


  nand
  g3360
  (
    n3105,
    n223,
    n2879,
    n417,
    n2185
  );


  nand
  g3361
  (
    n3096,
    n339,
    n281,
    n251,
    n2909
  );


  xor
  g3362
  (
    n3208,
    n2942,
    n389,
    n446,
    n435
  );


  nand
  g3363
  (
    n3206,
    n245,
    n2888,
    n396,
    n270
  );


  xor
  g3364
  (
    n3021,
    n453,
    n2460,
    n2869,
    n301
  );


  and
  g3365
  (
    n3317,
    n2679,
    n457,
    n250,
    n264
  );


  nand
  g3366
  (
    n3305,
    n2011,
    n2941,
    n2097,
    n2606
  );


  xor
  g3367
  (
    n3279,
    n2530,
    n2958,
    n2615,
    n2441
  );


  or
  g3368
  (
    n3033,
    n2895,
    n360,
    n483,
    n2914
  );


  nand
  g3369
  (
    n3041,
    n2412,
    n452,
    n2968,
    n2008
  );


  nand
  g3370
  (
    n3487,
    n373,
    n275,
    n2633,
    n2985
  );


  xnor
  g3371
  (
    n3147,
    n467,
    n363,
    n477,
    n2195
  );


  or
  g3372
  (
    n3238,
    n2887,
    n290,
    n2840,
    n403
  );


  xnor
  g3373
  (
    n3396,
    n2542,
    n2873,
    n2700,
    n2891
  );


  xor
  g3374
  (
    n3384,
    n2878,
    n365,
    n2450,
    n2702
  );


  nor
  g3375
  (
    n3164,
    n265,
    n2904,
    n2926,
    n2505
  );


  xnor
  g3376
  (
    n3508,
    n411,
    n433,
    n2963,
    n2454
  );


  nor
  g3377
  (
    n3609,
    n2976,
    n2087,
    n340,
    n489
  );


  nor
  g3378
  (
    n3002,
    n2948,
    n493,
    n395,
    n2065
  );


  or
  g3379
  (
    n3166,
    n236,
    n328,
    n2903,
    n2897
  );


  xnor
  g3380
  (
    n3146,
    n2865,
    n376,
    n2527,
    n486
  );


  xnor
  g3381
  (
    n2999,
    n462,
    n2952,
    n2380,
    n2189
  );


  xnor
  g3382
  (
    n3006,
    n2324,
    n414,
    n2262,
    n2665
  );


  or
  g3383
  (
    n3284,
    n2713,
    n310,
    n361,
    n2927
  );


  xor
  g3384
  (
    n3117,
    n2183,
    n2884,
    n2706,
    n2484
  );


  nand
  g3385
  (
    n3576,
    n333,
    n2663,
    n2871,
    n2500
  );


  or
  g3386
  (
    n3529,
    n2925,
    n2988,
    n235,
    n2875
  );


  nand
  g3387
  (
    n3323,
    n2970,
    n491,
    n2469,
    n2594
  );


  and
  g3388
  (
    n3299,
    n2845,
    n2962,
    n2874,
    n2598
  );


  or
  g3389
  (
    n3219,
    n2965,
    n276,
    n2482,
    n229
  );


  nor
  g3390
  (
    n3342,
    n389,
    n2870,
    n2425,
    n2682
  );


  nor
  g3391
  (
    n3275,
    n2064,
    n316,
    n230,
    n2026
  );


  xnor
  g3392
  (
    n3097,
    n254,
    n323,
    n2992,
    n2271
  );


  xnor
  g3393
  (
    n3567,
    n2986,
    n2181,
    n2883,
    n2921
  );


  nand
  g3394
  (
    n3579,
    n2203,
    n439,
    n2468,
    n2981
  );


  or
  g3395
  (
    n3614,
    n2868,
    n2985,
    n225,
    n416
  );


  and
  g3396
  (
    n3440,
    n2416,
    n379,
    n2570,
    n304
  );


  nor
  g3397
  (
    n3316,
    n432,
    n2267,
    n2333,
    n2335
  );


  nor
  g3398
  (
    n3205,
    n304,
    n2874,
    n2888,
    n2078
  );


  and
  g3399
  (
    n3365,
    n439,
    n269,
    n300,
    n290
  );


  or
  g3400
  (
    n3448,
    n2988,
    n2969,
    n302,
    n2141
  );


  nor
  g3401
  (
    n3393,
    n2857,
    n2303,
    n269,
    n349
  );


  and
  g3402
  (
    n3028,
    n2205,
    n412,
    n2528,
    n273
  );


  xor
  g3403
  (
    n3421,
    n2984,
    n2914,
    n336,
    n482
  );


  xnor
  g3404
  (
    n3634,
    n227,
    n2006,
    n266,
    n2895
  );


  xor
  g3405
  (
    n3622,
    n258,
    n452,
    n2711,
    n449
  );


  and
  g3406
  (
    n3046,
    n2449,
    n454,
    n2929,
    n268
  );


  nand
  g3407
  (
    n3007,
    n272,
    n2882,
    n2955,
    n2841
  );


  or
  g3408
  (
    n3465,
    n398,
    n2567,
    n2186,
    n287
  );


  nor
  g3409
  (
    n3420,
    n2993,
    n2070,
    n2042,
    n214
  );


  xor
  g3410
  (
    n3476,
    n348,
    n2188,
    n466,
    n2524
  );


  or
  g3411
  (
    n3490,
    n2708,
    n2613,
    n2885,
    n426
  );


  xnor
  g3412
  (
    n3056,
    n2168,
    n421,
    n473,
    n442
  );


  or
  g3413
  (
    n3581,
    n2132,
    n358,
    n340,
    n2687
  );


  or
  g3414
  (
    n3035,
    n469,
    n2864,
    n481,
    n2958
  );


  nand
  g3415
  (
    n3015,
    n2150,
    n2697,
    n309,
    n2957
  );


  or
  g3416
  (
    n3523,
    n424,
    n2442,
    n297,
    n2860
  );


  or
  g3417
  (
    n3544,
    n267,
    n492,
    n464,
    n305
  );


  or
  g3418
  (
    n3477,
    n443,
    n379,
    n462,
    n2907
  );


  xor
  g3419
  (
    n3080,
    n479,
    n372,
    n389,
    n482
  );


  xnor
  g3420
  (
    n3063,
    n2706,
    n494,
    n280,
    n2356
  );


  xnor
  g3421
  (
    n3352,
    n297,
    n241,
    n362,
    n284
  );


  and
  g3422
  (
    n3012,
    n2047,
    n2616,
    n460,
    n245
  );


  nor
  g3423
  (
    n3406,
    n337,
    n2649,
    n2904,
    n262
  );


  or
  g3424
  (
    n3047,
    n2878,
    n2859,
    n222,
    n2710
  );


  xnor
  g3425
  (
    n3204,
    n2322,
    n2589,
    n2694,
    n305
  );


  nand
  g3426
  (
    n3098,
    n2502,
    n2555,
    n386,
    n387
  );


  and
  g3427
  (
    n3030,
    n387,
    n406,
    n250,
    n2857
  );


  or
  g3428
  (
    n3419,
    n2928,
    n2967,
    n262,
    n391
  );


  or
  g3429
  (
    n3094,
    n374,
    n2880,
    n2547,
    n2534
  );


  xnor
  g3430
  (
    n3509,
    n224,
    n2684,
    n2310,
    n443
  );


  or
  g3431
  (
    n3502,
    n2678,
    n221,
    n256,
    n488
  );


  xor
  g3432
  (
    n3286,
    n405,
    n390,
    n2395,
    n2712
  );


  xor
  g3433
  (
    n3135,
    n2389,
    n2951,
    n497,
    n2919
  );


  or
  g3434
  (
    n3374,
    n356,
    n238,
    n2127,
    n2873
  );


  and
  g3435
  (
    n3446,
    n2907,
    n2917,
    n313,
    n2923
  );


  xnor
  g3436
  (
    n3397,
    n403,
    n1993,
    n366,
    n467
  );


  nor
  g3437
  (
    n3327,
    n388,
    n2115,
    n2696,
    n2862
  );


  and
  g3438
  (
    n3172,
    n2889,
    n2886,
    n2862,
    n213
  );


  nand
  g3439
  (
    n3402,
    n2557,
    n2927,
    n1998,
    n2576
  );


  or
  g3440
  (
    n3389,
    n2562,
    n2696,
    n412,
    n2345
  );


  or
  g3441
  (
    n3122,
    n368,
    n2953,
    n470,
    n320
  );


  nor
  g3442
  (
    n3413,
    n491,
    n394,
    n2886,
    n2892
  );


  nand
  g3443
  (
    n3182,
    n370,
    n482,
    n2942,
    n393
  );


  xnor
  g3444
  (
    n3129,
    n254,
    n2861,
    n2931,
    n229
  );


  xnor
  g3445
  (
    n3357,
    n449,
    n227,
    n2268,
    n218
  );


  nand
  g3446
  (
    n3392,
    n266,
    n293,
    n2062,
    n2975
  );


  xnor
  g3447
  (
    n3547,
    n326,
    n362,
    n334,
    n356
  );


  and
  g3448
  (
    n3556,
    n2362,
    n435,
    n2924,
    n2336
  );


  xnor
  g3449
  (
    n3190,
    n291,
    n2252,
    n2634,
    n317
  );


  nor
  g3450
  (
    n3034,
    n2152,
    n2946,
    n2842,
    n271
  );


  nand
  g3451
  (
    n3303,
    n345,
    n2666,
    n420,
    n410
  );


  nor
  g3452
  (
    n3531,
    n2327,
    n369,
    n383,
    n2411
  );


  xor
  g3453
  (
    n3337,
    n457,
    n2949,
    n294,
    n219
  );


  or
  g3454
  (
    n3301,
    n2328,
    n2845,
    n236,
    n405
  );


  nand
  g3455
  (
    n3424,
    n271,
    n365,
    n2536,
    n2364
  );


  nor
  g3456
  (
    n3210,
    n2918,
    n217,
    n344,
    n2916
  );


  nor
  g3457
  (
    n3599,
    n2697,
    n303,
    n2977,
    n2918
  );


  xor
  g3458
  (
    n3496,
    n2863,
    n2989,
    n432,
    n2144
  );


  xor
  g3459
  (
    n3090,
    n2164,
    n2670,
    n386,
    n225
  );


  xnor
  g3460
  (
    n3488,
    n2851,
    n2210,
    n240,
    n2838
  );


  xor
  g3461
  (
    n3116,
    n2403,
    n2701,
    n2569,
    n2300
  );


  xor
  g3462
  (
    n3071,
    n414,
    n416,
    n495,
    n2575
  );


  and
  g3463
  (
    n3283,
    n493,
    n2860,
    n2089,
    n2374
  );


  xnor
  g3464
  (
    n3526,
    n2429,
    n2434,
    n2668,
    n2944
  );


  and
  g3465
  (
    n3613,
    n328,
    n2928,
    n237,
    n479
  );


  and
  g3466
  (
    n3469,
    n418,
    n2922,
    n2930,
    n2948
  );


  nand
  g3467
  (
    n3368,
    n2952,
    n2478,
    n487,
    n2932
  );


  xor
  g3468
  (
    n3229,
    n223,
    n478,
    n2208,
    n2884
  );


  xor
  g3469
  (
    n3449,
    n2009,
    n2862,
    n461,
    n2858
  );


  nor
  g3470
  (
    n3329,
    n2641,
    n2163,
    n2707,
    n484
  );


  nand
  g3471
  (
    n3501,
    n2436,
    n2492,
    n279,
    n2928
  );


  xnor
  g3472
  (
    n3570,
    n2697,
    n2971,
    n2180,
    n2848
  );


  xor
  g3473
  (
    n3131,
    n235,
    n2710,
    n284,
    n356
  );


  xor
  g3474
  (
    n3385,
    n450,
    n311,
    n408,
    n2628
  );


  nor
  g3475
  (
    n3394,
    n246,
    n2286,
    n2456,
    n402
  );


  nand
  g3476
  (
    n3505,
    n413,
    n366,
    n2131,
    n2435
  );


  nor
  g3477
  (
    n3010,
    n2698,
    n322,
    n336,
    n460
  );


  xor
  g3478
  (
    n3485,
    n2351,
    n234,
    n2396,
    n496
  );


  and
  g3479
  (
    n3052,
    n396,
    n2276,
    n2462,
    n2713
  );


  nor
  g3480
  (
    n3016,
    n252,
    n458,
    n2885,
    n267
  );


  or
  g3481
  (
    n3333,
    n2341,
    n377,
    n347,
    n2600
  );


  xor
  g3482
  (
    n3474,
    n253,
    n1994,
    n2592,
    n332
  );


  or
  g3483
  (
    n3087,
    n217,
    n2919,
    n2986,
    n419
  );


  or
  g3484
  (
    n3480,
    n349,
    n353,
    n299,
    n2241
  );


  or
  g3485
  (
    n3625,
    n344,
    n2055,
    n2385,
    n358
  );


  nand
  g3486
  (
    n3222,
    n448,
    n2285,
    n2856,
    n2024
  );


  nand
  g3487
  (
    n3582,
    n2388,
    n2844,
    n492,
    n264
  );


  xnor
  g3488
  (
    n3407,
    n2331,
    n447,
    n2317,
    n2977
  );


  xnor
  g3489
  (
    n3126,
    n463,
    n2082,
    n2191,
    n261
  );


  and
  g3490
  (
    n3040,
    n477,
    n438,
    n365,
    n2551
  );


  xnor
  g3491
  (
    n3514,
    n220,
    n441,
    n2698,
    n230
  );


  xnor
  g3492
  (
    n2996,
    n2409,
    n2710,
    n2930,
    n2894
  );


  and
  g3493
  (
    n3188,
    n2422,
    n449,
    n2920,
    n2081
  );


  or
  g3494
  (
    n3319,
    n381,
    n2437,
    n2991,
    n2877
  );


  xnor
  g3495
  (
    n3271,
    n313,
    n2587,
    n2568,
    n422
  );


  nand
  g3496
  (
    n3612,
    n2013,
    n2245,
    n359,
    n245
  );


  nand
  g3497
  (
    n3551,
    n2553,
    n280,
    n403,
    n279
  );


  nor
  g3498
  (
    n3004,
    n2347,
    n366,
    n2980,
    n231
  );


  xnor
  g3499
  (
    n3537,
    n399,
    n2514,
    n2032,
    n455
  );


  nand
  g3500
  (
    n3549,
    n2877,
    n2516,
    n372,
    n2541
  );


  xor
  g3501
  (
    n3031,
    n2911,
    n301,
    n2160,
    n2607
  );


  xnor
  g3502
  (
    n3169,
    n272,
    n2706,
    n233,
    n2686
  );


  or
  g3503
  (
    n3192,
    n492,
    n451,
    n346,
    n2030
  );


  xnor
  g3504
  (
    n3311,
    n435,
    n310,
    n2860,
    n2614
  );


  and
  g3505
  (
    n3557,
    n393,
    n2925,
    n2854,
    n334
  );


  nor
  g3506
  (
    n3439,
    n2161,
    n2938,
    n342,
    n2675
  );


  nand
  g3507
  (
    n3067,
    n2839,
    n2841,
    n2710,
    n304
  );


  nand
  g3508
  (
    n3512,
    n2496,
    n2910,
    n2709,
    n238
  );


  or
  g3509
  (
    n3604,
    n384,
    n302,
    n2377,
    n296
  );


  nand
  g3510
  (
    n3289,
    n270,
    n332,
    n457,
    n2382
  );


  nand
  g3511
  (
    n3088,
    n254,
    n285,
    n2265,
    n2926
  );


  nand
  g3512
  (
    n3070,
    n450,
    n361,
    n2696,
    n416
  );


  nand
  g3513
  (
    n3332,
    n2622,
    n438,
    n374,
    n375
  );


  and
  g3514
  (
    n3489,
    n466,
    n2680,
    n351,
    n2313
  );


  or
  g3515
  (
    n3536,
    n2846,
    n476,
    n2554,
    n431
  );


  nor
  g3516
  (
    n3022,
    n2899,
    n275,
    n437,
    n2837
  );


  xor
  g3517
  (
    n3468,
    n2229,
    n461,
    n2012,
    n2865
  );


  nand
  g3518
  (
    n3338,
    n411,
    n2488,
    n2859,
    n2052
  );


  xnor
  g3519
  (
    n3285,
    n215,
    n2577,
    n2960,
    n294
  );


  or
  g3520
  (
    n3174,
    n2521,
    n2937,
    n383,
    n2966
  );


  xnor
  g3521
  (
    n3542,
    n346,
    n454,
    n352,
    n266
  );


  xor
  g3522
  (
    n3331,
    n470,
    n456,
    n2982,
    n2418
  );


  xnor
  g3523
  (
    n3417,
    n2870,
    n2989,
    n418
  );


  xnor
  g3524
  (
    n3362,
    n416,
    n287,
    n2094,
    n353
  );


  xnor
  g3525
  (
    n3309,
    n2507,
    n445,
    n2158,
    n2993
  );


  and
  g3526
  (
    n3467,
    n2950,
    n483,
    n2897,
    n2861
  );


  and
  g3527
  (
    n3108,
    n2549,
    n2698,
    n2694,
    n423
  );


  nor
  g3528
  (
    n3218,
    n414,
    n2093,
    n402,
    n444
  );


  and
  g3529
  (
    n3587,
    n324,
    n305,
    n2506,
    n2282
  );


  xnor
  g3530
  (
    n3605,
    n312,
    n2136,
    n352,
    n2539
  );


  nor
  g3531
  (
    n3506,
    n291,
    n453,
    n327,
    n337
  );


  and
  g3532
  (
    n3569,
    n228,
    n371,
    n355,
    n238
  );


  nor
  g3533
  (
    n3341,
    n2688,
    n442,
    n396,
    n2153
  );


  xnor
  g3534
  (
    n3154,
    n463,
    n2863,
    n2571,
    n2991
  );


  nor
  g3535
  (
    n3495,
    n2650,
    n2940,
    n2438,
    n361
  );


  nand
  g3536
  (
    n3157,
    n2859,
    n244,
    n218,
    n2461
  );


  nor
  g3537
  (
    n3562,
    n2954,
    n348,
    n2509,
    n256
  );


  xnor
  g3538
  (
    n3078,
    n2440,
    n2896,
    n316,
    n344
  );


  xnor
  g3539
  (
    n3081,
    n2051,
    n355,
    n2176,
    n2695
  );


  xor
  g3540
  (
    n2995,
    n2477,
    n409,
    n258,
    n318
  );


  nand
  g3541
  (
    n3627,
    n2938,
    n2961,
    n287,
    n2651
  );


  xor
  g3542
  (
    n3048,
    n368,
    n2540,
    n249,
    n439
  );


  xnor
  g3543
  (
    n3532,
    n2919,
    n2918,
    n299,
    n2846
  );


  xnor
  g3544
  (
    n3241,
    n442,
    n446,
    n216,
    n2986
  );


  xor
  g3545
  (
    n3429,
    n269,
    n429,
    n2840,
    n2872
  );


  and
  g3546
  (
    n3511,
    n447,
    n2593,
    n230,
    n356
  );


  and
  g3547
  (
    n3151,
    n2025,
    n2114,
    n2224,
    n2897
  );


  nor
  g3548
  (
    n3410,
    n2266,
    n2618,
    n2619,
    n494
  );


  nand
  g3549
  (
    n3263,
    n2558,
    n277,
    n283,
    n2308
  );


  xnor
  g3550
  (
    n3093,
    n244,
    n2982,
    n2893,
    n2947
  );


  and
  g3551
  (
    n3026,
    n392,
    n2432,
    n2391,
    n442
  );


  and
  g3552
  (
    n3464,
    n2309,
    n481,
    n2910,
    n2281
  );


  xnor
  g3553
  (
    n3388,
    n275,
    n2702,
    n2901,
    n2635
  );


  xnor
  g3554
  (
    n3563,
    n471,
    n2320,
    n2312,
    n223
  );


  nand
  g3555
  (
    n3470,
    n424,
    n446,
    n398,
    n2238
  );


  xnor
  g3556
  (
    n3602,
    n2360,
    n2217,
    n2969,
    n2868
  );


  nor
  g3557
  (
    n3554,
    n2381,
    n2909,
    n2848,
    n369
  );


  xnor
  g3558
  (
    n3520,
    n279,
    n436,
    n2903,
    n444
  );


  xnor
  g3559
  (
    n3391,
    n2972,
    n249,
    n2874,
    n370
  );


  xnor
  g3560
  (
    n3615,
    n440,
    n2291,
    n391,
    n298
  );


  xnor
  g3561
  (
    n3336,
    n2876,
    n2182,
    n357,
    n430
  );


  xnor
  g3562
  (
    n3032,
    n2871,
    n444,
    n2852,
    n417
  );


  nor
  g3563
  (
    n3163,
    n476,
    n447,
    n300,
    n2212
  );


  xor
  g3564
  (
    n3632,
    n382,
    n2219,
    n428,
    n2214
  );


  or
  g3565
  (
    n3340,
    n2992,
    n311,
    n362,
    n2060
  );


  nand
  g3566
  (
    n3018,
    n341,
    n2284,
    n336,
    n2264
  );


  xnor
  g3567
  (
    n3119,
    n375,
    n2959,
    n2472,
    n469
  );


  and
  g3568
  (
    n3312,
    n2321,
    n2501,
    n2625,
    n2981
  );


  or
  g3569
  (
    n3432,
    n463,
    n2595,
    n2165,
    n397
  );


  nor
  g3570
  (
    n3548,
    n2522,
    n2966,
    n2851,
    n2702
  );


  xnor
  g3571
  (
    n3445,
    n2708,
    n251,
    n363,
    n2090
  );


  nor
  g3572
  (
    n3103,
    n2674,
    n402,
    n2912,
    n424
  );


  xnor
  g3573
  (
    n3212,
    n258,
    n406,
    n2699,
    n344
  );


  nand
  g3574
  (
    n3355,
    n351,
    n2903,
    n2254,
    n2447
  );


  xor
  g3575
  (
    n3084,
    n432,
    n2339,
    n2108,
    n2709
  );


  nor
  g3576
  (
    n3624,
    n219,
    n2927,
    n412,
    n262
  );


  or
  g3577
  (
    n3525,
    n252,
    n297,
    n2939,
    n436
  );


  nand
  g3578
  (
    n3130,
    n269,
    n2955,
    n2841,
    n261
  );


  nand
  g3579
  (
    n3106,
    n2517,
    n283,
    n2086,
    n367
  );


  nor
  g3580
  (
    n3136,
    n2709,
    n387,
    n2305,
    n427
  );


  nand
  g3581
  (
    n3364,
    n2964,
    n2861,
    n2975,
    n2965
  );


  or
  g3582
  (
    n3504,
    n2848,
    n2640,
    n329,
    n346
  );


  xnor
  g3583
  (
    n3059,
    n2877,
    n2923,
    n2531,
    n288
  );


  xor
  g3584
  (
    n3585,
    n2692,
    n343,
    n2588,
    n428
  );


  or
  g3585
  (
    n3023,
    n351,
    n2001,
    n2960,
    n229
  );


  xor
  g3586
  (
    n3325,
    n260,
    n2867,
    n2979,
    n425
  );


  xnor
  g3587
  (
    n3109,
    n237,
    n2673,
    n2504,
    n489
  );


  nor
  g3588
  (
    n3633,
    n243,
    n2982,
    n227,
    n2146
  );


  nor
  g3589
  (
    n3527,
    n316,
    n2932,
    n311,
    n2711
  );


  and
  g3590
  (
    n3287,
    n2068,
    n2608,
    n2400,
    n2889
  );


  and
  g3591
  (
    n3171,
    n247,
    n2342,
    n315,
    n2981
  );


  nand
  g3592
  (
    n3360,
    n2104,
    n2623,
    n465,
    n2994
  );


  and
  g3593
  (
    n3173,
    n2711,
    n2413,
    n2056,
    n2704
  );


  xor
  g3594
  (
    n3491,
    n329,
    n2559,
    n2894,
    n431
  );


  nand
  g3595
  (
    n3233,
    n2892,
    n2886,
    n2873,
    n302
  );


  or
  g3596
  (
    n3555,
    n2134,
    n464,
    n2652,
    n2912
  );


  and
  g3597
  (
    n3110,
    n243,
    n259,
    n2920,
    n215
  );


  xnor
  g3598
  (
    n3221,
    n2119,
    n2552,
    n2848,
    n2355
  );


  and
  g3599
  (
    n3189,
    n2048,
    n2643,
    n2905,
    n2046
  );


  nand
  g3600
  (
    n3630,
    n306,
    n2143,
    n2681,
    n283
  );


  or
  g3601
  (
    n3517,
    n2890,
    n286,
    n2226,
    n2949
  );


  and
  g3602
  (
    n3700,
    n3504,
    n3545,
    n3304,
    n3592
  );


  nand
  g3603
  (
    n3838,
    n3631,
    n3533,
    n3287,
    n3616
  );


  xnor
  g3604
  (
    n3725,
    n3595,
    n3273,
    n3384,
    n3581
  );


  nand
  g3605
  (
    n3661,
    n3539,
    n3496,
    n3307,
    n3348
  );


  nand
  g3606
  (
    n3754,
    n3181,
    n3156,
    n3589,
    n3554
  );


  xnor
  g3607
  (
    n3641,
    n3337,
    n3600,
    n3532,
    n3548
  );


  nand
  g3608
  (
    n3640,
    n3448,
    n3301,
    n3244,
    n3441
  );


  nor
  g3609
  (
    n3844,
    n3590,
    n3323,
    n3513,
    n3254
  );


  or
  g3610
  (
    n3887,
    n3100,
    n3448,
    n3403,
    n3595
  );


  xnor
  g3611
  (
    n3884,
    n3552,
    n3556,
    n3192,
    n3432
  );


  nor
  g3612
  (
    n3852,
    n3071,
    n3233,
    n3370,
    n3013
  );


  nor
  g3613
  (
    n3660,
    n3597,
    n3351,
    n3618,
    n3385
  );


  xnor
  g3614
  (
    n3836,
    n3487,
    n3527,
    n3081,
    n3247
  );


  and
  g3615
  (
    n3752,
    n3486,
    n3526,
    n3535,
    n3214
  );


  xnor
  g3616
  (
    n3780,
    n3604,
    n3550,
    n3073,
    n3317
  );


  nand
  g3617
  (
    n3689,
    n3602,
    n3561,
    n3202,
    n3406
  );


  nand
  g3618
  (
    n3669,
    n3551,
    n3353,
    n3494,
    n3369
  );


  xor
  g3619
  (
    n3761,
    n3608,
    n3266,
    n3514,
    n3321
  );


  or
  g3620
  (
    n3901,
    n3477,
    n3239,
    n3397,
    n3560
  );


  nor
  g3621
  (
    n3924,
    n3597,
    n3185,
    n3278,
    n3428
  );


  nor
  g3622
  (
    n3648,
    n3180,
    n3567,
    n3481,
    n3599
  );


  nand
  g3623
  (
    n3853,
    n3568,
    n3559,
    n3186,
    n3253
  );


  xor
  g3624
  (
    n3849,
    n499,
    n3057,
    n3607,
    n3503
  );


  nor
  g3625
  (
    n3900,
    n3519,
    n3036,
    n3611,
    n3356
  );


  or
  g3626
  (
    n3772,
    n3471,
    n3584,
    n3617,
    n2725
  );


  or
  g3627
  (
    n3724,
    n3620,
    n3497,
    n3425,
    n3246
  );


  nor
  g3628
  (
    n3830,
    n3593,
    n3495,
    n3559,
    n3544
  );


  xor
  g3629
  (
    n3706,
    n3531,
    n3213,
    n498,
    n3024
  );


  or
  g3630
  (
    n3664,
    n3360,
    n3613,
    n3491,
    n3612
  );


  xnor
  g3631
  (
    n3855,
    n3513,
    n3501,
    n3055,
    n3533
  );


  nor
  g3632
  (
    n3825,
    n3328,
    n3578,
    n3506,
    n3618
  );


  nor
  g3633
  (
    n3680,
    n3524,
    n3487,
    n3518,
    n3409
  );


  nand
  g3634
  (
    n3771,
    n3325,
    n3493,
    n3167,
    n3546
  );


  and
  g3635
  (
    n3860,
    n3251,
    n3566,
    n3168,
    n3308
  );


  or
  g3636
  (
    n3883,
    n3441,
    n3068,
    n3303,
    n3079
  );


  nand
  g3637
  (
    n3691,
    n3174,
    n3623,
    n3550,
    n3512
  );


  nor
  g3638
  (
    n3877,
    n3556,
    n3442,
    n3437,
    n3573
  );


  or
  g3639
  (
    n3893,
    n3499,
    n3127,
    n3596,
    n3241
  );


  nand
  g3640
  (
    n3718,
    n3572,
    n3454,
    n3188,
    n3087
  );


  nand
  g3641
  (
    n3801,
    n3505,
    n3484,
    n3481,
    n3533
  );


  xnor
  g3642
  (
    n3815,
    n3524,
    n3570,
    n499,
    n3416
  );


  or
  g3643
  (
    n3828,
    n3632,
    n3059,
    n3105,
    n3436
  );


  nand
  g3644
  (
    n3760,
    n3231,
    n3103,
    n3634,
    n3283
  );


  nor
  g3645
  (
    n3834,
    n3494,
    n3495,
    n3234,
    n3530
  );


  nor
  g3646
  (
    n3927,
    n3506,
    n3512,
    n3630,
    n3064
  );


  nand
  g3647
  (
    n3788,
    n3533,
    n3104,
    n3596,
    n3135
  );


  and
  g3648
  (
    n3842,
    n3600,
    n3607,
    n3112,
    n3579
  );


  nand
  g3649
  (
    n3779,
    n3470,
    n3452,
    n3143,
    n3534
  );


  or
  g3650
  (
    n3687,
    n3200,
    n3621,
    n3487,
    n3570
  );


  xnor
  g3651
  (
    n3802,
    n3620,
    n3151,
    n3207,
    n3561
  );


  and
  g3652
  (
    n3890,
    n3074,
    n3377,
    n3540,
    n3561
  );


  or
  g3653
  (
    n3917,
    n3524,
    n3612,
    n3459,
    n3493
  );


  xnor
  g3654
  (
    n3821,
    n3183,
    n3521,
    n3612,
    n3224
  );


  or
  g3655
  (
    n3919,
    n3368,
    n3530,
    n3131,
    n3593
  );


  xor
  g3656
  (
    n3733,
    n3601,
    n3532,
    n3507,
    n3511
  );


  xor
  g3657
  (
    n3719,
    n3623,
    n3400,
    n3553,
    n3514
  );


  nand
  g3658
  (
    n3750,
    n3169,
    n3222,
    n3550,
    n3228
  );


  xor
  g3659
  (
    n3866,
    n3172,
    n3113,
    n3451,
    n3420
  );


  nor
  g3660
  (
    n3829,
    n3208,
    n3086,
    n3257,
    n3628
  );


  and
  g3661
  (
    n3874,
    n3538,
    n3426,
    n3373,
    n3025
  );


  and
  g3662
  (
    n3695,
    n3330,
    n3586,
    n3392,
    n3474
  );


  xnor
  g3663
  (
    n3932,
    n3542,
    n3314,
    n3546,
    n3510
  );


  nand
  g3664
  (
    n3651,
    n3277,
    n3509,
    n3033,
    n3413
  );


  nor
  g3665
  (
    n3694,
    n3546,
    n3285,
    n3477,
    n3608
  );


  and
  g3666
  (
    n3770,
    n3475,
    n3453,
    n3210,
    n3529
  );


  xnor
  g3667
  (
    n3746,
    n3219,
    n3245,
    n3609,
    n3503
  );


  xor
  g3668
  (
    n3872,
    n3342,
    n3572,
    n3489,
    n3440
  );


  and
  g3669
  (
    n3848,
    n3435,
    n3490,
    n3288,
    n3400
  );


  nor
  g3670
  (
    n3753,
    n3227,
    n3621,
    n3211,
    n3155
  );


  nor
  g3671
  (
    n3777,
    n3582,
    n3464,
    n3536,
    n3476
  );


  xor
  g3672
  (
    n3693,
    n3515,
    n3498,
    n3577,
    n3583
  );


  and
  g3673
  (
    n3726,
    n3132,
    n3520,
    n3498,
    n3028
  );


  or
  g3674
  (
    n3644,
    n3556,
    n3054,
    n3479,
    n3361
  );


  nor
  g3675
  (
    n3878,
    n3422,
    n3594,
    n3617,
    n3473
  );


  xor
  g3676
  (
    n3716,
    n3197,
    n3173,
    n3162,
    n3587
  );


  xor
  g3677
  (
    n3937,
    n3030,
    n3555,
    n3518,
    n3548
  );


  nor
  g3678
  (
    n3696,
    n3625,
    n3417,
    n3119,
    n3350
  );


  nor
  g3679
  (
    n3812,
    n3428,
    n3446,
    n3622,
    n3521
  );


  nand
  g3680
  (
    n3858,
    n3223,
    n3261,
    n3102,
    n3196
  );


  nor
  g3681
  (
    n3843,
    n3389,
    n3465,
    n3199,
    n3549
  );


  and
  g3682
  (
    n3906,
    n3443,
    n3098,
    n3620,
    n3165
  );


  or
  g3683
  (
    n3863,
    n3204,
    n3506,
    n3189,
    n3123
  );


  or
  g3684
  (
    n3810,
    n3499,
    n3494,
    n3577,
    n3534
  );


  or
  g3685
  (
    n3663,
    n3522,
    n2997,
    n3497,
    n3633
  );


  xor
  g3686
  (
    n3657,
    n3517,
    n3016,
    n3502,
    n3595
  );


  nor
  g3687
  (
    n3637,
    n3506,
    n3627,
    n3387,
    n3603
  );


  xor
  g3688
  (
    n3923,
    n3095,
    n3596,
    n3535,
    n3009
  );


  nand
  g3689
  (
    n3806,
    n3466,
    n3421,
    n3292,
    n3158
  );


  nand
  g3690
  (
    n3727,
    n3061,
    n3171,
    n3378,
    n3148
  );


  xor
  g3691
  (
    n3921,
    n3570,
    n3129,
    n3598,
    n3339
  );


  and
  g3692
  (
    n3655,
    n3495,
    n3053,
    n3601,
    n3121
  );


  and
  g3693
  (
    n3676,
    n3324,
    n3271,
    n3632,
    n3109
  );


  or
  g3694
  (
    n3915,
    n3332,
    n3456,
    n3541,
    n3116
  );


  nand
  g3695
  (
    n3930,
    n3610,
    n3606,
    n3355,
    n3581
  );


  nor
  g3696
  (
    n3736,
    n3599,
    n3110,
    n3576,
    n3489
  );


  or
  g3697
  (
    n3811,
    n3396,
    n3575,
    n3367,
    n3482
  );


  nand
  g3698
  (
    n3672,
    n3382,
    n3042,
    n3407,
    n3629
  );


  xor
  g3699
  (
    n3814,
    n3589,
    n3259,
    n3516,
    n3255
  );


  xor
  g3700
  (
    n3894,
    n2995,
    n3620,
    n3407,
    n3510
  );


  xor
  g3701
  (
    n3831,
    n3240,
    n3478,
    n3547,
    n3150
  );


  nand
  g3702
  (
    n3854,
    n3503,
    n3320,
    n3500,
    n3616
  );


  xor
  g3703
  (
    n3650,
    n3225,
    n3405,
    n3563,
    n3451
  );


  nand
  g3704
  (
    n3645,
    n3076,
    n3576,
    n3594,
    n3578
  );


  xor
  g3705
  (
    n3839,
    n3310,
    n3037,
    n3468,
    n3592
  );


  nand
  g3706
  (
    n3820,
    n3563,
    n3187,
    n3139,
    n3275
  );


  xnor
  g3707
  (
    n3705,
    n3358,
    n3221,
    n3464,
    n3438
  );


  xnor
  g3708
  (
    n3671,
    n3579,
    n3516,
    n3379,
    n3004
  );


  and
  g3709
  (
    n3833,
    n3408,
    n3521,
    n3366,
    n2998
  );


  or
  g3710
  (
    n3850,
    n3491,
    n3483,
    n3066,
    n3531
  );


  nor
  g3711
  (
    n3767,
    n3509,
    n3466,
    n3412,
    n3614
  );


  xnor
  g3712
  (
    n3816,
    n3284,
    n3418,
    n3164,
    n3546
  );


  xnor
  g3713
  (
    n3666,
    n3437,
    n3040,
    n3423,
    n3542
  );


  or
  g3714
  (
    n3879,
    n3576,
    n3545,
    n3035,
    n3478
  );


  and
  g3715
  (
    n3713,
    n3454,
    n3590,
    n3545,
    n3599
  );


  or
  g3716
  (
    n3766,
    n3409,
    n3487,
    n3163,
    n3463
  );


  nor
  g3717
  (
    n3668,
    n3041,
    n3039,
    n3526,
    n3497
  );


  and
  g3718
  (
    n3667,
    n3630,
    n3557,
    n3514,
    n3563
  );


  nor
  g3719
  (
    n3659,
    n3146,
    n3209,
    n3499,
    n3588
  );


  and
  g3720
  (
    n3907,
    n3508,
    n3302,
    n3631,
    n3352
  );


  xnor
  g3721
  (
    n3837,
    n3329,
    n3482,
    n3619,
    n3319
  );


  nand
  g3722
  (
    n3649,
    n3582,
    n3453,
    n3562,
    n3125
  );


  and
  g3723
  (
    n3643,
    n3590,
    n3427,
    n3522,
    n3520
  );


  or
  g3724
  (
    n3933,
    n3621,
    n3230,
    n3517,
    n3572
  );


  xor
  g3725
  (
    n3789,
    n3492,
    n3152,
    n3047,
    n3048
  );


  or
  g3726
  (
    n3805,
    n3458,
    n3580,
    n3134,
    n3364
  );


  nor
  g3727
  (
    n3679,
    n3628,
    n3500,
    n3516,
    n3607
  );


  nand
  g3728
  (
    n3795,
    n3263,
    n3517,
    n3235,
    n3443
  );


  or
  g3729
  (
    n3774,
    n3488,
    n3179,
    n3540,
    n3282
  );


  and
  g3730
  (
    n3797,
    n3408,
    n3490,
    n3614,
    n3549
  );


  xnor
  g3731
  (
    n3936,
    n3608,
    n3267,
    n3594,
    n3473
  );


  nor
  g3732
  (
    n3749,
    n3498,
    n3415,
    n3530,
    n3607
  );


  nor
  g3733
  (
    n3721,
    n3606,
    n3510,
    n3015,
    n2728
  );


  nor
  g3734
  (
    n3870,
    n3161,
    n3496,
    n3544,
    n3566
  );


  and
  g3735
  (
    n3756,
    n3170,
    n3294,
    n3333,
    n3518
  );


  and
  g3736
  (
    n3867,
    n3540,
    n3106,
    n3077,
    n3538
  );


  xor
  g3737
  (
    n3840,
    n3010,
    n3504,
    n3512,
    n3524
  );


  or
  g3738
  (
    n3819,
    n3560,
    n3615,
    n3584,
    n3606
  );


  xnor
  g3739
  (
    n3677,
    n3569,
    n3433,
    n3523,
    n3336
  );


  nand
  g3740
  (
    n3683,
    n3434,
    n3138,
    n3396,
    n3058
  );


  or
  g3741
  (
    n3684,
    n3511,
    n3029,
    n3584,
    n3565
  );


  nor
  g3742
  (
    n3757,
    n3398,
    n3019,
    n3394,
    n3477
  );


  nand
  g3743
  (
    n3741,
    n3562,
    n3525,
    n3427,
    n3531
  );


  and
  g3744
  (
    n3675,
    n498,
    n3327,
    n3479,
    n3440
  );


  or
  g3745
  (
    n3928,
    n3096,
    n3527,
    n3528,
    n3060
  );


  or
  g3746
  (
    n3781,
    n3450,
    n3141,
    n3519,
    n3627
  );


  nand
  g3747
  (
    n3856,
    n3532,
    n3520,
    n3515,
    n3507
  );


  and
  g3748
  (
    n3709,
    n3435,
    n3588,
    n3605,
    n3406
  );


  and
  g3749
  (
    n3737,
    n3574,
    n3218,
    n3547,
    n3564
  );


  nand
  g3750
  (
    n3886,
    n3537,
    n3611,
    n3031,
    n3346
  );


  xnor
  g3751
  (
    n3846,
    n3335,
    n3562,
    n3626,
    n3137
  );


  and
  g3752
  (
    n3739,
    n3462,
    n3529,
    n3600,
    n3553
  );


  or
  g3753
  (
    n3763,
    n3474,
    n3589,
    n3588,
    n3517
  );


  and
  g3754
  (
    n3796,
    n3272,
    n3411,
    n3515,
    n3585
  );


  and
  g3755
  (
    n3732,
    n3515,
    n3215,
    n3475,
    n3313
  );


  nand
  g3756
  (
    n3818,
    n3601,
    n3007,
    n3502,
    n3554
  );


  or
  g3757
  (
    n3734,
    n3625,
    n3126,
    n3547,
    n3479
  );


  and
  g3758
  (
    n3824,
    n3295,
    n3633,
    n3472,
    n3421
  );


  or
  g3759
  (
    n3686,
    n3484,
    n3488,
    n3338,
    n3566
  );


  nor
  g3760
  (
    n3782,
    n3590,
    n3001,
    n3536,
    n3615
  );


  nand
  g3761
  (
    n3873,
    n3264,
    n3120,
    n3232,
    n3386
  );


  or
  g3762
  (
    n3835,
    n3564,
    n3518,
    n3470,
    n3569
  );


  nand
  g3763
  (
    n3861,
    n498,
    n3628,
    n3498,
    n3492
  );


  and
  g3764
  (
    n3800,
    n3270,
    n3489,
    n3449,
    n3593
  );


  nand
  g3765
  (
    n3759,
    n3322,
    n3051,
    n3613,
    n3585
  );


  or
  g3766
  (
    n3722,
    n3122,
    n3497,
    n3501,
    n3402
  );


  xnor
  g3767
  (
    n3914,
    n3505,
    n3571,
    n3551,
    n3044
  );


  nand
  g3768
  (
    n3712,
    n499,
    n3554,
    n3492,
    n3229
  );


  xor
  g3769
  (
    n3707,
    n3595,
    n3565,
    n3416,
    n3099
  );


  nand
  g3770
  (
    n3784,
    n3575,
    n3147,
    n3523,
    n3447
  );


  xor
  g3771
  (
    n3783,
    n3483,
    n3080,
    n3444,
    n3291
  );


  nor
  g3772
  (
    n3794,
    n3374,
    n3262,
    n3012,
    n3594
  );


  nor
  g3773
  (
    n3717,
    n3268,
    n3456,
    n3558,
    n3598
  );


  or
  g3774
  (
    n3896,
    n3388,
    n3115,
    n3543,
    n3043
  );


  nand
  g3775
  (
    n3787,
    n3340,
    n3536,
    n3078,
    n3510
  );


  nand
  g3776
  (
    n3768,
    n3534,
    n3532,
    n3493,
    n3238
  );


  nor
  g3777
  (
    n3808,
    n3331,
    n3509,
    n3166,
    n3359
  );


  nand
  g3778
  (
    n3636,
    n3604,
    n3571,
    n3062,
    n3381
  );


  nor
  g3779
  (
    n3891,
    n3463,
    n3299,
    n3539,
    n3419
  );


  or
  g3780
  (
    n3869,
    n3050,
    n2727,
    n3468,
    n3457
  );


  or
  g3781
  (
    n3875,
    n3046,
    n3519,
    n3559,
    n3375
  );


  and
  g3782
  (
    n3888,
    n3496,
    n3571,
    n3417,
    n3501
  );


  or
  g3783
  (
    n3665,
    n3101,
    n3587,
    n3622,
    n3582
  );


  nand
  g3784
  (
    n3775,
    n3136,
    n3526,
    n2722,
    n3622
  );


  xnor
  g3785
  (
    n3735,
    n3484,
    n3216,
    n3469,
    n3633
  );


  or
  g3786
  (
    n3865,
    n3511,
    n3553,
    n3527,
    n3413
  );


  or
  g3787
  (
    n3925,
    n3606,
    n3391,
    n3508,
    n3422
  );


  or
  g3788
  (
    n3720,
    n3564,
    n3548,
    n3274,
    n3289
  );


  or
  g3789
  (
    n3868,
    n3142,
    n3558,
    n3410,
    n3513
  );


  or
  g3790
  (
    n3785,
    n3536,
    n3624,
    n3312,
    n3542
  );


  nand
  g3791
  (
    n3674,
    n3286,
    n3571,
    n3556,
    n3438
  );


  and
  g3792
  (
    n3807,
    n3618,
    n3111,
    n3555,
    n3535
  );


  nand
  g3793
  (
    n3744,
    n3550,
    n3011,
    n3612,
    n3433
  );


  nor
  g3794
  (
    n3857,
    n3380,
    n3494,
    n3582,
    n3567
  );


  xnor
  g3795
  (
    n3658,
    n3583,
    n3193,
    n3108,
    n3544
  );


  nor
  g3796
  (
    n3685,
    n3591,
    n3525,
    n3578,
    n3430
  );


  and
  g3797
  (
    n3703,
    n3528,
    n3619,
    n3610,
    n3032
  );


  xor
  g3798
  (
    n3692,
    n3557,
    n3538,
    n3618,
    n3585
  );


  or
  g3799
  (
    n3909,
    n3140,
    n3585,
    n3431,
    n3237
  );


  and
  g3800
  (
    n3897,
    n3423,
    n3083,
    n3347,
    n3415
  );


  nor
  g3801
  (
    n3714,
    n3194,
    n3570,
    n3411,
    n3572
  );


  or
  g3802
  (
    n3793,
    n3621,
    n3569,
    n3541,
    n3519
  );


  and
  g3803
  (
    n3698,
    n3243,
    n3602,
    n3471,
    n3090
  );


  xor
  g3804
  (
    n3798,
    n3118,
    n3491,
    n3020,
    n3226
  );


  or
  g3805
  (
    n3799,
    n3467,
    n3474,
    n3006,
    n3555
  );


  and
  g3806
  (
    n3690,
    n3130,
    n3613,
    n3567,
    n3027
  );


  xnor
  g3807
  (
    n3699,
    n3624,
    n3584,
    n3149,
    n3539
  );


  or
  g3808
  (
    n3646,
    n3520,
    n3341,
    n3501,
    n3124
  );


  nor
  g3809
  (
    n3702,
    n3002,
    n3509,
    n3603,
    n3157
  );


  xor
  g3810
  (
    n3769,
    n3442,
    n3507,
    n3575,
    n3480
  );


  xnor
  g3811
  (
    n3895,
    n3488,
    n3560,
    n3569,
    n3424
  );


  nand
  g3812
  (
    n3876,
    n3541,
    n3634,
    n3176,
    n3552
  );


  nand
  g3813
  (
    n3871,
    n3544,
    n3522,
    n3000,
    n3557
  );


  nand
  g3814
  (
    n3889,
    n3567,
    n3523,
    n3034,
    n3450
  );


  xnor
  g3815
  (
    n3728,
    n3481,
    n3298,
    n3260,
    n3601
  );


  xor
  g3816
  (
    n3885,
    n3499,
    n3623,
    n3465,
    n3628
  );


  xnor
  g3817
  (
    n3862,
    n3500,
    n3539,
    n3602,
    n3588
  );


  and
  g3818
  (
    n3790,
    n3092,
    n3613,
    n3486,
    n3085
  );


  xor
  g3819
  (
    n3851,
    n3489,
    n3583,
    n3589,
    n3605
  );


  xor
  g3820
  (
    n3786,
    n3371,
    n3554,
    n3484,
    n3529
  );


  xor
  g3821
  (
    n3704,
    n3005,
    n3383,
    n3398,
    n3178
  );


  xnor
  g3822
  (
    n3656,
    n3564,
    n3508,
    n3545,
    n3557
  );


  and
  g3823
  (
    n3826,
    n3608,
    n3537,
    n3630,
    n3279
  );


  nand
  g3824
  (
    n3653,
    n3300,
    n3290,
    n3587,
    n3581
  );


  or
  g3825
  (
    n3701,
    n2999,
    n3591,
    n3479,
    n3485
  );


  and
  g3826
  (
    n3881,
    n3580,
    n3568,
    n3281,
    n3587
  );


  xor
  g3827
  (
    n3708,
    n3558,
    n3603,
    n3114,
    n3491
  );


  nand
  g3828
  (
    n3710,
    n3446,
    n3551,
    n3558,
    n3619
  );


  or
  g3829
  (
    n3762,
    n3184,
    n3502,
    n3552,
    n3483
  );


  xnor
  g3830
  (
    n3642,
    n3349,
    n3252,
    n3609,
    n3372
  );


  xor
  g3831
  (
    n3755,
    n3611,
    n3568,
    n3038,
    n3297
  );


  nor
  g3832
  (
    n3731,
    n3551,
    n3610,
    n3633,
    n3203
  );


  or
  g3833
  (
    n3911,
    n3249,
    n2726,
    n3082,
    n3439
  );


  nand
  g3834
  (
    n3764,
    n3543,
    n3495,
    n3560,
    n3485
  );


  nor
  g3835
  (
    n3823,
    n3579,
    n3631,
    n3537,
    n3376
  );


  or
  g3836
  (
    n3723,
    n3476,
    n3469,
    n3296,
    n3599
  );


  nand
  g3837
  (
    n3792,
    n3424,
    n3504,
    n3014,
    n3531
  );


  xnor
  g3838
  (
    n3638,
    n3549,
    n3527,
    n3316,
    n3555
  );


  xor
  g3839
  (
    n3905,
    n3426,
    n3344,
    n3436,
    n3552
  );


  nand
  g3840
  (
    n3920,
    n3459,
    n3486,
    n3625,
    n3439
  );


  xor
  g3841
  (
    n3926,
    n3395,
    n3256,
    n3072,
    n3577
  );


  or
  g3842
  (
    n3832,
    n3429,
    n3021,
    n3580,
    n3159
  );


  nand
  g3843
  (
    n3934,
    n3547,
    n3505,
    n3575,
    n3553
  );


  xnor
  g3844
  (
    n3931,
    n3420,
    n3480,
    n3390,
    n3160
  );


  nand
  g3845
  (
    n3912,
    n3414,
    n3632,
    n3343,
    n3088
  );


  nand
  g3846
  (
    n3809,
    n3615,
    n3566,
    n3610,
    n3206
  );


  or
  g3847
  (
    n3813,
    n3485,
    n3627,
    n3528
  );


  nor
  g3848
  (
    n3859,
    n3250,
    n3490,
    n3521,
    n3586
  );


  or
  g3849
  (
    n3822,
    n3596,
    n3574,
    n3493,
    n3052
  );


  xor
  g3850
  (
    n3681,
    n3399,
    n3397,
    n3475,
    n3444
  );


  and
  g3851
  (
    n3899,
    n3403,
    n3107,
    n3175,
    n3619
  );


  xnor
  g3852
  (
    n3803,
    n3128,
    n3634,
    n3410,
    n3089
  );


  and
  g3853
  (
    n3910,
    n3591,
    n3154,
    n3220,
    n3309
  );


  nor
  g3854
  (
    n3635,
    n3631,
    n3445,
    n3075,
    n3432
  );


  nor
  g3855
  (
    n3929,
    n3461,
    n3191,
    n2996,
    n3622
  );


  nor
  g3856
  (
    n3730,
    n3614,
    n3529,
    n3455,
    n3056
  );


  xor
  g3857
  (
    n3904,
    n3492,
    n3363,
    n3565,
    n3429
  );


  nand
  g3858
  (
    n3697,
    n3609,
    n3507,
    n3018,
    n3602
  );


  xor
  g3859
  (
    n3776,
    n3217,
    n3198,
    n2723,
    n3481
  );


  nand
  g3860
  (
    n3748,
    n3093,
    n3212,
    n3530,
    n3583
  );


  xnor
  g3861
  (
    n3758,
    n3534,
    n3617,
    n3485,
    n3452
  );


  xnor
  g3862
  (
    n3715,
    n3404,
    n3586,
    n3461,
    n3460
  );


  nand
  g3863
  (
    n3841,
    n3543,
    n3434,
    n3626,
    n3412
  );


  or
  g3864
  (
    n3740,
    n3593,
    n3097,
    n3500,
    n3445
  );


  nand
  g3865
  (
    n3773,
    n3576,
    n3505,
    n3586,
    n3483
  );


  nor
  g3866
  (
    n3908,
    n3419,
    n3486,
    n3482,
    n3512
  );


  xnor
  g3867
  (
    n3678,
    n3504,
    n3293,
    n3063,
    n3117
  );


  xor
  g3868
  (
    n3662,
    n3626,
    n3045,
    n3627,
    n3458
  );


  or
  g3869
  (
    n3639,
    n2724,
    n3574,
    n3311,
    n3190
  );


  or
  g3870
  (
    n3711,
    n3592,
    n3525,
    n3455,
    n3091
  );


  xor
  g3871
  (
    n3688,
    n3488,
    n498,
    n3357,
    n3023
  );


  nand
  g3872
  (
    n3845,
    n3537,
    n3615,
    n3182,
    n3431
  );


  or
  g3873
  (
    n3922,
    n3543,
    n3145,
    n3548,
    n3144
  );


  xnor
  g3874
  (
    n3791,
    n3305,
    n3503,
    n3482,
    n3449
  );


  or
  g3875
  (
    n3738,
    n3605,
    n3473,
    n3604,
    n3563
  );


  xnor
  g3876
  (
    n3817,
    n3559,
    n3447,
    n3609,
    n3540
  );


  nand
  g3877
  (
    n3882,
    n3542,
    n3511,
    n3280,
    n3568
  );


  and
  g3878
  (
    n3898,
    n3549,
    n3393,
    n3632,
    n3265
  );


  and
  g3879
  (
    n3804,
    n3565,
    n3414,
    n3513,
    n3315
  );


  xnor
  g3880
  (
    n3743,
    n3094,
    n3573,
    n3629,
    n3133
  );


  or
  g3881
  (
    n3673,
    n3626,
    n3490,
    n3153,
    n3597
  );


  and
  g3882
  (
    n3903,
    n3269,
    n3508,
    n3069,
    n3616
  );


  and
  g3883
  (
    n3745,
    n3462,
    n3629,
    n3580,
    n3022
  );


  or
  g3884
  (
    n3751,
    n3017,
    n3201,
    n3236,
    n3354
  );


  xnor
  g3885
  (
    n3654,
    n3541,
    n3195,
    n3318,
    n3334
  );


  or
  g3886
  (
    n3647,
    n3405,
    n3616,
    n3526,
    n3523
  );


  xnor
  g3887
  (
    n3918,
    n3573,
    n3561,
    n3401,
    n3525
  );


  xnor
  g3888
  (
    n3778,
    n3579,
    n3276,
    n3502,
    n3478
  );


  nor
  g3889
  (
    n3902,
    n3604,
    n3003,
    n3248,
    n3472
  );


  or
  g3890
  (
    n3916,
    n3467,
    n3457,
    n3430,
    n3401
  );


  or
  g3891
  (
    n3847,
    n3399,
    n3630,
    n3026,
    n3365
  );


  nor
  g3892
  (
    n3765,
    n3404,
    n3538,
    n3578,
    n3597
  );


  xor
  g3893
  (
    n3682,
    n3480,
    n3522,
    n3535,
    n3425
  );


  nand
  g3894
  (
    n3880,
    n3476,
    n3617,
    n3008,
    n3345
  );


  xor
  g3895
  (
    n3827,
    n3603,
    n3496,
    n3362,
    n3402
  );


  and
  g3896
  (
    n3913,
    n3516,
    n3177,
    n3562,
    n3067
  );


  xor
  g3897
  (
    n3935,
    n3634,
    n3258,
    n3306,
    n3611
  );


  or
  g3898
  (
    n3670,
    n3460,
    n3592,
    n3623,
    n3624
  );


  xnor
  g3899
  (
    n3747,
    n3573,
    n3326,
    n3629,
    n3242
  );


  xor
  g3900
  (
    n3742,
    n3395,
    n3598,
    n3574,
    n3480
  );


  and
  g3901
  (
    n3729,
    n3591,
    n3418,
    n3600,
    n3605
  );


  and
  g3902
  (
    n3864,
    n3514,
    n3625,
    n3598,
    n3205
  );


  xor
  g3903
  (
    n3652,
    n3624,
    n3070,
    n3084,
    n3581
  );


  nand
  g3904
  (
    n3892,
    n3614,
    n3577,
    n3049,
    n3065
  );


  xnor
  g3905
  (
    n3984,
    n3813,
    n3852,
    n3663,
    n3773
  );


  or
  g3906
  (
    n3996,
    n3658,
    n3786,
    n3661,
    n3859
  );


  nor
  g3907
  (
    n3959,
    n3882,
    n3841,
    n3722,
    n3640
  );


  xor
  g3908
  (
    n3945,
    n3835,
    n3937,
    n3920,
    n3917
  );


  and
  g3909
  (
    n3970,
    n3654,
    n3667,
    n3862,
    n3838
  );


  or
  g3910
  (
    n3995,
    n3639,
    n3879,
    n3724,
    n3816
  );


  xor
  g3911
  (
    n3968,
    n3704,
    n3686,
    n3888,
    n3766
  );


  xor
  g3912
  (
    n3981,
    n3779,
    n3695,
    n3914,
    n3702
  );


  xnor
  g3913
  (
    n3973,
    n3815,
    n3865,
    n3897,
    n3713
  );


  and
  g3914
  (
    n3993,
    n3928,
    n3818,
    n3844,
    n3669
  );


  xor
  g3915
  (
    n3999,
    n3714,
    n3926,
    n3925,
    n3774
  );


  and
  g3916
  (
    n3942,
    n3834,
    n3740,
    n3636,
    n3902
  );


  nand
  g3917
  (
    n4004,
    n3797,
    n3670,
    n3689,
    n3730
  );


  xnor
  g3918
  (
    n3956,
    n3697,
    n3923,
    n3848,
    n3727
  );


  and
  g3919
  (
    n4000,
    n3668,
    n3742,
    n3770,
    n3906
  );


  xnor
  g3920
  (
    n3980,
    n3802,
    n3645,
    n3653,
    n3791
  );


  xor
  g3921
  (
    n4009,
    n3664,
    n3768,
    n3655,
    n3771
  );


  nand
  g3922
  (
    n3960,
    n3728,
    n3849,
    n3646,
    n3806
  );


  nor
  g3923
  (
    n3997,
    n3693,
    n3784,
    n3638,
    n3832
  );


  xnor
  g3924
  (
    n4007,
    n3793,
    n3935,
    n3691,
    n3800
  );


  nand
  g3925
  (
    n4001,
    n3873,
    n3796,
    n3681,
    n3703
  );


  nand
  g3926
  (
    n3947,
    n3680,
    n3687,
    n3885,
    n3764
  );


  nand
  g3927
  (
    n3976,
    n3843,
    n3666,
    n3899,
    n3783
  );


  nor
  g3928
  (
    n3990,
    n3876,
    n3828,
    n3720,
    n3812
  );


  nand
  g3929
  (
    n3946,
    n3734,
    n3694,
    n3860,
    n3708
  );


  nand
  g3930
  (
    n3986,
    n3787,
    n3679,
    n3912,
    n3830
  );


  or
  g3931
  (
    n3969,
    n3649,
    n3840,
    n3878,
    n3851
  );


  or
  g3932
  (
    n3983,
    n3678,
    n3706,
    n3934,
    n3656
  );


  and
  g3933
  (
    n3948,
    n3725,
    n3785,
    n3842,
    n3652
  );


  or
  g3934
  (
    n4006,
    n3880,
    n3677,
    n3753,
    n3765
  );


  xor
  g3935
  (
    n3998,
    n3814,
    n3748,
    n3836,
    n3870
  );


  and
  g3936
  (
    n3978,
    n3877,
    n3671,
    n3754,
    n3886
  );


  or
  g3937
  (
    n3940,
    n3905,
    n3891,
    n3864,
    n3858
  );


  nor
  g3938
  (
    n3963,
    n3745,
    n3867,
    n3769,
    n3821
  );


  xnor
  g3939
  (
    n3975,
    n3744,
    n3642,
    n3637,
    n3854
  );


  nand
  g3940
  (
    n3989,
    n3718,
    n3732,
    n3712,
    n3736
  );


  and
  g3941
  (
    n3951,
    n3916,
    n3807,
    n3889,
    n3756
  );


  xnor
  g3942
  (
    n3954,
    n3875,
    n3837,
    n3665,
    n3698
  );


  xnor
  g3943
  (
    n3961,
    n3781,
    n3651,
    n3696,
    n3672
  );


  xnor
  g3944
  (
    n3985,
    n3823,
    n3777,
    n499,
    n3760
  );


  and
  g3945
  (
    n3938,
    n3635,
    n3794,
    n3909,
    n3673
  );


  nor
  g3946
  (
    n3988,
    n3790,
    n3798,
    n3690,
    n3801
  );


  or
  g3947
  (
    n4003,
    n3758,
    n3692,
    n3737,
    n3921
  );


  and
  g3948
  (
    n3958,
    n3767,
    n3741,
    n3685,
    n3789
  );


  nor
  g3949
  (
    n4011,
    n3927,
    n3780,
    n3911,
    n3644
  );


  nor
  g3950
  (
    n3987,
    n3782,
    n3641,
    n3743,
    n3811
  );


  nor
  g3951
  (
    n3977,
    n3874,
    n3857,
    n3822,
    n3660
  );


  nor
  g3952
  (
    n3952,
    n3831,
    n3824,
    n3898,
    n3869
  );


  xnor
  g3953
  (
    n4005,
    n3717,
    n3825,
    n3775,
    n3861
  );


  or
  g3954
  (
    n3939,
    n3751,
    n3839,
    n3868,
    n3759
  );


  or
  g3955
  (
    n3991,
    n3711,
    n3804,
    n3731,
    n3762
  );


  nand
  g3956
  (
    n3966,
    n3729,
    n3772,
    n3715,
    n3872
  );


  xnor
  g3957
  (
    n3971,
    n3688,
    n3919,
    n3719,
    n3845
  );


  or
  g3958
  (
    n3962,
    n3819,
    n3805,
    n3659,
    n3795
  );


  xor
  g3959
  (
    n3943,
    n3750,
    n3846,
    n3932,
    n3827
  );


  nand
  g3960
  (
    n3964,
    n3710,
    n3908,
    n3735,
    n3709
  );


  xor
  g3961
  (
    n3974,
    n3778,
    n3643,
    n3915,
    n3931
  );


  xor
  g3962
  (
    n3953,
    n3896,
    n3829,
    n3817,
    n3674
  );


  xnor
  g3963
  (
    n4002,
    n3648,
    n3810,
    n3763,
    n3657
  );


  or
  g3964
  (
    n3994,
    n3833,
    n3746,
    n3647,
    n3929
  );


  or
  g3965
  (
    n3950,
    n3707,
    n3676,
    n3683,
    n3881
  );


  nand
  g3966
  (
    n3967,
    n3894,
    n3799,
    n3792,
    n3682
  );


  xnor
  g3967
  (
    n4010,
    n3757,
    n3863,
    n3705,
    n3884
  );


  xor
  g3968
  (
    n3979,
    n3887,
    n3721,
    n3856,
    n3776
  );


  nand
  g3969
  (
    n3957,
    n3871,
    n3904,
    n3895,
    n3903
  );


  xnor
  g3970
  (
    n4008,
    n3913,
    n3820,
    n3936,
    n3933
  );


  or
  g3971
  (
    n3965,
    n3699,
    n3701,
    n3922,
    n3738
  );


  and
  g3972
  (
    n3944,
    n3918,
    n3866,
    n3910,
    n3892
  );


  xnor
  g3973
  (
    n3949,
    n3749,
    n3924,
    n3803,
    n3733
  );


  and
  g3974
  (
    n4012,
    n3893,
    n3752,
    n3808,
    n3662
  );


  xnor
  g3975
  (
    n3941,
    n3853,
    n3723,
    n3700,
    n3901
  );


  and
  g3976
  (
    n3992,
    n3883,
    n3761,
    n3747,
    n3675
  );


  and
  g3977
  (
    n3955,
    n3847,
    n3788,
    n3809,
    n3684
  );


  and
  g3978
  (
    n3982,
    n3726,
    n3855,
    n3900,
    n3826
  );


  and
  g3979
  (
    n3972,
    n3850,
    n3930,
    n3755,
    n3890
  );


  xnor
  g3980
  (
    n4013,
    n3907,
    n3716,
    n3650,
    n3739
  );


  nand
  g3981
  (
    n4028,
    n3951,
    n3991,
    n4002,
    n3970
  );


  nor
  g3982
  (
    n4017,
    n3952,
    n3971,
    n4005,
    n3994
  );


  and
  g3983
  (
    n4020,
    n3939,
    n3992,
    n3954,
    n3963
  );


  xnor
  g3984
  (
    n4014,
    n3960,
    n3958,
    n3947,
    n3999
  );


  xor
  g3985
  (
    AntiSAT_key_wire,
    n3997,
    n3969,
    n3962,
    n4009
  );


  or
  g3986
  (
    n4016,
    n3959,
    n3979,
    n3946,
    n3938
  );


  nor
  g3987
  (
    n4031,
    n3983,
    n3974,
    n3989,
    n4013
  );


  xor
  g3988
  (
    n4032,
    n3957,
    n3986,
    n3984,
    n3973
  );


  and
  g3989
  (
    n4024,
    n3980,
    n3975,
    n3967,
    n3995
  );


  or
  g3990
  (
    n4026,
    n4004,
    n4003,
    n3978,
    n4008
  );


  xnor
  g3991
  (
    n4022,
    n4001,
    n3956,
    n3950,
    n3998
  );


  xnor
  g3992
  (
    n4029,
    n4007,
    n3977,
    n3988,
    n3945
  );


  xor
  g3993
  (
    n4025,
    n3941,
    n3940,
    n4006,
    n3955
  );


  nor
  g3994
  (
    n4015,
    n3968,
    n3981,
    n4010,
    n4011
  );


  xor
  g3995
  (
    n4021,
    n3948,
    n4012,
    n3972,
    n4000
  );


  or
  g3996
  (
    n4030,
    n3996,
    n3982,
    n3964,
    n3949
  );


  xor
  g3997
  (
    n4023,
    n3943,
    n3990,
    n3987,
    n3953
  );


  nand
  g3998
  (
    n4027,
    n3965,
    n3993,
    n3942,
    n3985
  );


  or
  g3999
  (
    n4019,
    n3976,
    n3966,
    n3961,
    n3944
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n4018,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

