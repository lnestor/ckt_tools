

module Stat_1387_39_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n1312,
  n1320,
  n1383,
  n1417,
  n1414,
  n1411,
  n1415,
  n1410,
  n1407,
  n1405,
  n1408,
  n1418,
  n1413,
  n1412,
  n1409,
  n1406,
  n1416,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1312;output n1320;output n1383;output n1417;output n1414;output n1411;output n1415;output n1410;output n1407;output n1405;output n1408;output n1418;output n1413;output n1412;output n1409;output n1406;output n1416;
  wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n138,
    n22
  );


  not
  g1
  (
    n66,
    n25
  );


  not
  g2
  (
    n104,
    n29
  );


  not
  g3
  (
    n111,
    n20
  );


  not
  g4
  (
    n98,
    n30
  );


  buf
  g5
  (
    n127,
    n31
  );


  buf
  g6
  (
    n88,
    n3
  );


  buf
  g7
  (
    n34,
    n12
  );


  buf
  g8
  (
    n140,
    n16
  );


  not
  g9
  (
    n42,
    n13
  );


  not
  g10
  (
    n96,
    n8
  );


  buf
  g11
  (
    KeyWire_0_10,
    n15
  );


  buf
  g12
  (
    n36,
    n1
  );


  not
  g13
  (
    n117,
    n14
  );


  not
  g14
  (
    n143,
    n4
  );


  buf
  g15
  (
    n99,
    n28
  );


  buf
  g16
  (
    n49,
    n6
  );


  not
  g17
  (
    n62,
    n23
  );


  buf
  g18
  (
    n78,
    n8
  );


  not
  g19
  (
    n68,
    n9
  );


  not
  g20
  (
    n131,
    n28
  );


  not
  g21
  (
    n75,
    n23
  );


  buf
  g22
  (
    n59,
    n21
  );


  buf
  g23
  (
    n112,
    n21
  );


  not
  g24
  (
    n125,
    n25
  );


  buf
  g25
  (
    n60,
    n26
  );


  not
  g26
  (
    n53,
    n10
  );


  not
  g27
  (
    n87,
    n20
  );


  not
  g28
  (
    n126,
    n7
  );


  buf
  g29
  (
    n82,
    n13
  );


  not
  g30
  (
    n50,
    n22
  );


  buf
  g31
  (
    n56,
    n19
  );


  buf
  g32
  (
    n85,
    n25
  );


  buf
  g33
  (
    n100,
    n9
  );


  buf
  g34
  (
    n101,
    n10
  );


  not
  g35
  (
    KeyWire_0_8,
    n3
  );


  not
  g36
  (
    n73,
    n17
  );


  buf
  g37
  (
    n128,
    n17
  );


  buf
  g38
  (
    n40,
    n14
  );


  buf
  g39
  (
    n84,
    n20
  );


  not
  g40
  (
    n48,
    n18
  );


  not
  g41
  (
    n135,
    n30
  );


  not
  g42
  (
    n141,
    n27
  );


  not
  g43
  (
    n77,
    n18
  );


  not
  g44
  (
    n136,
    n29
  );


  not
  g45
  (
    n121,
    n24
  );


  buf
  g46
  (
    n86,
    n5
  );


  buf
  g47
  (
    n145,
    n11
  );


  buf
  g48
  (
    n32,
    n3
  );


  not
  g49
  (
    n124,
    n31
  );


  not
  g50
  (
    n64,
    n23
  );


  buf
  g51
  (
    n132,
    n15
  );


  buf
  g52
  (
    n92,
    n11
  );


  not
  g53
  (
    n146,
    n4
  );


  buf
  g54
  (
    n103,
    n5
  );


  buf
  g55
  (
    n144,
    n30
  );


  not
  g56
  (
    n55,
    n1
  );


  not
  g57
  (
    n44,
    n29
  );


  buf
  g58
  (
    n47,
    n16
  );


  buf
  g59
  (
    n37,
    n27
  );


  buf
  g60
  (
    n150,
    n27
  );


  buf
  g61
  (
    n130,
    n17
  );


  not
  g62
  (
    n97,
    n9
  );


  buf
  g63
  (
    n129,
    n21
  );


  buf
  g64
  (
    n46,
    n26
  );


  not
  g65
  (
    n80,
    n13
  );


  not
  g66
  (
    n39,
    n2
  );


  not
  g67
  (
    n113,
    n19
  );


  buf
  g68
  (
    n133,
    n24
  );


  buf
  g69
  (
    n83,
    n1
  );


  buf
  g70
  (
    n57,
    n16
  );


  not
  g71
  (
    n79,
    n20
  );


  not
  g72
  (
    n148,
    n13
  );


  buf
  g73
  (
    n41,
    n3
  );


  buf
  g74
  (
    n94,
    n22
  );


  not
  g75
  (
    n106,
    n8
  );


  buf
  g76
  (
    n151,
    n7
  );


  buf
  g77
  (
    n115,
    n24
  );


  not
  g78
  (
    n76,
    n8
  );


  not
  g79
  (
    n43,
    n29
  );


  not
  g80
  (
    n38,
    n11
  );


  not
  g81
  (
    n137,
    n6
  );


  not
  g82
  (
    KeyWire_0_23,
    n17
  );


  not
  g83
  (
    n67,
    n10
  );


  buf
  g84
  (
    n45,
    n26
  );


  not
  g85
  (
    n54,
    n12
  );


  buf
  g86
  (
    n61,
    n31
  );


  buf
  g87
  (
    n119,
    n1
  );


  not
  g88
  (
    n102,
    n16
  );


  buf
  g89
  (
    n33,
    n30
  );


  buf
  g90
  (
    n95,
    n6
  );


  buf
  g91
  (
    n71,
    n24
  );


  buf
  g92
  (
    n93,
    n9
  );


  not
  g93
  (
    n153,
    n28
  );


  not
  g94
  (
    n110,
    n26
  );


  not
  g95
  (
    n74,
    n2
  );


  not
  g96
  (
    n35,
    n19
  );


  buf
  g97
  (
    n107,
    n19
  );


  not
  g98
  (
    n108,
    n14
  );


  not
  g99
  (
    n58,
    n22
  );


  not
  g100
  (
    n65,
    n15
  );


  not
  g101
  (
    n152,
    n2
  );


  buf
  g102
  (
    n122,
    n27
  );


  buf
  g103
  (
    n134,
    n7
  );


  not
  g104
  (
    n81,
    n2
  );


  not
  g105
  (
    n139,
    n11
  );


  buf
  g106
  (
    n155,
    n12
  );


  buf
  g107
  (
    n118,
    n31
  );


  not
  g108
  (
    n105,
    n4
  );


  not
  g109
  (
    n72,
    n6
  );


  not
  g110
  (
    n89,
    n18
  );


  not
  g111
  (
    n109,
    n5
  );


  not
  g112
  (
    n142,
    n18
  );


  not
  g113
  (
    n51,
    n14
  );


  not
  g114
  (
    n69,
    n28
  );


  buf
  g115
  (
    n154,
    n21
  );


  buf
  g116
  (
    n70,
    n4
  );


  buf
  g117
  (
    n147,
    n10
  );


  buf
  g118
  (
    n114,
    n7
  );


  buf
  g119
  (
    n116,
    n15
  );


  not
  g120
  (
    n90,
    n23
  );


  buf
  g121
  (
    n149,
    n5
  );


  not
  g122
  (
    n123,
    n12
  );


  buf
  g123
  (
    n91,
    n25
  );


  not
  g124
  (
    n425,
    n127
  );


  not
  g125
  (
    n199,
    n55
  );


  buf
  g126
  (
    n468,
    n38
  );


  not
  g127
  (
    n544,
    n68
  );


  buf
  g128
  (
    n497,
    n120
  );


  buf
  g129
  (
    n554,
    n83
  );


  not
  g130
  (
    n160,
    n82
  );


  not
  g131
  (
    n248,
    n34
  );


  buf
  g132
  (
    n326,
    n53
  );


  not
  g133
  (
    n435,
    n129
  );


  not
  g134
  (
    n266,
    n48
  );


  buf
  g135
  (
    n182,
    n94
  );


  not
  g136
  (
    n181,
    n107
  );


  buf
  g137
  (
    n277,
    n58
  );


  not
  g138
  (
    n189,
    n144
  );


  buf
  g139
  (
    n548,
    n144
  );


  buf
  g140
  (
    n178,
    n112
  );


  not
  g141
  (
    n247,
    n91
  );


  buf
  g142
  (
    n483,
    n38
  );


  not
  g143
  (
    n504,
    n34
  );


  buf
  g144
  (
    n562,
    n100
  );


  not
  g145
  (
    n542,
    n98
  );


  not
  g146
  (
    n180,
    n87
  );


  not
  g147
  (
    n228,
    n43
  );


  buf
  g148
  (
    n158,
    n46
  );


  buf
  g149
  (
    KeyWire_0_2,
    n97
  );


  not
  g150
  (
    n264,
    n52
  );


  buf
  g151
  (
    n231,
    n111
  );


  buf
  g152
  (
    n249,
    n35
  );


  not
  g153
  (
    n455,
    n102
  );


  buf
  g154
  (
    n293,
    n92
  );


  not
  g155
  (
    n357,
    n150
  );


  buf
  g156
  (
    n443,
    n51
  );


  not
  g157
  (
    n531,
    n151
  );


  not
  g158
  (
    n431,
    n108
  );


  not
  g159
  (
    n419,
    n102
  );


  buf
  g160
  (
    n543,
    n110
  );


  buf
  g161
  (
    n423,
    n98
  );


  buf
  g162
  (
    n446,
    n148
  );


  not
  g163
  (
    n209,
    n96
  );


  buf
  g164
  (
    n278,
    n137
  );


  buf
  g165
  (
    n371,
    n125
  );


  buf
  g166
  (
    n445,
    n122
  );


  not
  g167
  (
    n269,
    n64
  );


  buf
  g168
  (
    n167,
    n146
  );


  not
  g169
  (
    n476,
    n50
  );


  buf
  g170
  (
    n241,
    n41
  );


  buf
  g171
  (
    n456,
    n133
  );


  buf
  g172
  (
    n492,
    n69
  );


  buf
  g173
  (
    n349,
    n111
  );


  buf
  g174
  (
    n333,
    n69
  );


  not
  g175
  (
    n294,
    n113
  );


  buf
  g176
  (
    n232,
    n33
  );


  not
  g177
  (
    n533,
    n89
  );


  not
  g178
  (
    n442,
    n88
  );


  not
  g179
  (
    n321,
    n58
  );


  not
  g180
  (
    n496,
    n93
  );


  buf
  g181
  (
    n457,
    n147
  );


  buf
  g182
  (
    n210,
    n88
  );


  not
  g183
  (
    n522,
    n150
  );


  not
  g184
  (
    n283,
    n113
  );


  not
  g185
  (
    n545,
    n122
  );


  buf
  g186
  (
    n304,
    n71
  );


  buf
  g187
  (
    n424,
    n135
  );


  buf
  g188
  (
    n398,
    n77
  );


  not
  g189
  (
    n405,
    n114
  );


  buf
  g190
  (
    n203,
    n82
  );


  buf
  g191
  (
    n342,
    n150
  );


  not
  g192
  (
    n233,
    n130
  );


  buf
  g193
  (
    n460,
    n122
  );


  not
  g194
  (
    n478,
    n72
  );


  not
  g195
  (
    n156,
    n110
  );


  not
  g196
  (
    n380,
    n116
  );


  not
  g197
  (
    n348,
    n60
  );


  not
  g198
  (
    n253,
    n138
  );


  buf
  g199
  (
    n428,
    n63
  );


  not
  g200
  (
    KeyWire_0_30,
    n82
  );


  buf
  g201
  (
    n308,
    n140
  );


  not
  g202
  (
    n271,
    n63
  );


  buf
  g203
  (
    n353,
    n45
  );


  not
  g204
  (
    n316,
    n117
  );


  not
  g205
  (
    n179,
    n96
  );


  not
  g206
  (
    n299,
    n106
  );


  buf
  g207
  (
    n465,
    n38
  );


  not
  g208
  (
    n514,
    n47
  );


  buf
  g209
  (
    n450,
    n145
  );


  buf
  g210
  (
    n565,
    n130
  );


  not
  g211
  (
    n280,
    n146
  );


  buf
  g212
  (
    n307,
    n87
  );


  not
  g213
  (
    n251,
    n33
  );


  not
  g214
  (
    n461,
    n120
  );


  buf
  g215
  (
    n296,
    n42
  );


  not
  g216
  (
    n212,
    n36
  );


  not
  g217
  (
    n257,
    n44
  );


  buf
  g218
  (
    n218,
    n73
  );


  buf
  g219
  (
    n161,
    n42
  );


  buf
  g220
  (
    n555,
    n101
  );


  not
  g221
  (
    n281,
    n68
  );


  not
  g222
  (
    n370,
    n93
  );


  buf
  g223
  (
    n451,
    n33
  );


  buf
  g224
  (
    n394,
    n71
  );


  not
  g225
  (
    n183,
    n95
  );


  not
  g226
  (
    KeyWire_0_7,
    n118
  );


  buf
  g227
  (
    n332,
    n129
  );


  not
  g228
  (
    n235,
    n66
  );


  not
  g229
  (
    n368,
    n136
  );


  not
  g230
  (
    n305,
    n95
  );


  buf
  g231
  (
    n337,
    n84
  );


  not
  g232
  (
    n567,
    n67
  );


  not
  g233
  (
    n384,
    n146
  );


  not
  g234
  (
    n513,
    n116
  );


  buf
  g235
  (
    n426,
    n129
  );


  not
  g236
  (
    n577,
    n119
  );


  buf
  g237
  (
    n201,
    n101
  );


  not
  g238
  (
    n290,
    n89
  );


  buf
  g239
  (
    n434,
    n143
  );


  buf
  g240
  (
    n338,
    n35
  );


  not
  g241
  (
    n340,
    n90
  );


  not
  g242
  (
    n570,
    n43
  );


  buf
  g243
  (
    n331,
    n85
  );


  not
  g244
  (
    n314,
    n125
  );


  buf
  g245
  (
    n523,
    n68
  );


  not
  g246
  (
    n339,
    n71
  );


  buf
  g247
  (
    n335,
    n96
  );


  buf
  g248
  (
    n170,
    n131
  );


  not
  g249
  (
    n355,
    n117
  );


  buf
  g250
  (
    n345,
    n55
  );


  buf
  g251
  (
    n298,
    n121
  );


  not
  g252
  (
    n493,
    n141
  );


  not
  g253
  (
    n444,
    n128
  );


  buf
  g254
  (
    n250,
    n134
  );


  not
  g255
  (
    n206,
    n70
  );


  not
  g256
  (
    n500,
    n136
  );


  buf
  g257
  (
    n459,
    n145
  );


  not
  g258
  (
    n558,
    n149
  );


  buf
  g259
  (
    n323,
    n81
  );


  not
  g260
  (
    KeyWire_0_1,
    n106
  );


  not
  g261
  (
    n529,
    n118
  );


  buf
  g262
  (
    n341,
    n39
  );


  buf
  g263
  (
    n315,
    n92
  );


  not
  g264
  (
    n411,
    n144
  );


  buf
  g265
  (
    n470,
    n144
  );


  buf
  g266
  (
    n226,
    n149
  );


  not
  g267
  (
    n372,
    n101
  );


  not
  g268
  (
    n255,
    n49
  );


  buf
  g269
  (
    n552,
    n86
  );


  not
  g270
  (
    KeyWire_0_26,
    n54
  );


  buf
  g271
  (
    n524,
    n48
  );


  buf
  g272
  (
    n469,
    n41
  );


  buf
  g273
  (
    n288,
    n150
  );


  not
  g274
  (
    n268,
    n43
  );


  buf
  g275
  (
    n192,
    n81
  );


  buf
  g276
  (
    n361,
    n75
  );


  buf
  g277
  (
    n291,
    n99
  );


  not
  g278
  (
    n485,
    n36
  );


  not
  g279
  (
    n408,
    n65
  );


  not
  g280
  (
    n526,
    n42
  );


  not
  g281
  (
    KeyWire_0_17,
    n116
  );


  buf
  g282
  (
    n360,
    n85
  );


  buf
  g283
  (
    n213,
    n138
  );


  buf
  g284
  (
    n187,
    n37
  );


  buf
  g285
  (
    n244,
    n143
  );


  buf
  g286
  (
    n441,
    n124
  );


  buf
  g287
  (
    n193,
    n52
  );


  not
  g288
  (
    n534,
    n45
  );


  buf
  g289
  (
    n162,
    n51
  );


  buf
  g290
  (
    n184,
    n59
  );


  not
  g291
  (
    n303,
    n88
  );


  buf
  g292
  (
    n260,
    n103
  );


  not
  g293
  (
    n310,
    n44
  );


  not
  g294
  (
    n168,
    n107
  );


  buf
  g295
  (
    n172,
    n107
  );


  buf
  g296
  (
    n169,
    n35
  );


  not
  g297
  (
    n207,
    n112
  );


  not
  g298
  (
    n525,
    n57
  );


  not
  g299
  (
    n563,
    n87
  );


  buf
  g300
  (
    n225,
    n53
  );


  not
  g301
  (
    n490,
    n86
  );


  buf
  g302
  (
    n448,
    n127
  );


  not
  g303
  (
    n378,
    n70
  );


  buf
  g304
  (
    n252,
    n95
  );


  buf
  g305
  (
    n575,
    n37
  );


  not
  g306
  (
    n412,
    n151
  );


  not
  g307
  (
    n258,
    n115
  );


  buf
  g308
  (
    n373,
    n115
  );


  not
  g309
  (
    n388,
    n64
  );


  not
  g310
  (
    n363,
    n55
  );


  not
  g311
  (
    n163,
    n33
  );


  not
  g312
  (
    n479,
    n92
  );


  buf
  g313
  (
    n352,
    n130
  );


  buf
  g314
  (
    n275,
    n121
  );


  buf
  g315
  (
    n190,
    n91
  );


  not
  g316
  (
    n322,
    n132
  );


  not
  g317
  (
    n254,
    n119
  );


  not
  g318
  (
    n375,
    n123
  );


  buf
  g319
  (
    n503,
    n146
  );


  not
  g320
  (
    n477,
    n131
  );


  not
  g321
  (
    n417,
    n94
  );


  not
  g322
  (
    n272,
    n104
  );


  buf
  g323
  (
    n312,
    n54
  );


  not
  g324
  (
    n227,
    n133
  );


  buf
  g325
  (
    n392,
    n124
  );


  buf
  g326
  (
    n382,
    n56
  );


  buf
  g327
  (
    KeyWire_0_13,
    n123
  );


  buf
  g328
  (
    n367,
    n137
  );


  buf
  g329
  (
    n462,
    n46
  );


  not
  g330
  (
    n230,
    n80
  );


  not
  g331
  (
    n385,
    n141
  );


  not
  g332
  (
    n389,
    n120
  );


  buf
  g333
  (
    n236,
    n147
  );


  not
  g334
  (
    n471,
    n54
  );


  not
  g335
  (
    n166,
    n73
  );


  buf
  g336
  (
    n377,
    n60
  );


  buf
  g337
  (
    n520,
    n92
  );


  not
  g338
  (
    n211,
    n86
  );


  buf
  g339
  (
    n379,
    n50
  );


  not
  g340
  (
    n222,
    n147
  );


  not
  g341
  (
    n539,
    n99
  );


  buf
  g342
  (
    n505,
    n147
  );


  buf
  g343
  (
    n175,
    n94
  );


  buf
  g344
  (
    n430,
    n137
  );


  not
  g345
  (
    n506,
    n78
  );


  buf
  g346
  (
    n574,
    n126
  );


  buf
  g347
  (
    n157,
    n57
  );


  buf
  g348
  (
    n400,
    n67
  );


  not
  g349
  (
    n383,
    n151
  );


  not
  g350
  (
    n414,
    n72
  );


  buf
  g351
  (
    n559,
    n48
  );


  not
  g352
  (
    n320,
    n143
  );


  not
  g353
  (
    n200,
    n108
  );


  not
  g354
  (
    n437,
    n104
  );


  not
  g355
  (
    n540,
    n125
  );


  not
  g356
  (
    n202,
    n134
  );


  buf
  g357
  (
    n324,
    n148
  );


  buf
  g358
  (
    n495,
    n131
  );


  buf
  g359
  (
    n297,
    n41
  );


  buf
  g360
  (
    n510,
    n70
  );


  buf
  g361
  (
    n214,
    n44
  );


  buf
  g362
  (
    n420,
    n99
  );


  not
  g363
  (
    n220,
    n78
  );


  buf
  g364
  (
    n196,
    n102
  );


  not
  g365
  (
    n501,
    n115
  );


  not
  g366
  (
    n564,
    n99
  );


  not
  g367
  (
    n356,
    n40
  );


  buf
  g368
  (
    KeyWire_0_20,
    n39
  );


  not
  g369
  (
    KeyWire_0_24,
    n62
  );


  buf
  g370
  (
    n240,
    n128
  );


  not
  g371
  (
    n393,
    n65
  );


  buf
  g372
  (
    n334,
    n98
  );


  not
  g373
  (
    n343,
    n139
  );


  buf
  g374
  (
    n215,
    n78
  );


  buf
  g375
  (
    n229,
    n90
  );


  not
  g376
  (
    n482,
    n136
  );


  not
  g377
  (
    n458,
    n68
  );


  not
  g378
  (
    n480,
    n116
  );


  buf
  g379
  (
    n195,
    n81
  );


  buf
  g380
  (
    n481,
    n97
  );


  buf
  g381
  (
    n440,
    n100
  );


  buf
  g382
  (
    n286,
    n59
  );


  buf
  g383
  (
    n306,
    n49
  );


  buf
  g384
  (
    n366,
    n104
  );


  buf
  g385
  (
    n381,
    n108
  );


  buf
  g386
  (
    n511,
    n89
  );


  not
  g387
  (
    n535,
    n76
  );


  buf
  g388
  (
    n487,
    n105
  );


  not
  g389
  (
    n551,
    n101
  );


  buf
  g390
  (
    n566,
    n119
  );


  buf
  g391
  (
    n413,
    n97
  );


  buf
  g392
  (
    n568,
    n75
  );


  buf
  g393
  (
    n573,
    n121
  );


  buf
  g394
  (
    n197,
    n50
  );


  buf
  g395
  (
    n295,
    n94
  );


  not
  g396
  (
    n262,
    n46
  );


  buf
  g397
  (
    n365,
    n66
  );


  buf
  g398
  (
    n376,
    n115
  );


  buf
  g399
  (
    n464,
    n103
  );


  not
  g400
  (
    n289,
    n76
  );


  buf
  g401
  (
    n301,
    n54
  );


  not
  g402
  (
    n403,
    n47
  );


  not
  g403
  (
    n282,
    n113
  );


  not
  g404
  (
    n171,
    n142
  );


  buf
  g405
  (
    n354,
    n60
  );


  buf
  g406
  (
    n387,
    n83
  );


  buf
  g407
  (
    n530,
    n79
  );


  not
  g408
  (
    n317,
    n34
  );


  buf
  g409
  (
    n395,
    n103
  );


  not
  g410
  (
    n473,
    n78
  );


  buf
  g411
  (
    n313,
    n118
  );


  buf
  g412
  (
    n454,
    n87
  );


  not
  g413
  (
    n176,
    n80
  );


  not
  g414
  (
    n547,
    n139
  );


  not
  g415
  (
    n390,
    n45
  );


  buf
  g416
  (
    n261,
    n138
  );


  not
  g417
  (
    n409,
    n128
  );


  not
  g418
  (
    n300,
    n59
  );


  buf
  g419
  (
    n569,
    n74
  );


  not
  g420
  (
    n351,
    n75
  );


  not
  g421
  (
    n410,
    n47
  );


  not
  g422
  (
    n246,
    n49
  );


  buf
  g423
  (
    n242,
    n91
  );


  not
  g424
  (
    n452,
    n93
  );


  buf
  g425
  (
    n494,
    n32
  );


  buf
  g426
  (
    n188,
    n80
  );


  buf
  g427
  (
    n527,
    n126
  );


  buf
  g428
  (
    n362,
    n41
  );


  buf
  g429
  (
    n432,
    n137
  );


  not
  g430
  (
    n406,
    n74
  );


  not
  g431
  (
    n509,
    n110
  );


  buf
  g432
  (
    n475,
    n123
  );


  not
  g433
  (
    n364,
    n109
  );


  buf
  g434
  (
    KeyWire_0_9,
    n91
  );


  not
  g435
  (
    n401,
    n126
  );


  buf
  g436
  (
    n204,
    n148
  );


  buf
  g437
  (
    n499,
    n56
  );


  not
  g438
  (
    n402,
    n110
  );


  not
  g439
  (
    n541,
    n93
  );


  not
  g440
  (
    n359,
    n36
  );


  not
  g441
  (
    n416,
    n66
  );


  buf
  g442
  (
    n263,
    n102
  );


  buf
  g443
  (
    n498,
    n122
  );


  buf
  g444
  (
    n532,
    n140
  );


  buf
  g445
  (
    n234,
    n74
  );


  buf
  g446
  (
    n550,
    n145
  );


  not
  g447
  (
    n256,
    n112
  );


  not
  g448
  (
    n347,
    n105
  );


  buf
  g449
  (
    n274,
    n61
  );


  not
  g450
  (
    n186,
    n32
  );


  not
  g451
  (
    n327,
    n61
  );


  buf
  g452
  (
    n217,
    n148
  );


  buf
  g453
  (
    n546,
    n73
  );


  buf
  g454
  (
    n466,
    n53
  );


  not
  g455
  (
    n418,
    n149
  );


  buf
  g456
  (
    n515,
    n51
  );


  not
  g457
  (
    n336,
    n103
  );


  buf
  g458
  (
    n279,
    n90
  );


  not
  g459
  (
    n285,
    n151
  );


  buf
  g460
  (
    n194,
    n45
  );


  buf
  g461
  (
    n502,
    n64
  );


  buf
  g462
  (
    n284,
    n55
  );


  not
  g463
  (
    n512,
    n140
  );


  not
  g464
  (
    n407,
    n80
  );


  not
  g465
  (
    n521,
    n88
  );


  buf
  g466
  (
    n221,
    n58
  );


  not
  g467
  (
    n318,
    n32
  );


  buf
  g468
  (
    n427,
    n143
  );


  not
  g469
  (
    n404,
    n37
  );


  not
  g470
  (
    n287,
    n57
  );


  buf
  g471
  (
    n557,
    n90
  );


  not
  g472
  (
    n159,
    n139
  );


  not
  g473
  (
    n537,
    n40
  );


  buf
  g474
  (
    n191,
    n79
  );


  not
  g475
  (
    n164,
    n62
  );


  not
  g476
  (
    n549,
    n114
  );


  not
  g477
  (
    KeyWire_0_11,
    n109
  );


  not
  g478
  (
    n223,
    n138
  );


  buf
  g479
  (
    n536,
    n43
  );


  not
  g480
  (
    n238,
    n126
  );


  buf
  g481
  (
    n350,
    n85
  );


  not
  g482
  (
    n576,
    n48
  );


  not
  g483
  (
    n330,
    n111
  );


  not
  g484
  (
    n556,
    n52
  );


  buf
  g485
  (
    n358,
    n63
  );


  not
  g486
  (
    n489,
    n83
  );


  not
  g487
  (
    n369,
    n47
  );


  buf
  g488
  (
    n344,
    n114
  );


  not
  g489
  (
    n174,
    n89
  );


  buf
  g490
  (
    n463,
    n123
  );


  buf
  g491
  (
    n528,
    n109
  );


  buf
  g492
  (
    n518,
    n85
  );


  buf
  g493
  (
    n517,
    n134
  );


  not
  g494
  (
    n216,
    n76
  );


  buf
  g495
  (
    n519,
    n107
  );


  buf
  g496
  (
    n397,
    n39
  );


  buf
  g497
  (
    n173,
    n84
  );


  not
  g498
  (
    n325,
    n98
  );


  not
  g499
  (
    n422,
    n81
  );


  not
  g500
  (
    n453,
    n124
  );


  not
  g501
  (
    n399,
    n106
  );


  not
  g502
  (
    n433,
    n84
  );


  buf
  g503
  (
    n267,
    n59
  );


  buf
  g504
  (
    n270,
    n105
  );


  buf
  g505
  (
    n516,
    n60
  );


  buf
  g506
  (
    KeyWire_0_18,
    n79
  );


  buf
  g507
  (
    n208,
    n141
  );


  buf
  g508
  (
    n319,
    n77
  );


  buf
  g509
  (
    n438,
    n124
  );


  not
  g510
  (
    n538,
    n132
  );


  not
  g511
  (
    n436,
    n61
  );


  buf
  g512
  (
    n429,
    n51
  );


  buf
  g513
  (
    n292,
    n133
  );


  not
  g514
  (
    n259,
    n67
  );


  not
  g515
  (
    n177,
    n130
  );


  not
  g516
  (
    n484,
    n42
  );


  not
  g517
  (
    n467,
    n132
  );


  not
  g518
  (
    n449,
    n128
  );


  not
  g519
  (
    n571,
    n142
  );


  not
  g520
  (
    n265,
    n56
  );


  not
  g521
  (
    n311,
    n135
  );


  buf
  g522
  (
    n346,
    n40
  );


  not
  g523
  (
    n553,
    n82
  );


  buf
  g524
  (
    KeyWire_0_28,
    n64
  );


  not
  g525
  (
    n507,
    n69
  );


  xnor
  g526
  (
    n386,
    n83,
    n34
  );


  and
  g527
  (
    n165,
    n142,
    n77,
    n97,
    n127
  );


  or
  g528
  (
    n561,
    n65,
    n129,
    n62,
    n139
  );


  and
  g529
  (
    KeyWire_0_27,
    n96,
    n100,
    n44,
    n113
  );


  and
  g530
  (
    n239,
    n135,
    n39,
    n106,
    n132
  );


  or
  g531
  (
    n224,
    n121,
    n49,
    n77,
    n65
  );


  nor
  g532
  (
    n245,
    n117,
    n131,
    n69,
    n40
  );


  nand
  g533
  (
    n391,
    n35,
    n136,
    n149,
    n63
  );


  xnor
  g534
  (
    n474,
    n53,
    n36,
    n105,
    n119
  );


  nor
  g535
  (
    n488,
    n38,
    n73,
    n46,
    n118
  );


  nand
  g536
  (
    n421,
    n104,
    n76,
    n56,
    n84
  );


  xor
  g537
  (
    n329,
    n125,
    n133,
    n100,
    n74
  );


  nor
  g538
  (
    n198,
    n71,
    n57,
    n79,
    n75
  );


  xnor
  g539
  (
    n243,
    n70,
    n108,
    n32,
    n62
  );


  nor
  g540
  (
    n439,
    n72,
    n66,
    n120,
    n111
  );


  nor
  g541
  (
    n396,
    n127,
    n58,
    n61,
    n72
  );


  and
  g542
  (
    n486,
    n135,
    n145,
    n95,
    n67
  );


  or
  g543
  (
    n276,
    n134,
    n142,
    n117,
    n86
  );


  and
  g544
  (
    n447,
    n50,
    n140,
    n141,
    n37
  );


  nand
  g545
  (
    n508,
    n52,
    n112,
    n109,
    n114
  );


  not
  g546
  (
    n688,
    n314
  );


  not
  g547
  (
    n669,
    n170
  );


  not
  g548
  (
    n727,
    n308
  );


  buf
  g549
  (
    n739,
    n285
  );


  buf
  g550
  (
    KeyWire_0_0,
    n222
  );


  buf
  g551
  (
    n691,
    n274
  );


  buf
  g552
  (
    n623,
    n309
  );


  not
  g553
  (
    n648,
    n173
  );


  buf
  g554
  (
    n689,
    n303
  );


  buf
  g555
  (
    n663,
    n209
  );


  not
  g556
  (
    n625,
    n209
  );


  buf
  g557
  (
    n616,
    n251
  );


  not
  g558
  (
    n675,
    n347
  );


  not
  g559
  (
    n615,
    n169
  );


  not
  g560
  (
    n600,
    n287
  );


  not
  g561
  (
    n700,
    n184
  );


  not
  g562
  (
    n681,
    n286
  );


  not
  g563
  (
    n706,
    n173
  );


  not
  g564
  (
    n729,
    n222
  );


  not
  g565
  (
    n750,
    n330
  );


  buf
  g566
  (
    n581,
    n263
  );


  buf
  g567
  (
    n666,
    n264
  );


  buf
  g568
  (
    n762,
    n228
  );


  not
  g569
  (
    n670,
    n258
  );


  not
  g570
  (
    n715,
    n267
  );


  buf
  g571
  (
    n754,
    n235
  );


  not
  g572
  (
    n597,
    n348
  );


  not
  g573
  (
    n585,
    n313
  );


  not
  g574
  (
    n760,
    n291
  );


  not
  g575
  (
    n718,
    n199
  );


  buf
  g576
  (
    n653,
    n266
  );


  buf
  g577
  (
    n631,
    n349
  );


  buf
  g578
  (
    n723,
    n204
  );


  buf
  g579
  (
    n769,
    n223
  );


  not
  g580
  (
    n731,
    n273
  );


  buf
  g581
  (
    n752,
    n282
  );


  buf
  g582
  (
    n589,
    n215
  );


  buf
  g583
  (
    n733,
    n199
  );


  buf
  g584
  (
    n740,
    n331
  );


  buf
  g585
  (
    n599,
    n264
  );


  buf
  g586
  (
    n747,
    n300
  );


  not
  g587
  (
    n620,
    n270
  );


  not
  g588
  (
    n614,
    n240
  );


  buf
  g589
  (
    n743,
    n157
  );


  buf
  g590
  (
    n776,
    n351
  );


  not
  g591
  (
    n745,
    n162
  );


  buf
  g592
  (
    n696,
    n161
  );


  buf
  g593
  (
    n725,
    n249
  );


  not
  g594
  (
    n734,
    n342
  );


  buf
  g595
  (
    n596,
    n332
  );


  buf
  g596
  (
    n774,
    n200
  );


  buf
  g597
  (
    n621,
    n252
  );


  not
  g598
  (
    n661,
    n254
  );


  not
  g599
  (
    n652,
    n314
  );


  not
  g600
  (
    n682,
    n299
  );


  buf
  g601
  (
    n757,
    n333
  );


  buf
  g602
  (
    n645,
    n244
  );


  not
  g603
  (
    n741,
    n227
  );


  buf
  g604
  (
    n707,
    n318
  );


  buf
  g605
  (
    n618,
    n252
  );


  buf
  g606
  (
    n619,
    n335
  );


  not
  g607
  (
    n612,
    n185
  );


  not
  g608
  (
    n719,
    n343
  );


  not
  g609
  (
    n679,
    n305
  );


  not
  g610
  (
    KeyWire_0_25,
    n185
  );


  buf
  g611
  (
    n736,
    n307
  );


  buf
  g612
  (
    n654,
    n174
  );


  buf
  g613
  (
    n755,
    n319
  );


  not
  g614
  (
    n758,
    n242
  );


  buf
  g615
  (
    n698,
    n353
  );


  not
  g616
  (
    n678,
    n281
  );


  not
  g617
  (
    n632,
    n212
  );


  buf
  g618
  (
    n677,
    n166
  );


  not
  g619
  (
    n580,
    n337
  );


  buf
  g620
  (
    n629,
    n218
  );


  not
  g621
  (
    n703,
    n238
  );


  not
  g622
  (
    n628,
    n213
  );


  not
  g623
  (
    n694,
    n345
  );


  not
  g624
  (
    n642,
    n344
  );


  not
  g625
  (
    n668,
    n269
  );


  buf
  g626
  (
    n635,
    n334
  );


  not
  g627
  (
    KeyWire_0_12,
    n215
  );


  buf
  g628
  (
    n770,
    n329
  );


  buf
  g629
  (
    n686,
    n231
  );


  buf
  g630
  (
    n637,
    n266
  );


  not
  g631
  (
    n651,
    n187
  );


  not
  g632
  (
    n705,
    n217
  );


  not
  g633
  (
    n659,
    n262
  );


  not
  g634
  (
    n773,
    n355
  );


  not
  g635
  (
    n673,
    n354
  );


  buf
  g636
  (
    n605,
    n304
  );


  not
  g637
  (
    n609,
    n294
  );


  not
  g638
  (
    n601,
    n285
  );


  buf
  g639
  (
    n710,
    n188
  );


  not
  g640
  (
    n647,
    n168
  );


  buf
  g641
  (
    n712,
    n172
  );


  not
  g642
  (
    n685,
    n186
  );


  not
  g643
  (
    n713,
    n159
  );


  not
  g644
  (
    n656,
    n316
  );


  not
  g645
  (
    n708,
    n286
  );


  not
  g646
  (
    n704,
    n283
  );


  not
  g647
  (
    n626,
    n253
  );


  buf
  g648
  (
    n764,
    n338
  );


  not
  g649
  (
    n639,
    n326
  );


  buf
  g650
  (
    n594,
    n187
  );


  buf
  g651
  (
    n749,
    n310
  );


  not
  g652
  (
    n671,
    n191
  );


  not
  g653
  (
    n765,
    n164
  );


  buf
  g654
  (
    n697,
    n224
  );


  not
  g655
  (
    n606,
    n275
  );


  buf
  g656
  (
    n584,
    n256
  );


  not
  g657
  (
    n582,
    n302
  );


  not
  g658
  (
    n728,
    n304
  );


  buf
  g659
  (
    KeyWire_0_6,
    n271
  );


  buf
  g660
  (
    n683,
    n258
  );


  buf
  g661
  (
    n638,
    n254
  );


  not
  g662
  (
    n579,
    n290
  );


  not
  g663
  (
    n726,
    n292
  );


  not
  g664
  (
    n634,
    n325
  );


  not
  g665
  (
    n607,
    n214
  );


  buf
  g666
  (
    n735,
    n224
  );


  not
  g667
  (
    n768,
    n217
  );


  not
  g668
  (
    n650,
    n311
  );


  buf
  g669
  (
    n744,
    n246
  );


  buf
  g670
  (
    n717,
    n297
  );


  not
  g671
  (
    n640,
    n293
  );


  buf
  g672
  (
    n664,
    n196
  );


  not
  g673
  (
    n662,
    n207
  );


  buf
  g674
  (
    n593,
    n163
  );


  buf
  g675
  (
    n636,
    n346
  );


  buf
  g676
  (
    KeyWire_0_16,
    n317
  );


  buf
  g677
  (
    n687,
    n294
  );


  nand
  g678
  (
    n598,
    n282,
    n208
  );


  xnor
  g679
  (
    n595,
    n322,
    n165
  );


  xnor
  g680
  (
    n701,
    n219,
    n260,
    n295,
    n184
  );


  nand
  g681
  (
    n646,
    n177,
    n236,
    n339,
    n211
  );


  nand
  g682
  (
    n766,
    n348,
    n192,
    n234,
    n179
  );


  or
  g683
  (
    KeyWire_0_14,
    n298,
    n307,
    n165,
    n158
  );


  nand
  g684
  (
    n611,
    n245,
    n228,
    n158,
    n229
  );


  nor
  g685
  (
    n644,
    n189,
    n175,
    n318,
    n262
  );


  nand
  g686
  (
    n714,
    n268,
    n239,
    n316,
    n163
  );


  or
  g687
  (
    n603,
    n313,
    n226,
    n328,
    n181
  );


  and
  g688
  (
    n622,
    n347,
    n171,
    n168,
    n216
  );


  xor
  g689
  (
    n592,
    n240,
    n250,
    n161,
    n274
  );


  nor
  g690
  (
    n660,
    n351,
    n324,
    n279,
    n164
  );


  or
  g691
  (
    n587,
    n336,
    n269,
    n340,
    n334
  );


  and
  g692
  (
    n721,
    n194,
    n270,
    n261,
    n230
  );


  or
  g693
  (
    n630,
    n195,
    n201,
    n189,
    n331
  );


  xor
  g694
  (
    n617,
    n259,
    n238,
    n204,
    n169
  );


  xor
  g695
  (
    n655,
    n311,
    n225,
    n246,
    n273
  );


  xor
  g696
  (
    n742,
    n305,
    n292,
    n231,
    n247
  );


  nor
  g697
  (
    n583,
    n349,
    n179,
    n214,
    n284
  );


  and
  g698
  (
    n709,
    n181,
    n206,
    n172,
    n166
  );


  xor
  g699
  (
    n763,
    n248,
    n295,
    n308,
    n322
  );


  xor
  g700
  (
    n759,
    n345,
    n203,
    n263,
    n190
  );


  or
  g701
  (
    n658,
    n284,
    n265,
    n195,
    n355
  );


  nor
  g702
  (
    n676,
    n182,
    n194,
    n213,
    n244
  );


  and
  g703
  (
    n590,
    n210,
    n281,
    n156,
    n198
  );


  xor
  g704
  (
    KeyWire_0_29,
    n162,
    n177,
    n167,
    n200
  );


  xnor
  g705
  (
    n680,
    n324,
    n280,
    n206,
    n237
  );


  xnor
  g706
  (
    n772,
    n183,
    n293,
    n212,
    n336
  );


  nor
  g707
  (
    n756,
    n277,
    n191,
    n193,
    n216
  );


  and
  g708
  (
    n627,
    n291,
    n234,
    n288,
    n271
  );


  xor
  g709
  (
    n604,
    n352,
    n225,
    n190,
    n344
  );


  or
  g710
  (
    n722,
    n220,
    n340,
    n289,
    n174
  );


  and
  g711
  (
    n711,
    n339,
    n288,
    n253,
    n211
  );


  nor
  g712
  (
    n624,
    n188,
    n332,
    n256,
    n178
  );


  nor
  g713
  (
    n777,
    n198,
    n299,
    n242,
    n272
  );


  xnor
  g714
  (
    n716,
    n197,
    n277,
    n306
  );


  xnor
  g715
  (
    n730,
    n219,
    n241,
    n267,
    n278
  );


  xnor
  g716
  (
    n767,
    n160,
    n226,
    n283,
    n303
  );


  nand
  g717
  (
    n761,
    n327,
    n350,
    n223
  );


  nor
  g718
  (
    n633,
    n296,
    n300,
    n255,
    n180
  );


  nor
  g719
  (
    n695,
    n321,
    n272,
    n289,
    n193
  );


  xor
  g720
  (
    n649,
    n275,
    n248,
    n301,
    n325
  );


  and
  g721
  (
    n665,
    n328,
    n312,
    n342,
    n343
  );


  or
  g722
  (
    n732,
    n170,
    n280,
    n197,
    n297
  );


  nor
  g723
  (
    n591,
    n323,
    n320,
    n220,
    n233
  );


  xnor
  g724
  (
    n613,
    n176,
    n341,
    n210,
    n183
  );


  or
  g725
  (
    n748,
    n207,
    n320,
    n329,
    n180
  );


  xnor
  g726
  (
    n578,
    n221,
    n278,
    n250,
    n178
  );


  xnor
  g727
  (
    n657,
    n315,
    n243,
    n160,
    n255
  );


  nor
  g728
  (
    n751,
    n243,
    n235,
    n230,
    n327
  );


  nor
  g729
  (
    n684,
    n247,
    n186,
    n257,
    n205
  );


  nand
  g730
  (
    n690,
    n287,
    n249,
    n310,
    n171
  );


  nand
  g731
  (
    n608,
    n337,
    n296,
    n346,
    n201
  );


  xnor
  g732
  (
    n720,
    n290,
    n335,
    n317,
    n301
  );


  or
  g733
  (
    n643,
    n205,
    n239,
    n298,
    n354
  );


  nor
  g734
  (
    n737,
    n352,
    n309,
    n268,
    n323
  );


  and
  g735
  (
    n610,
    n338,
    n260,
    n236,
    n257
  );


  nor
  g736
  (
    n672,
    n203,
    n251,
    n202,
    n276
  );


  nand
  g737
  (
    n586,
    n229,
    n233,
    n319,
    n208
  );


  nor
  g738
  (
    n674,
    n202,
    n341,
    n245,
    n192
  );


  and
  g739
  (
    n692,
    n241,
    n326,
    n182,
    n156
  );


  and
  g740
  (
    n746,
    n302,
    n159,
    n265,
    n321
  );


  or
  g741
  (
    n699,
    n315,
    n232,
    n259,
    n279
  );


  and
  g742
  (
    n771,
    n176,
    n167,
    n312,
    n232
  );


  or
  g743
  (
    n667,
    n175,
    n237,
    n196,
    n218
  );


  or
  g744
  (
    n693,
    n261,
    n157,
    n227,
    n221
  );


  or
  g745
  (
    n641,
    n330,
    n333,
    n353,
    n276
  );


  not
  g746
  (
    n866,
    n390
  );


  buf
  g747
  (
    n806,
    n366
  );


  buf
  g748
  (
    n864,
    n421
  );


  not
  g749
  (
    n818,
    n632
  );


  buf
  g750
  (
    n787,
    n678
  );


  not
  g751
  (
    n782,
    n683
  );


  buf
  g752
  (
    n786,
    n423
  );


  buf
  g753
  (
    n832,
    n743
  );


  or
  g754
  (
    n871,
    n756,
    n697,
    n607,
    n629
  );


  and
  g755
  (
    n819,
    n646,
    n374,
    n430,
    n761
  );


  or
  g756
  (
    n820,
    n411,
    n365,
    n377,
    n692
  );


  and
  g757
  (
    n804,
    n734,
    n358,
    n676,
    n363
  );


  xnor
  g758
  (
    n794,
    n431,
    n435,
    n583,
    n653
  );


  nand
  g759
  (
    n858,
    n356,
    n400,
    n420,
    n762
  );


  xor
  g760
  (
    n783,
    n384,
    n392,
    n400,
    n387
  );


  xor
  g761
  (
    n838,
    n361,
    n730,
    n609,
    n382
  );


  and
  g762
  (
    n873,
    n394,
    n590,
    n429,
    n598
  );


  nor
  g763
  (
    n816,
    n397,
    n751,
    n402,
    n765
  );


  and
  g764
  (
    n853,
    n417,
    n735,
    n687,
    n406
  );


  xor
  g765
  (
    n843,
    n723,
    n580,
    n406,
    n766
  );


  xnor
  g766
  (
    n869,
    n699,
    n688,
    n388,
    n367
  );


  or
  g767
  (
    n854,
    n648,
    n373,
    n693,
    n635
  );


  nand
  g768
  (
    n827,
    n642,
    n720,
    n601,
    n746
  );


  nor
  g769
  (
    n835,
    n617,
    n368,
    n380,
    n433
  );


  or
  g770
  (
    n862,
    n395,
    n401,
    n435,
    n658
  );


  and
  g771
  (
    n793,
    n584,
    n373,
    n370,
    n423
  );


  nor
  g772
  (
    n792,
    n718,
    n602,
    n404,
    n733
  );


  nand
  g773
  (
    KeyWire_0_19,
    n690,
    n659,
    n424,
    n732
  );


  nand
  g774
  (
    n863,
    n611,
    n385,
    n403,
    n756
  );


  nand
  g775
  (
    n802,
    n389,
    n713,
    n633,
    n375
  );


  xnor
  g776
  (
    n789,
    n670,
    n766,
    n358,
    n432
  );


  xnor
  g777
  (
    n805,
    n739,
    n685,
    n428,
    n765
  );


  or
  g778
  (
    n855,
    n621,
    n405,
    n403,
    n631
  );


  or
  g779
  (
    n791,
    n694,
    n684,
    n737,
    n582
  );


  xnor
  g780
  (
    n859,
    n359,
    n421,
    n378,
    n744
  );


  or
  g781
  (
    n801,
    n395,
    n759,
    n589,
    n422
  );


  xnor
  g782
  (
    n861,
    n364,
    n715,
    n591,
    n387
  );


  nand
  g783
  (
    n876,
    n376,
    n360,
    n711,
    n615
  );


  or
  g784
  (
    n870,
    n754,
    n759,
    n357,
    n752
  );


  xor
  g785
  (
    n821,
    n764,
    n408,
    n657,
    n378
  );


  or
  g786
  (
    n825,
    n741,
    n665,
    n717,
    n691
  );


  nand
  g787
  (
    n829,
    n760,
    n647,
    n593,
    n592
  );


  or
  g788
  (
    n808,
    n651,
    n391,
    n605,
    n757
  );


  nor
  g789
  (
    n779,
    n702,
    n695,
    n414,
    n636
  );


  nor
  g790
  (
    n796,
    n396,
    n763,
    n587,
    n415
  );


  and
  g791
  (
    n851,
    n600,
    n639,
    n761,
    n418
  );


  xor
  g792
  (
    n844,
    n412,
    n751,
    n371,
    n705
  );


  or
  g793
  (
    n846,
    n614,
    n748,
    n622,
    n755
  );


  or
  g794
  (
    n840,
    n383,
    n357,
    n434,
    n426
  );


  nor
  g795
  (
    n809,
    n595,
    n757,
    n663,
    n381
  );


  xor
  g796
  (
    n795,
    n764,
    n579,
    n578,
    n418
  );


  and
  g797
  (
    n831,
    n411,
    n376,
    n727,
    n738
  );


  nand
  g798
  (
    n849,
    n638,
    n731,
    n362,
    n745
  );


  nand
  g799
  (
    n833,
    n425,
    n752,
    n366,
    n654
  );


  or
  g800
  (
    n815,
    n626,
    n655,
    n393,
    n425
  );


  nand
  g801
  (
    n812,
    n650,
    n640,
    n415,
    n669
  );


  or
  g802
  (
    n872,
    n384,
    n372,
    n382,
    n641
  );


  and
  g803
  (
    n822,
    n413,
    n408,
    n677,
    n405
  );


  and
  g804
  (
    n852,
    n399,
    n597,
    n586,
    n728
  );


  and
  g805
  (
    n860,
    n581,
    n666,
    n753,
    n763
  );


  nand
  g806
  (
    n807,
    n379,
    n672,
    n427,
    n383
  );


  xor
  g807
  (
    n857,
    n725,
    n392,
    n431,
    n414
  );


  xor
  g808
  (
    n830,
    n369,
    n394,
    n628,
    n625
  );


  xnor
  g809
  (
    n834,
    n767,
    n624,
    n645,
    n402
  );


  xnor
  g810
  (
    n790,
    n675,
    n767,
    n643,
    n668
  );


  and
  g811
  (
    n847,
    n374,
    n634,
    n682,
    n365
  );


  xnor
  g812
  (
    n813,
    n417,
    n627,
    n608,
    n644
  );


  nand
  g813
  (
    n814,
    n686,
    n721,
    n385,
    n612
  );


  nor
  g814
  (
    n837,
    n432,
    n710,
    n742,
    n719
  );


  xnor
  g815
  (
    n810,
    n398,
    n420,
    n372,
    n412
  );


  xor
  g816
  (
    n817,
    n360,
    n724,
    n390,
    n637
  );


  and
  g817
  (
    n875,
    n424,
    n413,
    n409,
    n410
  );


  and
  g818
  (
    n778,
    n398,
    n660,
    n429,
    n753
  );


  xnor
  g819
  (
    KeyWire_0_21,
    n613,
    n436,
    n661,
    n416
  );


  or
  g820
  (
    n800,
    n716,
    n698,
    n708,
    n391
  );


  nand
  g821
  (
    n865,
    n371,
    n434,
    n679,
    n393
  );


  nand
  g822
  (
    n799,
    n404,
    n616,
    n379,
    n388
  );


  and
  g823
  (
    n850,
    n736,
    n623,
    n416,
    n704
  );


  nor
  g824
  (
    n868,
    n620,
    n389,
    n758,
    n362
  );


  nand
  g825
  (
    n826,
    n422,
    n410,
    n755,
    n709
  );


  xnor
  g826
  (
    n785,
    n706,
    n437,
    n656,
    n696
  );


  nor
  g827
  (
    n811,
    n673,
    n437,
    n722,
    n428
  );


  nor
  g828
  (
    n797,
    n750,
    n407,
    n760,
    n649
  );


  xor
  g829
  (
    n784,
    n370,
    n762,
    n604,
    n369
  );


  nand
  g830
  (
    n824,
    n375,
    n380,
    n618,
    n681
  );


  or
  g831
  (
    n803,
    n606,
    n667,
    n754,
    n436
  );


  nand
  g832
  (
    n798,
    n610,
    n401,
    n368,
    n662
  );


  nor
  g833
  (
    n836,
    n356,
    n363,
    n700,
    n712
  );


  or
  g834
  (
    n780,
    n749,
    n361,
    n603,
    n701
  );


  or
  g835
  (
    n839,
    n433,
    n419,
    n427,
    n396
  );


  xnor
  g836
  (
    n842,
    n652,
    n364,
    n768,
    n619
  );


  and
  g837
  (
    n856,
    n707,
    n594,
    n367,
    n729
  );


  nand
  g838
  (
    n845,
    n630,
    n740,
    n399,
    n671
  );


  and
  g839
  (
    n788,
    n386,
    n359,
    n430,
    n426
  );


  xor
  g840
  (
    n823,
    n758,
    n419,
    n599,
    n680
  );


  xnor
  g841
  (
    n867,
    n407,
    n397,
    n726,
    n714
  );


  nand
  g842
  (
    n874,
    n585,
    n747,
    n689,
    n377
  );


  nand
  g843
  (
    n848,
    n381,
    n703,
    n674,
    n409
  );


  nor
  g844
  (
    n781,
    n664,
    n588,
    n596,
    n386
  );


  buf
  g845
  (
    n886,
    n778
  );


  not
  g846
  (
    n879,
    n787
  );


  nor
  g847
  (
    n878,
    n783,
    n781
  );


  and
  g848
  (
    n883,
    n784,
    n791,
    n786,
    n788
  );


  or
  g849
  (
    n882,
    n787,
    n791,
    n778,
    n782
  );


  nor
  g850
  (
    n884,
    n792,
    n792,
    n789,
    n790
  );


  xor
  g851
  (
    n880,
    n779,
    n793,
    n784,
    n785
  );


  and
  g852
  (
    n881,
    n789,
    n781,
    n782,
    n785
  );


  and
  g853
  (
    n885,
    n780,
    n783,
    n788,
    n793
  );


  nand
  g854
  (
    n877,
    n786,
    n780,
    n779,
    n790
  );


  xnor
  g855
  (
    n888,
    n880,
    n881,
    n883,
    n877
  );


  nand
  g856
  (
    n893,
    n878,
    n882,
    n881
  );


  nor
  g857
  (
    n887,
    n884,
    n880,
    n879
  );


  xor
  g858
  (
    n891,
    n878,
    n883,
    n884,
    n879
  );


  nor
  g859
  (
    KeyWire_0_4,
    n878,
    n883,
    n877,
    n882
  );


  xnor
  g860
  (
    n892,
    n880,
    n884,
    n877,
    n878
  );


  or
  g861
  (
    n894,
    n882,
    n881,
    n879
  );


  nand
  g862
  (
    n889,
    n877,
    n883,
    n884,
    n879
  );


  and
  g863
  (
    n902,
    n443,
    n441,
    n442,
    n447
  );


  nor
  g864
  (
    n901,
    n887,
    n449,
    n448
  );


  nor
  g865
  (
    n897,
    n446,
    n439,
    n891,
    n893
  );


  xnor
  g866
  (
    n896,
    n892,
    n440,
    n890,
    n888
  );


  nand
  g867
  (
    n899,
    n445,
    n447,
    n441,
    n438
  );


  and
  g868
  (
    n898,
    n440,
    n889,
    n438,
    n442
  );


  or
  g869
  (
    n895,
    n443,
    n444,
    n445,
    n893
  );


  nand
  g870
  (
    n900,
    n446,
    n439,
    n444,
    n448
  );


  buf
  g871
  (
    n929,
    n455
  );


  not
  g872
  (
    n912,
    n450
  );


  not
  g873
  (
    n917,
    n775
  );


  not
  g874
  (
    n928,
    n898
  );


  not
  g875
  (
    n922,
    n898
  );


  not
  g876
  (
    n915,
    n894
  );


  not
  g877
  (
    n904,
    n895
  );


  not
  g878
  (
    n924,
    n773
  );


  buf
  g879
  (
    n925,
    n901
  );


  not
  g880
  (
    n923,
    n899
  );


  and
  g881
  (
    n916,
    n798,
    n796
  );


  or
  g882
  (
    n903,
    n776,
    n453,
    n902,
    n899
  );


  xnor
  g883
  (
    n920,
    n896,
    n775,
    n902,
    n899
  );


  nand
  g884
  (
    n930,
    n896,
    n796,
    n900
  );


  nand
  g885
  (
    n921,
    n897,
    n895,
    n772,
    n774
  );


  and
  g886
  (
    n919,
    n774,
    n896,
    n770,
    n769
  );


  nor
  g887
  (
    n909,
    n777,
    n451,
    n454,
    n897
  );


  nor
  g888
  (
    n918,
    n799,
    n900,
    n795,
    n899
  );


  or
  g889
  (
    n905,
    n771,
    n456,
    n457,
    n901
  );


  nand
  g890
  (
    n906,
    n455,
    n795,
    n798,
    n794
  );


  xnor
  g891
  (
    n907,
    n898,
    n777,
    n452,
    n776
  );


  or
  g892
  (
    n926,
    n902,
    n457,
    n453,
    n797
  );


  or
  g893
  (
    n927,
    n771,
    n900,
    n894,
    n768
  );


  and
  g894
  (
    n911,
    n772,
    n450,
    n773,
    n901
  );


  nand
  g895
  (
    n913,
    n454,
    n898,
    n769,
    n896
  );


  xnor
  g896
  (
    n914,
    n794,
    n897,
    n451,
    n152
  );


  xnor
  g897
  (
    n910,
    n902,
    n452,
    n897,
    n770
  );


  nand
  g898
  (
    KeyWire_0_22,
    n797,
    n895,
    n456,
    n901
  );


  nand
  g899
  (
    n1007,
    n546,
    n831,
    n568,
    n918
  );


  xor
  g900
  (
    n956,
    n911,
    n903,
    n557,
    n478
  );


  and
  g901
  (
    n935,
    n467,
    n909,
    n921,
    n905
  );


  xor
  g902
  (
    n995,
    n562,
    n822,
    n491,
    n564
  );


  nand
  g903
  (
    n955,
    n559,
    n906,
    n903,
    n484
  );


  nor
  g904
  (
    n1021,
    n574,
    n805,
    n924,
    n503
  );


  and
  g905
  (
    n966,
    n498,
    n472,
    n538,
    n907
  );


  xor
  g906
  (
    n983,
    n806,
    n920,
    n473,
    n534
  );


  or
  g907
  (
    n1029,
    n919,
    n476,
    n530,
    n526
  );


  and
  g908
  (
    n954,
    n535,
    n569,
    n561,
    n918
  );


  nand
  g909
  (
    n1010,
    n528,
    n826,
    n832,
    n464
  );


  and
  g910
  (
    n981,
    n824,
    n916,
    n912,
    n905
  );


  or
  g911
  (
    n988,
    n550,
    n486,
    n914,
    n574
  );


  or
  g912
  (
    n968,
    n519,
    n561,
    n904,
    n825
  );


  nand
  g913
  (
    n992,
    n509,
    n527,
    n904,
    n501
  );


  nand
  g914
  (
    n982,
    n542,
    n816,
    n536,
    n516
  );


  nor
  g915
  (
    n1037,
    n827,
    n571,
    n805,
    n911
  );


  xor
  g916
  (
    n1020,
    n469,
    n568,
    n928,
    n483
  );


  nand
  g917
  (
    n959,
    n565,
    n559,
    n804,
    n906
  );


  nor
  g918
  (
    n1041,
    n523,
    n487,
    n562,
    n516
  );


  xor
  g919
  (
    n987,
    n570,
    n488,
    n912,
    n552
  );


  xnor
  g920
  (
    n964,
    n572,
    n926,
    n461,
    n922
  );


  nand
  g921
  (
    n996,
    n825,
    n803,
    n504,
    n480
  );


  xnor
  g922
  (
    n974,
    n574,
    n826,
    n930,
    n495
  );


  nand
  g923
  (
    n985,
    n507,
    n925,
    n475,
    n494
  );


  nor
  g924
  (
    n936,
    n533,
    n495,
    n490,
    n551
  );


  or
  g925
  (
    n1039,
    n549,
    n567,
    n508,
    n923
  );


  nor
  g926
  (
    n1013,
    n907,
    n917,
    n928,
    n489
  );


  or
  g927
  (
    n1027,
    n543,
    n513,
    n522,
    n925
  );


  nor
  g928
  (
    n1016,
    n553,
    n514,
    n806,
    n552
  );


  or
  g929
  (
    n975,
    n528,
    n925,
    n922,
    n926
  );


  nor
  g930
  (
    n943,
    n472,
    n501,
    n921,
    n831
  );


  xnor
  g931
  (
    n1006,
    n563,
    n920,
    n926,
    n478
  );


  or
  g932
  (
    n941,
    n517,
    n914,
    n512,
    n463
  );


  nand
  g933
  (
    n972,
    n511,
    n567,
    n919,
    n460
  );


  or
  g934
  (
    n997,
    n499,
    n560,
    n815,
    n801
  );


  xnor
  g935
  (
    n980,
    n916,
    n461,
    n928,
    n568
  );


  and
  g936
  (
    n932,
    n570,
    n527,
    n908,
    n812
  );


  nand
  g937
  (
    n979,
    n830,
    n927,
    n565,
    n575
  );


  and
  g938
  (
    n942,
    n484,
    n913,
    n531,
    n800
  );


  and
  g939
  (
    n1040,
    n811,
    n468,
    n918,
    n818
  );


  and
  g940
  (
    n1003,
    n908,
    n910,
    n808
  );


  or
  g941
  (
    n931,
    n497,
    n542,
    n914,
    n814
  );


  nor
  g942
  (
    n1038,
    n910,
    n565,
    n919,
    n813
  );


  or
  g943
  (
    n990,
    n820,
    n547,
    n485,
    n917
  );


  xnor
  g944
  (
    n971,
    n504,
    n923,
    n915
  );


  nor
  g945
  (
    n1036,
    n569,
    n556,
    n489,
    n908
  );


  xnor
  g946
  (
    n967,
    n930,
    n924,
    n814,
    n510
  );


  nand
  g947
  (
    n984,
    n917,
    n462,
    n829
  );


  xor
  g948
  (
    n960,
    n544,
    n502,
    n487,
    n498
  );


  or
  g949
  (
    n939,
    n493,
    n463,
    n560,
    n801
  );


  nor
  g950
  (
    n1015,
    n520,
    n912,
    n541,
    n471
  );


  xor
  g951
  (
    n1028,
    n906,
    n802,
    n482,
    n493
  );


  xnor
  g952
  (
    n953,
    n477,
    n930,
    n514,
    n518
  );


  or
  g953
  (
    n1008,
    n522,
    n548,
    n541,
    n515
  );


  xnor
  g954
  (
    n1042,
    n519,
    n474,
    n909,
    n828
  );


  nand
  g955
  (
    n962,
    n465,
    n914,
    n572,
    n921
  );


  xor
  g956
  (
    n998,
    n569,
    n563,
    n500,
    n821
  );


  xnor
  g957
  (
    n1017,
    n570,
    n488,
    n486,
    n471
  );


  xor
  g958
  (
    n938,
    n470,
    n567,
    n562,
    n816
  );


  nor
  g959
  (
    n961,
    n926,
    n909,
    n458,
    n919
  );


  nand
  g960
  (
    n1032,
    n523,
    n572,
    n566,
    n554
  );


  xnor
  g961
  (
    n973,
    n911,
    n492,
    n923,
    n483
  );


  xnor
  g962
  (
    n994,
    n813,
    n565,
    n479,
    n920
  );


  nor
  g963
  (
    n949,
    n561,
    n529,
    n808,
    n465
  );


  and
  g964
  (
    n937,
    n529,
    n819,
    n497,
    n517
  );


  and
  g965
  (
    n1000,
    n799,
    n570,
    n913,
    n927
  );


  xnor
  g966
  (
    n1031,
    n526,
    n555,
    n564,
    n807
  );


  and
  g967
  (
    n1035,
    n910,
    n467,
    n909,
    n502
  );


  xor
  g968
  (
    n965,
    n466,
    n573,
    n917,
    n800
  );


  nand
  g969
  (
    n947,
    n515,
    n548,
    n563,
    n525
  );


  nand
  g970
  (
    n999,
    n557,
    n930,
    n479,
    n821
  );


  nor
  g971
  (
    n978,
    n916,
    n513,
    n556,
    n507
  );


  nor
  g972
  (
    n989,
    n503,
    n531,
    n809,
    n485
  );


  and
  g973
  (
    n952,
    n820,
    n905,
    n929,
    n903
  );


  nand
  g974
  (
    n1030,
    n530,
    n540,
    n545,
    n815
  );


  nor
  g975
  (
    n1033,
    n532,
    n571,
    n913,
    n537
  );


  or
  g976
  (
    n986,
    n807,
    n532,
    n524,
    n929
  );


  xor
  g977
  (
    n1002,
    n823,
    n480,
    n560,
    n827
  );


  or
  g978
  (
    n1022,
    n920,
    n490,
    n491,
    n509
  );


  and
  g979
  (
    n1001,
    n505,
    n832,
    n810,
    n500
  );


  xnor
  g980
  (
    n969,
    n505,
    n521,
    n824,
    n496
  );


  xor
  g981
  (
    n1009,
    n822,
    n547,
    n907,
    n563
  );


  and
  g982
  (
    n993,
    n904,
    n575,
    n521,
    n460
  );


  xor
  g983
  (
    n991,
    n545,
    n462,
    n925,
    n918
  );


  and
  g984
  (
    n1012,
    n468,
    n496,
    n804,
    n575
  );


  xnor
  g985
  (
    n976,
    n568,
    n907,
    n903,
    n458
  );


  or
  g986
  (
    n958,
    n464,
    n569,
    n905,
    n573
  );


  xnor
  g987
  (
    n957,
    n912,
    n573,
    n553,
    n539
  );


  nor
  g988
  (
    n944,
    n817,
    n566,
    n533,
    n562
  );


  xor
  g989
  (
    n963,
    n474,
    n506,
    n566,
    n923
  );


  nor
  g990
  (
    n946,
    n564,
    n566,
    n904,
    n922
  );


  xor
  g991
  (
    n934,
    n492,
    n550,
    n508,
    n512
  );


  xor
  g992
  (
    n970,
    n506,
    n573,
    n823,
    n546
  );


  nor
  g993
  (
    n1023,
    n518,
    n833,
    n459,
    n470
  );


  xnor
  g994
  (
    n1004,
    n571,
    n524,
    n555,
    n499
  );


  or
  g995
  (
    n948,
    n906,
    n924,
    n544,
    n543
  );


  xnor
  g996
  (
    n940,
    n558,
    n929,
    n535,
    n473
  );


  and
  g997
  (
    n1018,
    n538,
    n572,
    n511,
    n466
  );


  xor
  g998
  (
    n1024,
    n476,
    n574,
    n561,
    n828
  );


  and
  g999
  (
    n1014,
    n567,
    n809,
    n475,
    n818
  );


  and
  g1000
  (
    n951,
    n481,
    n549,
    n927,
    n560
  );


  xnor
  g1001
  (
    n945,
    n803,
    n812,
    n575,
    n830
  );


  nand
  g1002
  (
    n1026,
    n817,
    n481,
    n554,
    n564
  );


  nand
  g1003
  (
    n933,
    n916,
    n819,
    n482,
    n927
  );


  or
  g1004
  (
    n1025,
    n520,
    n915,
    n477,
    n525
  );


  nand
  g1005
  (
    n950,
    n924,
    n928,
    n539,
    n510
  );


  xor
  g1006
  (
    n1019,
    n811,
    n908,
    n571,
    n534
  );


  xor
  g1007
  (
    n1005,
    n911,
    n810,
    n469,
    n921
  );


  and
  g1008
  (
    n1034,
    n913,
    n537,
    n802,
    n540
  );


  or
  g1009
  (
    n1011,
    n459,
    n494,
    n915,
    n929
  );


  and
  g1010
  (
    n977,
    n922,
    n536,
    n558,
    n551
  );


  buf
  g1011
  (
    n1050,
    n935
  );


  not
  g1012
  (
    n1045,
    n937
  );


  buf
  g1013
  (
    n1043,
    n933
  );


  buf
  g1014
  (
    n1047,
    n938
  );


  buf
  g1015
  (
    n1058,
    n936
  );


  buf
  g1016
  (
    n1056,
    n934
  );


  buf
  g1017
  (
    n1057,
    n931
  );


  buf
  g1018
  (
    n1053,
    n932
  );


  not
  g1019
  (
    n1048,
    n933
  );


  buf
  g1020
  (
    n1054,
    n937
  );


  buf
  g1021
  (
    n1052,
    n936
  );


  buf
  g1022
  (
    n1055,
    n932
  );


  not
  g1023
  (
    n1046,
    n934
  );


  buf
  g1024
  (
    n1049,
    n935
  );


  buf
  g1025
  (
    n1044,
    n938
  );


  not
  g1026
  (
    n1051,
    n931
  );


  not
  g1027
  (
    n1060,
    n1048
  );


  buf
  g1028
  (
    n1061,
    n1054
  );


  buf
  g1029
  (
    n1072,
    n1053
  );


  buf
  g1030
  (
    n1065,
    n1044
  );


  buf
  g1031
  (
    n1068,
    n1048
  );


  not
  g1032
  (
    n1073,
    n1053
  );


  xnor
  g1033
  (
    n1076,
    n1049,
    n1044
  );


  xor
  g1034
  (
    n1070,
    n1043,
    n1050,
    n1051,
    n1055
  );


  and
  g1035
  (
    n1064,
    n1046,
    n1044,
    n1056,
    n1054
  );


  xor
  g1036
  (
    n1075,
    n1048,
    n1053,
    n1052,
    n1043
  );


  or
  g1037
  (
    n1067,
    n1057,
    n1057,
    n1056,
    n1049
  );


  xor
  g1038
  (
    n1062,
    n1047,
    n1046,
    n1043,
    n1051
  );


  or
  g1039
  (
    n1077,
    n1052,
    n1047,
    n1054,
    n1050
  );


  xor
  g1040
  (
    n1063,
    n1057,
    n1054,
    n1043,
    n1047
  );


  nor
  g1041
  (
    n1074,
    n1049,
    n1045,
    n1055
  );


  nand
  g1042
  (
    n1071,
    n1056,
    n1056,
    n1045,
    n1050
  );


  nand
  g1043
  (
    n1078,
    n1045,
    n1052,
    n1047
  );


  xor
  g1044
  (
    n1066,
    n1055,
    n1050,
    n1049,
    n1051
  );


  and
  g1045
  (
    n1059,
    n1051,
    n1057,
    n1055,
    n1053
  );


  xor
  g1046
  (
    n1069,
    n1048,
    n1046,
    n1044
  );


  or
  g1047
  (
    n1093,
    n1070,
    n1060,
    n1066,
    n1061
  );


  xor
  g1048
  (
    n1090,
    n1060,
    n1062,
    n1065,
    n1072
  );


  xnor
  g1049
  (
    n1083,
    n1071,
    n1065,
    n1073,
    n1064
  );


  or
  g1050
  (
    n1084,
    n1063,
    n1061,
    n1074,
    n1073
  );


  xor
  g1051
  (
    n1079,
    n1065,
    n1067,
    n1063,
    n1059
  );


  nand
  g1052
  (
    n1085,
    n1064,
    n1066,
    n1062
  );


  or
  g1053
  (
    n1088,
    n1073,
    n1074,
    n1068,
    n1069
  );


  nand
  g1054
  (
    n1087,
    n1062,
    n1073,
    n1064,
    n1063
  );


  xnor
  g1055
  (
    n1092,
    n1071,
    n1069,
    n1061,
    n1062
  );


  and
  g1056
  (
    n1094,
    n1068,
    n1059
  );


  and
  g1057
  (
    n1081,
    n1070,
    n1072,
    n1068,
    n1069
  );


  and
  g1058
  (
    n1080,
    n1061,
    n1072,
    n1070,
    n1064
  );


  or
  g1059
  (
    n1089,
    n1071,
    n1074,
    n1069,
    n1060
  );


  xnor
  g1060
  (
    n1091,
    n1067,
    n1072,
    n1071,
    n1066
  );


  xor
  g1061
  (
    n1086,
    n1059,
    n1074,
    n1067,
    n1070
  );


  and
  g1062
  (
    n1082,
    n1063,
    n1060,
    n1067,
    n1065
  );


  not
  g1063
  (
    n1105,
    n1082
  );


  buf
  g1064
  (
    n1103,
    n1081
  );


  buf
  g1065
  (
    n1099,
    n1079
  );


  not
  g1066
  (
    n1095,
    n1079
  );


  buf
  g1067
  (
    n1102,
    n1081
  );


  buf
  g1068
  (
    n1109,
    n1079
  );


  buf
  g1069
  (
    n1110,
    n1081
  );


  buf
  g1070
  (
    n1097,
    n1080
  );


  not
  g1071
  (
    n1100,
    n1080
  );


  not
  g1072
  (
    n1096,
    n1082
  );


  buf
  g1073
  (
    n1108,
    n1081
  );


  not
  g1074
  (
    n1106,
    n1080
  );


  buf
  g1075
  (
    n1098,
    n1082
  );


  not
  g1076
  (
    n1101,
    n1082
  );


  buf
  g1077
  (
    n1107,
    n1079
  );


  not
  g1078
  (
    n1104,
    n1080
  );


  nor
  g1079
  (
    n1137,
    n1096,
    n956,
    n958,
    n959
  );


  xor
  g1080
  (
    n1111,
    n1109,
    n1110,
    n939,
    n941
  );


  xnor
  g1081
  (
    n1117,
    n946,
    n948,
    n954,
    n956
  );


  nor
  g1082
  (
    n1136,
    n1098,
    n940,
    n953,
    n943
  );


  xor
  g1083
  (
    n1116,
    n1099,
    n1098,
    n1102,
    n956
  );


  and
  g1084
  (
    n1123,
    n1104,
    n1095,
    n1096,
    n957
  );


  nor
  g1085
  (
    n1112,
    n1096,
    n955,
    n1109,
    n1102
  );


  xor
  g1086
  (
    n1114,
    n959,
    n945,
    n1103,
    n940
  );


  nand
  g1087
  (
    n1131,
    n1108,
    n1106,
    n1110,
    n950
  );


  or
  g1088
  (
    n1118,
    n952,
    n1105,
    n962,
    n961
  );


  and
  g1089
  (
    n1113,
    n1104,
    n958,
    n939,
    n1101
  );


  xnor
  g1090
  (
    n1120,
    n1104,
    n942,
    n947,
    n1103
  );


  or
  g1091
  (
    n1126,
    n947,
    n957,
    n958,
    n949
  );


  or
  g1092
  (
    KeyWire_0_31,
    n1103,
    n1101,
    n1099,
    n1110
  );


  xor
  g1093
  (
    n1139,
    n1108,
    n1106,
    n1107
  );


  nand
  g1094
  (
    n1115,
    n944,
    n952,
    n951,
    n961
  );


  nor
  g1095
  (
    n1121,
    n962,
    n950,
    n1097,
    n948
  );


  xnor
  g1096
  (
    n1135,
    n1100,
    n962,
    n1095,
    n954
  );


  and
  g1097
  (
    n1128,
    n1100,
    n1100,
    n1099,
    n960
  );


  xor
  g1098
  (
    n1119,
    n1108,
    n943,
    n942,
    n951
  );


  xnor
  g1099
  (
    n1140,
    n1097,
    n1107,
    n949,
    n957
  );


  or
  g1100
  (
    n1125,
    n1104,
    n1108,
    n959,
    n1095
  );


  nand
  g1101
  (
    n1127,
    n1098,
    n960,
    n1102
  );


  nand
  g1102
  (
    n1129,
    n946,
    n1097,
    n1106,
    n1107
  );


  xor
  g1103
  (
    n1132,
    n1099,
    n1105,
    n954,
    n1109
  );


  nand
  g1104
  (
    n1130,
    n1097,
    n1103,
    n1110,
    n961
  );


  xnor
  g1105
  (
    n1138,
    n955,
    n1102,
    n1101,
    n941
  );


  nand
  g1106
  (
    n1134,
    n1105,
    n1109,
    n1101,
    n1100
  );


  xor
  g1107
  (
    n1122,
    n945,
    n1106,
    n1098,
    n944
  );


  and
  g1108
  (
    n1133,
    n955,
    n1105,
    n953,
    n963
  );


  xnor
  g1109
  (
    n1141,
    n1133,
    n836,
    n1139,
    n1134
  );


  xnor
  g1110
  (
    n1148,
    n1129,
    n834,
    n1117,
    n1130
  );


  nand
  g1111
  (
    n1151,
    n1131,
    n1126,
    n1140,
    n1118
  );


  xnor
  g1112
  (
    n1150,
    n1134,
    n1140,
    n1138,
    n1124
  );


  nor
  g1113
  (
    n1147,
    n1131,
    n1123,
    n1124,
    n1122
  );


  and
  g1114
  (
    n1153,
    n1137,
    n1138,
    n1125,
    n1119
  );


  xor
  g1115
  (
    n1142,
    n1139,
    n836,
    n1115,
    n1130
  );


  xor
  g1116
  (
    n1143,
    n834,
    n1123,
    n1136,
    n1128
  );


  nor
  g1117
  (
    n1146,
    n1135,
    n835,
    n1127
  );


  xnor
  g1118
  (
    n1144,
    n1120,
    n1133,
    n1136,
    n1111
  );


  and
  g1119
  (
    n1152,
    n1121,
    n1127,
    n1112,
    n1137
  );


  and
  g1120
  (
    n1154,
    n1132,
    n1114,
    n1125,
    n1113
  );


  nor
  g1121
  (
    n1145,
    n1128,
    n833,
    n1129,
    n837
  );


  xor
  g1122
  (
    n1149,
    n1126,
    n1132,
    n1135,
    n1116
  );


  or
  g1123
  (
    n1159,
    n965,
    n965,
    n964,
    n1144
  );


  xor
  g1124
  (
    n1160,
    n1148,
    n1153,
    n1152,
    n1151
  );


  xor
  g1125
  (
    n1161,
    n1143,
    n965,
    n1145,
    n1142
  );


  xnor
  g1126
  (
    n1157,
    n967,
    n1149,
    n1147,
    n966
  );


  xnor
  g1127
  (
    n1155,
    n1146,
    n964,
    n967,
    n1150
  );


  nand
  g1128
  (
    n1156,
    n966,
    n1154,
    n963,
    n964
  );


  xor
  g1129
  (
    n1158,
    n967,
    n966,
    n963,
    n1141
  );


  not
  g1130
  (
    n1163,
    n1083
  );


  nor
  g1131
  (
    n1162,
    n1160,
    n969,
    n1087,
    n1086
  );


  xnor
  g1132
  (
    n1170,
    n1084,
    n969,
    n1158,
    n1160
  );


  xor
  g1133
  (
    n1172,
    n1155,
    n968,
    n1161,
    n1088
  );


  nand
  g1134
  (
    n1169,
    n1161,
    n968,
    n576,
    n1085
  );


  or
  g1135
  (
    n1171,
    n1083,
    n1159,
    n969
  );


  nand
  g1136
  (
    n1173,
    n1088,
    n1085,
    n1083
  );


  or
  g1137
  (
    n1175,
    n1087,
    n1156,
    n970
  );


  xor
  g1138
  (
    n1164,
    n1087,
    n1157,
    n1084,
    n1058
  );


  or
  g1139
  (
    n1168,
    n1058,
    n1084,
    n1085,
    n1086
  );


  nor
  g1140
  (
    n1167,
    n1087,
    n1158,
    n576,
    n1084
  );


  nand
  g1141
  (
    n1166,
    n1088,
    n1156,
    n968,
    n1058
  );


  or
  g1142
  (
    n1165,
    n1088,
    n1161,
    n1058,
    n1155
  );


  and
  g1143
  (
    n1174,
    n1086,
    n1086,
    n1157,
    n1083
  );


  not
  g1144
  (
    n1181,
    n1162
  );


  buf
  g1145
  (
    n1178,
    n1165
  );


  not
  g1146
  (
    n1180,
    n1162
  );


  not
  g1147
  (
    n1184,
    n1167
  );


  not
  g1148
  (
    n1179,
    n1164
  );


  not
  g1149
  (
    n1176,
    n1168
  );


  buf
  g1150
  (
    n1183,
    n1166
  );


  buf
  g1151
  (
    n1177,
    n1164
  );


  and
  g1152
  (
    n1182,
    n1167,
    n1166,
    n1169,
    n1165
  );


  nor
  g1153
  (
    n1185,
    n1169,
    n1168,
    n1163
  );


  and
  g1154
  (
    n1189,
    n1177,
    n1176,
    n1183,
    n1179
  );


  xor
  g1155
  (
    n1188,
    n1181,
    n1182,
    n1184
  );


  xnor
  g1156
  (
    n1186,
    n1183,
    n1181,
    n1177,
    n1178
  );


  nor
  g1157
  (
    n1187,
    n1178,
    n1180,
    n1179
  );


  buf
  g1158
  (
    n1197,
    n1187
  );


  buf
  g1159
  (
    n1193,
    n1189
  );


  buf
  g1160
  (
    n1191,
    n1187
  );


  not
  g1161
  (
    n1194,
    n1188
  );


  nand
  g1162
  (
    n1196,
    n1188,
    n1186
  );


  xor
  g1163
  (
    n1195,
    n970,
    n1189
  );


  nand
  g1164
  (
    n1192,
    n1187,
    n1186,
    n1188
  );


  and
  g1165
  (
    n1190,
    n971,
    n1188,
    n1189
  );


  nand
  g1166
  (
    n1203,
    n1194,
    n1195,
    n842,
    n1190
  );


  xor
  g1167
  (
    n1198,
    n843,
    n844,
    n972,
    n839
  );


  and
  g1168
  (
    n1199,
    n971,
    n973,
    n1197,
    n972
  );


  xnor
  g1169
  (
    n1205,
    n973,
    n840,
    n843
  );


  nand
  g1170
  (
    n1202,
    n1196,
    n841,
    n972,
    n973
  );


  or
  g1171
  (
    n1204,
    n838,
    n838,
    n837,
    n1193
  );


  xor
  g1172
  (
    n1200,
    n1191,
    n1192,
    n845,
    n839
  );


  and
  g1173
  (
    n1201,
    n844,
    n842,
    n841,
    n971
  );


  or
  g1174
  (
    n1215,
    n1200,
    n978,
    n975,
    n1199
  );


  and
  g1175
  (
    n1225,
    n975,
    n1173,
    n1089
  );


  nand
  g1176
  (
    n1208,
    n1090,
    n976,
    n1076,
    n1204
  );


  and
  g1177
  (
    n1216,
    n1172,
    n1200,
    n1205,
    n1090
  );


  and
  g1178
  (
    n1218,
    n852,
    n1170,
    n1198,
    n1200
  );


  xor
  g1179
  (
    n1207,
    n848,
    n1171,
    n1075,
    n850
  );


  xor
  g1180
  (
    n1210,
    n1205,
    n1198,
    n1203,
    n1204
  );


  or
  g1181
  (
    n1228,
    n1202,
    n847,
    n1090,
    n851
  );


  nor
  g1182
  (
    n1224,
    n1199,
    n1203,
    n1172,
    n846
  );


  nand
  g1183
  (
    n1221,
    n1078,
    n1078,
    n852,
    n850
  );


  and
  g1184
  (
    n1222,
    n847,
    n1205,
    n848,
    n1202
  );


  and
  g1185
  (
    n1206,
    n849,
    n978,
    n1089,
    n979
  );


  xor
  g1186
  (
    n1213,
    n1201,
    n1077,
    n851
  );


  nand
  g1187
  (
    n1223,
    n1078,
    n845,
    n1201,
    n1199
  );


  xnor
  g1188
  (
    n1211,
    n1202,
    n849,
    n1201,
    n1077
  );


  xnor
  g1189
  (
    n1229,
    n1202,
    n1076,
    n1205,
    n1075
  );


  and
  g1190
  (
    n1214,
    n978,
    n976,
    n1089,
    n1203
  );


  and
  g1191
  (
    n1212,
    n1203,
    n1200,
    n976,
    n1201
  );


  nor
  g1192
  (
    n1217,
    n977,
    n974,
    n1199,
    n1075
  );


  and
  g1193
  (
    n1227,
    n974,
    n1204,
    n978,
    n977
  );


  and
  g1194
  (
    n1226,
    n1170,
    n1076,
    n1204
  );


  xor
  g1195
  (
    n1219,
    n1171,
    n1075,
    n1077,
    n846
  );


  nand
  g1196
  (
    n1209,
    n1089,
    n977,
    n1090,
    n1198
  );


  nor
  g1197
  (
    n1220,
    n975,
    n1198,
    n974,
    n1078
  );


  xnor
  g1198
  (
    n1293,
    n997,
    n1018,
    n1006,
    n1223
  );


  or
  g1199
  (
    n1242,
    n1013,
    n1007,
    n1218,
    n979
  );


  xnor
  g1200
  (
    n1299,
    n979,
    n993,
    n1011,
    n1215
  );


  xor
  g1201
  (
    n1256,
    n983,
    n998,
    n1210,
    n1206
  );


  nand
  g1202
  (
    n1286,
    n1228,
    n1032,
    n1026,
    n1018
  );


  nand
  g1203
  (
    n1235,
    n990,
    n1216,
    n987,
    n981
  );


  nand
  g1204
  (
    n1245,
    n986,
    n1009,
    n154,
    n987
  );


  nand
  g1205
  (
    KeyWire_0_15,
    n1007,
    n1208,
    n154,
    n981
  );


  and
  g1206
  (
    n1272,
    n990,
    n152,
    n1031,
    n1221
  );


  or
  g1207
  (
    n1306,
    n1215,
    n1024,
    n1000,
    n1028
  );


  xnor
  g1208
  (
    n1249,
    n1225,
    n1214,
    n980,
    n1028
  );


  nor
  g1209
  (
    n1304,
    n1222,
    n1006,
    n1022,
    n1219
  );


  nor
  g1210
  (
    n1284,
    n1223,
    n1014,
    n988,
    n1013
  );


  and
  g1211
  (
    n1311,
    n1030,
    n1227,
    n1021,
    n999
  );


  xnor
  g1212
  (
    n1240,
    n1217,
    n1223,
    n1006,
    n1218
  );


  xnor
  g1213
  (
    n1310,
    n1023,
    n1219,
    n1227,
    n1006
  );


  nor
  g1214
  (
    n1232,
    n1207,
    n1212,
    n1213,
    n1024
  );


  or
  g1215
  (
    n1263,
    n1010,
    n1210,
    n1014,
    n1216
  );


  and
  g1216
  (
    n1257,
    n1217,
    n1020,
    n997,
    n154
  );


  and
  g1217
  (
    n1296,
    n983,
    n1016,
    n1213,
    n1029
  );


  and
  g1218
  (
    n1271,
    n1218,
    n1030,
    n1013,
    n994
  );


  nor
  g1219
  (
    n1231,
    n1010,
    n1229,
    n1018,
    n1022
  );


  xor
  g1220
  (
    n1307,
    n1220,
    n988,
    n991
  );


  or
  g1221
  (
    n1251,
    n1023,
    n1225,
    n1017,
    n993
  );


  nand
  g1222
  (
    n1241,
    n1032,
    n1216,
    n1011
  );


  nor
  g1223
  (
    n1267,
    n1013,
    n1005,
    n1211,
    n1030
  );


  nor
  g1224
  (
    n1280,
    n1021,
    n990,
    n1004,
    n1026
  );


  nor
  g1225
  (
    n1278,
    n1207,
    n982,
    n1008,
    n984
  );


  nor
  g1226
  (
    n1260,
    n1213,
    n1214,
    n1024,
    n1032
  );


  nor
  g1227
  (
    n1301,
    n984,
    n1022,
    n1212,
    n1211
  );


  and
  g1228
  (
    n1233,
    n982,
    n998,
    n1033,
    n1023
  );


  xor
  g1229
  (
    n1253,
    n1025,
    n992,
    n996,
    n998
  );


  or
  g1230
  (
    n1289,
    n1017,
    n988,
    n982,
    n1031
  );


  or
  g1231
  (
    n1236,
    n1222,
    n1003,
    n1027,
    n991
  );


  xor
  g1232
  (
    n1277,
    n1008,
    n1021,
    n995,
    n1025
  );


  and
  g1233
  (
    n1302,
    n1015,
    n990,
    n1009,
    n1029
  );


  and
  g1234
  (
    n1287,
    n1028,
    n1009,
    n1209,
    n1031
  );


  and
  g1235
  (
    n1292,
    n1008,
    n1213,
    n153,
    n992
  );


  and
  g1236
  (
    n1230,
    n989,
    n991,
    n1025,
    n1005
  );


  nor
  g1237
  (
    n1308,
    n1001,
    n1033,
    n989,
    n1019
  );


  nand
  g1238
  (
    n1276,
    n1224,
    n1027,
    n1219,
    n1209
  );


  or
  g1239
  (
    n1261,
    n986,
    n1207,
    n152,
    n1004
  );


  nand
  g1240
  (
    n1294,
    n1018,
    n1003,
    n988,
    n1002
  );


  xor
  g1241
  (
    n1275,
    n1227,
    n989,
    n1031,
    n985
  );


  and
  g1242
  (
    n1274,
    n1034,
    n1002,
    n1212,
    n1209
  );


  and
  g1243
  (
    n1266,
    n1026,
    n1028,
    n993,
    n982
  );


  nand
  g1244
  (
    n1244,
    n996,
    n1016,
    n1218,
    n1227
  );


  nand
  g1245
  (
    n1262,
    n1005,
    n985,
    n998,
    n1225
  );


  or
  g1246
  (
    n1234,
    n1001,
    n1010,
    n1229,
    n1228
  );


  xnor
  g1247
  (
    n1298,
    n1002,
    n1221,
    n1034,
    n1014
  );


  nor
  g1248
  (
    n1259,
    n1208,
    n1011,
    n1026,
    n1220
  );


  or
  g1249
  (
    n1297,
    n1016,
    n1229,
    n1224,
    n987
  );


  nand
  g1250
  (
    n1264,
    n999,
    n1030,
    n1000,
    n1017
  );


  nor
  g1251
  (
    n1300,
    n1214,
    n1209,
    n1221,
    n999
  );


  and
  g1252
  (
    n1237,
    n1210,
    n1020,
    n1208,
    n1029
  );


  or
  g1253
  (
    n1243,
    n981,
    n995,
    n980,
    n997
  );


  and
  g1254
  (
    n1290,
    n1207,
    n992,
    n980,
    n1023
  );


  and
  g1255
  (
    n1258,
    n1215,
    n1027,
    n1000,
    n1009
  );


  or
  g1256
  (
    n1254,
    n1029,
    n1007,
    n1220,
    n1226
  );


  or
  g1257
  (
    n1295,
    n1020,
    n994,
    n153,
    n1004
  );


  and
  g1258
  (
    n1248,
    n1229,
    n1215,
    n1024,
    n1033
  );


  and
  g1259
  (
    n1270,
    n1217,
    n979,
    n1021,
    n1001
  );


  xnor
  g1260
  (
    n1283,
    n1206,
    n981,
    n1210,
    n1217
  );


  and
  g1261
  (
    n1303,
    n1003,
    n1007,
    n1225,
    n1010
  );


  xnor
  g1262
  (
    n1238,
    n1015,
    n985,
    n1000
  );


  or
  g1263
  (
    n1291,
    n1015,
    n1012,
    n992,
    n999
  );


  nand
  g1264
  (
    n1281,
    n1022,
    n1034,
    n1224,
    n1219
  );


  nor
  g1265
  (
    n1239,
    n983,
    n1017,
    n1206,
    n153
  );


  xor
  g1266
  (
    n1255,
    n1228,
    n1011,
    n1002,
    n1211
  );


  xor
  g1267
  (
    n1250,
    n1008,
    n1220,
    n153,
    n1020
  );


  nor
  g1268
  (
    n1282,
    n997,
    n1003,
    n980,
    n1226
  );


  or
  g1269
  (
    n1252,
    n1226,
    n1033,
    n1019,
    n1222
  );


  nand
  g1270
  (
    n1285,
    n1214,
    n1224,
    n987,
    n984
  );


  xor
  g1271
  (
    n1247,
    n1012,
    n1211,
    n986,
    n984
  );


  xor
  g1272
  (
    n1269,
    n1019,
    n1012,
    n1025,
    n1004
  );


  xnor
  g1273
  (
    n1246,
    n1206,
    n1221,
    n995,
    n1222
  );


  xnor
  g1274
  (
    n1273,
    n1208,
    n996,
    n983,
    n1027
  );


  nand
  g1275
  (
    n1305,
    n1001,
    n986,
    n1014,
    n1019
  );


  nor
  g1276
  (
    n1288,
    n1226,
    n989,
    n996,
    n1212
  );


  nor
  g1277
  (
    n1309,
    n1015,
    n1223,
    n995,
    n994
  );


  nor
  g1278
  (
    n1265,
    n994,
    n152,
    n1032,
    n1016
  );


  nor
  g1279
  (
    n1268,
    n1012,
    n1005,
    n993,
    n1228
  );


  not
  g1280
  (
    n1316,
    n1233
  );


  not
  g1281
  (
    n1317,
    n1238
  );


  not
  g1282
  (
    n1315,
    n1232
  );


  and
  g1283
  (
    n1313,
    n1231,
    n1239,
    n1240
  );


  or
  g1284
  (
    n1314,
    n1236,
    n1230,
    n1237
  );


  xor
  g1285
  (
    n1312,
    n1241,
    n1235,
    n1234
  );


  xnor
  g1286
  (
    n1318,
    n1314,
    n1316,
    n1315,
    n1313
  );


  xnor
  g1287
  (
    n1321,
    n855,
    n854,
    n857
  );


  and
  g1288
  (
    n1320,
    n853,
    n855,
    n1318,
    n856
  );


  or
  g1289
  (
    n1319,
    n856,
    n1318,
    n853
  );


  xnor
  g1290
  (
    n1323,
    n858,
    n858,
    n857,
    n1321
  );


  nand
  g1291
  (
    n1322,
    n885,
    n1320,
    n859
  );


  not
  g1292
  (
    n1328,
    n860
  );


  not
  g1293
  (
    n1327,
    n1323
  );


  nor
  g1294
  (
    n1326,
    n1322,
    n860
  );


  or
  g1295
  (
    n1324,
    n1243,
    n861,
    n862
  );


  nand
  g1296
  (
    n1329,
    n1244,
    n1323
  );


  nand
  g1297
  (
    n1325,
    n1322,
    n1242,
    n862,
    n863
  );


  xnor
  g1298
  (
    n1334,
    n869,
    n1175,
    n1326,
    n1037
  );


  xnor
  g1299
  (
    KeyWire_0_5,
    n869,
    n1094,
    n863,
    n1329
  );


  or
  g1300
  (
    n1348,
    n1038,
    n1324,
    n1036,
    n1035
  );


  xor
  g1301
  (
    n1333,
    n1328,
    n1324,
    n1326,
    n1037
  );


  xor
  g1302
  (
    n1342,
    n867,
    n871,
    n1174,
    n1035
  );


  xor
  g1303
  (
    n1349,
    n1091,
    n870,
    n1094,
    n1327
  );


  xor
  g1304
  (
    n1339,
    n866,
    n865,
    n1091
  );


  nor
  g1305
  (
    n1343,
    n1328,
    n1094,
    n865,
    n1092
  );


  nand
  g1306
  (
    n1330,
    n1327,
    n1174,
    n1324,
    n1091
  );


  and
  g1307
  (
    n1337,
    n1185,
    n1185,
    n864,
    n1034
  );


  xnor
  g1308
  (
    n1335,
    n1175,
    n1036,
    n1326,
    n1324
  );


  xor
  g1309
  (
    n1340,
    n1037,
    n1329,
    n1094,
    n1326
  );


  nand
  g1310
  (
    n1332,
    n1327,
    n1093,
    n1036
  );


  xnor
  g1311
  (
    n1345,
    n870,
    n866,
    n1093,
    n868
  );


  and
  g1312
  (
    n1338,
    n1035,
    n1092,
    n864,
    n1329
  );


  xnor
  g1313
  (
    n1336,
    n1325,
    n1327,
    n1184,
    n1093
  );


  nand
  g1314
  (
    n1331,
    n1317,
    n1035,
    n1092,
    n1325
  );


  and
  g1315
  (
    n1347,
    n1328,
    n1328,
    n1092,
    n1175
  );


  nand
  g1316
  (
    KeyWire_0_3,
    n1037,
    n1325,
    n1036
  );


  xor
  g1317
  (
    n1344,
    n1329,
    n868,
    n867,
    n1038
  );


  nor
  g1318
  (
    n1372,
    n1332,
    n1273,
    n1330,
    n1341
  );


  and
  g1319
  (
    n1361,
    n1346,
    n1310,
    n1255,
    n1348
  );


  or
  g1320
  (
    n1379,
    n1254,
    n1348,
    n1295,
    n1266
  );


  xor
  g1321
  (
    n1358,
    n1249,
    n1348,
    n1299,
    n1349
  );


  xor
  g1322
  (
    n1373,
    n155,
    n155,
    n1253,
    n1248
  );


  and
  g1323
  (
    n1362,
    n1311,
    n1291,
    n1257,
    n1247
  );


  nand
  g1324
  (
    n1376,
    n1284,
    n1301,
    n1331,
    n1280
  );


  xor
  g1325
  (
    n1378,
    n1348,
    n1300,
    n1306,
    n1279
  );


  or
  g1326
  (
    n1357,
    n1343,
    n1334,
    n1272,
    n1285
  );


  or
  g1327
  (
    n1366,
    n1332,
    n1245,
    n1267,
    n1333
  );


  xnor
  g1328
  (
    n1371,
    n1343,
    n1263,
    n1337,
    n1344
  );


  or
  g1329
  (
    n1355,
    n1345,
    n1341,
    n1278,
    n1305
  );


  and
  g1330
  (
    n1377,
    n1336,
    n1270,
    n1333,
    n1338
  );


  xnor
  g1331
  (
    n1356,
    n1275,
    n1262,
    n1271,
    n1261
  );


  and
  g1332
  (
    n1352,
    n1290,
    n1256,
    n1277,
    n1298
  );


  xor
  g1333
  (
    n1351,
    n1308,
    n1251,
    n1260,
    n1265
  );


  nand
  g1334
  (
    n1375,
    n1347,
    n1264,
    n1346,
    n1340
  );


  or
  g1335
  (
    n1370,
    n154,
    n1338,
    n1342,
    n1281
  );


  nor
  g1336
  (
    n1368,
    n1347,
    n1335,
    n1269
  );


  nor
  g1337
  (
    n1359,
    n1246,
    n1288,
    n1292,
    n1304
  );


  nor
  g1338
  (
    n1363,
    n1349,
    n1345,
    n1294,
    n155
  );


  nor
  g1339
  (
    n1354,
    n1336,
    n1282,
    n1289,
    n1259
  );


  xnor
  g1340
  (
    n1353,
    n1340,
    n1337,
    n1349,
    n1344
  );


  xor
  g1341
  (
    n1360,
    n1334,
    n1330,
    n1286,
    n1258
  );


  or
  g1342
  (
    n1364,
    n1302,
    n1342,
    n1331,
    n1346
  );


  nor
  g1343
  (
    n1350,
    n155,
    n1347,
    n1293,
    n1283
  );


  xor
  g1344
  (
    n1374,
    n1274,
    n1347,
    n1307,
    n1287
  );


  xor
  g1345
  (
    n1369,
    n1346,
    n1303,
    n1296,
    n1349
  );


  xor
  g1346
  (
    n1365,
    n1339,
    n1252,
    n1268,
    n1250
  );


  or
  g1347
  (
    n1367,
    n1339,
    n1309,
    n1297,
    n1276
  );


  buf
  g1348
  (
    n1382,
    n1353
  );


  not
  g1349
  (
    n1381,
    n1354
  );


  buf
  g1350
  (
    n1384,
    n1350
  );


  buf
  g1351
  (
    n1380,
    n1351
  );


  buf
  g1352
  (
    n1383,
    n1352
  );


  xor
  g1353
  (
    n1386,
    n1381,
    n576,
    n1382,
    n1384
  );


  or
  g1354
  (
    n1385,
    n577,
    n577,
    n576,
    n1383
  );


  not
  g1355
  (
    n1390,
    n1386
  );


  not
  g1356
  (
    n1389,
    n1385
  );


  not
  g1357
  (
    n1387,
    n1386
  );


  buf
  g1358
  (
    n1388,
    n1385
  );


  and
  g1359
  (
    n1391,
    n1388,
    n1387,
    n1389
  );


  and
  g1360
  (
    n1392,
    n1388,
    n871,
    n1390
  );


  nand
  g1361
  (
    n1393,
    n577,
    n577,
    n1392,
    n1391
  );


  buf
  g1362
  (
    n1394,
    n1393
  );


  and
  g1363
  (
    n1395,
    n873,
    n872,
    n1394
  );


  xnor
  g1364
  (
    n1396,
    n872,
    n872,
    n873,
    n1394
  );


  or
  g1365
  (
    n1402,
    n885,
    n1396,
    n1362,
    n1395
  );


  nor
  g1366
  (
    n1397,
    n886,
    n1395,
    n1358,
    n1396
  );


  nor
  g1367
  (
    n1398,
    n1039,
    n1359,
    n1038,
    n1040
  );


  nor
  g1368
  (
    n1401,
    n1040,
    n1039,
    n885,
    n1356
  );


  xor
  g1369
  (
    n1399,
    n886,
    n1355,
    n885,
    n1039
  );


  and
  g1370
  (
    n1403,
    n1396,
    n886,
    n1040,
    n1357
  );


  xnor
  g1371
  (
    n1404,
    n886,
    n1396,
    n1360,
    n1361
  );


  nor
  g1372
  (
    n1400,
    n1038,
    n1395,
    n1039
  );


  nand
  g1373
  (
    n1416,
    n874,
    n1401,
    n875,
    n1371
  );


  or
  g1374
  (
    n1414,
    n1369,
    n873,
    n875,
    n876
  );


  and
  g1375
  (
    n1406,
    n1377,
    n875,
    n1042,
    n873
  );


  and
  g1376
  (
    n1408,
    n1399,
    n1376,
    n1041,
    n1042
  );


  or
  g1377
  (
    n1409,
    n1041,
    n876,
    n1399,
    n1379
  );


  and
  g1378
  (
    n1413,
    n1400,
    n1403,
    n1404,
    n1372
  );


  xnor
  g1379
  (
    n1412,
    n874,
    n1041,
    n1367,
    n1374
  );


  nor
  g1380
  (
    n1405,
    n1364,
    n1403,
    n1040,
    n875
  );


  nor
  g1381
  (
    n1407,
    n1373,
    n1042,
    n1400,
    n1366
  );


  xor
  g1382
  (
    n1418,
    n1397,
    n1401,
    n1370,
    n1365
  );


  xnor
  g1383
  (
    n1415,
    n1398,
    n874,
    n876
  );


  nor
  g1384
  (
    n1417,
    n1042,
    n1368,
    n1363,
    n1398
  );


  nor
  g1385
  (
    n1411,
    n1375,
    n1402,
    n1041
  );


  xnor
  g1386
  (
    n1410,
    n1404,
    n876,
    n1397,
    n1378
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n724,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n560,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n472,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1346,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n890,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1341,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n702,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n273,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n120,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n237,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n63,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n219,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n588,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n328,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n775,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1279,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n738,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n302,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n309,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n828,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n205,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n841,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n908,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n52,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n374,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n753,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n415,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n185,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n491,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n602,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n572,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1124,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

