

module Stat_1071_333
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n45,
  n46,
  n47,
  n48,
  n49,
  n50,
  n51,
  n52,
  n358,
  n361,
  n340,
  n360,
  n355,
  n345,
  n338,
  n362,
  n356,
  n335,
  n353,
  n359,
  n354,
  n1004,
  n1070,
  n1059,
  n1056,
  n1053,
  n1060,
  n1062,
  n1057,
  n1052,
  n1071,
  n1072,
  n1058,
  n1055,
  n1073,
  n1065,
  n1061,
  n1074,
  n1063,
  n1114,
  n1092,
  n1093,
  n1107,
  n1102,
  n1113,
  n1105,
  n1120,
  n1094,
  n1121,
  n1098,
  n1104,
  n1116,
  n1101,
  n1112,
  n1119,
  n1097,
  n1118,
  n1110,
  n1103,
  n1095,
  n1123,
  n1100,
  n1117,
  n1111,
  n1109,
  n1099,
  n1096,
  n1106,
  n1115,
  n1108,
  n1122,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63,
  keyIn_0_64,
  keyIn_0_65,
  keyIn_0_66,
  keyIn_0_67,
  keyIn_0_68,
  keyIn_0_69,
  keyIn_0_70,
  keyIn_0_71,
  keyIn_0_72,
  keyIn_0_73,
  keyIn_0_74,
  keyIn_0_75,
  keyIn_0_76,
  keyIn_0_77,
  keyIn_0_78,
  keyIn_0_79,
  keyIn_0_80,
  keyIn_0_81,
  keyIn_0_82,
  keyIn_0_83,
  keyIn_0_84,
  keyIn_0_85,
  keyIn_0_86,
  keyIn_0_87,
  keyIn_0_88,
  keyIn_0_89,
  keyIn_0_90,
  keyIn_0_91,
  keyIn_0_92,
  keyIn_0_93,
  keyIn_0_94,
  keyIn_0_95,
  keyIn_0_96,
  keyIn_0_97,
  keyIn_0_98,
  keyIn_0_99,
  keyIn_0_100,
  keyIn_0_101,
  keyIn_0_102,
  keyIn_0_103
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input n40;input n41;input n42;input n43;input n44;input n45;input n46;input n47;input n48;input n49;input n50;input n51;input n52;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;input keyIn_0_64;input keyIn_0_65;input keyIn_0_66;input keyIn_0_67;input keyIn_0_68;input keyIn_0_69;input keyIn_0_70;input keyIn_0_71;input keyIn_0_72;input keyIn_0_73;input keyIn_0_74;input keyIn_0_75;input keyIn_0_76;input keyIn_0_77;input keyIn_0_78;input keyIn_0_79;input keyIn_0_80;input keyIn_0_81;input keyIn_0_82;input keyIn_0_83;input keyIn_0_84;input keyIn_0_85;input keyIn_0_86;input keyIn_0_87;input keyIn_0_88;input keyIn_0_89;input keyIn_0_90;input keyIn_0_91;input keyIn_0_92;input keyIn_0_93;input keyIn_0_94;input keyIn_0_95;input keyIn_0_96;input keyIn_0_97;input keyIn_0_98;input keyIn_0_99;input keyIn_0_100;input keyIn_0_101;input keyIn_0_102;input keyIn_0_103;
  output n358;output n361;output n340;output n360;output n355;output n345;output n338;output n362;output n356;output n335;output n353;output n359;output n354;output n1004;output n1070;output n1059;output n1056;output n1053;output n1060;output n1062;output n1057;output n1052;output n1071;output n1072;output n1058;output n1055;output n1073;output n1065;output n1061;output n1074;output n1063;output n1114;output n1092;output n1093;output n1107;output n1102;output n1113;output n1105;output n1120;output n1094;output n1121;output n1098;output n1104;output n1116;output n1101;output n1112;output n1119;output n1097;output n1118;output n1110;output n1103;output n1095;output n1123;output n1100;output n1117;output n1111;output n1109;output n1099;output n1096;output n1106;output n1115;output n1108;output n1122;
  wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n336;wire n337;wire n339;wire n341;wire n342;wire n343;wire n344;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n357;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1054;wire n1064;wire n1066;wire n1067;wire n1068;wire n1069;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire g_input_0_32;wire gbar_input_0_32;wire g_input_0_33;wire gbar_input_0_33;wire g_input_0_34;wire gbar_input_0_34;wire g_input_0_35;wire gbar_input_0_35;wire g_input_0_36;wire gbar_input_0_36;wire g_input_0_37;wire gbar_input_0_37;wire g_input_0_38;wire gbar_input_0_38;wire g_input_0_39;wire gbar_input_0_39;wire g_input_0_40;wire gbar_input_0_40;wire g_input_0_41;wire gbar_input_0_41;wire g_input_0_42;wire gbar_input_0_42;wire g_input_0_43;wire gbar_input_0_43;wire g_input_0_44;wire gbar_input_0_44;wire g_input_0_45;wire gbar_input_0_45;wire g_input_0_46;wire gbar_input_0_46;wire g_input_0_47;wire gbar_input_0_47;wire g_input_0_48;wire gbar_input_0_48;wire g_input_0_49;wire gbar_input_0_49;wire g_input_0_50;wire gbar_input_0_50;wire g_input_0_51;wire gbar_input_0_51;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n81,
    n21
  );


  buf
  g1
  (
    n90,
    n34
  );


  not
  g2
  (
    n186,
    n17
  );


  not
  g3
  (
    n131,
    n27
  );


  not
  g4
  (
    n86,
    n43
  );


  buf
  g5
  (
    n75,
    n35
  );


  buf
  g6
  (
    n165,
    n23
  );


  not
  g7
  (
    n118,
    n37
  );


  buf
  g8
  (
    n132,
    n7
  );


  not
  g9
  (
    n217,
    n41
  );


  buf
  g10
  (
    n91,
    n12
  );


  buf
  g11
  (
    n202,
    n15
  );


  buf
  g12
  (
    n181,
    n33
  );


  buf
  g13
  (
    n155,
    n38
  );


  not
  g14
  (
    n211,
    n17
  );


  buf
  g15
  (
    n56,
    n9
  );


  not
  g16
  (
    n218,
    n46
  );


  not
  g17
  (
    n92,
    n28
  );


  not
  g18
  (
    n177,
    n20
  );


  not
  g19
  (
    n68,
    n27
  );


  not
  g20
  (
    n224,
    n22
  );


  not
  g21
  (
    n144,
    n31
  );


  not
  g22
  (
    n72,
    n16
  );


  not
  g23
  (
    n191,
    n12
  );


  not
  g24
  (
    n120,
    n41
  );


  not
  g25
  (
    n114,
    n17
  );


  not
  g26
  (
    n125,
    n22
  );


  not
  g27
  (
    n149,
    n16
  );


  not
  g28
  (
    n195,
    n41
  );


  buf
  g29
  (
    n167,
    n28
  );


  not
  g30
  (
    n89,
    n34
  );


  not
  g31
  (
    n99,
    n9
  );


  buf
  g32
  (
    n200,
    n42
  );


  buf
  g33
  (
    n94,
    n12
  );


  buf
  g34
  (
    n219,
    n29
  );


  not
  g35
  (
    n112,
    n30
  );


  buf
  g36
  (
    n123,
    n13
  );


  buf
  g37
  (
    n192,
    n31
  );


  not
  g38
  (
    n142,
    n4
  );


  not
  g39
  (
    n166,
    n19
  );


  not
  g40
  (
    n203,
    n4
  );


  not
  g41
  (
    n110,
    n5
  );


  not
  g42
  (
    n184,
    n13
  );


  buf
  g43
  (
    n170,
    n23
  );


  buf
  g44
  (
    n182,
    n18
  );


  not
  g45
  (
    n204,
    n32
  );


  not
  g46
  (
    n162,
    n22
  );


  buf
  g47
  (
    n158,
    n40
  );


  not
  g48
  (
    n199,
    n45
  );


  buf
  g49
  (
    n117,
    n23
  );


  not
  g50
  (
    n226,
    n14
  );


  not
  g51
  (
    n212,
    n42
  );


  buf
  g52
  (
    n65,
    n44
  );


  not
  g53
  (
    n220,
    n35
  );


  buf
  g54
  (
    n208,
    n28
  );


  not
  g55
  (
    n95,
    n47
  );


  not
  g56
  (
    n221,
    n39
  );


  not
  g57
  (
    n126,
    n46
  );


  buf
  g58
  (
    n135,
    n26
  );


  buf
  g59
  (
    n215,
    n18
  );


  buf
  g60
  (
    n105,
    n35
  );


  buf
  g61
  (
    n97,
    n1
  );


  not
  g62
  (
    n148,
    n33
  );


  buf
  g63
  (
    n57,
    n7
  );


  not
  g64
  (
    n156,
    n3
  );


  buf
  g65
  (
    n185,
    n43
  );


  not
  g66
  (
    n160,
    n7
  );


  buf
  g67
  (
    n150,
    n11
  );


  not
  g68
  (
    n139,
    n38
  );


  not
  g69
  (
    n198,
    n25
  );


  not
  g70
  (
    n61,
    n27
  );


  not
  g71
  (
    n84,
    n46
  );


  buf
  g72
  (
    n128,
    n23
  );


  not
  g73
  (
    n79,
    n31
  );


  not
  g74
  (
    n176,
    n9
  );


  not
  g75
  (
    n67,
    n26
  );


  not
  g76
  (
    n141,
    n14
  );


  buf
  g77
  (
    n136,
    n36
  );


  buf
  g78
  (
    n80,
    n1
  );


  buf
  g79
  (
    n146,
    n22
  );


  not
  g80
  (
    n213,
    n24
  );


  not
  g81
  (
    n122,
    n10
  );


  buf
  g82
  (
    n71,
    n6
  );


  not
  g83
  (
    n133,
    n5
  );


  buf
  g84
  (
    n147,
    n34
  );


  buf
  g85
  (
    n164,
    n40
  );


  buf
  g86
  (
    n154,
    n15
  );


  not
  g87
  (
    n109,
    n39
  );


  buf
  g88
  (
    n77,
    n44
  );


  buf
  g89
  (
    n159,
    n33
  );


  buf
  g90
  (
    n207,
    n16
  );


  not
  g91
  (
    n223,
    n18
  );


  buf
  g92
  (
    n174,
    n40
  );


  buf
  g93
  (
    n124,
    n24
  );


  not
  g94
  (
    n87,
    n36
  );


  buf
  g95
  (
    n60,
    n42
  );


  buf
  g96
  (
    n134,
    n39
  );


  not
  g97
  (
    n111,
    n15
  );


  not
  g98
  (
    n169,
    n3
  );


  buf
  g99
  (
    n93,
    n10
  );


  not
  g100
  (
    n188,
    n18
  );


  not
  g101
  (
    n103,
    n19
  );


  buf
  g102
  (
    n121,
    n20
  );


  not
  g103
  (
    n171,
    n32
  );


  buf
  g104
  (
    n113,
    n29
  );


  buf
  g105
  (
    n64,
    n20
  );


  not
  g106
  (
    n145,
    n6
  );


  buf
  g107
  (
    n173,
    n20
  );


  buf
  g108
  (
    n175,
    n33
  );


  buf
  g109
  (
    n54,
    n8
  );


  buf
  g110
  (
    n201,
    n32
  );


  not
  g111
  (
    n225,
    n10
  );


  not
  g112
  (
    n190,
    n8
  );


  not
  g113
  (
    n197,
    n36
  );


  not
  g114
  (
    n107,
    n37
  );


  buf
  g115
  (
    n62,
    n7
  );


  buf
  g116
  (
    n161,
    n25
  );


  buf
  g117
  (
    n116,
    n44
  );


  buf
  g118
  (
    n83,
    n43
  );


  not
  g119
  (
    n108,
    n40
  );


  not
  g120
  (
    n187,
    n21
  );


  not
  g121
  (
    n88,
    n47
  );


  not
  g122
  (
    n63,
    n31
  );


  not
  g123
  (
    n209,
    n38
  );


  buf
  g124
  (
    n193,
    n45
  );


  buf
  g125
  (
    n101,
    n28
  );


  buf
  g126
  (
    n102,
    n43
  );


  not
  g127
  (
    n82,
    n30
  );


  not
  g128
  (
    n196,
    n11
  );


  buf
  g129
  (
    n153,
    n14
  );


  buf
  g130
  (
    n168,
    n24
  );


  buf
  g131
  (
    n106,
    n16
  );


  not
  g132
  (
    n73,
    n30
  );


  buf
  g133
  (
    n127,
    n45
  );


  buf
  g134
  (
    n157,
    n12
  );


  buf
  g135
  (
    n137,
    n32
  );


  not
  g136
  (
    n172,
    n19
  );


  not
  g137
  (
    n189,
    n13
  );


  buf
  g138
  (
    n138,
    n36
  );


  not
  g139
  (
    n98,
    n21
  );


  buf
  g140
  (
    n163,
    n46
  );


  buf
  g141
  (
    n70,
    n26
  );


  buf
  g142
  (
    n222,
    n25
  );


  not
  g143
  (
    n151,
    n29
  );


  buf
  g144
  (
    n74,
    n41
  );


  buf
  g145
  (
    n69,
    n24
  );


  not
  g146
  (
    n104,
    n2
  );


  buf
  g147
  (
    n119,
    n9
  );


  not
  g148
  (
    n85,
    n10
  );


  not
  g149
  (
    n115,
    n15
  );


  buf
  g150
  (
    n55,
    n2
  );


  buf
  g151
  (
    n205,
    n26
  );


  buf
  g152
  (
    n58,
    n39
  );


  buf
  g153
  (
    n78,
    n14
  );


  not
  g154
  (
    n129,
    n44
  );


  buf
  g155
  (
    n214,
    n8
  );


  buf
  g156
  (
    n53,
    n37
  );


  buf
  g157
  (
    n76,
    n29
  );


  buf
  g158
  (
    n100,
    n11
  );


  buf
  g159
  (
    n210,
    n35
  );


  not
  g160
  (
    n194,
    n19
  );


  buf
  g161
  (
    n66,
    n42
  );


  not
  g162
  (
    n206,
    n25
  );


  not
  g163
  (
    n143,
    n11
  );


  not
  g164
  (
    n152,
    n45
  );


  buf
  g165
  (
    n178,
    n38
  );


  buf
  g166
  (
    n183,
    n8
  );


  buf
  g167
  (
    n216,
    n13
  );


  buf
  g168
  (
    n130,
    n34
  );


  not
  g169
  (
    n180,
    n37
  );


  not
  g170
  (
    n96,
    n30
  );


  not
  g171
  (
    n59,
    n21
  );


  buf
  g172
  (
    n140,
    n27
  );


  not
  g173
  (
    n179,
    n17
  );


  buf
  g174
  (
    n314,
    n124
  );


  not
  g175
  (
    n301,
    n121
  );


  buf
  g176
  (
    n229,
    n115
  );


  not
  g177
  (
    n275,
    n71
  );


  buf
  g178
  (
    n296,
    n72
  );


  buf
  g179
  (
    n298,
    n92
  );


  buf
  g180
  (
    n260,
    n106
  );


  buf
  g181
  (
    n268,
    n90
  );


  not
  g182
  (
    n321,
    n110
  );


  buf
  g183
  (
    n323,
    n95
  );


  not
  g184
  (
    n262,
    n120
  );


  not
  g185
  (
    n292,
    n65
  );


  buf
  g186
  (
    n289,
    n87
  );


  buf
  g187
  (
    n315,
    n68
  );


  buf
  g188
  (
    n249,
    n56
  );


  not
  g189
  (
    n228,
    n91
  );


  buf
  g190
  (
    n310,
    n74
  );


  buf
  g191
  (
    n328,
    n83
  );


  buf
  g192
  (
    n251,
    n89
  );


  buf
  g193
  (
    n320,
    n113
  );


  not
  g194
  (
    n239,
    n91
  );


  buf
  g195
  (
    n243,
    n95
  );


  not
  g196
  (
    n317,
    n63
  );


  not
  g197
  (
    n327,
    n92
  );


  buf
  g198
  (
    n253,
    n55
  );


  buf
  g199
  (
    n306,
    n58
  );


  buf
  g200
  (
    n265,
    n103
  );


  buf
  g201
  (
    n311,
    n98
  );


  not
  g202
  (
    n264,
    n122
  );


  not
  g203
  (
    n333,
    n66
  );


  buf
  g204
  (
    n303,
    n79
  );


  not
  g205
  (
    n281,
    n104
  );


  not
  g206
  (
    n242,
    n107
  );


  buf
  g207
  (
    n330,
    n57
  );


  not
  g208
  (
    n284,
    n105
  );


  buf
  g209
  (
    n259,
    n100
  );


  not
  g210
  (
    n304,
    n96
  );


  not
  g211
  (
    n232,
    n111
  );


  not
  g212
  (
    n250,
    n119
  );


  not
  g213
  (
    n270,
    n60
  );


  not
  g214
  (
    n247,
    n125
  );


  not
  g215
  (
    n231,
    n93
  );


  buf
  g216
  (
    n300,
    n73
  );


  not
  g217
  (
    n322,
    n102
  );


  not
  g218
  (
    n291,
    n64
  );


  buf
  g219
  (
    n316,
    n116
  );


  not
  g220
  (
    n263,
    n90
  );


  buf
  g221
  (
    n278,
    n89
  );


  buf
  g222
  (
    n283,
    n107
  );


  buf
  g223
  (
    n288,
    n87
  );


  buf
  g224
  (
    n332,
    n76
  );


  not
  g225
  (
    n257,
    n114
  );


  not
  g226
  (
    n307,
    n67
  );


  not
  g227
  (
    n318,
    n93
  );


  buf
  g228
  (
    n258,
    n112
  );


  not
  g229
  (
    n240,
    n80
  );


  buf
  g230
  (
    n234,
    n99
  );


  not
  g231
  (
    n256,
    n84
  );


  buf
  g232
  (
    n241,
    n113
  );


  not
  g233
  (
    n293,
    n88
  );


  not
  g234
  (
    n227,
    n88
  );


  not
  g235
  (
    n271,
    n105
  );


  not
  g236
  (
    n277,
    n81
  );


  buf
  g237
  (
    n269,
    n69
  );


  not
  g238
  (
    n309,
    n59
  );


  not
  g239
  (
    n313,
    n94
  );


  buf
  g240
  (
    n329,
    n75
  );


  buf
  g241
  (
    n245,
    n77
  );


  buf
  g242
  (
    n308,
    n125
  );


  buf
  g243
  (
    n286,
    n101
  );


  not
  g244
  (
    n324,
    n122
  );


  buf
  g245
  (
    n236,
    n121
  );


  buf
  g246
  (
    n279,
    n61
  );


  not
  g247
  (
    n266,
    n123
  );


  not
  g248
  (
    n326,
    n114
  );


  not
  g249
  (
    n261,
    n70
  );


  buf
  g250
  (
    n312,
    n96
  );


  not
  g251
  (
    n287,
    n62
  );


  buf
  g252
  (
    n297,
    n117
  );


  not
  g253
  (
    n280,
    n119
  );


  buf
  g254
  (
    n274,
    n94
  );


  not
  g255
  (
    n267,
    n106
  );


  not
  g256
  (
    n273,
    n110
  );


  buf
  g257
  (
    n255,
    n116
  );


  not
  g258
  (
    n299,
    n126
  );


  not
  g259
  (
    n325,
    n54
  );


  buf
  g260
  (
    n248,
    n120
  );


  buf
  g261
  (
    n331,
    n97
  );


  not
  g262
  (
    n302,
    n98
  );


  buf
  g263
  (
    n246,
    n118
  );


  buf
  g264
  (
    n238,
    n109
  );


  not
  g265
  (
    n334,
    n53
  );


  buf
  g266
  (
    n254,
    n78
  );


  not
  g267
  (
    n285,
    n123
  );


  buf
  g268
  (
    n295,
    n102
  );


  not
  g269
  (
    n244,
    n101
  );


  buf
  g270
  (
    n272,
    n111
  );


  buf
  g271
  (
    n252,
    n109
  );


  not
  g272
  (
    n230,
    n100
  );


  buf
  g273
  (
    n305,
    n117
  );


  not
  g274
  (
    n290,
    n124
  );


  not
  g275
  (
    n282,
    n97
  );


  not
  g276
  (
    n237,
    n86
  );


  not
  g277
  (
    n235,
    n115
  );


  not
  g278
  (
    n294,
    n99
  );


  buf
  g279
  (
    n276,
    n85
  );


  xnor
  g280
  (
    n233,
    n108,
    n118,
    n112
  );


  nand
  g281
  (
    n319,
    n103,
    n104,
    n108,
    n82
  );


  nor
  g282
  (
    n353,
    n230,
    n127
  );


  nand
  g283
  (
    n359,
    n289,
    n257,
    n240,
    n275
  );


  nor
  g284
  (
    n339,
    n251,
    n273,
    n242,
    n255
  );


  nor
  g285
  (
    n362,
    n303,
    n295,
    n282,
    n228
  );


  or
  g286
  (
    n340,
    n262,
    n235,
    n284,
    n247
  );


  nor
  g287
  (
    n360,
    n241,
    n298,
    n261,
    n297
  );


  nor
  g288
  (
    n355,
    n266,
    n290,
    n319,
    n278
  );


  nor
  g289
  (
    n337,
    n129,
    n271,
    n128,
    n311
  );


  and
  g290
  (
    n348,
    n283,
    n329,
    n310,
    n236
  );


  and
  g291
  (
    n346,
    n245,
    n127,
    n288,
    n231
  );


  xnor
  g292
  (
    n357,
    n299,
    n321,
    n291,
    n252
  );


  nor
  g293
  (
    n352,
    n307,
    n277,
    n269,
    n272
  );


  xor
  g294
  (
    n341,
    n315,
    n300,
    n265,
    n246
  );


  nor
  g295
  (
    n344,
    n227,
    n332,
    n293,
    n243
  );


  and
  g296
  (
    n350,
    n233,
    n308,
    n260,
    n232
  );


  and
  g297
  (
    n356,
    n274,
    n287,
    n258,
    n314
  );


  xnor
  g298
  (
    n361,
    n254,
    n267,
    n305,
    n244
  );


  nor
  g299
  (
    n354,
    n229,
    n280,
    n325,
    n238
  );


  xor
  g300
  (
    n349,
    n126,
    n323,
    n302,
    n306
  );


  or
  g301
  (
    n342,
    n322,
    n237,
    n256,
    n263
  );


  xor
  g302
  (
    n338,
    n320,
    n264,
    n253,
    n285
  );


  and
  g303
  (
    n336,
    n249,
    n309,
    n270,
    n331
  );


  xor
  g304
  (
    n358,
    n334,
    n318,
    n276,
    n286
  );


  nor
  g305
  (
    n347,
    n326,
    n301,
    n294,
    n328
  );


  or
  g306
  (
    n363,
    n248,
    n317,
    n279,
    n312
  );


  or
  g307
  (
    n343,
    n313,
    n330,
    n259,
    n268
  );


  nor
  g308
  (
    n335,
    n234,
    n333,
    n128,
    n296
  );


  xnor
  g309
  (
    n345,
    n250,
    n292,
    n316,
    n239
  );


  xor
  g310
  (
    n351,
    n281,
    n304,
    n327,
    n324
  );


  buf
  g311
  (
    n368,
    n49
  );


  not
  g312
  (
    n372,
    n51
  );


  not
  g313
  (
    n370,
    n358
  );


  not
  g314
  (
    n365,
    n356
  );


  buf
  g315
  (
    n367,
    n50
  );


  xor
  g316
  (
    n375,
    n50,
    n351
  );


  xnor
  g317
  (
    n374,
    n48,
    n49
  );


  xnor
  g318
  (
    n364,
    n48,
    n47,
    n348
  );


  nor
  g319
  (
    n376,
    n48,
    n360,
    n359
  );


  nand
  g320
  (
    n371,
    n354,
    n50
  );


  xor
  g321
  (
    n369,
    n350,
    n355,
    n352
  );


  xnor
  g322
  (
    n366,
    n357,
    n47,
    n353
  );


  and
  g323
  (
    n373,
    n49,
    n349,
    n48
  );


  xnor
  g324
  (
    n387,
    n140,
    n366,
    n365
  );


  or
  g325
  (
    n385,
    n144,
    n140,
    n143,
    n137
  );


  nor
  g326
  (
    n388,
    n133,
    n132,
    n135,
    n367
  );


  and
  g327
  (
    n383,
    n132,
    n142,
    n143,
    n366
  );


  nor
  g328
  (
    n379,
    n365,
    n136,
    n129,
    n146
  );


  nor
  g329
  (
    n386,
    n145,
    n364,
    n131
  );


  and
  g330
  (
    n380,
    n144,
    n146,
    n138,
    n133
  );


  nand
  g331
  (
    n382,
    n139,
    n134,
    n366,
    n135
  );


  nand
  g332
  (
    n381,
    n130,
    n139,
    n142,
    n136
  );


  or
  g333
  (
    n378,
    n147,
    n131,
    n366,
    n367
  );


  and
  g334
  (
    n384,
    n134,
    n145,
    n137,
    n130
  );


  or
  g335
  (
    n377,
    n365,
    n141,
    n138
  );


  buf
  g336
  (
    n391,
    n379
  );


  not
  g337
  (
    n393,
    n380
  );


  not
  g338
  (
    n398,
    n377
  );


  not
  g339
  (
    n397,
    n378
  );


  not
  g340
  (
    n392,
    n378
  );


  buf
  g341
  (
    n396,
    n381
  );


  not
  g342
  (
    n390,
    n379
  );


  not
  g343
  (
    n395,
    n381
  );


  not
  g344
  (
    n389,
    n380
  );


  buf
  g345
  (
    n394,
    n377
  );


  buf
  g346
  (
    n400,
    n362
  );


  not
  g347
  (
    n401,
    n392
  );


  buf
  g348
  (
    n402,
    n361
  );


  and
  g349
  (
    n399,
    n389,
    n390,
    n391
  );


  buf
  g350
  (
    n406,
    n400
  );


  not
  g351
  (
    n408,
    n399
  );


  not
  g352
  (
    n409,
    n400
  );


  buf
  g353
  (
    n404,
    n401
  );


  not
  g354
  (
    n405,
    n400
  );


  not
  g355
  (
    n407,
    n399
  );


  not
  g356
  (
    n412,
    n399
  );


  not
  g357
  (
    n403,
    n400
  );


  buf
  g358
  (
    n411,
    n401
  );


  buf
  g359
  (
    n410,
    n399
  );


  not
  g360
  (
    n414,
    n406
  );


  buf
  g361
  (
    n422,
    n404
  );


  buf
  g362
  (
    n418,
    n385
  );


  not
  g363
  (
    n417,
    n404
  );


  buf
  g364
  (
    n425,
    n403
  );


  not
  g365
  (
    n427,
    n403
  );


  not
  g366
  (
    n419,
    n403
  );


  buf
  g367
  (
    n426,
    n383
  );


  not
  g368
  (
    n415,
    n405
  );


  buf
  g369
  (
    n421,
    n403
  );


  buf
  g370
  (
    n420,
    n406
  );


  not
  g371
  (
    n413,
    n404
  );


  nand
  g372
  (
    n424,
    n404,
    n386,
    n384,
    n382
  );


  xnor
  g373
  (
    n416,
    n385,
    n405,
    n406
  );


  nor
  g374
  (
    n423,
    n383,
    n382,
    n405,
    n384
  );


  nor
  g375
  (
    n436,
    n163,
    n157,
    n156,
    n153
  );


  and
  g376
  (
    n428,
    n151,
    n164,
    n152,
    n158
  );


  nand
  g377
  (
    n431,
    n150,
    n155,
    n413,
    n152
  );


  xnor
  g378
  (
    n435,
    n396,
    n166,
    n162
  );


  xor
  g379
  (
    n434,
    n163,
    n150,
    n414,
    n147
  );


  nand
  g380
  (
    n432,
    n416,
    n413,
    n414,
    n167
  );


  nor
  g381
  (
    n444,
    n161,
    n168,
    n169,
    n413
  );


  nand
  g382
  (
    n430,
    n393,
    n168,
    n416,
    n414
  );


  nand
  g383
  (
    n440,
    n154,
    n157,
    n415
  );


  and
  g384
  (
    n443,
    n415,
    n149,
    n395
  );


  xnor
  g385
  (
    n439,
    n165,
    n161,
    n414,
    n167
  );


  xor
  g386
  (
    n442,
    n159,
    n166,
    n160,
    n154
  );


  xnor
  g387
  (
    n429,
    n148,
    n151,
    n413,
    n165
  );


  nor
  g388
  (
    n437,
    n416,
    n155,
    n160,
    n417
  );


  xor
  g389
  (
    n433,
    n394,
    n415,
    n153,
    n416
  );


  nand
  g390
  (
    n441,
    n398,
    n148,
    n164,
    n158
  );


  nand
  g391
  (
    n438,
    n159,
    n156,
    n169,
    n397
  );


  buf
  g392
  (
    n446,
    n433
  );


  buf
  g393
  (
    n475,
    n428
  );


  buf
  g394
  (
    n470,
    n429
  );


  not
  g395
  (
    n458,
    n436
  );


  buf
  g396
  (
    n467,
    n429
  );


  not
  g397
  (
    n468,
    n433
  );


  not
  g398
  (
    n478,
    n435
  );


  not
  g399
  (
    n469,
    n431
  );


  not
  g400
  (
    n454,
    n429
  );


  buf
  g401
  (
    n471,
    n430
  );


  not
  g402
  (
    n453,
    n430
  );


  buf
  g403
  (
    n449,
    n434
  );


  buf
  g404
  (
    n477,
    n434
  );


  buf
  g405
  (
    n474,
    n432
  );


  buf
  g406
  (
    n447,
    n435
  );


  not
  g407
  (
    n462,
    n434
  );


  buf
  g408
  (
    n455,
    n433
  );


  buf
  g409
  (
    n459,
    n430
  );


  not
  g410
  (
    n460,
    n431
  );


  buf
  g411
  (
    n451,
    n401
  );


  buf
  g412
  (
    n448,
    n437
  );


  not
  g413
  (
    n464,
    n432
  );


  buf
  g414
  (
    n476,
    n436
  );


  buf
  g415
  (
    n473,
    n432
  );


  buf
  g416
  (
    n456,
    n431
  );


  not
  g417
  (
    n457,
    n401
  );


  buf
  g418
  (
    n465,
    n402
  );


  buf
  g419
  (
    n445,
    n431
  );


  not
  g420
  (
    n472,
    n436
  );


  not
  g421
  (
    n463,
    n402
  );


  buf
  g422
  (
    n452,
    n429
  );


  not
  g423
  (
    n466,
    n402
  );


  xnor
  g424
  (
    n461,
    n430,
    n435,
    n433,
    n402
  );


  nand
  g425
  (
    n450,
    n435,
    n436,
    n432,
    n434
  );


  not
  g426
  (
    n492,
    n460
  );


  buf
  g427
  (
    n527,
    n472
  );


  not
  g428
  (
    n522,
    n453
  );


  not
  g429
  (
    n520,
    n462
  );


  not
  g430
  (
    n521,
    n412
  );


  buf
  g431
  (
    n496,
    n477
  );


  buf
  g432
  (
    n533,
    n476
  );


  buf
  g433
  (
    n497,
    n452
  );


  buf
  g434
  (
    n498,
    n463
  );


  buf
  g435
  (
    n529,
    n412
  );


  buf
  g436
  (
    n495,
    n475
  );


  buf
  g437
  (
    n547,
    n474
  );


  not
  g438
  (
    n534,
    n412
  );


  not
  g439
  (
    n523,
    n410
  );


  not
  g440
  (
    n516,
    n455
  );


  not
  g441
  (
    n532,
    n463
  );


  buf
  g442
  (
    n511,
    n466
  );


  buf
  g443
  (
    n528,
    n451
  );


  not
  g444
  (
    n526,
    n451
  );


  buf
  g445
  (
    n517,
    n464
  );


  buf
  g446
  (
    n513,
    n458
  );


  not
  g447
  (
    n536,
    n409
  );


  buf
  g448
  (
    n530,
    n412
  );


  buf
  g449
  (
    n524,
    n407
  );


  not
  g450
  (
    n509,
    n467
  );


  buf
  g451
  (
    n518,
    n445
  );


  not
  g452
  (
    n546,
    n454
  );


  not
  g453
  (
    n541,
    n407
  );


  not
  g454
  (
    n525,
    n448
  );


  buf
  g455
  (
    n499,
    n457
  );


  not
  g456
  (
    n484,
    n478
  );


  buf
  g457
  (
    n551,
    n462
  );


  buf
  g458
  (
    n481,
    n447
  );


  buf
  g459
  (
    n488,
    n468
  );


  not
  g460
  (
    n543,
    n453
  );


  buf
  g461
  (
    n480,
    n409
  );


  buf
  g462
  (
    n519,
    n408
  );


  not
  g463
  (
    n505,
    n469
  );


  not
  g464
  (
    n504,
    n473
  );


  buf
  g465
  (
    n507,
    n446
  );


  buf
  g466
  (
    n514,
    n471
  );


  not
  g467
  (
    n539,
    n410
  );


  not
  g468
  (
    n549,
    n470
  );


  not
  g469
  (
    n537,
    n410
  );


  buf
  g470
  (
    n502,
    n410
  );


  not
  g471
  (
    n506,
    n458
  );


  buf
  g472
  (
    n500,
    n469
  );


  buf
  g473
  (
    n487,
    n457
  );


  not
  g474
  (
    n503,
    n472
  );


  buf
  g475
  (
    n508,
    n452
  );


  not
  g476
  (
    n485,
    n411
  );


  buf
  g477
  (
    n512,
    n411
  );


  not
  g478
  (
    n479,
    n467
  );


  not
  g479
  (
    n542,
    n406
  );


  not
  g480
  (
    n515,
    n476
  );


  buf
  g481
  (
    n548,
    n459
  );


  buf
  g482
  (
    n491,
    n465
  );


  buf
  g483
  (
    n540,
    n408
  );


  not
  g484
  (
    n486,
    n468
  );


  buf
  g485
  (
    n494,
    n461
  );


  not
  g486
  (
    n531,
    n409
  );


  not
  g487
  (
    n483,
    n477
  );


  buf
  g488
  (
    n510,
    n476
  );


  not
  g489
  (
    n482,
    n475
  );


  nor
  g490
  (
    n490,
    n409,
    n478
  );


  xor
  g491
  (
    n489,
    n408,
    n454,
    n411,
    n456
  );


  xnor
  g492
  (
    n493,
    n466,
    n464,
    n407,
    n470
  );


  or
  g493
  (
    n535,
    n477,
    n447,
    n411,
    n449
  );


  nor
  g494
  (
    n550,
    n460,
    n474,
    n450
  );


  nand
  g495
  (
    n538,
    n478,
    n465,
    n473,
    n477
  );


  nand
  g496
  (
    n545,
    n476,
    n445,
    n446,
    n459
  );


  and
  g497
  (
    n544,
    n407,
    n449,
    n461,
    n455
  );


  xor
  g498
  (
    n501,
    n408,
    n456,
    n471,
    n448
  );


  buf
  g499
  (
    n679,
    n374
  );


  not
  g500
  (
    n583,
    n525
  );


  not
  g501
  (
    n556,
    n506
  );


  buf
  g502
  (
    n736,
    n504
  );


  buf
  g503
  (
    n669,
    n371
  );


  not
  g504
  (
    n690,
    n488
  );


  not
  g505
  (
    n732,
    n502
  );


  not
  g506
  (
    n589,
    n372
  );


  buf
  g507
  (
    n705,
    n424
  );


  not
  g508
  (
    n668,
    n421
  );


  not
  g509
  (
    n594,
    n522
  );


  buf
  g510
  (
    n597,
    n419
  );


  not
  g511
  (
    n622,
    n486
  );


  buf
  g512
  (
    n579,
    n489
  );


  not
  g513
  (
    n581,
    n512
  );


  not
  g514
  (
    n719,
    n523
  );


  not
  g515
  (
    n708,
    n518
  );


  buf
  g516
  (
    n649,
    n370
  );


  not
  g517
  (
    n704,
    n417
  );


  buf
  g518
  (
    n738,
    n523
  );


  buf
  g519
  (
    n667,
    n367
  );


  not
  g520
  (
    n695,
    n524
  );


  buf
  g521
  (
    n559,
    n486
  );


  buf
  g522
  (
    n701,
    n425
  );


  buf
  g523
  (
    n682,
    n482
  );


  buf
  g524
  (
    n663,
    n498
  );


  not
  g525
  (
    n716,
    n369
  );


  buf
  g526
  (
    n595,
    n516
  );


  buf
  g527
  (
    n647,
    n485
  );


  buf
  g528
  (
    n602,
    n482
  );


  buf
  g529
  (
    n606,
    n525
  );


  not
  g530
  (
    n684,
    n51
  );


  not
  g531
  (
    n591,
    n514
  );


  not
  g532
  (
    n554,
    n515
  );


  buf
  g533
  (
    n672,
    n484
  );


  not
  g534
  (
    n697,
    n499
  );


  buf
  g535
  (
    n648,
    n483
  );


  not
  g536
  (
    n607,
    n507
  );


  buf
  g537
  (
    n747,
    n508
  );


  not
  g538
  (
    n592,
    n521
  );


  buf
  g539
  (
    n702,
    n514
  );


  not
  g540
  (
    n557,
    n512
  );


  not
  g541
  (
    n715,
    n485
  );


  buf
  g542
  (
    n694,
    n507
  );


  not
  g543
  (
    n641,
    n375
  );


  not
  g544
  (
    n588,
    n523
  );


  buf
  g545
  (
    n689,
    n505
  );


  buf
  g546
  (
    n656,
    n500
  );


  not
  g547
  (
    n565,
    n526
  );


  buf
  g548
  (
    n662,
    n503
  );


  not
  g549
  (
    n564,
    n525
  );


  not
  g550
  (
    n692,
    n505
  );


  not
  g551
  (
    n745,
    n370
  );


  not
  g552
  (
    n660,
    n495
  );


  buf
  g553
  (
    n568,
    n483
  );


  buf
  g554
  (
    n670,
    n504
  );


  buf
  g555
  (
    n737,
    n513
  );


  not
  g556
  (
    n561,
    n513
  );


  not
  g557
  (
    n643,
    n374
  );


  buf
  g558
  (
    n610,
    n427
  );


  buf
  g559
  (
    n553,
    n482
  );


  buf
  g560
  (
    n612,
    n519
  );


  not
  g561
  (
    n666,
    n512
  );


  not
  g562
  (
    n638,
    n526
  );


  not
  g563
  (
    n603,
    n417
  );


  not
  g564
  (
    n575,
    n487
  );


  not
  g565
  (
    n582,
    n371
  );


  not
  g566
  (
    n664,
    n519
  );


  not
  g567
  (
    n744,
    n506
  );


  buf
  g568
  (
    n584,
    n512
  );


  not
  g569
  (
    n593,
    n495
  );


  buf
  g570
  (
    n713,
    n523
  );


  buf
  g571
  (
    n628,
    n424
  );


  not
  g572
  (
    n632,
    n510
  );


  not
  g573
  (
    n640,
    n524
  );


  not
  g574
  (
    n609,
    n494
  );


  buf
  g575
  (
    n634,
    n370
  );


  not
  g576
  (
    n650,
    n514
  );


  not
  g577
  (
    n717,
    n521
  );


  not
  g578
  (
    n600,
    n527
  );


  not
  g579
  (
    n636,
    n422
  );


  not
  g580
  (
    n631,
    n492
  );


  not
  g581
  (
    n651,
    n486
  );


  buf
  g582
  (
    n611,
    n374
  );


  buf
  g583
  (
    n659,
    n479
  );


  buf
  g584
  (
    n567,
    n479
  );


  buf
  g585
  (
    n635,
    n368
  );


  not
  g586
  (
    n637,
    n420
  );


  not
  g587
  (
    n680,
    n484
  );


  not
  g588
  (
    n729,
    n423
  );


  not
  g589
  (
    n639,
    n484
  );


  not
  g590
  (
    n574,
    n503
  );


  not
  g591
  (
    n566,
    n491
  );


  not
  g592
  (
    n655,
    n524
  );


  not
  g593
  (
    n723,
    n498
  );


  buf
  g594
  (
    n601,
    n499
  );


  buf
  g595
  (
    n552,
    n424
  );


  not
  g596
  (
    n710,
    n490
  );


  buf
  g597
  (
    n709,
    n425
  );


  buf
  g598
  (
    n590,
    n487
  );


  buf
  g599
  (
    n735,
    n480
  );


  not
  g600
  (
    n731,
    n518
  );


  not
  g601
  (
    n645,
    n517
  );


  buf
  g602
  (
    n742,
    n498
  );


  not
  g603
  (
    n586,
    n481
  );


  not
  g604
  (
    n711,
    n502
  );


  buf
  g605
  (
    n569,
    n368
  );


  buf
  g606
  (
    n617,
    n373
  );


  not
  g607
  (
    n573,
    n421
  );


  buf
  g608
  (
    n726,
    n491
  );


  not
  g609
  (
    n571,
    n496
  );


  buf
  g610
  (
    n703,
    n480
  );


  buf
  g611
  (
    n721,
    n485
  );


  buf
  g612
  (
    n707,
    n423
  );


  buf
  g613
  (
    n678,
    n375
  );


  buf
  g614
  (
    n706,
    n490
  );


  not
  g615
  (
    n741,
    n504
  );


  not
  g616
  (
    n728,
    n511
  );


  not
  g617
  (
    n677,
    n501
  );


  buf
  g618
  (
    n654,
    n488
  );


  not
  g619
  (
    n714,
    n499
  );


  buf
  g620
  (
    n691,
    n422
  );


  not
  g621
  (
    n587,
    n516
  );


  not
  g622
  (
    n646,
    n521
  );


  not
  g623
  (
    n657,
    n518
  );


  not
  g624
  (
    n661,
    n418
  );


  buf
  g625
  (
    n696,
    n418
  );


  not
  g626
  (
    n621,
    n506
  );


  not
  g627
  (
    n577,
    n500
  );


  buf
  g628
  (
    n722,
    n509
  );


  not
  g629
  (
    n739,
    n503
  );


  buf
  g630
  (
    n720,
    n527
  );


  buf
  g631
  (
    n683,
    n498
  );


  buf
  g632
  (
    n674,
    n490
  );


  buf
  g633
  (
    n626,
    n516
  );


  not
  g634
  (
    n743,
    n419
  );


  buf
  g635
  (
    n576,
    n522
  );


  buf
  g636
  (
    n693,
    n509
  );


  buf
  g637
  (
    n700,
    n481
  );


  buf
  g638
  (
    n653,
    n495
  );


  not
  g639
  (
    n624,
    n497
  );


  not
  g640
  (
    n676,
    n501
  );


  not
  g641
  (
    n604,
    n426
  );


  not
  g642
  (
    n681,
    n526
  );


  buf
  g643
  (
    n699,
    n369
  );


  buf
  g644
  (
    n608,
    n525
  );


  buf
  g645
  (
    n652,
    n519
  );


  not
  g646
  (
    n630,
    n504
  );


  not
  g647
  (
    n614,
    n492
  );


  not
  g648
  (
    n616,
    n516
  );


  not
  g649
  (
    n740,
    n502
  );


  not
  g650
  (
    n688,
    n491
  );


  buf
  g651
  (
    n633,
    n493
  );


  not
  g652
  (
    n727,
    n426
  );


  not
  g653
  (
    n733,
    n509
  );


  buf
  g654
  (
    n725,
    n519
  );


  buf
  g655
  (
    n734,
    n421
  );


  buf
  g656
  (
    n730,
    n427
  );


  buf
  g657
  (
    n686,
    n483
  );


  buf
  g658
  (
    n665,
    n510
  );


  not
  g659
  (
    n599,
    n511
  );


  not
  g660
  (
    n625,
    n493
  );


  buf
  g661
  (
    n555,
    n499
  );


  buf
  g662
  (
    n558,
    n375
  );


  buf
  g663
  (
    n642,
    n508
  );


  buf
  g664
  (
    n658,
    n488
  );


  buf
  g665
  (
    n580,
    n372
  );


  not
  g666
  (
    n629,
    n495
  );


  not
  g667
  (
    n644,
    n368
  );


  buf
  g668
  (
    n578,
    n522
  );


  nor
  g669
  (
    n746,
    n487,
    n487,
    n505,
    n501
  );


  xor
  g670
  (
    n675,
    n518,
    n421,
    n493,
    n484
  );


  nand
  g671
  (
    n619,
    n419,
    n520,
    n508,
    n506
  );


  nor
  g672
  (
    n687,
    n372,
    n427,
    n502,
    n492
  );


  and
  g673
  (
    n718,
    n481,
    n522,
    n427,
    n510
  );


  xnor
  g674
  (
    n724,
    n486,
    n520,
    n524,
    n420
  );


  xnor
  g675
  (
    n671,
    n493,
    n371,
    n425,
    n419
  );


  xor
  g676
  (
    n605,
    n526,
    n510,
    n485,
    n491
  );


  nor
  g677
  (
    n623,
    n511,
    n511,
    n501,
    n517
  );


  xor
  g678
  (
    n615,
    n503,
    n515,
    n423,
    n418
  );


  xor
  g679
  (
    n712,
    n497,
    n521,
    n368,
    n492
  );


  nand
  g680
  (
    n618,
    n508,
    n370,
    n488,
    n509
  );


  and
  g681
  (
    n620,
    n424,
    n373,
    n507,
    n482
  );


  xnor
  g682
  (
    n563,
    n517,
    n496,
    n515,
    n373
  );


  xor
  g683
  (
    n585,
    n423,
    n514,
    n479,
    n494
  );


  xnor
  g684
  (
    n685,
    n520,
    n527,
    n417,
    n422
  );


  xor
  g685
  (
    n698,
    n489,
    n372,
    n527,
    n497
  );


  xnor
  g686
  (
    n570,
    n373,
    n418,
    n479,
    n481
  );


  nor
  g687
  (
    n596,
    n489,
    n515,
    n500,
    n367
  );


  and
  g688
  (
    n562,
    n513,
    n507,
    n489,
    n490
  );


  nand
  g689
  (
    n572,
    n480,
    n420,
    n425,
    n375
  );


  nor
  g690
  (
    n673,
    n494,
    n497,
    n369,
    n420
  );


  or
  g691
  (
    n560,
    n513,
    n422,
    n505,
    n426
  );


  and
  g692
  (
    n598,
    n520,
    n496,
    n500
  );


  xor
  g693
  (
    n627,
    n369,
    n517,
    n494,
    n426
  );


  nand
  g694
  (
    n613,
    n374,
    n480,
    n371,
    n483
  );


  buf
  g695
  (
    n748,
    n556
  );


  not
  g696
  (
    n753,
    n552
  );


  not
  g697
  (
    n749,
    n555
  );


  not
  g698
  (
    n751,
    n557
  );


  not
  g699
  (
    n754,
    n553
  );


  and
  g700
  (
    n750,
    n552,
    n554,
    n556
  );


  nor
  g701
  (
    n752,
    n557,
    n555,
    n553,
    n554
  );


  not
  g702
  (
    n761,
    n561
  );


  nor
  g703
  (
    n762,
    n564,
    n748,
    n562
  );


  or
  g704
  (
    n755,
    n558,
    n753,
    n566,
    n750
  );


  nand
  g705
  (
    n757,
    n752,
    n478,
    n564,
    n565
  );


  nor
  g706
  (
    n759,
    n563,
    n559,
    n562,
    n565
  );


  xor
  g707
  (
    n756,
    n560,
    n563,
    n754,
    n561
  );


  and
  g708
  (
    n760,
    n170,
    n560,
    n559,
    n558
  );


  nor
  g709
  (
    n758,
    n566,
    n751,
    n749,
    n754
  );


  xnor
  g710
  (
    n791,
    n538,
    n541,
    n551,
    n542
  );


  xor
  g711
  (
    n780,
    n544,
    n543,
    n529,
    n539
  );


  nor
  g712
  (
    n764,
    n759,
    n755,
    n533,
    n535
  );


  xnor
  g713
  (
    n766,
    n758,
    n539,
    n550,
    n551
  );


  nand
  g714
  (
    n786,
    n761,
    n534,
    n536,
    n539
  );


  xor
  g715
  (
    n788,
    n755,
    n757,
    n529,
    n538
  );


  xor
  g716
  (
    n768,
    n760,
    n550,
    n545,
    n759
  );


  xnor
  g717
  (
    n785,
    n548,
    n545,
    n536,
    n538
  );


  xnor
  g718
  (
    n763,
    n547,
    n755,
    n530,
    n535
  );


  nand
  g719
  (
    n772,
    n534,
    n546,
    n544,
    n759
  );


  or
  g720
  (
    n783,
    n548,
    n756,
    n541
  );


  and
  g721
  (
    n767,
    n543,
    n756,
    n544,
    n530
  );


  and
  g722
  (
    n787,
    n543,
    n528,
    n760,
    n762
  );


  or
  g723
  (
    n776,
    n757,
    n540,
    n543,
    n551
  );


  nor
  g724
  (
    n765,
    n535,
    n540,
    n545,
    n528
  );


  xor
  g725
  (
    n774,
    n529,
    n549,
    n542,
    n537
  );


  or
  g726
  (
    n770,
    n762,
    n548,
    n547,
    n758
  );


  nor
  g727
  (
    n781,
    n531,
    n762,
    n542,
    n540
  );


  and
  g728
  (
    n775,
    n761,
    n756,
    n528,
    n546
  );


  and
  g729
  (
    n784,
    n547,
    n544,
    n755,
    n546
  );


  and
  g730
  (
    n779,
    n550,
    n528,
    n761
  );


  xor
  g731
  (
    n773,
    n538,
    n530,
    n535,
    n551
  );


  nand
  g732
  (
    n794,
    n760,
    n757,
    n541,
    n547
  );


  and
  g733
  (
    n771,
    n529,
    n534,
    n542,
    n545
  );


  xnor
  g734
  (
    n793,
    n536,
    n537,
    n532,
    n533
  );


  or
  g735
  (
    n778,
    n533,
    n762,
    n758,
    n757
  );


  xnor
  g736
  (
    n782,
    n532,
    n534,
    n531
  );


  xor
  g737
  (
    n792,
    n531,
    n530,
    n760,
    n532
  );


  xnor
  g738
  (
    n789,
    n537,
    n541,
    n549,
    n536
  );


  nand
  g739
  (
    n790,
    n550,
    n759,
    n532,
    n533
  );


  or
  g740
  (
    n777,
    n758,
    n539,
    n546,
    n549
  );


  nor
  g741
  (
    n769,
    n537,
    n549,
    n548,
    n540
  );


  not
  g742
  (
    n810,
    n780
  );


  buf
  g743
  (
    n801,
    n570
  );


  buf
  g744
  (
    n814,
    n568
  );


  not
  g745
  (
    n804,
    n569
  );


  buf
  g746
  (
    n796,
    n766
  );


  not
  g747
  (
    n809,
    n773
  );


  buf
  g748
  (
    n808,
    n764
  );


  buf
  g749
  (
    n813,
    n779
  );


  not
  g750
  (
    n795,
    n780
  );


  not
  g751
  (
    n798,
    n778
  );


  not
  g752
  (
    n812,
    n765
  );


  not
  g753
  (
    n797,
    n569
  );


  not
  g754
  (
    n802,
    n567
  );


  not
  g755
  (
    n803,
    n567
  );


  not
  g756
  (
    n811,
    n568
  );


  not
  g757
  (
    n805,
    n767
  );


  buf
  g758
  (
    n799,
    n781
  );


  not
  g759
  (
    n806,
    n768
  );


  xor
  g760
  (
    n800,
    n777,
    n770
  );


  nor
  g761
  (
    n807,
    n763,
    n771,
    n769,
    n772
  );


  nor
  g762
  (
    n815,
    n774,
    n775,
    n776,
    n779
  );


  xnor
  g763
  (
    n820,
    n171,
    n212,
    n196,
    n800
  );


  xnor
  g764
  (
    n853,
    n797,
    n796,
    n191
  );


  and
  g765
  (
    n847,
    n215,
    n193,
    n206
  );


  xor
  g766
  (
    n838,
    n174,
    n203,
    n216,
    n795
  );


  xor
  g767
  (
    n842,
    n799,
    n575,
    n800,
    n796
  );


  nand
  g768
  (
    n849,
    n216,
    n185,
    n173,
    n573
  );


  nor
  g769
  (
    n827,
    n217,
    n804,
    n226,
    n225
  );


  nor
  g770
  (
    n817,
    n207,
    n191,
    n209,
    n176
  );


  nand
  g771
  (
    n856,
    n571,
    n795,
    n192,
    n179
  );


  xor
  g772
  (
    n816,
    n223,
    n204,
    n209,
    n193
  );


  xor
  g773
  (
    n852,
    n183,
    n201,
    n204,
    n197
  );


  or
  g774
  (
    n846,
    n184,
    n210,
    n219,
    n187
  );


  xor
  g775
  (
    n841,
    n182,
    n798,
    n217,
    n223
  );


  nor
  g776
  (
    n843,
    n179,
    n576,
    n186,
    n220
  );


  and
  g777
  (
    n833,
    n180,
    n805,
    n226,
    n804
  );


  and
  g778
  (
    n826,
    n800,
    n207,
    n225,
    n574
  );


  nor
  g779
  (
    n857,
    n796,
    n214,
    n181,
    n196
  );


  nand
  g780
  (
    n854,
    n577,
    n214,
    n799,
    n194
  );


  nor
  g781
  (
    n850,
    n213,
    n186,
    n202,
    n578
  );


  nor
  g782
  (
    n819,
    n195,
    n208,
    n804,
    n220
  );


  nand
  g783
  (
    n845,
    n570,
    n195,
    n221,
    n175
  );


  and
  g784
  (
    n823,
    n218,
    n575,
    n572,
    n221
  );


  or
  g785
  (
    n839,
    n797,
    n571,
    n218,
    n574
  );


  xor
  g786
  (
    n822,
    n205,
    n801,
    n188
  );


  and
  g787
  (
    n837,
    n198,
    n177,
    n170,
    n224
  );


  nor
  g788
  (
    n818,
    n181,
    n212,
    n172,
    n798
  );


  xnor
  g789
  (
    n825,
    n798,
    n222,
    n803,
    n573
  );


  and
  g790
  (
    n832,
    n802,
    n205,
    n219,
    n190
  );


  or
  g791
  (
    n831,
    n199,
    n189,
    n187,
    n201
  );


  nand
  g792
  (
    n844,
    n199,
    n211,
    n215,
    n801
  );


  xor
  g793
  (
    n855,
    n178,
    n224,
    n797,
    n184
  );


  and
  g794
  (
    n828,
    n176,
    n222,
    n572,
    n194
  );


  or
  g795
  (
    n858,
    n211,
    n797,
    n803,
    n802
  );


  xnor
  g796
  (
    n829,
    n175,
    n171,
    n182,
    n801
  );


  and
  g797
  (
    n840,
    n803,
    n197,
    n208,
    n189
  );


  or
  g798
  (
    n821,
    n210,
    n803,
    n576,
    n795
  );


  nor
  g799
  (
    n836,
    n802,
    n190,
    n178,
    n577
  );


  or
  g800
  (
    n835,
    n798,
    n200,
    n802
  );


  nor
  g801
  (
    n834,
    n174,
    n173,
    n801,
    n198
  );


  or
  g802
  (
    n848,
    n795,
    n800,
    n172,
    n799
  );


  xnor
  g803
  (
    n824,
    n202,
    n192,
    n177,
    n180
  );


  nand
  g804
  (
    n851,
    n185,
    n805,
    n183,
    n203
  );


  xor
  g805
  (
    n830,
    n213,
    n805,
    n804,
    n799
  );


  buf
  g806
  (
    n863,
    n819
  );


  buf
  g807
  (
    n859,
    n828
  );


  not
  g808
  (
    n861,
    n822
  );


  buf
  g809
  (
    n862,
    n817
  );


  buf
  g810
  (
    n860,
    n51
  );


  xnor
  g811
  (
    n866,
    n827,
    n52,
    n826
  );


  nor
  g812
  (
    n864,
    n818,
    n816,
    n825,
    n821
  );


  xnor
  g813
  (
    n865,
    n824,
    n823,
    n51,
    n820
  );


  and
  g814
  (
    n871,
    n579,
    n860,
    n863,
    n792
  );


  xnor
  g815
  (
    n874,
    n794,
    n861,
    n782
  );


  nor
  g816
  (
    n873,
    n794,
    n792,
    n793,
    n784
  );


  nor
  g817
  (
    n870,
    n785,
    n783,
    n790,
    n863
  );


  xor
  g818
  (
    n872,
    n862,
    n859,
    n788,
    n789
  );


  xor
  g819
  (
    n869,
    n786,
    n793,
    n781,
    n784
  );


  or
  g820
  (
    n875,
    n860,
    n859,
    n791,
    n787
  );


  or
  g821
  (
    n867,
    n788,
    n791,
    n862,
    n789
  );


  nor
  g822
  (
    n868,
    n787,
    n785,
    n861,
    n578
  );


  and
  g823
  (
    n876,
    n579,
    n790,
    n786,
    n783
  );


  xnor
  g824
  (
    n888,
    n814,
    n870,
    n583,
    n875
  );


  nor
  g825
  (
    n887,
    n806,
    n585,
    n813,
    n808
  );


  nand
  g826
  (
    n878,
    n809,
    n876,
    n807,
    n814
  );


  nor
  g827
  (
    n893,
    n873,
    n811,
    n812,
    n809
  );


  and
  g828
  (
    n882,
    n584,
    n586,
    n815
  );


  nor
  g829
  (
    n889,
    n585,
    n868,
    n813
  );


  xnor
  g830
  (
    n883,
    n580,
    n807,
    n869,
    n876
  );


  nand
  g831
  (
    n886,
    n815,
    n811,
    n874,
    n867
  );


  nor
  g832
  (
    n881,
    n810,
    n810,
    n815,
    n808
  );


  xor
  g833
  (
    n890,
    n809,
    n875,
    n874,
    n807
  );


  or
  g834
  (
    n880,
    n810,
    n814,
    n582,
    n807
  );


  xor
  g835
  (
    n885,
    n872,
    n580,
    n805,
    n871
  );


  and
  g836
  (
    n879,
    n806,
    n873,
    n581,
    n871
  );


  nor
  g837
  (
    n892,
    n808,
    n808,
    n582,
    n869
  );


  nand
  g838
  (
    n877,
    n583,
    n812,
    n810
  );


  or
  g839
  (
    n891,
    n811,
    n581,
    n806,
    n813
  );


  and
  g840
  (
    n884,
    n870,
    n584,
    n809,
    n814
  );


  xnor
  g841
  (
    n894,
    n872,
    n812,
    n811,
    n806
  );


  nor
  g842
  (
    n921,
    n882,
    n598,
    n596,
    n884
  );


  or
  g843
  (
    n943,
    n656,
    n879,
    n659
  );


  nand
  g844
  (
    n932,
    n847,
    n625,
    n631,
    n637
  );


  xor
  g845
  (
    n896,
    n620,
    n609,
    n832,
    n660
  );


  and
  g846
  (
    n942,
    n625,
    n888,
    n635,
    n894
  );


  nand
  g847
  (
    n908,
    n617,
    n663,
    n590,
    n636
  );


  xnor
  g848
  (
    n945,
    n650,
    n892,
    n669,
    n656
  );


  nor
  g849
  (
    n963,
    n889,
    n884,
    n586,
    n599
  );


  xnor
  g850
  (
    n901,
    n631,
    n661,
    n880,
    n842
  );


  and
  g851
  (
    n922,
    n880,
    n657,
    n605,
    n626
  );


  xnor
  g852
  (
    n931,
    n632,
    n882,
    n619,
    n603
  );


  xnor
  g853
  (
    n937,
    n587,
    n649,
    n668,
    n597
  );


  and
  g854
  (
    n903,
    n597,
    n890,
    n637,
    n883
  );


  or
  g855
  (
    n965,
    n604,
    n880,
    n611,
    n881
  );


  and
  g856
  (
    n899,
    n670,
    n851,
    n622,
    n882
  );


  xor
  g857
  (
    n957,
    n830,
    n659,
    n652,
    n878
  );


  xor
  g858
  (
    n898,
    n881,
    n651,
    n878,
    n890
  );


  or
  g859
  (
    n920,
    n894,
    n837,
    n600,
    n886
  );


  and
  g860
  (
    n948,
    n833,
    n593,
    n849,
    n630
  );


  nand
  g861
  (
    n952,
    n849,
    n642,
    n622,
    n893
  );


  nand
  g862
  (
    n918,
    n601,
    n885,
    n612,
    n610
  );


  nand
  g863
  (
    n900,
    n846,
    n852,
    n626,
    n666
  );


  nor
  g864
  (
    n964,
    n606,
    n592,
    n588,
    n621
  );


  xor
  g865
  (
    n905,
    n884,
    n891,
    n646,
    n605
  );


  xnor
  g866
  (
    n930,
    n891,
    n665,
    n877,
    n842
  );


  nand
  g867
  (
    n923,
    n623,
    n669,
    n643,
    n640
  );


  nor
  g868
  (
    n949,
    n654,
    n604,
    n594,
    n613
  );


  and
  g869
  (
    n958,
    n607,
    n628,
    n632,
    n655
  );


  xnor
  g870
  (
    n929,
    n840,
    n846,
    n589,
    n606
  );


  or
  g871
  (
    n961,
    n608,
    n848,
    n850,
    n645
  );


  nand
  g872
  (
    n924,
    n589,
    n641,
    n613,
    n834
  );


  xor
  g873
  (
    n928,
    n841,
    n829,
    n616,
    n591
  );


  and
  g874
  (
    n950,
    n599,
    n612,
    n661,
    n630
  );


  nand
  g875
  (
    n960,
    n835,
    n670,
    n624,
    n843
  );


  or
  g876
  (
    n966,
    n633,
    n884,
    n878,
    n837
  );


  or
  g877
  (
    n935,
    n590,
    n840,
    n648,
    n608
  );


  xor
  g878
  (
    n944,
    n888,
    n634,
    n838,
    n835
  );


  xnor
  g879
  (
    n959,
    n614,
    n883,
    n587,
    n888
  );


  xor
  g880
  (
    n940,
    n880,
    n618,
    n892
  );


  nor
  g881
  (
    n946,
    n651,
    n894,
    n889,
    n847
  );


  xnor
  g882
  (
    n912,
    n883,
    n643,
    n641,
    n607
  );


  or
  g883
  (
    n926,
    n595,
    n889,
    n891,
    n666
  );


  nand
  g884
  (
    n915,
    n640,
    n636,
    n893,
    n885
  );


  and
  g885
  (
    n925,
    n662,
    n883,
    n600,
    n592
  );


  nand
  g886
  (
    n910,
    n639,
    n644,
    n629,
    n619
  );


  or
  g887
  (
    n941,
    n888,
    n617,
    n658,
    n645
  );


  and
  g888
  (
    n916,
    n646,
    n634,
    n653,
    n844
  );


  or
  g889
  (
    n954,
    n887,
    n594,
    n662,
    n881
  );


  and
  g890
  (
    n953,
    n664,
    n660,
    n596,
    n879
  );


  nand
  g891
  (
    n936,
    n602,
    n887,
    n663,
    n603
  );


  or
  g892
  (
    n927,
    n839,
    n650,
    n892,
    n618
  );


  or
  g893
  (
    n938,
    n602,
    n621,
    n639,
    n889
  );


  xor
  g894
  (
    n933,
    n610,
    n667,
    n629
  );


  xor
  g895
  (
    n895,
    n886,
    n839,
    n593,
    n668
  );


  nor
  g896
  (
    n934,
    n615,
    n638,
    n623,
    n614
  );


  nand
  g897
  (
    n939,
    n653,
    n893,
    n624,
    n894
  );


  nand
  g898
  (
    n907,
    n655,
    n627,
    n595,
    n845
  );


  nand
  g899
  (
    n897,
    n834,
    n890,
    n844,
    n601
  );


  xor
  g900
  (
    n955,
    n620,
    n628,
    n654,
    n881
  );


  nor
  g901
  (
    n962,
    n588,
    n887,
    n879,
    n882
  );


  nor
  g902
  (
    n902,
    n836,
    n635,
    n886,
    n831
  );


  xor
  g903
  (
    n919,
    n885,
    n838,
    n831,
    n609
  );


  nor
  g904
  (
    n956,
    n648,
    n833,
    n611,
    n843
  );


  nor
  g905
  (
    n917,
    n633,
    n845,
    n644,
    n591
  );


  and
  g906
  (
    n947,
    n598,
    n878,
    n830,
    n638
  );


  nand
  g907
  (
    n951,
    n848,
    n657,
    n649,
    n877
  );


  xnor
  g908
  (
    n906,
    n851,
    n665,
    n877,
    n829
  );


  and
  g909
  (
    n909,
    n658,
    n647,
    n885,
    n615
  );


  nand
  g910
  (
    n913,
    n877,
    n647,
    n891,
    n850
  );


  and
  g911
  (
    n914,
    n616,
    n890,
    n832,
    n841
  );


  xor
  g912
  (
    n904,
    n836,
    n627,
    n887,
    n652
  );


  xnor
  g913
  (
    n911,
    n664,
    n893,
    n642,
    n886
  );


  buf
  g914
  (
    n990,
    n898
  );


  not
  g915
  (
    n972,
    n900
  );


  not
  g916
  (
    n967,
    n918
  );


  buf
  g917
  (
    n974,
    n916
  );


  buf
  g918
  (
    n975,
    n912
  );


  not
  g919
  (
    n991,
    n917
  );


  not
  g920
  (
    n988,
    n922
  );


  buf
  g921
  (
    n977,
    n914
  );


  buf
  g922
  (
    n982,
    n906
  );


  not
  g923
  (
    n968,
    n903
  );


  buf
  g924
  (
    n978,
    n899
  );


  buf
  g925
  (
    n970,
    n919
  );


  buf
  g926
  (
    n969,
    n897
  );


  buf
  g927
  (
    n987,
    n907
  );


  not
  g928
  (
    n994,
    n913
  );


  not
  g929
  (
    n980,
    n910
  );


  not
  g930
  (
    n986,
    n904
  );


  not
  g931
  (
    n973,
    n908
  );


  buf
  g932
  (
    n983,
    n901
  );


  buf
  g933
  (
    n976,
    n902
  );


  buf
  g934
  (
    n985,
    n896
  );


  buf
  g935
  (
    n984,
    n915
  );


  buf
  g936
  (
    n981,
    n905
  );


  not
  g937
  (
    n993,
    n895
  );


  not
  g938
  (
    n989,
    n909
  );


  buf
  g939
  (
    n971,
    n911
  );


  buf
  g940
  (
    n979,
    n920
  );


  buf
  g941
  (
    n992,
    n921
  );


  xor
  g942
  (
    AntiSAT_key_wire,
    n970,
    n982,
    n441,
    n437
  );


  or
  g943
  (
    n1007,
    n387,
    n438,
    n439,
    n437
  );


  or
  g944
  (
    n1002,
    n441,
    n443,
    n967,
    n439
  );


  xor
  g945
  (
    n1009,
    n438,
    n994,
    n442
  );


  nor
  g946
  (
    n997,
    n440,
    n439,
    n443,
    n444
  );


  xor
  g947
  (
    n1012,
    n974,
    n989,
    n986,
    n981
  );


  xor
  g948
  (
    n999,
    n993,
    n972,
    n439,
    n437
  );


  and
  g949
  (
    n1003,
    n991,
    n442,
    n976,
    n444
  );


  or
  g950
  (
    n1005,
    n442,
    n968,
    n388,
    n985
  );


  nor
  g951
  (
    n1006,
    n988,
    n991,
    n984,
    n388
  );


  xnor
  g952
  (
    n996,
    n438,
    n441,
    n977,
    n993
  );


  xnor
  g953
  (
    n995,
    n992,
    n969,
    n443,
    n990
  );


  nor
  g954
  (
    n998,
    n973,
    n978,
    n983,
    n438
  );


  or
  g955
  (
    n1001,
    n992,
    n979,
    n987,
    n923
  );


  nor
  g956
  (
    n1011,
    n440,
    n994,
    n989,
    n386
  );


  xnor
  g957
  (
    n1010,
    n387,
    n975,
    n443,
    n671
  );


  nor
  g958
  (
    n1000,
    n671,
    n444,
    n980,
    n440
  );


  xor
  g959
  (
    n1008,
    n440,
    n971,
    n441,
    n990
  );


  xor
  g960
  (
    n1023,
    n1006,
    n855,
    n1001,
    n376
  );


  or
  g961
  (
    n1013,
    n856,
    n855,
    n927,
    n940
  );


  xnor
  g962
  (
    n1016,
    n933,
    n376,
    n931,
    n924
  );


  xnor
  g963
  (
    n1025,
    n998,
    n997,
    n852,
    n1008
  );


  nand
  g964
  (
    n1015,
    n1003,
    n929,
    n376
  );


  and
  g965
  (
    n1021,
    n935,
    n853,
    n363,
    n947
  );


  nand
  g966
  (
    n1020,
    n856,
    n925,
    n936,
    n854
  );


  and
  g967
  (
    n1022,
    n1007,
    n943,
    n854,
    n1002
  );


  or
  g968
  (
    n1018,
    n937,
    n945,
    n672,
    n996
  );


  or
  g969
  (
    n1024,
    n942,
    n939,
    n1009,
    n1000
  );


  nor
  g970
  (
    n1017,
    n938,
    n932,
    n672,
    n946
  );


  nand
  g971
  (
    n1026,
    n857,
    n999,
    n944,
    n928
  );


  nand
  g972
  (
    n1014,
    n941,
    n1004,
    n948,
    n1005
  );


  nand
  g973
  (
    n1019,
    n930,
    n934,
    n853,
    n926
  );


  xnor
  g974
  (
    n1027,
    n959,
    n1014,
    n960,
    n954
  );


  xnor
  g975
  (
    n1030,
    n1013,
    n956,
    n950,
    n1014
  );


  xor
  g976
  (
    n1028,
    n952,
    n1013,
    n949,
    n953
  );


  xor
  g977
  (
    n1029,
    n951,
    n955,
    n957,
    n958
  );


  not
  g978
  (
    n1034,
    n1028
  );


  buf
  g979
  (
    n1033,
    n673
  );


  xnor
  g980
  (
    n1031,
    n674,
    n673
  );


  nor
  g981
  (
    n1032,
    n674,
    n1027
  );


  not
  g982
  (
    n1045,
    n866
  );


  buf
  g983
  (
    n1050,
    n52
  );


  buf
  g984
  (
    n1038,
    n388
  );


  buf
  g985
  (
    n1037,
    n1033
  );


  buf
  g986
  (
    n1035,
    n858
  );


  and
  g987
  (
    n1046,
    n866,
    n961,
    n1033
  );


  and
  g988
  (
    n1041,
    n866,
    n1032,
    n388,
    n1034
  );


  xnor
  g989
  (
    n1047,
    n1031,
    n865,
    n1010
  );


  xnor
  g990
  (
    n1040,
    n963,
    n858,
    n864,
    n1012
  );


  xnor
  g991
  (
    n1048,
    n1031,
    n865,
    n864,
    n52
  );


  nor
  g992
  (
    n1044,
    n1034,
    n965,
    n1032,
    n864
  );


  xor
  g993
  (
    n1042,
    n863,
    n1033,
    n964
  );


  xor
  g994
  (
    n1036,
    n1034,
    n857,
    n962,
    n1031
  );


  nand
  g995
  (
    n1043,
    n444,
    n1031,
    n1032,
    n1011
  );


  or
  g996
  (
    n1049,
    n1032,
    n52,
    n1034,
    n863
  );


  nor
  g997
  (
    n1039,
    n866,
    n865,
    n966,
    n864
  );


  or
  g998
  (
    n1061,
    n1043,
    n690,
    n682
  );


  xor
  g999
  (
    n1074,
    n1035,
    n1018,
    n1026,
    n1022
  );


  xor
  g1000
  (
    n1054,
    n676,
    n1042,
    n1020,
    n677
  );


  xnor
  g1001
  (
    n1053,
    n1025,
    n685,
    n1021,
    n1044
  );


  nand
  g1002
  (
    n1057,
    n1019,
    n1044,
    n1049,
    n1020
  );


  nand
  g1003
  (
    n1051,
    n680,
    n1050,
    n682
  );


  nor
  g1004
  (
    n1065,
    n681,
    n1018,
    n1025,
    n1047
  );


  xnor
  g1005
  (
    n1058,
    n1020,
    n683,
    n686,
    n1024
  );


  xnor
  g1006
  (
    n1067,
    n1020,
    n676,
    n686,
    n1017
  );


  or
  g1007
  (
    n1068,
    n689,
    n1017,
    n1025,
    n675
  );


  or
  g1008
  (
    n1066,
    n679,
    n1026,
    n1023,
    n1038
  );


  nand
  g1009
  (
    n1052,
    n1025,
    n1046,
    n1048,
    n1024
  );


  nand
  g1010
  (
    n1060,
    n1024,
    n1021,
    n1022
  );


  and
  g1011
  (
    n1064,
    n1015,
    n683,
    n1023,
    n1049
  );


  xnor
  g1012
  (
    n1070,
    n687,
    n1019,
    n1015,
    n1023
  );


  or
  g1013
  (
    n1062,
    n1037,
    n1021,
    n689,
    n688
  );


  or
  g1014
  (
    n1072,
    n1040,
    n1047,
    n1023,
    n679
  );


  or
  g1015
  (
    n1056,
    n677,
    n1043,
    n1016,
    n1045
  );


  nor
  g1016
  (
    n1055,
    n691,
    n1026,
    n684,
    n688
  );


  or
  g1017
  (
    n1069,
    n1048,
    n685,
    n1026,
    n678
  );


  nand
  g1018
  (
    n1059,
    n684,
    n1021,
    n1022,
    n1036
  );


  nand
  g1019
  (
    n1063,
    n691,
    n681,
    n687,
    n675
  );


  xnor
  g1020
  (
    n1071,
    n1041,
    n1016,
    n1024,
    n1039
  );


  and
  g1021
  (
    n1073,
    n1046,
    n678,
    n1045,
    n680
  );


  nand
  g1022
  (
    n1075,
    n693,
    n695,
    n1029,
    n1028
  );


  nand
  g1023
  (
    n1077,
    n1072,
    n1030,
    n1028,
    n696
  );


  xor
  g1024
  (
    n1076,
    n693,
    n1074,
    n1030,
    n1071
  );


  xnor
  g1025
  (
    n1081,
    n1073,
    n694,
    n692,
    n695
  );


  or
  g1026
  (
    n1080,
    n1069,
    n694,
    n692,
    n1028
  );


  nor
  g1027
  (
    n1079,
    n1030,
    n1030,
    n1070,
    n696
  );


  xnor
  g1028
  (
    n1078,
    n1068,
    n1029
  );


  not
  g1029
  (
    n1083,
    n1075
  );


  not
  g1030
  (
    n1082,
    n1075
  );


  xor
  g1031
  (
    n1091,
    n702,
    n707,
    n1082,
    n705
  );


  nor
  g1032
  (
    n1087,
    n700,
    n1083,
    n701,
    n704
  );


  or
  g1033
  (
    n1088,
    n698,
    n704,
    n701,
    n699
  );


  and
  g1034
  (
    n1086,
    n1083,
    n1082,
    n706
  );


  nand
  g1035
  (
    n1085,
    n700,
    n707,
    n697,
    n699
  );


  nand
  g1036
  (
    n1084,
    n708,
    n703,
    n697
  );


  and
  g1037
  (
    n1089,
    n702,
    n1082,
    n708,
    n705
  );


  or
  g1038
  (
    n1090,
    n698,
    n706,
    n1083
  );


  xnor
  g1039
  (
    n1110,
    n1085,
    n712,
    n741,
    n1090
  );


  and
  g1040
  (
    n1103,
    n729,
    n718,
    n736,
    n745
  );


  nand
  g1041
  (
    n1092,
    n1085,
    n732,
    n731,
    n1076
  );


  xnor
  g1042
  (
    n1111,
    n745,
    n719,
    n1081,
    n1078
  );


  xor
  g1043
  (
    n1100,
    n1078,
    n746,
    n747,
    n1091
  );


  nor
  g1044
  (
    n1112,
    n746,
    n1081,
    n727,
    n738
  );


  nor
  g1045
  (
    n1105,
    n712,
    n735,
    n1085,
    n1077
  );


  xnor
  g1046
  (
    n1114,
    n711,
    n711,
    n1086,
    n729
  );


  or
  g1047
  (
    n1119,
    n1088,
    n715,
    n1084
  );


  xnor
  g1048
  (
    n1106,
    n717,
    n740,
    n1089,
    n731
  );


  nand
  g1049
  (
    n1104,
    n1087,
    n1091,
    n1089,
    n1084
  );


  or
  g1050
  (
    n1120,
    n1086,
    n1080,
    n737,
    n747
  );


  xnor
  g1051
  (
    n1109,
    n718,
    n710,
    n744
  );


  or
  g1052
  (
    n1122,
    n728,
    n733,
    n1086
  );


  xor
  g1053
  (
    n1097,
    n742,
    n713,
    n734,
    n730
  );


  xnor
  g1054
  (
    n1101,
    n717,
    n1091,
    n716,
    n724
  );


  xnor
  g1055
  (
    n1094,
    n1091,
    n726,
    n734,
    n1077
  );


  nand
  g1056
  (
    n1116,
    n1076,
    n742,
    n730,
    n728
  );


  xor
  g1057
  (
    n1115,
    n1089,
    n741,
    n721,
    n1090
  );


  xnor
  g1058
  (
    n1118,
    n1088,
    n716,
    n723,
    n714
  );


  xor
  g1059
  (
    n1095,
    n1087,
    n1086,
    n1081,
    n710
  );


  and
  g1060
  (
    n1096,
    n721,
    n713,
    n738,
    n1090
  );


  and
  g1061
  (
    n1098,
    n719,
    n743,
    n1079
  );


  or
  g1062
  (
    n1108,
    n709,
    n714,
    n720,
    n1085
  );


  nor
  g1063
  (
    n1107,
    n746,
    n724,
    n723,
    n737
  );


  or
  g1064
  (
    n1123,
    n722,
    n740,
    n735,
    n732
  );


  or
  g1065
  (
    n1113,
    n722,
    n1084,
    n746,
    n747
  );


  or
  g1066
  (
    n1102,
    n1080,
    n743,
    n747,
    n720
  );


  and
  g1067
  (
    n1121,
    n1087,
    n736,
    n1089,
    n1090
  );


  xnor
  g1068
  (
    n1099,
    n715,
    n739,
    n1087,
    n725
  );


  xor
  g1069
  (
    n1093,
    n1088,
    n727,
    n726,
    n709
  );


  xnor
  g1070
  (
    n1117,
    n1088,
    n725,
    n739,
    n1081
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_0,
    keyIn_0_52,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_1,
    keyIn_0_53,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_2,
    keyIn_0_54,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_3,
    keyIn_0_55,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_4,
    keyIn_0_56,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_5,
    keyIn_0_57,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_6,
    keyIn_0_58,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_7,
    keyIn_0_59,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_8,
    keyIn_0_60,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_9,
    keyIn_0_61,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_10,
    keyIn_0_62,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_11,
    keyIn_0_63,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_64
  (
    gbar_input_0_12,
    keyIn_0_64,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_65
  (
    gbar_input_0_13,
    keyIn_0_65,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_66
  (
    gbar_input_0_14,
    keyIn_0_66,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_67
  (
    gbar_input_0_15,
    keyIn_0_67,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_68
  (
    gbar_input_0_16,
    keyIn_0_68,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_69
  (
    gbar_input_0_17,
    keyIn_0_69,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_70
  (
    gbar_input_0_18,
    keyIn_0_70,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_71
  (
    gbar_input_0_19,
    keyIn_0_71,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_72
  (
    gbar_input_0_20,
    keyIn_0_72,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_73
  (
    gbar_input_0_21,
    keyIn_0_73,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_74
  (
    gbar_input_0_22,
    keyIn_0_74,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_75
  (
    gbar_input_0_23,
    keyIn_0_75,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_76
  (
    gbar_input_0_24,
    keyIn_0_76,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_77
  (
    gbar_input_0_25,
    keyIn_0_77,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_78
  (
    gbar_input_0_26,
    keyIn_0_78,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_79
  (
    gbar_input_0_27,
    keyIn_0_79,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_80
  (
    gbar_input_0_28,
    keyIn_0_80,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_81
  (
    gbar_input_0_29,
    keyIn_0_81,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_82
  (
    gbar_input_0_30,
    keyIn_0_82,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_83
  (
    gbar_input_0_31,
    keyIn_0_83,
    n32
  );


  xor
  KeyPIGate_0_32
  (
    g_input_0_32,
    keyIn_0_32,
    n33
  );


  xor
  KeyPIGate_0_84
  (
    gbar_input_0_32,
    keyIn_0_84,
    n33
  );


  xor
  KeyPIGate_0_33
  (
    g_input_0_33,
    keyIn_0_33,
    n34
  );


  xor
  KeyPIGate_0_85
  (
    gbar_input_0_33,
    keyIn_0_85,
    n34
  );


  xor
  KeyPIGate_0_34
  (
    g_input_0_34,
    keyIn_0_34,
    n35
  );


  xor
  KeyPIGate_0_86
  (
    gbar_input_0_34,
    keyIn_0_86,
    n35
  );


  xor
  KeyPIGate_0_35
  (
    g_input_0_35,
    keyIn_0_35,
    n36
  );


  xor
  KeyPIGate_0_87
  (
    gbar_input_0_35,
    keyIn_0_87,
    n36
  );


  xor
  KeyPIGate_0_36
  (
    g_input_0_36,
    keyIn_0_36,
    n37
  );


  xor
  KeyPIGate_0_88
  (
    gbar_input_0_36,
    keyIn_0_88,
    n37
  );


  xor
  KeyPIGate_0_37
  (
    g_input_0_37,
    keyIn_0_37,
    n38
  );


  xor
  KeyPIGate_0_89
  (
    gbar_input_0_37,
    keyIn_0_89,
    n38
  );


  xor
  KeyPIGate_0_38
  (
    g_input_0_38,
    keyIn_0_38,
    n39
  );


  xor
  KeyPIGate_0_90
  (
    gbar_input_0_38,
    keyIn_0_90,
    n39
  );


  xor
  KeyPIGate_0_39
  (
    g_input_0_39,
    keyIn_0_39,
    n40
  );


  xor
  KeyPIGate_0_91
  (
    gbar_input_0_39,
    keyIn_0_91,
    n40
  );


  xor
  KeyPIGate_0_40
  (
    g_input_0_40,
    keyIn_0_40,
    n41
  );


  xor
  KeyPIGate_0_92
  (
    gbar_input_0_40,
    keyIn_0_92,
    n41
  );


  xor
  KeyPIGate_0_41
  (
    g_input_0_41,
    keyIn_0_41,
    n42
  );


  xor
  KeyPIGate_0_93
  (
    gbar_input_0_41,
    keyIn_0_93,
    n42
  );


  xor
  KeyPIGate_0_42
  (
    g_input_0_42,
    keyIn_0_42,
    n43
  );


  xor
  KeyPIGate_0_94
  (
    gbar_input_0_42,
    keyIn_0_94,
    n43
  );


  xor
  KeyPIGate_0_43
  (
    g_input_0_43,
    keyIn_0_43,
    n44
  );


  xor
  KeyPIGate_0_95
  (
    gbar_input_0_43,
    keyIn_0_95,
    n44
  );


  xor
  KeyPIGate_0_44
  (
    g_input_0_44,
    keyIn_0_44,
    n45
  );


  xor
  KeyPIGate_0_96
  (
    gbar_input_0_44,
    keyIn_0_96,
    n45
  );


  xor
  KeyPIGate_0_45
  (
    g_input_0_45,
    keyIn_0_45,
    n46
  );


  xor
  KeyPIGate_0_97
  (
    gbar_input_0_45,
    keyIn_0_97,
    n46
  );


  xor
  KeyPIGate_0_46
  (
    g_input_0_46,
    keyIn_0_46,
    n47
  );


  xor
  KeyPIGate_0_98
  (
    gbar_input_0_46,
    keyIn_0_98,
    n47
  );


  xor
  KeyPIGate_0_47
  (
    g_input_0_47,
    keyIn_0_47,
    n48
  );


  xor
  KeyPIGate_0_99
  (
    gbar_input_0_47,
    keyIn_0_99,
    n48
  );


  xor
  KeyPIGate_0_48
  (
    g_input_0_48,
    keyIn_0_48,
    n49
  );


  xor
  KeyPIGate_0_100
  (
    gbar_input_0_48,
    keyIn_0_100,
    n49
  );


  xor
  KeyPIGate_0_49
  (
    g_input_0_49,
    keyIn_0_49,
    n50
  );


  xor
  KeyPIGate_0_101
  (
    gbar_input_0_49,
    keyIn_0_101,
    n50
  );


  xor
  KeyPIGate_0_50
  (
    g_input_0_50,
    keyIn_0_50,
    n51
  );


  xor
  KeyPIGate_0_102
  (
    gbar_input_0_50,
    keyIn_0_102,
    n51
  );


  xor
  KeyPIGate_0_51
  (
    g_input_0_51,
    keyIn_0_51,
    n52
  );


  xor
  KeyPIGate_0_103
  (
    gbar_input_0_51,
    keyIn_0_103,
    n52
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31,
    g_input_0_32,
    g_input_0_33,
    g_input_0_34,
    g_input_0_35,
    g_input_0_36,
    g_input_0_37,
    g_input_0_38,
    g_input_0_39,
    g_input_0_40,
    g_input_0_41,
    g_input_0_42,
    g_input_0_43,
    g_input_0_44,
    g_input_0_45,
    g_input_0_46,
    g_input_0_47,
    g_input_0_48,
    g_input_0_49,
    g_input_0_50,
    g_input_0_51
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31,
    gbar_input_0_32,
    gbar_input_0_33,
    gbar_input_0_34,
    gbar_input_0_35,
    gbar_input_0_36,
    gbar_input_0_37,
    gbar_input_0_38,
    gbar_input_0_39,
    gbar_input_0_40,
    gbar_input_0_41,
    gbar_input_0_42,
    gbar_input_0_43,
    gbar_input_0_44,
    gbar_input_0_45,
    gbar_input_0_46,
    gbar_input_0_47,
    gbar_input_0_48,
    gbar_input_0_49,
    gbar_input_0_50,
    gbar_input_0_51
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n1004,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

