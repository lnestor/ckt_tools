

module Stat_1426_22_3
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n566,
  n580,
  n570,
  n588,
  n582,
  n587,
  n572,
  n571,
  n584,
  n585,
  n586,
  n577,
  n565,
  n564,
  n1451,
  n1446,
  n1448,
  n1450,
  n1449,
  n1447,
  n1444,
  n1445
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n566;output n580;output n570;output n588;output n582;output n587;output n572;output n571;output n584;output n585;output n586;output n577;output n565;output n564;output n1451;output n1446;output n1448;output n1450;output n1449;output n1447;output n1444;output n1445;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n567;wire n568;wire n569;wire n573;wire n574;wire n575;wire n576;wire n578;wire n579;wire n581;wire n583;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  buf
  g0
  (
    n73,
    n18
  );


  not
  g1
  (
    n62,
    n11
  );


  not
  g2
  (
    n116,
    n10
  );


  not
  g3
  (
    n108,
    n23
  );


  not
  g4
  (
    n29,
    n23
  );


  not
  g5
  (
    n122,
    n14
  );


  buf
  g6
  (
    n106,
    n21
  );


  buf
  g7
  (
    n68,
    n3
  );


  buf
  g8
  (
    n51,
    n16
  );


  buf
  g9
  (
    n102,
    n5
  );


  buf
  g10
  (
    n100,
    n20
  );


  not
  g11
  (
    n47,
    n4
  );


  buf
  g12
  (
    n82,
    n25
  );


  not
  g13
  (
    n52,
    n18
  );


  buf
  g14
  (
    n53,
    n25
  );


  buf
  g15
  (
    KeyWire_0_10,
    n9
  );


  buf
  g16
  (
    n75,
    n21
  );


  buf
  g17
  (
    n84,
    n11
  );


  buf
  g18
  (
    n77,
    n14
  );


  buf
  g19
  (
    n44,
    n4
  );


  buf
  g20
  (
    n87,
    n2
  );


  buf
  g21
  (
    n37,
    n5
  );


  not
  g22
  (
    n54,
    n7
  );


  buf
  g23
  (
    n70,
    n9
  );


  not
  g24
  (
    n40,
    n2
  );


  not
  g25
  (
    n121,
    n21
  );


  not
  g26
  (
    n115,
    n16
  );


  buf
  g27
  (
    n98,
    n10
  );


  not
  g28
  (
    n72,
    n7
  );


  buf
  g29
  (
    n34,
    n4
  );


  not
  g30
  (
    n113,
    n17
  );


  not
  g31
  (
    n120,
    n19
  );


  buf
  g32
  (
    n86,
    n15
  );


  not
  g33
  (
    n55,
    n1
  );


  not
  g34
  (
    n32,
    n18
  );


  buf
  g35
  (
    n78,
    n14
  );


  not
  g36
  (
    n110,
    n22
  );


  not
  g37
  (
    n63,
    n1
  );


  buf
  g38
  (
    n83,
    n15
  );


  buf
  g39
  (
    n26,
    n6
  );


  not
  g40
  (
    n27,
    n21
  );


  not
  g41
  (
    n80,
    n10
  );


  not
  g42
  (
    n69,
    n5
  );


  not
  g43
  (
    n124,
    n19
  );


  not
  g44
  (
    n58,
    n4
  );


  not
  g45
  (
    n88,
    n7
  );


  buf
  g46
  (
    n125,
    n23
  );


  buf
  g47
  (
    n90,
    n16
  );


  not
  g48
  (
    n71,
    n3
  );


  buf
  g49
  (
    n96,
    n3
  );


  buf
  g50
  (
    n101,
    n22
  );


  not
  g51
  (
    n109,
    n8
  );


  buf
  g52
  (
    n45,
    n9
  );


  not
  g53
  (
    n38,
    n19
  );


  not
  g54
  (
    n65,
    n15
  );


  not
  g55
  (
    n57,
    n24
  );


  not
  g56
  (
    n111,
    n2
  );


  not
  g57
  (
    n93,
    n24
  );


  not
  g58
  (
    n60,
    n12
  );


  not
  g59
  (
    n81,
    n24
  );


  not
  g60
  (
    n107,
    n11
  );


  not
  g61
  (
    n36,
    n17
  );


  not
  g62
  (
    n33,
    n12
  );


  not
  g63
  (
    n66,
    n9
  );


  not
  g64
  (
    n28,
    n12
  );


  buf
  g65
  (
    n31,
    n1
  );


  not
  g66
  (
    n91,
    n13
  );


  buf
  g67
  (
    n117,
    n5
  );


  not
  g68
  (
    n105,
    n11
  );


  buf
  g69
  (
    n74,
    n13
  );


  not
  g70
  (
    n97,
    n6
  );


  buf
  g71
  (
    n56,
    n3
  );


  buf
  g72
  (
    n94,
    n2
  );


  not
  g73
  (
    n99,
    n6
  );


  buf
  g74
  (
    n76,
    n14
  );


  buf
  g75
  (
    n79,
    n10
  );


  buf
  g76
  (
    n85,
    n7
  );


  buf
  g77
  (
    n64,
    n16
  );


  buf
  g78
  (
    n112,
    n22
  );


  buf
  g79
  (
    n119,
    n13
  );


  buf
  g80
  (
    n30,
    n20
  );


  not
  g81
  (
    n46,
    n24
  );


  buf
  g82
  (
    n95,
    n18
  );


  buf
  g83
  (
    n42,
    n1
  );


  not
  g84
  (
    n49,
    n17
  );


  not
  g85
  (
    n123,
    n23
  );


  buf
  g86
  (
    n118,
    n19
  );


  buf
  g87
  (
    KeyWire_0_2,
    n12
  );


  not
  g88
  (
    n104,
    n6
  );


  buf
  g89
  (
    n103,
    n22
  );


  not
  g90
  (
    n35,
    n8
  );


  buf
  g91
  (
    n48,
    n17
  );


  buf
  g92
  (
    n39,
    n15
  );


  buf
  g93
  (
    n43,
    n25
  );


  not
  g94
  (
    n114,
    n8
  );


  buf
  g95
  (
    n61,
    n25
  );


  not
  g96
  (
    n67,
    n8
  );


  buf
  g97
  (
    n41,
    n20
  );


  buf
  g98
  (
    n92,
    n20
  );


  buf
  g99
  (
    n50,
    n13
  );


  not
  g100
  (
    n193,
    n91
  );


  not
  g101
  (
    n152,
    n124
  );


  not
  g102
  (
    n129,
    n66
  );


  not
  g103
  (
    n134,
    n75
  );


  buf
  g104
  (
    n159,
    n36
  );


  buf
  g105
  (
    n203,
    n36
  );


  buf
  g106
  (
    n163,
    n67
  );


  buf
  g107
  (
    n138,
    n39
  );


  buf
  g108
  (
    n149,
    n67
  );


  not
  g109
  (
    n237,
    n44
  );


  not
  g110
  (
    n166,
    n77
  );


  buf
  g111
  (
    n183,
    n27
  );


  not
  g112
  (
    n180,
    n118
  );


  not
  g113
  (
    n214,
    n108
  );


  buf
  g114
  (
    n228,
    n34
  );


  not
  g115
  (
    n208,
    n78
  );


  buf
  g116
  (
    n215,
    n34
  );


  buf
  g117
  (
    n241,
    n37
  );


  not
  g118
  (
    n187,
    n81
  );


  buf
  g119
  (
    n195,
    n98
  );


  buf
  g120
  (
    n229,
    n101
  );


  not
  g121
  (
    n133,
    n96
  );


  buf
  g122
  (
    n179,
    n82
  );


  buf
  g123
  (
    n234,
    n41
  );


  buf
  g124
  (
    n168,
    n111
  );


  not
  g125
  (
    n258,
    n26
  );


  not
  g126
  (
    n225,
    n84
  );


  buf
  g127
  (
    n142,
    n48
  );


  buf
  g128
  (
    n233,
    n97
  );


  not
  g129
  (
    n167,
    n43
  );


  buf
  g130
  (
    n242,
    n71
  );


  buf
  g131
  (
    n252,
    n40
  );


  not
  g132
  (
    n217,
    n73
  );


  not
  g133
  (
    n197,
    n123
  );


  buf
  g134
  (
    n137,
    n125
  );


  buf
  g135
  (
    n169,
    n40
  );


  not
  g136
  (
    n190,
    n37
  );


  buf
  g137
  (
    n249,
    n115
  );


  not
  g138
  (
    n223,
    n78
  );


  buf
  g139
  (
    n143,
    n71
  );


  buf
  g140
  (
    n165,
    n124
  );


  not
  g141
  (
    n236,
    n122
  );


  buf
  g142
  (
    n256,
    n105
  );


  not
  g143
  (
    n262,
    n76
  );


  buf
  g144
  (
    n182,
    n75
  );


  not
  g145
  (
    n186,
    n120
  );


  buf
  g146
  (
    n191,
    n124
  );


  buf
  g147
  (
    n176,
    n119
  );


  and
  g148
  (
    n254,
    n123,
    n120
  );


  xor
  g149
  (
    n220,
    n35,
    n29
  );


  xor
  g150
  (
    n181,
    n81,
    n119,
    n93,
    n92
  );


  xor
  g151
  (
    n170,
    n102,
    n45,
    n77,
    n62
  );


  and
  g152
  (
    n157,
    n70,
    n38,
    n32
  );


  nor
  g153
  (
    n243,
    n52,
    n104,
    n116,
    n57
  );


  nand
  g154
  (
    n216,
    n55,
    n99,
    n82,
    n121
  );


  or
  g155
  (
    n206,
    n81,
    n62,
    n98,
    n65
  );


  or
  g156
  (
    n148,
    n73,
    n28,
    n48,
    n37
  );


  and
  g157
  (
    n257,
    n124,
    n121,
    n106,
    n107
  );


  and
  g158
  (
    n199,
    n103,
    n47,
    n42,
    n91
  );


  or
  g159
  (
    n255,
    n32,
    n112,
    n104,
    n59
  );


  nor
  g160
  (
    n218,
    n59,
    n105,
    n28,
    n69
  );


  nand
  g161
  (
    n146,
    n53,
    n69,
    n82,
    n83
  );


  xnor
  g162
  (
    n158,
    n95,
    n47,
    n99,
    n48
  );


  xor
  g163
  (
    n156,
    n81,
    n54,
    n107,
    n31
  );


  xnor
  g164
  (
    n202,
    n29,
    n92,
    n112,
    n49
  );


  nand
  g165
  (
    n160,
    n46,
    n44,
    n78,
    n65
  );


  xnor
  g166
  (
    n147,
    n63,
    n94,
    n67,
    n33
  );


  and
  g167
  (
    n232,
    n68,
    n40,
    n62,
    n109
  );


  nor
  g168
  (
    n161,
    n38,
    n68,
    n58,
    n47
  );


  xor
  g169
  (
    n230,
    n85,
    n58,
    n101,
    n59
  );


  or
  g170
  (
    n200,
    n53,
    n108,
    n70,
    n35
  );


  xnor
  g171
  (
    n194,
    n56,
    n41,
    n100,
    n97
  );


  and
  g172
  (
    n178,
    n55,
    n84,
    n54,
    n112
  );


  xor
  g173
  (
    n185,
    n105,
    n52,
    n74,
    n35
  );


  xor
  g174
  (
    n189,
    n95,
    n105,
    n76,
    n67
  );


  xor
  g175
  (
    n177,
    n38,
    n114,
    n50,
    n107
  );


  nor
  g176
  (
    n150,
    n46,
    n36,
    n97,
    n99
  );


  xnor
  g177
  (
    n204,
    n62,
    n97,
    n88,
    n83
  );


  or
  g178
  (
    n201,
    n43,
    n74,
    n103,
    n46
  );


  xor
  g179
  (
    n126,
    n84,
    n26,
    n45,
    n65
  );


  xor
  g180
  (
    n198,
    n94,
    n87,
    n56,
    n42
  );


  xnor
  g181
  (
    n211,
    n65,
    n64,
    n49,
    n70
  );


  xnor
  g182
  (
    n131,
    n27,
    n30,
    n33,
    n28
  );


  nor
  g183
  (
    n132,
    n76,
    n90,
    n87,
    n96
  );


  xor
  g184
  (
    n196,
    n39,
    n84,
    n85,
    n94
  );


  xor
  g185
  (
    n184,
    n54,
    n27,
    n61,
    n119
  );


  nand
  g186
  (
    n136,
    n90,
    n42,
    n72,
    n86
  );


  xnor
  g187
  (
    n227,
    n44,
    n125,
    n85,
    n86
  );


  or
  g188
  (
    n238,
    n125,
    n117,
    n89,
    n63
  );


  and
  g189
  (
    n154,
    n117,
    n55,
    n53,
    n101
  );


  or
  g190
  (
    n250,
    n94,
    n71,
    n113,
    n111
  );


  xnor
  g191
  (
    n128,
    n106,
    n101,
    n95,
    n107
  );


  nand
  g192
  (
    n192,
    n51,
    n117,
    n119,
    n28
  );


  nand
  g193
  (
    n153,
    n96,
    n104,
    n30,
    n43
  );


  nand
  g194
  (
    n210,
    n52,
    n100,
    n41,
    n115
  );


  nor
  g195
  (
    n219,
    n92,
    n118,
    n122,
    n47
  );


  and
  g196
  (
    n248,
    n59,
    n52,
    n34,
    n79
  );


  and
  g197
  (
    n239,
    n80,
    n122,
    n120,
    n61
  );


  xor
  g198
  (
    n144,
    n108,
    n43,
    n111,
    n39
  );


  nand
  g199
  (
    n226,
    n111,
    n80,
    n102
  );


  nand
  g200
  (
    n173,
    n56,
    n64,
    n85,
    n75
  );


  or
  g201
  (
    n205,
    n93,
    n66,
    n30,
    n63
  );


  and
  g202
  (
    n175,
    n90,
    n39,
    n118,
    n79
  );


  nor
  g203
  (
    n140,
    n51,
    n32,
    n83,
    n46
  );


  nor
  g204
  (
    n259,
    n113,
    n70,
    n61,
    n110
  );


  nand
  g205
  (
    n253,
    n121,
    n40,
    n29,
    n123
  );


  nand
  g206
  (
    n139,
    n109,
    n72,
    n49,
    n114
  );


  and
  g207
  (
    n127,
    n51,
    n102,
    n26,
    n77
  );


  or
  g208
  (
    n246,
    n31,
    n116,
    n75,
    n76
  );


  or
  g209
  (
    n174,
    n63,
    n95,
    n56,
    n112
  );


  and
  g210
  (
    n240,
    n87,
    n123,
    n89,
    n50
  );


  xor
  g211
  (
    n155,
    n58,
    n27,
    n106,
    n83
  );


  or
  g212
  (
    n222,
    n69,
    n103,
    n86,
    n115
  );


  xnor
  g213
  (
    n235,
    n33,
    n78,
    n98,
    n66
  );


  xnor
  g214
  (
    n135,
    n50,
    n44,
    n79,
    n114
  );


  and
  g215
  (
    n244,
    n60,
    n72,
    n45,
    n96
  );


  xor
  g216
  (
    n209,
    n36,
    n30,
    n116,
    n61
  );


  or
  g217
  (
    n245,
    n60,
    n64,
    n68,
    n80
  );


  nand
  g218
  (
    n172,
    n117,
    n33,
    n31
  );


  xor
  g219
  (
    n162,
    n58,
    n53,
    n73,
    n66
  );


  nand
  g220
  (
    n151,
    n93,
    n89,
    n48,
    n42
  );


  nand
  g221
  (
    n231,
    n89,
    n79,
    n26,
    n103
  );


  nor
  g222
  (
    n261,
    n125,
    n32,
    n88,
    n109
  );


  nor
  g223
  (
    n188,
    n34,
    n113,
    n45,
    n102
  );


  or
  g224
  (
    n224,
    n122,
    n41,
    n88,
    n55
  );


  nand
  g225
  (
    n212,
    n57,
    n115,
    n72,
    n71
  );


  and
  g226
  (
    n221,
    n57,
    n108,
    n64,
    n116
  );


  and
  g227
  (
    n171,
    n91,
    n74,
    n100,
    n29
  );


  or
  g228
  (
    n213,
    n109,
    n74,
    n37,
    n86
  );


  and
  g229
  (
    n130,
    n104,
    n77,
    n106,
    n110
  );


  xnor
  g230
  (
    n247,
    n99,
    n51,
    n69,
    n98
  );


  and
  g231
  (
    n207,
    n87,
    n120,
    n93,
    n60
  );


  and
  g232
  (
    n145,
    n35,
    n91,
    n73,
    n114
  );


  and
  g233
  (
    n164,
    n54,
    n57,
    n68,
    n121
  );


  or
  g234
  (
    n141,
    n49,
    n118,
    n110,
    n60
  );


  or
  g235
  (
    n251,
    n88,
    n110,
    n82,
    n100
  );


  nor
  g236
  (
    n260,
    n113,
    n50,
    n90,
    n92
  );


  buf
  g237
  (
    n285,
    n168
  );


  not
  g238
  (
    n264,
    n136
  );


  buf
  g239
  (
    n281,
    n156
  );


  not
  g240
  (
    n284,
    n161
  );


  not
  g241
  (
    n266,
    n181
  );


  buf
  g242
  (
    n273,
    n167
  );


  buf
  g243
  (
    n283,
    n147
  );


  buf
  g244
  (
    n279,
    n174
  );


  not
  g245
  (
    n280,
    n148
  );


  buf
  g246
  (
    n267,
    n164
  );


  buf
  g247
  (
    n268,
    n163
  );


  buf
  g248
  (
    n282,
    n137
  );


  not
  g249
  (
    n263,
    n138
  );


  buf
  g250
  (
    n288,
    n151
  );


  not
  g251
  (
    n287,
    n177
  );


  buf
  g252
  (
    n275,
    n175
  );


  not
  g253
  (
    n286,
    n165
  );


  not
  g254
  (
    n274,
    n129
  );


  xor
  g255
  (
    n269,
    n127,
    n170
  );


  nand
  g256
  (
    n272,
    n173,
    n128,
    n153,
    n141
  );


  xor
  g257
  (
    n278,
    n176,
    n134,
    n139,
    n152
  );


  or
  g258
  (
    n270,
    n130,
    n132,
    n166,
    n169
  );


  xnor
  g259
  (
    n289,
    n154,
    n135,
    n149,
    n144
  );


  nor
  g260
  (
    n290,
    n140,
    n155,
    n133,
    n142
  );


  xnor
  g261
  (
    n265,
    n126,
    n143,
    n160,
    n178
  );


  xor
  g262
  (
    n277,
    n131,
    n179,
    n146,
    n158
  );


  nand
  g263
  (
    n271,
    n172,
    n162,
    n150,
    n180
  );


  nand
  g264
  (
    n276,
    n157,
    n145,
    n171,
    n159
  );


  not
  g265
  (
    n304,
    n282
  );


  not
  g266
  (
    n293,
    n275
  );


  not
  g267
  (
    n321,
    n279
  );


  buf
  g268
  (
    n320,
    n281
  );


  not
  g269
  (
    n314,
    n273
  );


  not
  g270
  (
    n317,
    n269
  );


  buf
  g271
  (
    n309,
    n268
  );


  not
  g272
  (
    n300,
    n283
  );


  buf
  g273
  (
    n307,
    n277
  );


  buf
  g274
  (
    n318,
    n276
  );


  buf
  g275
  (
    n316,
    n281
  );


  buf
  g276
  (
    n291,
    n271
  );


  buf
  g277
  (
    n302,
    n283
  );


  not
  g278
  (
    n322,
    n284
  );


  not
  g279
  (
    n305,
    n281
  );


  buf
  g280
  (
    n296,
    n281
  );


  not
  g281
  (
    n310,
    n274
  );


  not
  g282
  (
    n306,
    n263
  );


  buf
  g283
  (
    n292,
    n272
  );


  buf
  g284
  (
    n319,
    n283
  );


  buf
  g285
  (
    n297,
    n278
  );


  not
  g286
  (
    n315,
    n266
  );


  not
  g287
  (
    n311,
    n282
  );


  buf
  g288
  (
    n298,
    n282
  );


  not
  g289
  (
    n295,
    n270
  );


  buf
  g290
  (
    n303,
    n264
  );


  not
  g291
  (
    n312,
    n283
  );


  buf
  g292
  (
    n308,
    n267
  );


  buf
  g293
  (
    n299,
    n282
  );


  buf
  g294
  (
    n301,
    n280
  );


  buf
  g295
  (
    n294,
    n284
  );


  buf
  g296
  (
    n313,
    n265
  );


  not
  g297
  (
    n365,
    n318
  );


  buf
  g298
  (
    n430,
    n292
  );


  buf
  g299
  (
    n397,
    n304
  );


  buf
  g300
  (
    n390,
    n300
  );


  not
  g301
  (
    n413,
    n303
  );


  not
  g302
  (
    n352,
    n308
  );


  not
  g303
  (
    n331,
    n316
  );


  not
  g304
  (
    n429,
    n314
  );


  buf
  g305
  (
    n363,
    n307
  );


  not
  g306
  (
    n404,
    n317
  );


  not
  g307
  (
    n392,
    n308
  );


  buf
  g308
  (
    n376,
    n296
  );


  not
  g309
  (
    n423,
    n302
  );


  buf
  g310
  (
    n426,
    n293
  );


  not
  g311
  (
    n444,
    n306
  );


  not
  g312
  (
    n389,
    n305
  );


  not
  g313
  (
    n326,
    n291
  );


  not
  g314
  (
    n338,
    n300
  );


  buf
  g315
  (
    n417,
    n311
  );


  buf
  g316
  (
    n373,
    n309
  );


  buf
  g317
  (
    n341,
    n322
  );


  not
  g318
  (
    n327,
    n313
  );


  not
  g319
  (
    n324,
    n317
  );


  not
  g320
  (
    n437,
    n295
  );


  buf
  g321
  (
    n332,
    n315
  );


  buf
  g322
  (
    n328,
    n293
  );


  not
  g323
  (
    n408,
    n299
  );


  buf
  g324
  (
    n371,
    n314
  );


  buf
  g325
  (
    n435,
    n318
  );


  buf
  g326
  (
    n368,
    n312
  );


  not
  g327
  (
    n353,
    n305
  );


  buf
  g328
  (
    n386,
    n297
  );


  buf
  g329
  (
    n336,
    n295
  );


  not
  g330
  (
    n391,
    n315
  );


  not
  g331
  (
    n401,
    n299
  );


  not
  g332
  (
    n334,
    n297
  );


  not
  g333
  (
    n337,
    n315
  );


  buf
  g334
  (
    n323,
    n320
  );


  buf
  g335
  (
    n333,
    n312
  );


  buf
  g336
  (
    n395,
    n303
  );


  not
  g337
  (
    n406,
    n297
  );


  not
  g338
  (
    n346,
    n321
  );


  not
  g339
  (
    n424,
    n305
  );


  not
  g340
  (
    n385,
    n305
  );


  not
  g341
  (
    n340,
    n320
  );


  not
  g342
  (
    n374,
    n311
  );


  not
  g343
  (
    n440,
    n301
  );


  buf
  g344
  (
    n358,
    n295
  );


  not
  g345
  (
    n414,
    n321
  );


  not
  g346
  (
    n416,
    n319
  );


  buf
  g347
  (
    n428,
    n312
  );


  buf
  g348
  (
    n402,
    n321
  );


  buf
  g349
  (
    n394,
    n306
  );


  buf
  g350
  (
    n356,
    n298
  );


  buf
  g351
  (
    n357,
    n293
  );


  not
  g352
  (
    n359,
    n313
  );


  buf
  g353
  (
    n396,
    n296
  );


  buf
  g354
  (
    n375,
    n294
  );


  not
  g355
  (
    n329,
    n313
  );


  buf
  g356
  (
    n364,
    n314
  );


  not
  g357
  (
    n432,
    n303
  );


  not
  g358
  (
    n399,
    n292
  );


  not
  g359
  (
    n398,
    n320
  );


  buf
  g360
  (
    n403,
    n316
  );


  buf
  g361
  (
    n438,
    n318
  );


  buf
  g362
  (
    n382,
    n306
  );


  buf
  g363
  (
    n427,
    n307
  );


  buf
  g364
  (
    n409,
    n312
  );


  buf
  g365
  (
    n446,
    n307
  );


  buf
  g366
  (
    n445,
    n302
  );


  buf
  g367
  (
    n367,
    n294
  );


  buf
  g368
  (
    n342,
    n313
  );


  not
  g369
  (
    n348,
    n300
  );


  not
  g370
  (
    n441,
    n318
  );


  not
  g371
  (
    n379,
    n317
  );


  not
  g372
  (
    n443,
    n309
  );


  buf
  g373
  (
    n330,
    n304
  );


  buf
  g374
  (
    n354,
    n309
  );


  buf
  g375
  (
    n349,
    n307
  );


  buf
  g376
  (
    n422,
    n298
  );


  not
  g377
  (
    n378,
    n299
  );


  buf
  g378
  (
    n344,
    n291
  );


  not
  g379
  (
    n347,
    n322
  );


  buf
  g380
  (
    n339,
    n319
  );


  not
  g381
  (
    n405,
    n309
  );


  not
  g382
  (
    n425,
    n321
  );


  buf
  g383
  (
    n418,
    n315
  );


  not
  g384
  (
    n433,
    n302
  );


  not
  g385
  (
    n345,
    n308
  );


  buf
  g386
  (
    n370,
    n292
  );


  not
  g387
  (
    n335,
    n304
  );


  buf
  g388
  (
    n420,
    n319
  );


  buf
  g389
  (
    n372,
    n304
  );


  buf
  g390
  (
    n442,
    n308
  );


  not
  g391
  (
    n351,
    n311
  );


  buf
  g392
  (
    n419,
    n319
  );


  not
  g393
  (
    n384,
    n301
  );


  not
  g394
  (
    n439,
    n317
  );


  buf
  g395
  (
    n380,
    n314
  );


  not
  g396
  (
    n400,
    n295
  );


  buf
  g397
  (
    n431,
    n310
  );


  buf
  g398
  (
    n369,
    n310
  );


  not
  g399
  (
    n343,
    n294
  );


  buf
  g400
  (
    n436,
    n310
  );


  not
  g401
  (
    n393,
    n299
  );


  buf
  g402
  (
    n366,
    n291
  );


  not
  g403
  (
    n387,
    n298
  );


  buf
  g404
  (
    n355,
    n292
  );


  buf
  g405
  (
    n360,
    n310
  );


  buf
  g406
  (
    n412,
    n316
  );


  buf
  g407
  (
    n381,
    n297
  );


  buf
  g408
  (
    n383,
    n296
  );


  not
  g409
  (
    n325,
    n298
  );


  not
  g410
  (
    n434,
    n301
  );


  not
  g411
  (
    n421,
    n311
  );


  buf
  g412
  (
    n362,
    n302
  );


  buf
  g413
  (
    n415,
    n293
  );


  not
  g414
  (
    n361,
    n306
  );


  buf
  g415
  (
    n411,
    n300
  );


  buf
  g416
  (
    n388,
    n294
  );


  buf
  g417
  (
    n407,
    n303
  );


  not
  g418
  (
    n350,
    n316
  );


  buf
  g419
  (
    n377,
    n320
  );


  and
  g420
  (
    n410,
    n301,
    n322,
    n296,
    n291
  );


  xnor
  g421
  (
    n470,
    n413,
    n377,
    n358,
    n427
  );


  xor
  g422
  (
    n450,
    n353,
    n415,
    n366,
    n382
  );


  nand
  g423
  (
    n455,
    n437,
    n428,
    n423,
    n414
  );


  xor
  g424
  (
    n495,
    n346,
    n401,
    n425,
    n383
  );


  or
  g425
  (
    n521,
    n379,
    n408,
    n358
  );


  nor
  g426
  (
    n474,
    n439,
    n440,
    n414,
    n362
  );


  or
  g427
  (
    n452,
    n358,
    n388,
    n384,
    n408
  );


  xor
  g428
  (
    n483,
    n400,
    n422,
    n435,
    n410
  );


  nand
  g429
  (
    n541,
    n381,
    n426,
    n395,
    n386
  );


  nand
  g430
  (
    n537,
    n443,
    n365,
    n440,
    n352
  );


  nand
  g431
  (
    n510,
    n407,
    n396,
    n413,
    n427
  );


  or
  g432
  (
    n525,
    n385,
    n405,
    n438,
    n337
  );


  nand
  g433
  (
    n466,
    n376,
    n384,
    n370
  );


  nor
  g434
  (
    n538,
    n401,
    n372,
    n427,
    n444
  );


  nor
  g435
  (
    n486,
    n403,
    n390,
    n369,
    n405
  );


  nand
  g436
  (
    n475,
    n392,
    n330,
    n364,
    n413
  );


  or
  g437
  (
    n494,
    n364,
    n364,
    n371,
    n441
  );


  and
  g438
  (
    n447,
    n323,
    n416,
    n398,
    n338
  );


  and
  g439
  (
    n531,
    n404,
    n376,
    n395,
    n367
  );


  nor
  g440
  (
    n454,
    n406,
    n397,
    n372,
    n379
  );


  nand
  g441
  (
    n448,
    n412,
    n423,
    n374,
    n414
  );


  or
  g442
  (
    n496,
    n435,
    n433,
    n392,
    n387
  );


  xor
  g443
  (
    n497,
    n444,
    n393,
    n392,
    n420
  );


  xor
  g444
  (
    KeyWire_0_14,
    n379,
    n404,
    n359,
    n387
  );


  xor
  g445
  (
    n457,
    n415,
    n444,
    n401,
    n354
  );


  nand
  g446
  (
    n453,
    n393,
    n387,
    n396,
    n421
  );


  or
  g447
  (
    n514,
    n399,
    n421,
    n342,
    n429
  );


  xor
  g448
  (
    n482,
    n392,
    n410,
    n419,
    n434
  );


  nand
  g449
  (
    n463,
    n439,
    n407,
    n336,
    n404
  );


  and
  g450
  (
    n503,
    n380,
    n433,
    n422,
    n406
  );


  and
  g451
  (
    n504,
    n357,
    n324,
    n437,
    n402
  );


  or
  g452
  (
    n468,
    n372,
    n378,
    n432,
    n403
  );


  nand
  g453
  (
    n508,
    n325,
    n383,
    n384,
    n444
  );


  nand
  g454
  (
    n520,
    n375,
    n416,
    n347,
    n417
  );


  xor
  g455
  (
    n459,
    n339,
    n388,
    n403,
    n439
  );


  nand
  g456
  (
    n485,
    n375,
    n418,
    n360,
    n387
  );


  nor
  g457
  (
    n501,
    n397,
    n363,
    n358,
    n417
  );


  and
  g458
  (
    n534,
    n374,
    n377,
    n430,
    n367
  );


  nand
  g459
  (
    n490,
    n403,
    n396,
    n359,
    n432
  );


  xnor
  g460
  (
    n458,
    n431,
    n443,
    n382,
    n359
  );


  or
  g461
  (
    n479,
    n442,
    n442,
    n405,
    n368
  );


  nor
  g462
  (
    n505,
    n397,
    n414,
    n355,
    n390
  );


  xnor
  g463
  (
    n513,
    n417,
    n362,
    n367,
    n397
  );


  nand
  g464
  (
    n500,
    n369,
    n409,
    n360,
    n381
  );


  xor
  g465
  (
    n539,
    n370,
    n390,
    n422,
    n349
  );


  xor
  g466
  (
    n542,
    n361,
    n419,
    n409,
    n416
  );


  nand
  g467
  (
    n488,
    n380,
    n417,
    n443,
    n385
  );


  xor
  g468
  (
    n465,
    n445,
    n419,
    n361,
    n381
  );


  nand
  g469
  (
    n530,
    n362,
    n369,
    n370,
    n421
  );


  and
  g470
  (
    n516,
    n441,
    n429,
    n438,
    n386
  );


  or
  g471
  (
    n492,
    n340,
    n424,
    n394,
    n334
  );


  and
  g472
  (
    n543,
    n378,
    n359,
    n411,
    n436
  );


  nand
  g473
  (
    n527,
    n366,
    n436,
    n333,
    n415
  );


  and
  g474
  (
    KeyWire_0_7,
    n383,
    n332,
    n415,
    n380
  );


  xor
  g475
  (
    n461,
    n329,
    n366,
    n382,
    n398
  );


  or
  g476
  (
    n491,
    n365,
    n430,
    n348,
    n369
  );


  or
  g477
  (
    n507,
    n378,
    n434,
    n326,
    n370
  );


  xnor
  g478
  (
    n469,
    n426,
    n371,
    n436,
    n411
  );


  nand
  g479
  (
    n518,
    n423,
    n365,
    n434,
    n350
  );


  or
  g480
  (
    n472,
    n425,
    n396,
    n418,
    n423
  );


  xnor
  g481
  (
    n489,
    n363,
    n394,
    n391,
    n401
  );


  nor
  g482
  (
    n467,
    n373,
    n328,
    n344,
    n430
  );


  or
  g483
  (
    n477,
    n341,
    n428,
    n399,
    n365
  );


  nor
  g484
  (
    n519,
    n412,
    n437,
    n393,
    n388
  );


  xnor
  g485
  (
    n523,
    n363,
    n366,
    n362,
    n411
  );


  nand
  g486
  (
    n502,
    n436,
    n439,
    n390,
    n398
  );


  nand
  g487
  (
    n451,
    n391,
    n445,
    n419,
    n383
  );


  or
  g488
  (
    n540,
    n375,
    n368,
    n378,
    n400
  );


  or
  g489
  (
    n478,
    n405,
    n406,
    n343,
    n400
  );


  xnor
  g490
  (
    n528,
    n409,
    n389,
    n371,
    n446
  );


  xnor
  g491
  (
    n498,
    n424,
    n368,
    n428,
    n331
  );


  xnor
  g492
  (
    n529,
    n430,
    n399,
    n386,
    n429
  );


  nand
  g493
  (
    n517,
    n385,
    n356,
    n373,
    n402
  );


  nand
  g494
  (
    n456,
    n407,
    n361,
    n433,
    n368
  );


  xnor
  g495
  (
    n512,
    n425,
    n382,
    n442,
    n407
  );


  xnor
  g496
  (
    n522,
    n379,
    n393,
    n389
  );


  nand
  g497
  (
    n462,
    n431,
    n432,
    n424,
    n410
  );


  nor
  g498
  (
    n493,
    n374,
    n435,
    n429,
    n440
  );


  xor
  g499
  (
    n536,
    n400,
    n432,
    n438,
    n377
  );


  xnor
  g500
  (
    n481,
    n437,
    n373,
    n351,
    n361
  );


  or
  g501
  (
    n526,
    n420,
    n442,
    n418,
    n435
  );


  xor
  g502
  (
    n535,
    n406,
    n364,
    n360,
    n394
  );


  and
  g503
  (
    n471,
    n371,
    n376,
    n381,
    n345
  );


  nand
  g504
  (
    n533,
    n395,
    n399,
    n398,
    n380
  );


  or
  g505
  (
    n480,
    n385,
    n440,
    n413,
    n409
  );


  nand
  g506
  (
    n499,
    n360,
    n394,
    n408,
    n426
  );


  nand
  g507
  (
    n464,
    n441,
    n402,
    n431,
    n375
  );


  and
  g508
  (
    n506,
    n412,
    n445,
    n420
  );


  and
  g509
  (
    n476,
    n388,
    n427,
    n424,
    n363
  );


  xor
  g510
  (
    n487,
    n391,
    n386,
    n373,
    n374
  );


  xnor
  g511
  (
    n524,
    n335,
    n418,
    n428,
    n389
  );


  and
  g512
  (
    n509,
    n411,
    n433,
    n425,
    n327
  );


  or
  g513
  (
    n515,
    n416,
    n404,
    n395,
    n421
  );


  or
  g514
  (
    n484,
    n402,
    n438,
    n422,
    n372
  );


  xor
  g515
  (
    n473,
    n391,
    n445,
    n412,
    n431
  );


  or
  g516
  (
    n449,
    n443,
    n367,
    n441,
    n377
  );


  and
  g517
  (
    n511,
    n434,
    n376,
    n410,
    n426
  );


  not
  g518
  (
    n544,
    n464
  );


  buf
  g519
  (
    n548,
    n453
  );


  nand
  g520
  (
    n546,
    n449,
    n451
  );


  xnor
  g521
  (
    n545,
    n457,
    n447,
    n459,
    n461
  );


  nand
  g522
  (
    n549,
    n456,
    n452,
    n454,
    n463
  );


  nor
  g523
  (
    n547,
    n448,
    n455,
    n462,
    n466
  );


  xnor
  g524
  (
    n550,
    n450,
    n458,
    n460,
    n465
  );


  not
  g525
  (
    n557,
    n547
  );


  not
  g526
  (
    n558,
    n545
  );


  not
  g527
  (
    n552,
    n550
  );


  not
  g528
  (
    n556,
    n285
  );


  not
  g529
  (
    n560,
    n546
  );


  not
  g530
  (
    n559,
    n548
  );


  not
  g531
  (
    n551,
    n550
  );


  nor
  g532
  (
    n553,
    n549,
    n285,
    n550
  );


  xnor
  g533
  (
    n554,
    n285,
    n544,
    n284
  );


  nand
  g534
  (
    n555,
    n550,
    n285,
    n286
  );


  not
  g535
  (
    n564,
    n554
  );


  buf
  g536
  (
    n567,
    n556
  );


  buf
  g537
  (
    n574,
    n480
  );


  not
  g538
  (
    n563,
    n556
  );


  buf
  g539
  (
    n585,
    n476
  );


  buf
  g540
  (
    n575,
    n555
  );


  buf
  g541
  (
    n581,
    n554
  );


  not
  g542
  (
    n577,
    n555
  );


  not
  g543
  (
    n588,
    n477
  );


  not
  g544
  (
    n579,
    n552
  );


  not
  g545
  (
    n583,
    n551
  );


  not
  g546
  (
    n587,
    n551
  );


  not
  g547
  (
    n580,
    n485
  );


  not
  g548
  (
    n562,
    n557
  );


  buf
  g549
  (
    n584,
    n558
  );


  buf
  g550
  (
    n578,
    n553
  );


  not
  g551
  (
    n570,
    n482
  );


  not
  g552
  (
    n589,
    n469
  );


  not
  g553
  (
    n586,
    n555
  );


  buf
  g554
  (
    n573,
    n475
  );


  buf
  g555
  (
    n582,
    n553
  );


  buf
  g556
  (
    n565,
    n556
  );


  not
  g557
  (
    n568,
    n483
  );


  xnor
  g558
  (
    n571,
    n553,
    n484,
    n555
  );


  and
  g559
  (
    n561,
    n473,
    n557,
    n553,
    n474
  );


  xnor
  g560
  (
    n576,
    n557,
    n552,
    n558,
    n478
  );


  nor
  g561
  (
    n569,
    n467,
    n479,
    n481,
    n472
  );


  xor
  g562
  (
    n566,
    n552,
    n554,
    n486
  );


  or
  g563
  (
    n572,
    n468,
    n556,
    n470,
    n551
  );


  nand
  g564
  (
    n590,
    n552,
    n471,
    n551,
    n557
  );


  not
  g565
  (
    n592,
    n487
  );


  nand
  g566
  (
    n591,
    n575,
    n576,
    n577
  );


  or
  g567
  (
    n593,
    n489,
    n488,
    n490,
    n591
  );


  nand
  g568
  (
    n595,
    n494,
    n492,
    n593,
    n493
  );


  xnor
  g569
  (
    n594,
    n593,
    n491,
    n495,
    n496
  );


  xnor
  g570
  (
    n601,
    n498,
    n503
  );


  nor
  g571
  (
    n600,
    n508,
    n504,
    n501,
    n594
  );


  and
  g572
  (
    n599,
    n446,
    n595,
    n594,
    n505
  );


  or
  g573
  (
    n597,
    n511,
    n509,
    n595,
    n499
  );


  xor
  g574
  (
    n596,
    n497,
    n446,
    n595,
    n506
  );


  nor
  g575
  (
    KeyWire_0_13,
    n446,
    n500,
    n512,
    n594
  );


  or
  g576
  (
    n602,
    n507,
    n595,
    n510,
    n502
  );


  not
  g577
  (
    n612,
    n599
  );


  not
  g578
  (
    n609,
    n598
  );


  not
  g579
  (
    n608,
    n600
  );


  not
  g580
  (
    n607,
    n600
  );


  not
  g581
  (
    n603,
    n599
  );


  not
  g582
  (
    n604,
    n600
  );


  not
  g583
  (
    n605,
    n601
  );


  not
  g584
  (
    n610,
    n597
  );


  buf
  g585
  (
    n606,
    n600
  );


  buf
  g586
  (
    n611,
    n596
  );


  not
  g587
  (
    n632,
    n592
  );


  not
  g588
  (
    n630,
    n579
  );


  buf
  g589
  (
    n625,
    n606
  );


  buf
  g590
  (
    n644,
    n612
  );


  buf
  g591
  (
    n616,
    n607
  );


  buf
  g592
  (
    n648,
    n611
  );


  not
  g593
  (
    n622,
    n182
  );


  not
  g594
  (
    n633,
    n608
  );


  buf
  g595
  (
    n638,
    n606
  );


  not
  g596
  (
    n636,
    n581
  );


  not
  g597
  (
    n641,
    n517
  );


  buf
  g598
  (
    n650,
    n610
  );


  not
  g599
  (
    n620,
    n580
  );


  buf
  g600
  (
    n629,
    n608
  );


  not
  g601
  (
    n628,
    n185
  );


  not
  g602
  (
    n640,
    n612
  );


  buf
  g603
  (
    n621,
    n612
  );


  buf
  g604
  (
    n634,
    n183
  );


  buf
  g605
  (
    n646,
    n604
  );


  buf
  g606
  (
    n615,
    n604
  );


  not
  g607
  (
    n649,
    n607
  );


  not
  g608
  (
    n626,
    n186
  );


  buf
  g609
  (
    n627,
    n611
  );


  not
  g610
  (
    n623,
    n184
  );


  buf
  g611
  (
    n645,
    n516
  );


  not
  g612
  (
    n637,
    n609
  );


  not
  g613
  (
    n643,
    n608
  );


  buf
  g614
  (
    n624,
    n609
  );


  buf
  g615
  (
    n651,
    n603
  );


  not
  g616
  (
    n639,
    n605
  );


  not
  g617
  (
    n619,
    n604
  );


  buf
  g618
  (
    n614,
    n605
  );


  not
  g619
  (
    n635,
    n187
  );


  not
  g620
  (
    n652,
    n610
  );


  nand
  g621
  (
    n631,
    n603,
    n611
  );


  and
  g622
  (
    n647,
    n513,
    n515,
    n605,
    n603
  );


  nand
  g623
  (
    n617,
    n608,
    n578,
    n603,
    n609
  );


  and
  g624
  (
    n613,
    n610,
    n612,
    n607,
    n606
  );


  xor
  g625
  (
    n642,
    n609,
    n604,
    n514,
    n610
  );


  or
  g626
  (
    n618,
    n606,
    n605,
    n611,
    n607
  );


  buf
  g627
  (
    n740,
    n619
  );


  buf
  g628
  (
    n683,
    n615
  );


  not
  g629
  (
    n694,
    n634
  );


  buf
  g630
  (
    n664,
    n640
  );


  buf
  g631
  (
    n773,
    n613
  );


  buf
  g632
  (
    n761,
    n652
  );


  buf
  g633
  (
    n791,
    n633
  );


  buf
  g634
  (
    n778,
    n632
  );


  buf
  g635
  (
    n794,
    n616
  );


  buf
  g636
  (
    n726,
    n645
  );


  buf
  g637
  (
    n688,
    n630
  );


  buf
  g638
  (
    n687,
    n633
  );


  buf
  g639
  (
    n789,
    n618
  );


  buf
  g640
  (
    n722,
    n651
  );


  not
  g641
  (
    n777,
    n624
  );


  not
  g642
  (
    n654,
    n652
  );


  not
  g643
  (
    n732,
    n629
  );


  buf
  g644
  (
    n690,
    n651
  );


  not
  g645
  (
    n719,
    n629
  );


  not
  g646
  (
    n710,
    n643
  );


  not
  g647
  (
    n769,
    n560
  );


  buf
  g648
  (
    n700,
    n621
  );


  buf
  g649
  (
    n781,
    n617
  );


  buf
  g650
  (
    n768,
    n625
  );


  buf
  g651
  (
    n691,
    n626
  );


  not
  g652
  (
    n783,
    n645
  );


  not
  g653
  (
    n747,
    n646
  );


  buf
  g654
  (
    n727,
    n618
  );


  not
  g655
  (
    n699,
    n613
  );


  not
  g656
  (
    n717,
    n631
  );


  not
  g657
  (
    n704,
    n622
  );


  buf
  g658
  (
    n698,
    n619
  );


  buf
  g659
  (
    n657,
    n632
  );


  buf
  g660
  (
    n674,
    n634
  );


  not
  g661
  (
    n729,
    n639
  );


  buf
  g662
  (
    n714,
    n620
  );


  not
  g663
  (
    n779,
    n633
  );


  buf
  g664
  (
    n749,
    n638
  );


  not
  g665
  (
    n667,
    n635
  );


  buf
  g666
  (
    n798,
    n625
  );


  not
  g667
  (
    n757,
    n286
  );


  not
  g668
  (
    n712,
    n643
  );


  buf
  g669
  (
    n684,
    n519
  );


  not
  g670
  (
    n662,
    n647
  );


  not
  g671
  (
    n663,
    n651
  );


  buf
  g672
  (
    n668,
    n628
  );


  not
  g673
  (
    n739,
    n643
  );


  buf
  g674
  (
    n692,
    n619
  );


  not
  g675
  (
    n800,
    n621
  );


  buf
  g676
  (
    n795,
    n647
  );


  not
  g677
  (
    n750,
    n639
  );


  not
  g678
  (
    n788,
    n646
  );


  not
  g679
  (
    n774,
    n619
  );


  not
  g680
  (
    n659,
    n644
  );


  not
  g681
  (
    n803,
    n650
  );


  not
  g682
  (
    n810,
    n617
  );


  buf
  g683
  (
    n790,
    n642
  );


  buf
  g684
  (
    n708,
    n627
  );


  not
  g685
  (
    n755,
    n622
  );


  buf
  g686
  (
    n758,
    n616
  );


  buf
  g687
  (
    n707,
    n624
  );


  buf
  g688
  (
    n745,
    n621
  );


  buf
  g689
  (
    n679,
    n629
  );


  buf
  g690
  (
    n706,
    n614
  );


  not
  g691
  (
    n793,
    n630
  );


  not
  g692
  (
    n665,
    n624
  );


  buf
  g693
  (
    n693,
    n558
  );


  buf
  g694
  (
    n780,
    n637
  );


  not
  g695
  (
    n762,
    n636
  );


  buf
  g696
  (
    n709,
    n627
  );


  not
  g697
  (
    n723,
    n622
  );


  buf
  g698
  (
    n799,
    n646
  );


  buf
  g699
  (
    n785,
    n559
  );


  buf
  g700
  (
    n660,
    n647
  );


  not
  g701
  (
    n801,
    n620
  );


  buf
  g702
  (
    n735,
    n637
  );


  buf
  g703
  (
    n812,
    n649
  );


  buf
  g704
  (
    n697,
    n623
  );


  not
  g705
  (
    n796,
    n633
  );


  not
  g706
  (
    n711,
    n621
  );


  buf
  g707
  (
    n753,
    n630
  );


  not
  g708
  (
    n678,
    n559
  );


  not
  g709
  (
    n720,
    n648
  );


  not
  g710
  (
    n696,
    n636
  );


  not
  g711
  (
    n731,
    n642
  );


  not
  g712
  (
    n737,
    n560
  );


  not
  g713
  (
    n682,
    n635
  );


  not
  g714
  (
    n686,
    n649
  );


  not
  g715
  (
    n772,
    n649
  );


  not
  g716
  (
    n724,
    n627
  );


  not
  g717
  (
    n666,
    n558
  );


  not
  g718
  (
    n701,
    n648
  );


  buf
  g719
  (
    n669,
    n614
  );


  buf
  g720
  (
    n658,
    n641
  );


  not
  g721
  (
    n656,
    n650
  );


  buf
  g722
  (
    n765,
    n618
  );


  not
  g723
  (
    n681,
    n648
  );


  buf
  g724
  (
    n743,
    n638
  );


  buf
  g725
  (
    n677,
    n617
  );


  not
  g726
  (
    n797,
    n631
  );


  buf
  g727
  (
    n759,
    n286
  );


  not
  g728
  (
    n738,
    n642
  );


  buf
  g729
  (
    n786,
    n638
  );


  buf
  g730
  (
    n672,
    n622
  );


  buf
  g731
  (
    n752,
    n640
  );


  buf
  g732
  (
    n775,
    n643
  );


  not
  g733
  (
    n728,
    n520
  );


  buf
  g734
  (
    n661,
    n646
  );


  buf
  g735
  (
    n676,
    n642
  );


  buf
  g736
  (
    n760,
    n632
  );


  not
  g737
  (
    n806,
    n615
  );


  not
  g738
  (
    n689,
    n628
  );


  buf
  g739
  (
    n736,
    n650
  );


  not
  g740
  (
    n811,
    n614
  );


  buf
  g741
  (
    n716,
    n620
  );


  not
  g742
  (
    n804,
    n640
  );


  not
  g743
  (
    n766,
    n614
  );


  buf
  g744
  (
    n721,
    n639
  );


  not
  g745
  (
    n733,
    n640
  );


  buf
  g746
  (
    n809,
    n560
  );


  buf
  g747
  (
    n705,
    n634
  );


  not
  g748
  (
    n754,
    n626
  );


  not
  g749
  (
    n653,
    n634
  );


  not
  g750
  (
    n746,
    n635
  );


  not
  g751
  (
    n807,
    n613
  );


  buf
  g752
  (
    n770,
    n651
  );


  buf
  g753
  (
    n742,
    n648
  );


  buf
  g754
  (
    n784,
    n625
  );


  not
  g755
  (
    n808,
    n623
  );


  buf
  g756
  (
    n802,
    n620
  );


  not
  g757
  (
    n805,
    n645
  );


  buf
  g758
  (
    n764,
    n624
  );


  buf
  g759
  (
    n776,
    n645
  );


  not
  g760
  (
    n787,
    n627
  );


  not
  g761
  (
    n671,
    n628
  );


  not
  g762
  (
    n741,
    n628
  );


  not
  g763
  (
    n756,
    n639
  );


  not
  g764
  (
    n744,
    n637
  );


  not
  g765
  (
    n675,
    n625
  );


  buf
  g766
  (
    n748,
    n636
  );


  buf
  g767
  (
    n713,
    n644
  );


  buf
  g768
  (
    n702,
    n521
  );


  not
  g769
  (
    n725,
    n649
  );


  not
  g770
  (
    n792,
    n615
  );


  not
  g771
  (
    n680,
    n635
  );


  buf
  g772
  (
    n767,
    n626
  );


  buf
  g773
  (
    n715,
    n641
  );


  not
  g774
  (
    n685,
    n647
  );


  not
  g775
  (
    n751,
    n636
  );


  not
  g776
  (
    n730,
    n652
  );


  buf
  g777
  (
    n670,
    n632
  );


  buf
  g778
  (
    n695,
    n613
  );


  buf
  g779
  (
    n734,
    n616
  );


  not
  g780
  (
    n718,
    n518
  );


  nand
  g781
  (
    n782,
    n629,
    n641
  );


  xnor
  g782
  (
    n763,
    n652,
    n630,
    n626,
    n616
  );


  or
  g783
  (
    n703,
    n623,
    n644,
    n637,
    n617
  );


  xnor
  g784
  (
    n655,
    n615,
    n638,
    n644,
    n618
  );


  xor
  g785
  (
    n673,
    n650,
    n559,
    n560
  );


  xor
  g786
  (
    n771,
    n623,
    n631,
    n641
  );


  not
  g787
  (
    n896,
    n788
  );


  buf
  g788
  (
    n1124,
    n716
  );


  not
  g789
  (
    n1078,
    n779
  );


  buf
  g790
  (
    n931,
    n736
  );


  not
  g791
  (
    n1019,
    n752
  );


  buf
  g792
  (
    n1069,
    n684
  );


  buf
  g793
  (
    n842,
    n783
  );


  not
  g794
  (
    n893,
    n678
  );


  not
  g795
  (
    n948,
    n672
  );


  not
  g796
  (
    n1140,
    n796
  );


  not
  g797
  (
    n972,
    n801
  );


  not
  g798
  (
    n1029,
    n687
  );


  buf
  g799
  (
    n933,
    n704
  );


  buf
  g800
  (
    n1012,
    n720
  );


  buf
  g801
  (
    n1064,
    n684
  );


  buf
  g802
  (
    n846,
    n782
  );


  not
  g803
  (
    n992,
    n668
  );


  not
  g804
  (
    n1000,
    n791
  );


  not
  g805
  (
    n814,
    n804
  );


  buf
  g806
  (
    n864,
    n751
  );


  not
  g807
  (
    n1110,
    n585
  );


  buf
  g808
  (
    n1093,
    n755
  );


  not
  g809
  (
    n1005,
    n671
  );


  not
  g810
  (
    n1159,
    n658
  );


  not
  g811
  (
    n901,
    n669
  );


  buf
  g812
  (
    n899,
    n775
  );


  buf
  g813
  (
    n924,
    n707
  );


  not
  g814
  (
    n1022,
    n801
  );


  not
  g815
  (
    n835,
    n706
  );


  not
  g816
  (
    n998,
    n794
  );


  not
  g817
  (
    n1130,
    n717
  );


  not
  g818
  (
    n848,
    n660
  );


  buf
  g819
  (
    n1041,
    n757
  );


  buf
  g820
  (
    n1166,
    n799
  );


  buf
  g821
  (
    n973,
    n791
  );


  not
  g822
  (
    n1091,
    n746
  );


  not
  g823
  (
    n851,
    n800
  );


  not
  g824
  (
    n1087,
    n788
  );


  not
  g825
  (
    n963,
    n737
  );


  not
  g826
  (
    n831,
    n721
  );


  not
  g827
  (
    n859,
    n688
  );


  buf
  g828
  (
    n919,
    n776
  );


  buf
  g829
  (
    n1073,
    n744
  );


  buf
  g830
  (
    n985,
    n673
  );


  not
  g831
  (
    n904,
    n808
  );


  not
  g832
  (
    n849,
    n689
  );


  not
  g833
  (
    KeyWire_0_8,
    n654
  );


  buf
  g834
  (
    n1056,
    n657
  );


  buf
  g835
  (
    n894,
    n701
  );


  not
  g836
  (
    n1102,
    n671
  );


  not
  g837
  (
    n921,
    n743
  );


  buf
  g838
  (
    n1082,
    n693
  );


  buf
  g839
  (
    n950,
    n761
  );


  buf
  g840
  (
    n1085,
    n670
  );


  not
  g841
  (
    n856,
    n793
  );


  not
  g842
  (
    n1151,
    n785
  );


  buf
  g843
  (
    n881,
    n763
  );


  not
  g844
  (
    n1126,
    n683
  );


  buf
  g845
  (
    n861,
    n670
  );


  not
  g846
  (
    n857,
    n761
  );


  not
  g847
  (
    n1074,
    n742
  );


  not
  g848
  (
    n1043,
    n753
  );


  not
  g849
  (
    n883,
    n672
  );


  buf
  g850
  (
    n957,
    n695
  );


  buf
  g851
  (
    n1128,
    n800
  );


  not
  g852
  (
    n836,
    n773
  );


  not
  g853
  (
    n913,
    n684
  );


  buf
  g854
  (
    n1112,
    n713
  );


  buf
  g855
  (
    n874,
    n792
  );


  not
  g856
  (
    n932,
    n701
  );


  buf
  g857
  (
    n886,
    n727
  );


  not
  g858
  (
    n915,
    n687
  );


  not
  g859
  (
    n1032,
    n804
  );


  buf
  g860
  (
    n1115,
    n802
  );


  not
  g861
  (
    n1161,
    n793
  );


  not
  g862
  (
    n1123,
    n798
  );


  buf
  g863
  (
    n995,
    n785
  );


  buf
  g864
  (
    n1081,
    n797
  );


  not
  g865
  (
    n863,
    n811
  );


  buf
  g866
  (
    n960,
    n721
  );


  not
  g867
  (
    n1158,
    n653
  );


  buf
  g868
  (
    n1153,
    n687
  );


  buf
  g869
  (
    n1173,
    n695
  );


  buf
  g870
  (
    n865,
    n653
  );


  buf
  g871
  (
    n1125,
    n756
  );


  buf
  g872
  (
    n1040,
    n740
  );


  buf
  g873
  (
    n1059,
    n709
  );


  buf
  g874
  (
    n1108,
    n702
  );


  buf
  g875
  (
    n838,
    n741
  );


  not
  g876
  (
    n912,
    n758
  );


  not
  g877
  (
    n1095,
    n670
  );


  buf
  g878
  (
    n970,
    n784
  );


  buf
  g879
  (
    n996,
    n655
  );


  buf
  g880
  (
    n1016,
    n673
  );


  not
  g881
  (
    n1097,
    n724
  );


  buf
  g882
  (
    n1172,
    n662
  );


  buf
  g883
  (
    n1046,
    n730
  );


  not
  g884
  (
    n939,
    n765
  );


  buf
  g885
  (
    n1044,
    n679
  );


  buf
  g886
  (
    n860,
    n660
  );


  buf
  g887
  (
    n1028,
    n762
  );


  buf
  g888
  (
    n887,
    n752
  );


  not
  g889
  (
    n1023,
    n743
  );


  not
  g890
  (
    n1114,
    n771
  );


  not
  g891
  (
    n1024,
    n798
  );


  buf
  g892
  (
    n1035,
    n786
  );


  buf
  g893
  (
    n1111,
    n666
  );


  not
  g894
  (
    n1065,
    n664
  );


  buf
  g895
  (
    n1120,
    n755
  );


  buf
  g896
  (
    n1163,
    n744
  );


  not
  g897
  (
    n1047,
    n737
  );


  buf
  g898
  (
    n934,
    n799
  );


  not
  g899
  (
    n815,
    n699
  );


  buf
  g900
  (
    n1026,
    n809
  );


  not
  g901
  (
    n920,
    n688
  );


  buf
  g902
  (
    n890,
    n659
  );


  buf
  g903
  (
    n1058,
    n746
  );


  buf
  g904
  (
    n971,
    n750
  );


  buf
  g905
  (
    n1094,
    n746
  );


  not
  g906
  (
    n1086,
    n760
  );


  buf
  g907
  (
    n850,
    n742
  );


  not
  g908
  (
    n952,
    n717
  );


  buf
  g909
  (
    n1122,
    n752
  );


  not
  g910
  (
    n1021,
    n664
  );


  buf
  g911
  (
    KeyWire_0_11,
    n588
  );


  buf
  g912
  (
    n1015,
    n673
  );


  buf
  g913
  (
    n882,
    n799
  );


  buf
  g914
  (
    n956,
    n728
  );


  not
  g915
  (
    n844,
    n782
  );


  not
  g916
  (
    n928,
    n680
  );


  buf
  g917
  (
    n898,
    n788
  );


  not
  g918
  (
    n823,
    n740
  );


  buf
  g919
  (
    n1017,
    n669
  );


  not
  g920
  (
    n1066,
    n674
  );


  buf
  g921
  (
    n1090,
    n715
  );


  buf
  g922
  (
    n945,
    n736
  );


  buf
  g923
  (
    n897,
    n808
  );


  not
  g924
  (
    n1175,
    n778
  );


  not
  g925
  (
    n822,
    n770
  );


  not
  g926
  (
    n1170,
    n798
  );


  buf
  g927
  (
    n941,
    n736
  );


  not
  g928
  (
    n983,
    n793
  );


  buf
  g929
  (
    n1062,
    n807
  );


  buf
  g930
  (
    n988,
    n747
  );


  not
  g931
  (
    n978,
    n653
  );


  not
  g932
  (
    n869,
    n810
  );


  buf
  g933
  (
    n1155,
    n778
  );


  buf
  g934
  (
    n1063,
    n703
  );


  not
  g935
  (
    n976,
    n777
  );


  buf
  g936
  (
    n830,
    n741
  );


  buf
  g937
  (
    n969,
    n759
  );


  not
  g938
  (
    n914,
    n760
  );


  buf
  g939
  (
    n930,
    n781
  );


  not
  g940
  (
    n1011,
    n666
  );


  not
  g941
  (
    n1092,
    n702
  );


  not
  g942
  (
    n1051,
    n697
  );


  not
  g943
  (
    n1137,
    n797
  );


  not
  g944
  (
    n1077,
    n725
  );


  not
  g945
  (
    n1060,
    n717
  );


  buf
  g946
  (
    n1160,
    n681
  );


  buf
  g947
  (
    n958,
    n719
  );


  buf
  g948
  (
    n1099,
    n722
  );


  not
  g949
  (
    n1080,
    n729
  );


  buf
  g950
  (
    n1118,
    n783
  );


  buf
  g951
  (
    n959,
    n772
  );


  not
  g952
  (
    n949,
    n765
  );


  not
  g953
  (
    n974,
    n706
  );


  not
  g954
  (
    n1003,
    n779
  );


  buf
  g955
  (
    n1142,
    n749
  );


  buf
  g956
  (
    n878,
    n655
  );


  not
  g957
  (
    n824,
    n717
  );


  not
  g958
  (
    n910,
    n704
  );


  buf
  g959
  (
    n876,
    n765
  );


  buf
  g960
  (
    n975,
    n688
  );


  not
  g961
  (
    n1138,
    n708
  );


  not
  g962
  (
    n1018,
    n791
  );


  not
  g963
  (
    n862,
    n685
  );


  buf
  g964
  (
    n1105,
    n769
  );


  not
  g965
  (
    n1149,
    n754
  );


  buf
  g966
  (
    n1054,
    n658
  );


  not
  g967
  (
    n1079,
    n658
  );


  buf
  g968
  (
    n923,
    n689
  );


  not
  g969
  (
    n1042,
    n703
  );


  buf
  g970
  (
    n967,
    n775
  );


  not
  g971
  (
    n946,
    n664
  );


  buf
  g972
  (
    n1014,
    n734
  );


  not
  g973
  (
    n922,
    n771
  );


  not
  g974
  (
    KeyWire_0_6,
    n668
  );


  not
  g975
  (
    n903,
    n803
  );


  not
  g976
  (
    n937,
    n756
  );


  buf
  g977
  (
    n1167,
    n790
  );


  not
  g978
  (
    n905,
    n801
  );


  not
  g979
  (
    n1169,
    n674
  );


  buf
  g980
  (
    n1107,
    n812
  );


  not
  g981
  (
    n1031,
    n680
  );


  buf
  g982
  (
    n880,
    n770
  );


  not
  g983
  (
    n936,
    n655
  );


  not
  g984
  (
    n1050,
    n682
  );


  not
  g985
  (
    n942,
    n770
  );


  not
  g986
  (
    n895,
    n781
  );


  not
  g987
  (
    n833,
    n794
  );


  buf
  g988
  (
    n858,
    n694
  );


  not
  g989
  (
    n840,
    n661
  );


  buf
  g990
  (
    n940,
    n801
  );


  buf
  g991
  (
    n917,
    n766
  );


  buf
  g992
  (
    n1098,
    n716
  );


  not
  g993
  (
    n1157,
    n698
  );


  not
  g994
  (
    n944,
    n704
  );


  buf
  g995
  (
    n1165,
    n762
  );


  not
  g996
  (
    n1036,
    n809
  );


  not
  g997
  (
    n1001,
    n747
  );


  not
  g998
  (
    n1076,
    n683
  );


  not
  g999
  (
    n1052,
    n660
  );


  not
  g1000
  (
    n1144,
    n776
  );


  not
  g1001
  (
    n891,
    n771
  );


  not
  g1002
  (
    n1141,
    n757
  );


  buf
  g1003
  (
    n1057,
    n710
  );


  not
  g1004
  (
    n871,
    n666
  );


  not
  g1005
  (
    n906,
    n807
  );


  buf
  g1006
  (
    n1129,
    n655
  );


  buf
  g1007
  (
    n885,
    n697
  );


  buf
  g1008
  (
    n1103,
    n766
  );


  not
  g1009
  (
    n935,
    n763
  );


  buf
  g1010
  (
    n1034,
    n734
  );


  not
  g1011
  (
    n1174,
    n733
  );


  not
  g1012
  (
    n926,
    n733
  );


  buf
  g1013
  (
    n816,
    n761
  );


  buf
  g1014
  (
    n927,
    n705
  );


  not
  g1015
  (
    n1020,
    n737
  );


  buf
  g1016
  (
    n1045,
    n745
  );


  buf
  g1017
  (
    n1131,
    n668
  );


  buf
  g1018
  (
    n909,
    n692
  );


  buf
  g1019
  (
    n854,
    n804
  );


  buf
  g1020
  (
    n834,
    n724
  );


  buf
  g1021
  (
    n821,
    n762
  );


  not
  g1022
  (
    n889,
    n683
  );


  not
  g1023
  (
    n986,
    n667
  );


  not
  g1024
  (
    n820,
    n729
  );


  buf
  g1025
  (
    n1089,
    n730
  );


  not
  g1026
  (
    n827,
    n784
  );


  not
  g1027
  (
    n868,
    n736
  );


  buf
  g1028
  (
    n1096,
    n772
  );


  not
  g1029
  (
    n1006,
    n762
  );


  not
  g1030
  (
    n1101,
    n733
  );


  not
  g1031
  (
    n1171,
    n745
  );


  buf
  g1032
  (
    n1104,
    n789
  );


  not
  g1033
  (
    n1106,
    n735
  );


  buf
  g1034
  (
    n1061,
    n802
  );


  buf
  g1035
  (
    n875,
    n735
  );


  not
  g1036
  (
    n938,
    n670
  );


  not
  g1037
  (
    n1004,
    n774
  );


  buf
  g1038
  (
    n1025,
    n711
  );


  not
  g1039
  (
    n843,
    n795
  );


  not
  g1040
  (
    n1154,
    n732
  );


  buf
  g1041
  (
    n994,
    n716
  );


  buf
  g1042
  (
    n1119,
    n710
  );


  not
  g1043
  (
    n1168,
    n719
  );


  buf
  g1044
  (
    n987,
    n738
  );


  buf
  g1045
  (
    n872,
    n749
  );


  not
  g1046
  (
    n1135,
    n696
  );


  not
  g1047
  (
    n817,
    n792
  );


  buf
  g1048
  (
    n837,
    n691
  );


  buf
  g1049
  (
    n911,
    n686
  );


  not
  g1050
  (
    n1109,
    n748
  );


  not
  g1051
  (
    n993,
    n738
  );


  not
  g1052
  (
    n1027,
    n724
  );


  buf
  g1053
  (
    n908,
    n653
  );


  buf
  g1054
  (
    n1147,
    n691
  );


  not
  g1055
  (
    n1146,
    n777
  );


  and
  g1056
  (
    n1164,
    n718,
    n727,
    n690,
    n742
  );


  xor
  g1057
  (
    n982,
    n700,
    n723,
    n786,
    n729
  );


  or
  g1058
  (
    n1176,
    n673,
    n675,
    n790,
    n812
  );


  nand
  g1059
  (
    n818,
    n708,
    n757,
    n720,
    n777
  );


  and
  g1060
  (
    n1037,
    n582,
    n693,
    n698,
    n714
  );


  nand
  g1061
  (
    n888,
    n726,
    n690,
    n728,
    n792
  );


  xnor
  g1062
  (
    n990,
    n785,
    n731,
    n734,
    n690
  );


  and
  g1063
  (
    n1053,
    n773,
    n735,
    n739,
    n696
  );


  or
  g1064
  (
    n991,
    n711,
    n741,
    n712,
    n743
  );


  nor
  g1065
  (
    n1071,
    n695,
    n584,
    n677,
    n699
  );


  and
  g1066
  (
    n1152,
    n750,
    n680,
    n698,
    n672
  );


  and
  g1067
  (
    n955,
    n719,
    n686,
    n767,
    n674
  );


  xnor
  g1068
  (
    n1116,
    n740,
    n758,
    n772,
    n682
  );


  or
  g1069
  (
    n1121,
    n689,
    n777,
    n750,
    n773
  );


  xor
  g1070
  (
    n1117,
    n812,
    n719,
    n782,
    n764
  );


  or
  g1071
  (
    n839,
    n795,
    n662,
    n767,
    n751
  );


  or
  g1072
  (
    n947,
    n703,
    n742,
    n810,
    n767
  );


  or
  g1073
  (
    n813,
    n667,
    n753,
    n714,
    n773
  );


  or
  g1074
  (
    n826,
    n808,
    n796,
    n665,
    n787
  );


  and
  g1075
  (
    n966,
    n682,
    n794,
    n805,
    n731
  );


  nor
  g1076
  (
    n1150,
    n709,
    n769,
    n779,
    n664
  );


  and
  g1077
  (
    n847,
    n701,
    n715,
    n676,
    n780
  );


  xor
  g1078
  (
    n1088,
    n699,
    n656,
    n659,
    n769
  );


  nor
  g1079
  (
    KeyWire_0_9,
    n756,
    n725,
    n793,
    n715
  );


  xnor
  g1080
  (
    n925,
    n795,
    n764,
    n700,
    n787
  );


  and
  g1081
  (
    n929,
    n810,
    n707,
    n751,
    n695
  );


  and
  g1082
  (
    n841,
    n677,
    n811,
    n709,
    n766
  );


  nor
  g1083
  (
    n961,
    n680,
    n660,
    n749,
    n754
  );


  xor
  g1084
  (
    n852,
    n759,
    n678,
    n755,
    n694
  );


  or
  g1085
  (
    n902,
    n741,
    n668,
    n656,
    n722
  );


  nand
  g1086
  (
    n953,
    n693,
    n676,
    n671,
    n696
  );


  xor
  g1087
  (
    n980,
    n797,
    n718,
    n720,
    n702
  );


  nand
  g1088
  (
    n845,
    n774,
    n775,
    n661,
    n812
  );


  nand
  g1089
  (
    n866,
    n789,
    n775,
    n778,
    n722
  );


  xnor
  g1090
  (
    n1083,
    n654,
    n657,
    n662,
    n687
  );


  xor
  g1091
  (
    n828,
    n669,
    n718,
    n781,
    n711
  );


  and
  g1092
  (
    n1048,
    n796,
    n806,
    n685
  );


  or
  g1093
  (
    n855,
    n694,
    n808,
    n807,
    n803
  );


  xor
  g1094
  (
    n1145,
    n745,
    n804,
    n689,
    n803
  );


  nor
  g1095
  (
    n884,
    n768,
    n789,
    n729,
    n787
  );


  xor
  g1096
  (
    n977,
    n688,
    n656,
    n734,
    n726
  );


  and
  g1097
  (
    n1156,
    n785,
    n764,
    n758,
    n710
  );


  xnor
  g1098
  (
    n951,
    n810,
    n765,
    n676,
    n748
  );


  and
  g1099
  (
    n1013,
    n713,
    n739,
    n716,
    n730
  );


  nor
  g1100
  (
    n962,
    n760,
    n656,
    n795,
    n737
  );


  xor
  g1101
  (
    n1139,
    n798,
    n784,
    n754,
    n686
  );


  xor
  g1102
  (
    n1113,
    n738,
    n774,
    n704,
    n780
  );


  nand
  g1103
  (
    n877,
    n709,
    n731,
    n693,
    n771
  );


  xor
  g1104
  (
    n907,
    n783,
    n679,
    n697,
    n665
  );


  or
  g1105
  (
    n965,
    n700,
    n675,
    n802,
    n725
  );


  xor
  g1106
  (
    n1049,
    n677,
    n728,
    n705,
    n747
  );


  or
  g1107
  (
    n1068,
    n663,
    n755,
    n781,
    n686
  );


  nand
  g1108
  (
    n999,
    n713,
    n745,
    n714,
    n683
  );


  or
  g1109
  (
    n1070,
    n724,
    n790,
    n789,
    n705
  );


  nand
  g1110
  (
    n832,
    n799,
    n732,
    n710,
    n730
  );


  nand
  g1111
  (
    n954,
    n692,
    n672,
    n685,
    n726
  );


  xnor
  g1112
  (
    n1134,
    n692,
    n791,
    n794,
    n654
  );


  or
  g1113
  (
    n1133,
    n727,
    n750,
    n731,
    n770
  );


  xor
  g1114
  (
    n870,
    n746,
    n772,
    n768,
    n764
  );


  nor
  g1115
  (
    n1143,
    n749,
    n714,
    n769,
    n780
  );


  xor
  g1116
  (
    n1002,
    n723,
    n757,
    n809,
    n587
  );


  xnor
  g1117
  (
    n968,
    n788,
    n759,
    n696,
    n728
  );


  nand
  g1118
  (
    n943,
    n786,
    n684,
    n677,
    n657
  );


  or
  g1119
  (
    n892,
    n590,
    n752,
    n805,
    n679
  );


  and
  g1120
  (
    n918,
    n721,
    n758,
    n760,
    n766
  );


  and
  g1121
  (
    n964,
    n691,
    n733,
    n682,
    n721
  );


  nand
  g1122
  (
    n1010,
    n661,
    n748,
    n751,
    n763
  );


  nor
  g1123
  (
    n979,
    n807,
    n701,
    n705,
    n800
  );


  xnor
  g1124
  (
    n1067,
    n711,
    n727,
    n666,
    n665
  );


  nand
  g1125
  (
    n997,
    n759,
    n663,
    n792,
    n722
  );


  xor
  g1126
  (
    n1030,
    n756,
    n723,
    n661,
    n796
  );


  and
  g1127
  (
    n1100,
    n589,
    n658,
    n783,
    n671
  );


  nor
  g1128
  (
    n867,
    n586,
    n694,
    n806,
    n738
  );


  or
  g1129
  (
    n984,
    n708,
    n702,
    n713,
    n806
  );


  xnor
  g1130
  (
    n1038,
    n663,
    n681,
    n778,
    n712
  );


  xor
  g1131
  (
    n1162,
    n659,
    n691,
    n662,
    n800
  );


  nor
  g1132
  (
    n1039,
    n690,
    n667,
    n726,
    n739
  );


  nand
  g1133
  (
    n981,
    n681,
    n739,
    n700,
    n703
  );


  or
  g1134
  (
    n1008,
    n692,
    n753,
    n707,
    n802
  );


  xnor
  g1135
  (
    n916,
    n809,
    n743,
    n787,
    n708
  );


  and
  g1136
  (
    n825,
    n723,
    n748,
    n754,
    n678
  );


  xnor
  g1137
  (
    n1075,
    n707,
    n675,
    n753,
    n761
  );


  nor
  g1138
  (
    n819,
    n676,
    n681,
    n744,
    n712
  );


  nor
  g1139
  (
    n1033,
    n674,
    n697,
    n776,
    n811
  );


  xnor
  g1140
  (
    n1132,
    n675,
    n779,
    n583,
    n803
  );


  nor
  g1141
  (
    n829,
    n768,
    n790,
    n732,
    n720
  );


  xor
  g1142
  (
    n1127,
    n747,
    n732,
    n805,
    n718
  );


  xor
  g1143
  (
    n1009,
    n712,
    n665,
    n784,
    n805
  );


  nand
  g1144
  (
    n1084,
    n774,
    n811,
    n706,
    n654
  );


  and
  g1145
  (
    n873,
    n679,
    n782,
    n768,
    n698
  );


  or
  g1146
  (
    n879,
    n667,
    n699,
    n725,
    n763
  );


  and
  g1147
  (
    n900,
    n663,
    n744,
    n786,
    n678
  );


  xor
  g1148
  (
    n1136,
    n776,
    n740,
    n659,
    n780
  );


  xor
  g1149
  (
    n1007,
    n706,
    n767,
    n657,
    n669
  );


  or
  g1150
  (
    n1072,
    n797,
    n735,
    n715,
    n685
  );


  nor
  g1151
  (
    n1242,
    n864,
    n1150,
    n897,
    n959
  );


  and
  g1152
  (
    KeyWire_0_4,
    n955,
    n1152,
    n1118,
    n1081
  );


  nand
  g1153
  (
    n1216,
    n1142,
    n983,
    n1085,
    n1160
  );


  or
  g1154
  (
    n1210,
    n881,
    n1117,
    n987,
    n831
  );


  nor
  g1155
  (
    n1220,
    n840,
    n835,
    n813,
    n997
  );


  nor
  g1156
  (
    n1235,
    n1091,
    n1073,
    n1070,
    n1068
  );


  and
  g1157
  (
    n1187,
    n850,
    n922,
    n1128,
    n940
  );


  nand
  g1158
  (
    n1192,
    n989,
    n925,
    n1138,
    n1054
  );


  nand
  g1159
  (
    n1260,
    n1082,
    n1129,
    n976,
    n1037
  );


  xor
  g1160
  (
    n1199,
    n1069,
    n885,
    n820,
    n1063
  );


  and
  g1161
  (
    n1270,
    n1016,
    n843,
    n1131,
    n601
  );


  and
  g1162
  (
    n1268,
    n969,
    n1042,
    n1161,
    n1155
  );


  nor
  g1163
  (
    n1182,
    n1130,
    n1076,
    n602,
    n848
  );


  or
  g1164
  (
    n1258,
    n960,
    n1014,
    n846,
    n839
  );


  nor
  g1165
  (
    n1236,
    n878,
    n1109,
    n952,
    n931
  );


  nand
  g1166
  (
    n1196,
    n823,
    n904,
    n944,
    n1162
  );


  and
  g1167
  (
    n1257,
    n1028,
    n893,
    n1088,
    n817
  );


  xnor
  g1168
  (
    n1185,
    n965,
    n819,
    n1079,
    n1001
  );


  xnor
  g1169
  (
    n1265,
    n837,
    n1163,
    n1030,
    n981
  );


  and
  g1170
  (
    n1239,
    n915,
    n1004,
    n1172,
    n1046
  );


  and
  g1171
  (
    n1225,
    n1043,
    n1025,
    n876,
    n1159
  );


  nand
  g1172
  (
    n1205,
    n891,
    n1021,
    n845,
    n1115
  );


  xor
  g1173
  (
    n1263,
    n1036,
    n886,
    n941,
    n936
  );


  and
  g1174
  (
    n1238,
    n1062,
    n911,
    n814,
    n1114
  );


  nand
  g1175
  (
    n1219,
    n1158,
    n1059,
    n1169,
    n870
  );


  or
  g1176
  (
    n1234,
    n921,
    n1136,
    n1065,
    n1072
  );


  and
  g1177
  (
    n1211,
    n907,
    n896,
    n1090,
    n1007
  );


  xor
  g1178
  (
    n1206,
    n834,
    n958,
    n1003,
    n1168
  );


  or
  g1179
  (
    n1197,
    n1011,
    n868,
    n1047,
    n1051
  );


  xor
  g1180
  (
    n1198,
    n929,
    n1145,
    n1008,
    n1040
  );


  xnor
  g1181
  (
    n1256,
    n1024,
    n1074,
    n1071,
    n949
  );


  nand
  g1182
  (
    n1223,
    n1092,
    n1015,
    n950,
    n1122
  );


  xnor
  g1183
  (
    n1233,
    n1141,
    n889,
    n903,
    n832
  );


  and
  g1184
  (
    n1246,
    n880,
    n866,
    n1018,
    n979
  );


  xor
  g1185
  (
    n1227,
    n1013,
    n875,
    n930,
    n900
  );


  nand
  g1186
  (
    n1221,
    n895,
    n838,
    n1098,
    n1107
  );


  or
  g1187
  (
    n1255,
    n1053,
    n905,
    n995,
    n522
  );


  xnor
  g1188
  (
    n1241,
    n602,
    n964,
    n914,
    n1166
  );


  xnor
  g1189
  (
    n1253,
    n934,
    n1135,
    n924,
    n888
  );


  xor
  g1190
  (
    n1231,
    n1097,
    n829,
    n1012,
    n1119
  );


  xnor
  g1191
  (
    n1217,
    n1056,
    n999,
    n1151,
    n827
  );


  xnor
  g1192
  (
    n1190,
    n1019,
    n1064,
    n894,
    n1132
  );


  xnor
  g1193
  (
    n1224,
    n816,
    n974,
    n1144,
    n1087
  );


  xor
  g1194
  (
    n1191,
    n1017,
    n1066,
    n1113,
    n991
  );


  xnor
  g1195
  (
    n1267,
    n1038,
    n986,
    n928,
    n1105
  );


  nor
  g1196
  (
    n1248,
    n871,
    n1165,
    n908,
    n1124
  );


  nand
  g1197
  (
    n1208,
    n917,
    n1026,
    n988,
    n1020
  );


  xor
  g1198
  (
    n1202,
    n1041,
    n882,
    n1174,
    n1078
  );


  nor
  g1199
  (
    n1230,
    n1034,
    n948,
    n1148,
    n856
  );


  xnor
  g1200
  (
    n1226,
    n978,
    n828,
    n927,
    n1133
  );


  nand
  g1201
  (
    n1245,
    n970,
    n1104,
    n935,
    n971
  );


  xnor
  g1202
  (
    n1249,
    n1127,
    n1173,
    n910,
    n1057
  );


  or
  g1203
  (
    n1215,
    n975,
    n869,
    n860,
    n1149
  );


  nand
  g1204
  (
    n1247,
    n1022,
    n902,
    n932,
    n602
  );


  or
  g1205
  (
    n1181,
    n883,
    n1045,
    n526,
    n1075
  );


  nor
  g1206
  (
    n1200,
    n879,
    n1094,
    n909,
    n1083
  );


  xnor
  g1207
  (
    n1232,
    n1171,
    n601,
    n1033,
    n873
  );


  xor
  g1208
  (
    n1203,
    n1099,
    n1061,
    n858,
    n1146
  );


  xnor
  g1209
  (
    n1264,
    n939,
    n874,
    n946,
    n992
  );


  and
  g1210
  (
    n1240,
    n825,
    n867,
    n1050,
    n1067
  );


  nor
  g1211
  (
    n1212,
    n977,
    n1111,
    n890,
    n1137
  );


  and
  g1212
  (
    n1195,
    n826,
    n1058,
    n945,
    n822
  );


  and
  g1213
  (
    n1207,
    n899,
    n525,
    n1010,
    n865
  );


  or
  g1214
  (
    n1201,
    n523,
    n877,
    n901,
    n1153
  );


  xnor
  g1215
  (
    n1259,
    n962,
    n824,
    n851,
    n1120
  );


  and
  g1216
  (
    n1229,
    n957,
    n967,
    n1006,
    n953
  );


  xnor
  g1217
  (
    n1237,
    n980,
    n815,
    n1123,
    n1005
  );


  and
  g1218
  (
    n1183,
    n859,
    n1035,
    n887,
    n1103
  );


  xnor
  g1219
  (
    n1177,
    n963,
    n1032,
    n861,
    n972
  );


  nor
  g1220
  (
    n1184,
    n1170,
    n990,
    n1009,
    n1101
  );


  or
  g1221
  (
    n1261,
    n884,
    n1089,
    n1125,
    n993
  );


  xnor
  g1222
  (
    n1252,
    n1084,
    n961,
    n601,
    n818
  );


  nor
  g1223
  (
    n1180,
    n1112,
    n1139,
    n951,
    n1077
  );


  nor
  g1224
  (
    n1186,
    n1167,
    n1044,
    n1096,
    n872
  );


  nor
  g1225
  (
    n1213,
    n855,
    n1023,
    n1140,
    n923
  );


  xnor
  g1226
  (
    n1262,
    n1086,
    n892,
    n842,
    n933
  );


  xor
  g1227
  (
    n1243,
    n926,
    n898,
    n906,
    n1156
  );


  nand
  g1228
  (
    n1222,
    n849,
    n857,
    n984,
    n985
  );


  xnor
  g1229
  (
    n1194,
    n1027,
    n821,
    n524,
    n1100
  );


  nor
  g1230
  (
    n1204,
    n847,
    n1126,
    n1121,
    n1000
  );


  nand
  g1231
  (
    n1209,
    n937,
    n1080,
    n1029,
    n916
  );


  xor
  g1232
  (
    n1266,
    n994,
    n982,
    n836,
    n919
  );


  xor
  g1233
  (
    n1193,
    n954,
    n1108,
    n998,
    n1134
  );


  or
  g1234
  (
    n1269,
    n1052,
    n833,
    n1102,
    n966
  );


  nand
  g1235
  (
    n1254,
    n1106,
    n1055,
    n956,
    n1060
  );


  nor
  g1236
  (
    n1251,
    n942,
    n1143,
    n1031,
    n1116
  );


  xnor
  g1237
  (
    n1214,
    n852,
    n854,
    n1175,
    n1049
  );


  xor
  g1238
  (
    n1188,
    n862,
    n920,
    n1164,
    n1157
  );


  or
  g1239
  (
    n1218,
    n1147,
    n1176,
    n943,
    n1110
  );


  and
  g1240
  (
    n1179,
    n938,
    n1048,
    n947,
    n973
  );


  nand
  g1241
  (
    n1250,
    n602,
    n853,
    n830,
    n1095
  );


  nand
  g1242
  (
    n1244,
    n912,
    n1093,
    n913,
    n863
  );


  and
  g1243
  (
    n1178,
    n1154,
    n918,
    n1039,
    n844
  );


  nor
  g1244
  (
    n1189,
    n841,
    n968,
    n1002,
    n996
  );


  not
  g1245
  (
    n1285,
    n1187
  );


  not
  g1246
  (
    n1275,
    n1228
  );


  buf
  g1247
  (
    n1314,
    n1216
  );


  buf
  g1248
  (
    n1311,
    n1229
  );


  not
  g1249
  (
    n1327,
    n1225
  );


  buf
  g1250
  (
    n1326,
    n1194
  );


  not
  g1251
  (
    n1301,
    n1183
  );


  not
  g1252
  (
    n1283,
    n1227
  );


  not
  g1253
  (
    n1273,
    n1179
  );


  buf
  g1254
  (
    n1286,
    n1195
  );


  buf
  g1255
  (
    n1320,
    n1201
  );


  not
  g1256
  (
    n1293,
    n1184
  );


  buf
  g1257
  (
    n1303,
    n1181
  );


  buf
  g1258
  (
    n1281,
    n1197
  );


  not
  g1259
  (
    n1296,
    n1214
  );


  buf
  g1260
  (
    n1294,
    n1186
  );


  not
  g1261
  (
    n1290,
    n1212
  );


  buf
  g1262
  (
    n1304,
    n1218
  );


  not
  g1263
  (
    n1277,
    n1204
  );


  not
  g1264
  (
    n1278,
    n1196
  );


  not
  g1265
  (
    n1315,
    n1198
  );


  buf
  g1266
  (
    n1292,
    n1232
  );


  not
  g1267
  (
    n1302,
    n1223
  );


  buf
  g1268
  (
    n1310,
    n1222
  );


  not
  g1269
  (
    n1305,
    n1219
  );


  buf
  g1270
  (
    n1280,
    n1211
  );


  buf
  g1271
  (
    n1298,
    n1189
  );


  buf
  g1272
  (
    n1282,
    n1185
  );


  buf
  g1273
  (
    n1312,
    n1192
  );


  buf
  g1274
  (
    n1317,
    n1217
  );


  buf
  g1275
  (
    n1291,
    n1206
  );


  buf
  g1276
  (
    n1288,
    n1188
  );


  buf
  g1277
  (
    n1325,
    n1203
  );


  not
  g1278
  (
    n1309,
    n1226
  );


  buf
  g1279
  (
    n1284,
    n1199
  );


  buf
  g1280
  (
    n1289,
    n1191
  );


  buf
  g1281
  (
    n1274,
    n1221
  );


  buf
  g1282
  (
    n1322,
    n1200
  );


  buf
  g1283
  (
    n1318,
    n1224
  );


  not
  g1284
  (
    n1287,
    n1177
  );


  not
  g1285
  (
    n1272,
    n1178
  );


  not
  g1286
  (
    n1328,
    n1210
  );


  buf
  g1287
  (
    n1316,
    n1202
  );


  not
  g1288
  (
    n1308,
    n1190
  );


  buf
  g1289
  (
    n1297,
    n1205
  );


  not
  g1290
  (
    n1300,
    n1220
  );


  buf
  g1291
  (
    n1279,
    n1182
  );


  not
  g1292
  (
    n1306,
    n1180
  );


  buf
  g1293
  (
    n1323,
    n1230
  );


  not
  g1294
  (
    n1271,
    n1208
  );


  buf
  g1295
  (
    n1276,
    n1209
  );


  not
  g1296
  (
    n1295,
    n1207
  );


  not
  g1297
  (
    n1313,
    n1231
  );


  not
  g1298
  (
    n1299,
    n1233
  );


  buf
  g1299
  (
    n1321,
    n1234
  );


  buf
  g1300
  (
    n1319,
    n1193
  );


  buf
  g1301
  (
    n1307,
    n1215
  );


  buf
  g1302
  (
    n1324,
    n1213
  );


  nand
  g1303
  (
    n1356,
    n1238,
    n1301,
    n1316
  );


  nand
  g1304
  (
    n1384,
    n1298,
    n242,
    n1318,
    n1276
  );


  xor
  g1305
  (
    KeyWire_0_3,
    n194,
    n248,
    n1314,
    n235
  );


  xnor
  g1306
  (
    n1380,
    n189,
    n1241,
    n1297,
    n1272
  );


  xnor
  g1307
  (
    n1381,
    n1325,
    n1248,
    n1286,
    n1273
  );


  nor
  g1308
  (
    n1397,
    n1321,
    n1298,
    n238,
    n1296
  );


  xnor
  g1309
  (
    n1360,
    n200,
    n1275,
    n1327,
    n1325
  );


  nand
  g1310
  (
    n1402,
    n1324,
    n1312,
    n1302,
    n1291
  );


  nor
  g1311
  (
    n1372,
    n1287,
    n1288,
    n1304,
    n1235
  );


  nand
  g1312
  (
    n1379,
    n239,
    n206,
    n1320,
    n218
  );


  nand
  g1313
  (
    n1370,
    n1307,
    n1322,
    n209,
    n528
  );


  nor
  g1314
  (
    n1339,
    n1328,
    n229,
    n247,
    n1284
  );


  xnor
  g1315
  (
    KeyWire_0_1,
    n205,
    n1246,
    n1322,
    n1283
  );


  xor
  g1316
  (
    n1338,
    n1245,
    n1317,
    n220,
    n1318
  );


  and
  g1317
  (
    n1364,
    n1300,
    n1249,
    n1323,
    n1299
  );


  and
  g1318
  (
    n1368,
    n1310,
    n1292,
    n1247,
    n1283
  );


  or
  g1319
  (
    n1378,
    n1323,
    n1277,
    n1282,
    n1275
  );


  xnor
  g1320
  (
    n1382,
    n1327,
    n1312,
    n1303
  );


  xnor
  g1321
  (
    n1399,
    n208,
    n258,
    n1274,
    n1276
  );


  nand
  g1322
  (
    n1351,
    n201,
    n1326,
    n533,
    n1297
  );


  xor
  g1323
  (
    n1391,
    n210,
    n1311,
    n1244,
    n226
  );


  and
  g1324
  (
    n1407,
    n214,
    n224,
    n1299,
    n211
  );


  nand
  g1325
  (
    n1373,
    n1289,
    n1289,
    n1277,
    n1272
  );


  or
  g1326
  (
    n1371,
    n215,
    n1304,
    n1281,
    n1319
  );


  or
  g1327
  (
    n1350,
    n1285,
    n1328,
    n1302,
    n233
  );


  or
  g1328
  (
    KeyWire_0_12,
    n1281,
    n1317,
    n1315,
    n1278
  );


  nor
  g1329
  (
    n1376,
    n190,
    n257,
    n1297,
    n1271
  );


  or
  g1330
  (
    n1359,
    n1305,
    n262,
    n532,
    n1278
  );


  xnor
  g1331
  (
    n1357,
    n1314,
    n1293,
    n1279,
    n228
  );


  xnor
  g1332
  (
    n1404,
    n1316,
    n199,
    n223,
    n1325
  );


  xnor
  g1333
  (
    n1366,
    n1286,
    n1324,
    n1314,
    n1298
  );


  and
  g1334
  (
    n1358,
    n216,
    n1315,
    n1294,
    n1283
  );


  xnor
  g1335
  (
    n1395,
    n1236,
    n1317,
    n1328,
    n195
  );


  and
  g1336
  (
    n1401,
    n1274,
    n1308,
    n1327,
    n1326
  );


  xnor
  g1337
  (
    n1353,
    n1307,
    n1275,
    n1294,
    n1305
  );


  and
  g1338
  (
    n1335,
    n243,
    n227,
    n1291,
    n1313
  );


  xnor
  g1339
  (
    n1329,
    n251,
    n1290,
    n1321,
    n1279
  );


  xor
  g1340
  (
    n1396,
    n236,
    n1324,
    n1271,
    n221
  );


  or
  g1341
  (
    n1405,
    n1305,
    n1287,
    n1308,
    n1309
  );


  xnor
  g1342
  (
    n1403,
    n212,
    n1313,
    n1323,
    n1271
  );


  nand
  g1343
  (
    n1400,
    n1313,
    n531,
    n1290,
    n198
  );


  xor
  g1344
  (
    n1365,
    n1318,
    n1306,
    n231,
    n1303
  );


  xor
  g1345
  (
    n1340,
    n1304,
    n1283,
    n1274,
    n1284
  );


  or
  g1346
  (
    n1394,
    n1292,
    n535,
    n1316,
    n261
  );


  xnor
  g1347
  (
    n1342,
    n1281,
    n1243,
    n256,
    n1306
  );


  nand
  g1348
  (
    n1333,
    n1242,
    n1306,
    n1303,
    n1278
  );


  and
  g1349
  (
    n1387,
    n249,
    n1325,
    n1299,
    n219
  );


  xor
  g1350
  (
    KeyWire_0_15,
    n1296,
    n322,
    n1324,
    n1312
  );


  nor
  g1351
  (
    n1410,
    n1327,
    n245,
    n1297,
    n202
  );


  xor
  g1352
  (
    n1385,
    n1309,
    n193,
    n197,
    n244
  );


  or
  g1353
  (
    n1388,
    n1272,
    n1240,
    n1301,
    n1311
  );


  xor
  g1354
  (
    n1383,
    n1319,
    n1296,
    n1285,
    n1289
  );


  nand
  g1355
  (
    n1336,
    n1307,
    n1280,
    n1322,
    n1308
  );


  nand
  g1356
  (
    n1331,
    n1290,
    n1293,
    n1307,
    n1301
  );


  nand
  g1357
  (
    n1346,
    n1309,
    n1271,
    n534,
    n260
  );


  and
  g1358
  (
    n1392,
    n1288,
    n213,
    n1273,
    n1319
  );


  xor
  g1359
  (
    n1367,
    n234,
    n1320,
    n1276,
    n1306
  );


  or
  g1360
  (
    n1408,
    n230,
    n1280,
    n1302,
    n1293
  );


  and
  g1361
  (
    n1409,
    n1298,
    n1294,
    n1302,
    n1295
  );


  nor
  g1362
  (
    KeyWire_0_5,
    n1311,
    n1276,
    n1304,
    n1279
  );


  xnor
  g1363
  (
    n1386,
    n1313,
    n222,
    n252,
    n1292
  );


  nand
  g1364
  (
    n1377,
    n1287,
    n1299,
    n1293,
    n1301
  );


  or
  g1365
  (
    n1332,
    n250,
    n1290,
    n1315,
    n529
  );


  nor
  g1366
  (
    n1389,
    n1280,
    n1280,
    n1326,
    n1300
  );


  nor
  g1367
  (
    n1345,
    n241,
    n1323,
    n1291,
    n1295
  );


  xor
  g1368
  (
    n1374,
    n217,
    n1295,
    n530,
    n1310
  );


  xor
  g1369
  (
    n1390,
    n1310,
    n1288,
    n225,
    n207
  );


  and
  g1370
  (
    n1341,
    n1321,
    n259,
    n1284,
    n1322
  );


  nor
  g1371
  (
    n1352,
    n1320,
    n1278,
    n204,
    n1291
  );


  xor
  g1372
  (
    n1348,
    n1309,
    n1279,
    n232,
    n1282
  );


  xor
  g1373
  (
    n1362,
    n196,
    n240,
    n1310,
    n1318
  );


  nor
  g1374
  (
    n1354,
    n253,
    n1321,
    n1294,
    n1315
  );


  nor
  g1375
  (
    n1398,
    n1311,
    n1285,
    n1300,
    n255
  );


  nor
  g1376
  (
    n1393,
    n1274,
    n1282,
    n1272,
    n1287
  );


  nor
  g1377
  (
    n1369,
    n1326,
    n254,
    n1288,
    n1285
  );


  nand
  g1378
  (
    n1347,
    n1281,
    n1296,
    n1286,
    n1277
  );


  nor
  g1379
  (
    n1330,
    n1303,
    n1308,
    n1320,
    n1305
  );


  and
  g1380
  (
    n1349,
    n1273,
    n1292,
    n1237,
    n203
  );


  xor
  g1381
  (
    n1344,
    n1317,
    n527,
    n1300,
    n246
  );


  nor
  g1382
  (
    n1411,
    n1277,
    n1314,
    n237,
    n1284
  );


  xnor
  g1383
  (
    n1406,
    n1319,
    n191,
    n1295,
    n1275
  );


  nor
  g1384
  (
    n1343,
    n192,
    n1286,
    n1328,
    n1239
  );


  nor
  g1385
  (
    n1363,
    n188,
    n1282,
    n1289,
    n1273
  );


  xnor
  g1386
  (
    n1437,
    n1368,
    n542,
    n1406,
    n1336
  );


  or
  g1387
  (
    n1419,
    n537,
    n1357,
    n1258,
    n290
  );


  xnor
  g1388
  (
    n1443,
    n1399,
    n1385,
    n1265,
    n1361
  );


  nand
  g1389
  (
    n1414,
    n290,
    n1330,
    n1261,
    n1411
  );


  nor
  g1390
  (
    n1431,
    n289,
    n1251,
    n1268,
    n1374
  );


  nand
  g1391
  (
    n1435,
    n1253,
    n1388,
    n1255,
    n1404
  );


  and
  g1392
  (
    n1428,
    n1262,
    n1354,
    n1379,
    n1386
  );


  nor
  g1393
  (
    n1433,
    n1337,
    n1376,
    n1398,
    n1334
  );


  or
  g1394
  (
    n1427,
    n1343,
    n1256,
    n1393,
    n1392
  );


  nand
  g1395
  (
    n1439,
    n1400,
    n287,
    n1329,
    n1333
  );


  or
  g1396
  (
    n1430,
    n287,
    n1341,
    n1391,
    n1367
  );


  and
  g1397
  (
    n1416,
    n1356,
    n539,
    n1364,
    n1401
  );


  nor
  g1398
  (
    n1415,
    n1397,
    n1410,
    n1335,
    n540
  );


  nor
  g1399
  (
    KeyWire_0_0,
    n1377,
    n1381,
    n1409,
    n1380
  );


  and
  g1400
  (
    n1429,
    n1366,
    n1396,
    n1344,
    n1370
  );


  xor
  g1401
  (
    n1424,
    n1359,
    n1353,
    n1263,
    n290
  );


  and
  g1402
  (
    n1413,
    n1346,
    n1362,
    n1378,
    n1383
  );


  nand
  g1403
  (
    n1434,
    n538,
    n1270,
    n1365,
    n1347
  );


  xnor
  g1404
  (
    n1442,
    n1259,
    n289,
    n1338,
    n287
  );


  and
  g1405
  (
    n1420,
    n290,
    n1363,
    n1349,
    n541
  );


  nand
  g1406
  (
    n1421,
    n1267,
    n1394,
    n1340,
    n1369
  );


  nor
  g1407
  (
    n1412,
    n1339,
    n1250,
    n1375,
    n289
  );


  nor
  g1408
  (
    n1436,
    n1373,
    n1348,
    n1389,
    n288
  );


  xnor
  g1409
  (
    n1418,
    n1372,
    n1358,
    n288,
    n1350
  );


  nand
  g1410
  (
    n1441,
    n1331,
    n1352,
    n1254,
    n1387
  );


  xor
  g1411
  (
    n1423,
    n1264,
    n1382,
    n1390,
    n536
  );


  or
  g1412
  (
    n1432,
    n1371,
    n1269,
    n288,
    n1266
  );


  nand
  g1413
  (
    n1422,
    n1260,
    n1252,
    n1402,
    n543
  );


  or
  g1414
  (
    n1425,
    n1407,
    n288,
    n1384,
    n1257
  );


  xor
  g1415
  (
    n1438,
    n289,
    n1395,
    n287,
    n1355
  );


  or
  g1416
  (
    n1440,
    n1408,
    n1403,
    n1360,
    n1351
  );


  or
  g1417
  (
    n1426,
    n1342,
    n1405,
    n1332,
    n1345
  );


  xnor
  g1418
  (
    n1445,
    n1431,
    n1430,
    n1437,
    n1425
  );


  xor
  g1419
  (
    n1451,
    n1414,
    n1429,
    n1441,
    n1424
  );


  xnor
  g1420
  (
    n1449,
    n1439,
    n1433,
    n1427,
    n1421
  );


  nor
  g1421
  (
    n1444,
    n1442,
    n1420,
    n1419,
    n1418
  );


  xor
  g1422
  (
    n1450,
    n1438,
    n1422,
    n1415,
    n1412
  );


  xor
  g1423
  (
    n1447,
    n1434,
    n1413,
    n1432,
    n1443
  );


  xor
  g1424
  (
    n1446,
    n1416,
    n1423,
    n1436,
    n1428
  );


  and
  g1425
  (
    n1448,
    n1417,
    n1426,
    n1440,
    n1435
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1417,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1361,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n59,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1334,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1228,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1355,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1055,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n460,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n989,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1148,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n89,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n853,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1337,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n598,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n532,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1375,
    KeyNOTWire_0_15
  );


endmodule


