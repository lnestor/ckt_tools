// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_2540_401 written by SynthGen on 2021/05/24 19:47:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_2540_401 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44,
 n940, n933, n939, n937, n926, n932, n938, n925,
 n935, n936, n931, n930, n929, n934, n2453, n2482,
 n2525, n2526, n2523, n2524, n2521, n2557, n2581, n2580,
 n2570, n2579, n2553, n2559, n2584, n2573, n2571, n2558,
 n2577, n2562, n2572, n2560, n2569, n2576, n2568, n2567,
 n2564, n2574, n2583, n2561, n2554, n2563, n2582, n2555,
 n2575, n2566, n2578, n2556, n2565);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44;

output n940, n933, n939, n937, n926, n932, n938, n925,
 n935, n936, n931, n930, n929, n934, n2453, n2482,
 n2525, n2526, n2523, n2524, n2521, n2557, n2581, n2580,
 n2570, n2579, n2553, n2559, n2584, n2573, n2571, n2558,
 n2577, n2562, n2572, n2560, n2569, n2576, n2568, n2567,
 n2564, n2574, n2583, n2561, n2554, n2563, n2582, n2555,
 n2575, n2566, n2578, n2556, n2565;

wire n45, n46, n47, n48, n49, n50, n51, n52,
 n53, n54, n55, n56, n57, n58, n59, n60,
 n61, n62, n63, n64, n65, n66, n67, n68,
 n69, n70, n71, n72, n73, n74, n75, n76,
 n77, n78, n79, n80, n81, n82, n83, n84,
 n85, n86, n87, n88, n89, n90, n91, n92,
 n93, n94, n95, n96, n97, n98, n99, n100,
 n101, n102, n103, n104, n105, n106, n107, n108,
 n109, n110, n111, n112, n113, n114, n115, n116,
 n117, n118, n119, n120, n121, n122, n123, n124,
 n125, n126, n127, n128, n129, n130, n131, n132,
 n133, n134, n135, n136, n137, n138, n139, n140,
 n141, n142, n143, n144, n145, n146, n147, n148,
 n149, n150, n151, n152, n153, n154, n155, n156,
 n157, n158, n159, n160, n161, n162, n163, n164,
 n165, n166, n167, n168, n169, n170, n171, n172,
 n173, n174, n175, n176, n177, n178, n179, n180,
 n181, n182, n183, n184, n185, n186, n187, n188,
 n189, n190, n191, n192, n193, n194, n195, n196,
 n197, n198, n199, n200, n201, n202, n203, n204,
 n205, n206, n207, n208, n209, n210, n211, n212,
 n213, n214, n215, n216, n217, n218, n219, n220,
 n221, n222, n223, n224, n225, n226, n227, n228,
 n229, n230, n231, n232, n233, n234, n235, n236,
 n237, n238, n239, n240, n241, n242, n243, n244,
 n245, n246, n247, n248, n249, n250, n251, n252,
 n253, n254, n255, n256, n257, n258, n259, n260,
 n261, n262, n263, n264, n265, n266, n267, n268,
 n269, n270, n271, n272, n273, n274, n275, n276,
 n277, n278, n279, n280, n281, n282, n283, n284,
 n285, n286, n287, n288, n289, n290, n291, n292,
 n293, n294, n295, n296, n297, n298, n299, n300,
 n301, n302, n303, n304, n305, n306, n307, n308,
 n309, n310, n311, n312, n313, n314, n315, n316,
 n317, n318, n319, n320, n321, n322, n323, n324,
 n325, n326, n327, n328, n329, n330, n331, n332,
 n333, n334, n335, n336, n337, n338, n339, n340,
 n341, n342, n343, n344, n345, n346, n347, n348,
 n349, n350, n351, n352, n353, n354, n355, n356,
 n357, n358, n359, n360, n361, n362, n363, n364,
 n365, n366, n367, n368, n369, n370, n371, n372,
 n373, n374, n375, n376, n377, n378, n379, n380,
 n381, n382, n383, n384, n385, n386, n387, n388,
 n389, n390, n391, n392, n393, n394, n395, n396,
 n397, n398, n399, n400, n401, n402, n403, n404,
 n405, n406, n407, n408, n409, n410, n411, n412,
 n413, n414, n415, n416, n417, n418, n419, n420,
 n421, n422, n423, n424, n425, n426, n427, n428,
 n429, n430, n431, n432, n433, n434, n435, n436,
 n437, n438, n439, n440, n441, n442, n443, n444,
 n445, n446, n447, n448, n449, n450, n451, n452,
 n453, n454, n455, n456, n457, n458, n459, n460,
 n461, n462, n463, n464, n465, n466, n467, n468,
 n469, n470, n471, n472, n473, n474, n475, n476,
 n477, n478, n479, n480, n481, n482, n483, n484,
 n485, n486, n487, n488, n489, n490, n491, n492,
 n493, n494, n495, n496, n497, n498, n499, n500,
 n501, n502, n503, n504, n505, n506, n507, n508,
 n509, n510, n511, n512, n513, n514, n515, n516,
 n517, n518, n519, n520, n521, n522, n523, n524,
 n525, n526, n527, n528, n529, n530, n531, n532,
 n533, n534, n535, n536, n537, n538, n539, n540,
 n541, n542, n543, n544, n545, n546, n547, n548,
 n549, n550, n551, n552, n553, n554, n555, n556,
 n557, n558, n559, n560, n561, n562, n563, n564,
 n565, n566, n567, n568, n569, n570, n571, n572,
 n573, n574, n575, n576, n577, n578, n579, n580,
 n581, n582, n583, n584, n585, n586, n587, n588,
 n589, n590, n591, n592, n593, n594, n595, n596,
 n597, n598, n599, n600, n601, n602, n603, n604,
 n605, n606, n607, n608, n609, n610, n611, n612,
 n613, n614, n615, n616, n617, n618, n619, n620,
 n621, n622, n623, n624, n625, n626, n627, n628,
 n629, n630, n631, n632, n633, n634, n635, n636,
 n637, n638, n639, n640, n641, n642, n643, n644,
 n645, n646, n647, n648, n649, n650, n651, n652,
 n653, n654, n655, n656, n657, n658, n659, n660,
 n661, n662, n663, n664, n665, n666, n667, n668,
 n669, n670, n671, n672, n673, n674, n675, n676,
 n677, n678, n679, n680, n681, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n758, n759, n760, n761, n762, n763, n764,
 n765, n766, n767, n768, n769, n770, n771, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n865, n866, n867, n868,
 n869, n870, n871, n872, n873, n874, n875, n876,
 n877, n878, n879, n880, n881, n882, n883, n884,
 n885, n886, n887, n888, n889, n890, n891, n892,
 n893, n894, n895, n896, n897, n898, n899, n900,
 n901, n902, n903, n904, n905, n906, n907, n908,
 n909, n910, n911, n912, n913, n914, n915, n916,
 n917, n918, n919, n920, n921, n922, n923, n924,
 n927, n928, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
 n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
 n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
 n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
 n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
 n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
 n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
 n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
 n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
 n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
 n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
 n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
 n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
 n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
 n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
 n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
 n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
 n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
 n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
 n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
 n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
 n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
 n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
 n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
 n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
 n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
 n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
 n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
 n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
 n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
 n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
 n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
 n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
 n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
 n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
 n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
 n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
 n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
 n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
 n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
 n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
 n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
 n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
 n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
 n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
 n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
 n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
 n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
 n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
 n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
 n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
 n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
 n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
 n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
 n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
 n2451, n2452, n2454, n2455, n2456, n2457, n2458, n2459,
 n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
 n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
 n2476, n2477, n2478, n2479, n2480, n2481, n2483, n2484,
 n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
 n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
 n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
 n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
 n2517, n2518, n2519, n2520, n2522, n2527, n2528, n2529,
 n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
 n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
 n2546, n2547, n2548, n2549, n2550, n2551, n2552;

buf  g0 (n206, n33);
not  g1 (n174, n33);
buf  g2 (n53, n4);
not  g3 (n186, n24);
not  g4 (n175, n19);
not  g5 (n69, n39);
not  g6 (n161, n15);
buf  g7 (n201, n39);
buf  g8 (n97, n15);
not  g9 (n103, n23);
buf  g10 (n105, n35);
not  g11 (n200, n26);
not  g12 (n57, n29);
buf  g13 (n124, n3);
buf  g14 (n156, n34);
not  g15 (n169, n6);
not  g16 (n157, n4);
buf  g17 (n94, n35);
not  g18 (n195, n42);
not  g19 (n77, n12);
not  g20 (n134, n36);
buf  g21 (n179, n12);
not  g22 (n80, n22);
buf  g23 (n145, n7);
not  g24 (n135, n44);
not  g25 (n99, n23);
buf  g26 (n146, n31);
not  g27 (n55, n8);
not  g28 (n81, n14);
not  g29 (n207, n10);
buf  g30 (n108, n23);
buf  g31 (n216, n5);
not  g32 (n117, n35);
buf  g33 (n164, n18);
buf  g34 (n180, n19);
not  g35 (n190, n11);
not  g36 (n49, n41);
not  g37 (n59, n20);
not  g38 (n155, n25);
buf  g39 (n126, n11);
buf  g40 (n88, n39);
buf  g41 (n170, n27);
buf  g42 (n107, n14);
buf  g43 (n65, n2);
buf  g44 (n106, n10);
not  g45 (n158, n17);
not  g46 (n139, n43);
not  g47 (n220, n8);
buf  g48 (n79, n9);
buf  g49 (n178, n36);
not  g50 (n185, n38);
buf  g51 (n149, n38);
not  g52 (n148, n8);
not  g53 (n151, n20);
not  g54 (n188, n31);
buf  g55 (n165, n17);
buf  g56 (n93, n41);
not  g57 (n120, n40);
buf  g58 (n127, n22);
buf  g59 (n109, n10);
not  g60 (n172, n33);
buf  g61 (n160, n26);
buf  g62 (n152, n40);
not  g63 (n154, n13);
not  g64 (n136, n6);
buf  g65 (n193, n19);
buf  g66 (n219, n17);
buf  g67 (n52, n11);
buf  g68 (n202, n9);
buf  g69 (n75, n16);
not  g70 (n101, n21);
not  g71 (n47, n34);
buf  g72 (n64, n8);
buf  g73 (n67, n14);
buf  g74 (n138, n43);
buf  g75 (n153, n25);
not  g76 (n45, n10);
not  g77 (n144, n44);
buf  g78 (n111, n19);
buf  g79 (n210, n18);
buf  g80 (n192, n15);
buf  g81 (n209, n7);
buf  g82 (n159, n32);
buf  g83 (n184, n38);
buf  g84 (n114, n6);
not  g85 (n133, n24);
not  g86 (n68, n21);
buf  g87 (n205, n25);
not  g88 (n62, n13);
buf  g89 (n95, n44);
buf  g90 (n168, n24);
not  g91 (n96, n35);
buf  g92 (n87, n1);
buf  g93 (n183, n18);
buf  g94 (n167, n29);
buf  g95 (n121, n41);
buf  g96 (n171, n4);
buf  g97 (n91, n5);
not  g98 (n177, n16);
not  g99 (n66, n44);
buf  g100 (n83, n21);
buf  g101 (n70, n2);
not  g102 (n60, n28);
buf  g103 (n58, n41);
buf  g104 (n74, n30);
buf  g105 (n50, n37);
buf  g106 (n173, n26);
not  g107 (n214, n39);
buf  g108 (n213, n40);
buf  g109 (n181, n42);
not  g110 (n56, n36);
not  g111 (n76, n11);
buf  g112 (n182, n13);
not  g113 (n116, n22);
buf  g114 (n54, n9);
buf  g115 (n208, n1);
not  g116 (n51, n23);
not  g117 (n166, n3);
buf  g118 (n85, n42);
buf  g119 (n217, n40);
buf  g120 (n199, n43);
not  g121 (n46, n15);
not  g122 (n113, n20);
buf  g123 (n78, n43);
not  g124 (n176, n1);
buf  g125 (n131, n2);
not  g126 (n84, n3);
not  g127 (n82, n30);
buf  g128 (n72, n27);
not  g129 (n204, n34);
buf  g130 (n104, n37);
not  g131 (n128, n7);
buf  g132 (n129, n32);
not  g133 (n141, n4);
not  g134 (n102, n29);
not  g135 (n147, n12);
buf  g136 (n163, n30);
buf  g137 (n196, n36);
not  g138 (n90, n38);
not  g139 (n197, n21);
not  g140 (n137, n20);
not  g141 (n118, n16);
buf  g142 (n140, n28);
buf  g143 (n86, n18);
not  g144 (n73, n9);
buf  g145 (n189, n7);
buf  g146 (n122, n26);
not  g147 (n119, n3);
buf  g148 (n130, n28);
buf  g149 (n71, n16);
buf  g150 (n194, n17);
buf  g151 (n100, n32);
not  g152 (n48, n27);
buf  g153 (n92, n24);
not  g154 (n211, n33);
not  g155 (n150, n34);
buf  g156 (n198, n14);
not  g157 (n63, n37);
buf  g158 (n212, n31);
not  g159 (n203, n32);
buf  g160 (n162, n37);
buf  g161 (n89, n27);
not  g162 (n123, n6);
buf  g163 (n215, n25);
not  g164 (n218, n13);
buf  g165 (n112, n12);
not  g166 (n132, n5);
buf  g167 (n125, n28);
not  g168 (n98, n2);
not  g169 (n115, n42);
buf  g170 (n110, n31);
not  g171 (n142, n29);
not  g172 (n191, n30);
buf  g173 (n187, n5);
not  g174 (n61, n22);
not  g175 (n143, n1);
not  g176 (n779, n125);
not  g177 (n431, n102);
buf  g178 (n577, n133);
buf  g179 (n556, n194);
not  g180 (n870, n101);
not  g181 (n254, n59);
not  g182 (n402, n176);
buf  g183 (n253, n178);
not  g184 (n524, n157);
buf  g185 (n643, n70);
buf  g186 (n889, n209);
not  g187 (n351, n86);
not  g188 (n799, n179);
not  g189 (n442, n158);
not  g190 (n589, n48);
not  g191 (n644, n152);
buf  g192 (n356, n170);
not  g193 (n774, n171);
buf  g194 (n624, n71);
buf  g195 (n848, n54);
not  g196 (n382, n182);
buf  g197 (n464, n100);
not  g198 (n626, n56);
buf  g199 (n830, n126);
buf  g200 (n560, n140);
not  g201 (n623, n167);
buf  g202 (n318, n200);
buf  g203 (n581, n76);
not  g204 (n437, n60);
not  g205 (n653, n98);
buf  g206 (n518, n77);
buf  g207 (n855, n86);
not  g208 (n270, n146);
not  g209 (n882, n52);
not  g210 (n311, n81);
buf  g211 (n479, n220);
buf  g212 (n233, n53);
buf  g213 (n664, n89);
buf  g214 (n591, n143);
not  g215 (n923, n85);
buf  g216 (n618, n170);
buf  g217 (n521, n197);
buf  g218 (n338, n70);
buf  g219 (n661, n101);
not  g220 (n527, n205);
not  g221 (n459, n168);
buf  g222 (n497, n99);
buf  g223 (n597, n94);
not  g224 (n908, n85);
not  g225 (n328, n73);
not  g226 (n612, n63);
buf  g227 (n826, n161);
not  g228 (n852, n218);
buf  g229 (n388, n164);
buf  g230 (n666, n45);
buf  g231 (n236, n219);
not  g232 (n372, n183);
buf  g233 (n821, n104);
not  g234 (n566, n214);
not  g235 (n361, n198);
not  g236 (n456, n83);
not  g237 (n244, n83);
not  g238 (n801, n140);
not  g239 (n829, n174);
not  g240 (n895, n47);
not  g241 (n691, n46);
buf  g242 (n627, n51);
buf  g243 (n711, n88);
buf  g244 (n505, n158);
not  g245 (n540, n96);
buf  g246 (n645, n175);
buf  g247 (n400, n79);
buf  g248 (n884, n104);
buf  g249 (n632, n53);
buf  g250 (n559, n169);
not  g251 (n552, n194);
buf  g252 (n547, n81);
buf  g253 (n381, n86);
not  g254 (n704, n217);
buf  g255 (n648, n57);
not  g256 (n256, n204);
buf  g257 (n782, n219);
buf  g258 (n385, n60);
not  g259 (n708, n193);
buf  g260 (n777, n197);
buf  g261 (n323, n72);
not  g262 (n823, n164);
not  g263 (n384, n191);
buf  g264 (n430, n82);
buf  g265 (n657, n67);
buf  g266 (n476, n142);
buf  g267 (n449, n106);
buf  g268 (n322, n93);
buf  g269 (n425, n50);
buf  g270 (n592, n184);
buf  g271 (n865, n177);
not  g272 (n825, n182);
not  g273 (n668, n71);
buf  g274 (n802, n210);
not  g275 (n791, n216);
buf  g276 (n881, n80);
not  g277 (n788, n132);
not  g278 (n488, n118);
buf  g279 (n490, n127);
not  g280 (n421, n84);
not  g281 (n371, n161);
not  g282 (n506, n103);
not  g283 (n586, n220);
buf  g284 (n780, n187);
not  g285 (n611, n81);
buf  g286 (n641, n149);
buf  g287 (n733, n92);
buf  g288 (n416, n94);
buf  g289 (n266, n207);
not  g290 (n501, n84);
not  g291 (n575, n48);
buf  g292 (n580, n186);
not  g293 (n241, n55);
buf  g294 (n740, n73);
not  g295 (n271, n163);
buf  g296 (n637, n123);
buf  g297 (n665, n155);
buf  g298 (n463, n216);
not  g299 (n550, n149);
not  g300 (n346, n55);
not  g301 (n427, n201);
not  g302 (n681, n106);
buf  g303 (n498, n85);
not  g304 (n485, n109);
buf  g305 (n594, n180);
buf  g306 (n838, n133);
buf  g307 (n538, n200);
buf  g308 (n806, n63);
buf  g309 (n844, n187);
buf  g310 (n869, n165);
not  g311 (n370, n66);
not  g312 (n342, n103);
buf  g313 (n707, n47);
not  g314 (n755, n87);
not  g315 (n878, n63);
buf  g316 (n794, n151);
not  g317 (n900, n185);
buf  g318 (n348, n54);
buf  g319 (n268, n167);
buf  g320 (n763, n208);
buf  g321 (n819, n200);
buf  g322 (n365, n108);
not  g323 (n354, n195);
not  g324 (n562, n100);
buf  g325 (n746, n99);
not  g326 (n689, n145);
not  g327 (n719, n196);
buf  g328 (n533, n52);
not  g329 (n724, n213);
not  g330 (n451, n53);
not  g331 (n263, n153);
buf  g332 (n678, n189);
not  g333 (n636, n56);
not  g334 (n658, n209);
not  g335 (n810, n115);
buf  g336 (n532, n214);
buf  g337 (n894, n49);
buf  g338 (n410, n117);
buf  g339 (n396, n188);
buf  g340 (n906, n58);
not  g341 (n325, n134);
not  g342 (n745, n140);
not  g343 (n567, n99);
not  g344 (n776, n82);
not  g345 (n863, n67);
not  g346 (n907, n116);
buf  g347 (n287, n212);
buf  g348 (n602, n168);
buf  g349 (n883, n71);
not  g350 (n734, n152);
not  g351 (n903, n195);
buf  g352 (n548, n138);
not  g353 (n500, n189);
not  g354 (n234, n71);
buf  g355 (n748, n171);
not  g356 (n596, n87);
buf  g357 (n905, n105);
not  g358 (n625, n121);
not  g359 (n327, n164);
buf  g360 (n433, n208);
not  g361 (n712, n115);
not  g362 (n670, n88);
not  g363 (n753, n55);
not  g364 (n549, n215);
not  g365 (n605, n80);
not  g366 (n687, n75);
buf  g367 (n909, n175);
buf  g368 (n457, n59);
buf  g369 (n230, n72);
buf  g370 (n887, n60);
not  g371 (n781, n176);
buf  g372 (n474, n141);
not  g373 (n531, n145);
buf  g374 (n555, n145);
buf  g375 (n293, n215);
not  g376 (n279, n188);
not  g377 (n335, n50);
not  g378 (n713, n183);
buf  g379 (n699, n139);
buf  g380 (n743, n215);
buf  g381 (n758, n141);
buf  g382 (n303, n211);
buf  g383 (n697, n203);
not  g384 (n873, n159);
not  g385 (n890, n179);
buf  g386 (n285, n165);
buf  g387 (n647, n191);
buf  g388 (n579, n129);
not  g389 (n493, n201);
not  g390 (n248, n96);
buf  g391 (n675, n75);
buf  g392 (n616, n148);
not  g393 (n920, n138);
not  g394 (n496, n127);
buf  g395 (n423, n64);
not  g396 (n811, n82);
buf  g397 (n332, n165);
buf  g398 (n409, n82);
buf  g399 (n642, n181);
buf  g400 (n470, n186);
not  g401 (n720, n192);
buf  g402 (n911, n109);
not  g403 (n314, n68);
not  g404 (n320, n113);
buf  g405 (n854, n157);
not  g406 (n761, n174);
not  g407 (n840, n168);
not  g408 (n765, n120);
buf  g409 (n558, n62);
not  g410 (n366, n48);
buf  g411 (n390, n182);
buf  g412 (n565, n144);
buf  g413 (n759, n113);
buf  g414 (n630, n114);
not  g415 (n570, n52);
buf  g416 (n918, n151);
not  g417 (n585, n159);
not  g418 (n462, n147);
not  g419 (n897, n217);
not  g420 (n526, n93);
buf  g421 (n688, n132);
buf  g422 (n291, n148);
not  g423 (n917, n129);
not  g424 (n726, n183);
not  g425 (n814, n122);
not  g426 (n730, n79);
not  g427 (n676, n108);
buf  g428 (n795, n106);
not  g429 (n617, n163);
buf  g430 (n387, n206);
buf  g431 (n503, n182);
buf  g432 (n242, n198);
buf  g433 (n283, n119);
buf  g434 (n329, n208);
buf  g435 (n317, n199);
not  g436 (n252, n130);
not  g437 (n334, n65);
buf  g438 (n709, n197);
buf  g439 (n672, n47);
not  g440 (n715, n136);
buf  g441 (n249, n126);
not  g442 (n614, n55);
not  g443 (n340, n59);
not  g444 (n921, n50);
buf  g445 (n621, n147);
not  g446 (n478, n62);
buf  g447 (n404, n169);
not  g448 (n519, n74);
not  g449 (n834, n73);
not  g450 (n510, n61);
not  g451 (n640, n138);
buf  g452 (n770, n154);
not  g453 (n523, n137);
not  g454 (n288, n104);
not  g455 (n495, n207);
buf  g456 (n662, n70);
not  g457 (n359, n49);
not  g458 (n835, n213);
not  g459 (n245, n216);
buf  g460 (n888, n131);
not  g461 (n786, n173);
not  g462 (n696, n210);
buf  g463 (n654, n95);
not  g464 (n871, n75);
buf  g465 (n259, n168);
not  g466 (n362, n172);
buf  g467 (n557, n131);
buf  g468 (n480, n48);
buf  g469 (n729, n87);
not  g470 (n435, n73);
buf  g471 (n635, n180);
buf  g472 (n899, n101);
not  g473 (n751, n123);
buf  g474 (n756, n119);
buf  g475 (n564, n205);
not  g476 (n659, n104);
buf  g477 (n492, n187);
buf  g478 (n828, n136);
buf  g479 (n554, n170);
buf  g480 (n536, n61);
buf  g481 (n639, n109);
buf  g482 (n469, n97);
not  g483 (n284, n167);
buf  g484 (n764, n112);
buf  g485 (n273, n214);
not  g486 (n376, n200);
buf  g487 (n880, n181);
not  g488 (n842, n75);
buf  g489 (n484, n204);
buf  g490 (n534, n126);
not  g491 (n750, n157);
buf  g492 (n595, n91);
buf  g493 (n299, n151);
buf  g494 (n649, n164);
not  g495 (n762, n173);
not  g496 (n238, n141);
not  g497 (n336, n202);
not  g498 (n499, n115);
not  g499 (n778, n118);
buf  g500 (n491, n143);
not  g501 (n306, n83);
buf  g502 (n913, n155);
buf  g503 (n584, n120);
not  g504 (n267, n45);
not  g505 (n784, n72);
buf  g506 (n783, n57);
not  g507 (n403, n85);
buf  g508 (n282, n74);
buf  g509 (n298, n163);
not  g510 (n374, n215);
not  g511 (n415, n100);
buf  g512 (n448, n64);
buf  g513 (n467, n203);
buf  g514 (n544, n68);
buf  g515 (n603, n185);
buf  g516 (n789, n155);
not  g517 (n805, n177);
not  g518 (n693, n197);
not  g519 (n465, n63);
buf  g520 (n773, n188);
buf  g521 (n702, n172);
not  g522 (n680, n51);
not  g523 (n551, n84);
not  g524 (n700, n149);
buf  g525 (n766, n179);
not  g526 (n772, n190);
not  g527 (n226, n84);
not  g528 (n522, n95);
not  g529 (n604, n91);
buf  g530 (n578, n146);
not  g531 (n669, n125);
not  g532 (n486, n190);
not  g533 (n331, n207);
buf  g534 (n915, n112);
buf  g535 (n429, n144);
buf  g536 (n414, n134);
not  g537 (n378, n133);
buf  g538 (n235, n122);
buf  g539 (n258, n132);
not  g540 (n877, n111);
buf  g541 (n228, n122);
not  g542 (n754, n94);
buf  g543 (n651, n132);
not  g544 (n695, n46);
not  g545 (n481, n142);
buf  g546 (n296, n125);
buf  g547 (n598, n201);
not  g548 (n512, n169);
not  g549 (n701, n66);
not  g550 (n265, n119);
not  g551 (n922, n120);
buf  g552 (n817, n177);
not  g553 (n418, n78);
buf  g554 (n309, n80);
buf  g555 (n790, n51);
not  g556 (n482, n66);
buf  g557 (n793, n89);
buf  g558 (n326, n96);
not  g559 (n399, n181);
buf  g560 (n816, n128);
buf  g561 (n694, n118);
not  g562 (n760, n174);
not  g563 (n721, n97);
not  g564 (n441, n195);
buf  g565 (n440, n136);
buf  g566 (n407, n86);
not  g567 (n477, n188);
not  g568 (n568, n191);
buf  g569 (n910, n61);
not  g570 (n690, n176);
not  g571 (n445, n165);
not  g572 (n472, n134);
buf  g573 (n247, n95);
buf  g574 (n833, n100);
not  g575 (n898, n193);
buf  g576 (n847, n206);
buf  g577 (n798, n156);
not  g578 (n892, n107);
buf  g579 (n367, n64);
buf  g580 (n237, n76);
buf  g581 (n741, n114);
buf  g582 (n785, n184);
buf  g583 (n227, n147);
not  g584 (n674, n169);
not  g585 (n804, n159);
not  g586 (n861, n64);
not  g587 (n858, n139);
not  g588 (n539, n166);
not  g589 (n722, n98);
not  g590 (n446, n107);
buf  g591 (n357, n160);
not  g592 (n737, n78);
not  g593 (n671, n123);
not  g594 (n269, n68);
buf  g595 (n358, n199);
not  g596 (n677, n56);
not  g597 (n364, n202);
not  g598 (n633, n49);
buf  g599 (n638, n162);
buf  g600 (n800, n192);
not  g601 (n412, n90);
buf  g602 (n663, n152);
buf  g603 (n321, n116);
not  g604 (n885, n126);
not  g605 (n489, n208);
not  g606 (n525, n51);
buf  g607 (n386, n119);
not  g608 (n432, n108);
not  g609 (n276, n212);
not  g610 (n593, n91);
buf  g611 (n839, n202);
not  g612 (n347, n191);
not  g613 (n901, n130);
buf  g614 (n406, n151);
buf  g615 (n319, n128);
buf  g616 (n822, n130);
not  g617 (n391, n149);
not  g618 (n727, n220);
buf  g619 (n808, n76);
not  g620 (n454, n74);
buf  g621 (n243, n66);
buf  g622 (n812, n184);
not  g623 (n514, n158);
buf  g624 (n373, n88);
not  g625 (n608, n62);
buf  g626 (n845, n120);
not  g627 (n610, n83);
buf  g628 (n535, n199);
buf  g629 (n606, n56);
buf  g630 (n316, n178);
not  g631 (n718, n203);
buf  g632 (n458, n190);
not  g633 (n893, n156);
buf  g634 (n511, n45);
not  g635 (n389, n105);
not  g636 (n420, n58);
not  g637 (n260, n217);
buf  g638 (n221, n72);
not  g639 (n424, n102);
not  g640 (n301, n87);
buf  g641 (n286, n212);
buf  g642 (n582, n113);
buf  g643 (n857, n98);
buf  g644 (n747, n144);
buf  g645 (n428, n118);
not  g646 (n815, n47);
not  g647 (n600, n160);
not  g648 (n613, n65);
buf  g649 (n652, n65);
buf  g650 (n588, n111);
not  g651 (n343, n124);
not  g652 (n629, n127);
buf  g653 (n239, n124);
not  g654 (n601, n213);
not  g655 (n487, n115);
not  g656 (n300, n57);
not  g657 (n703, n74);
not  g658 (n546, n198);
buf  g659 (n914, n198);
buf  g660 (n438, n194);
buf  g661 (n820, n181);
buf  g662 (n450, n144);
not  g663 (n257, n163);
buf  g664 (n561, n99);
buf  g665 (n516, n219);
not  g666 (n660, n136);
not  g667 (n609, n205);
buf  g668 (n867, n187);
buf  g669 (n509, n117);
not  g670 (n728, n97);
not  g671 (n723, n219);
buf  g672 (n836, n220);
not  g673 (n411, n199);
not  g674 (n813, n186);
buf  g675 (n231, n79);
buf  g676 (n818, n107);
not  g677 (n380, n121);
not  g678 (n471, n159);
buf  g679 (n422, n138);
not  g680 (n856, n111);
buf  g681 (n650, n210);
buf  g682 (n307, n141);
buf  g683 (n573, n192);
not  g684 (n732, n69);
not  g685 (n655, n173);
buf  g686 (n851, n171);
buf  g687 (n792, n171);
buf  g688 (n731, n79);
buf  g689 (n530, n93);
not  g690 (n912, n117);
buf  g691 (n305, n58);
buf  g692 (n902, n112);
buf  g693 (n853, n150);
buf  g694 (n809, n94);
not  g695 (n513, n54);
buf  g696 (n543, n90);
not  g697 (n735, n150);
buf  g698 (n916, n93);
buf  g699 (n872, n78);
buf  g700 (n736, n209);
not  g701 (n308, n175);
not  g702 (n686, n196);
buf  g703 (n345, n114);
buf  g704 (n904, n175);
not  g705 (n274, n123);
not  g706 (n831, n192);
buf  g707 (n222, n77);
not  g708 (n744, n166);
buf  g709 (n864, n189);
buf  g710 (n483, n92);
not  g711 (n698, n140);
buf  g712 (n607, n69);
not  g713 (n824, n97);
not  g714 (n837, n166);
buf  g715 (n827, n46);
buf  g716 (n310, n76);
buf  g717 (n769, n217);
not  g718 (n599, n162);
buf  g719 (n896, n112);
buf  g720 (n290, n194);
not  g721 (n859, n189);
not  g722 (n355, n213);
buf  g723 (n504, n113);
buf  g724 (n466, n210);
buf  g725 (n280, n203);
not  g726 (n710, n67);
not  g727 (n443, n90);
not  g728 (n537, n161);
not  g729 (n297, n110);
buf  g730 (n807, n124);
not  g731 (n225, n129);
not  g732 (n337, n162);
not  g733 (n375, n135);
buf  g734 (n520, n176);
not  g735 (n344, n135);
not  g736 (n460, n205);
buf  g737 (n315, n206);
buf  g738 (n405, n185);
not  g739 (n545, n160);
buf  g740 (n368, n178);
buf  g741 (n393, n135);
not  g742 (n352, n110);
buf  g743 (n379, n90);
not  g744 (n333, n161);
not  g745 (n574, n125);
not  g746 (n294, n172);
not  g747 (n563, n172);
not  g748 (n330, n214);
not  g749 (n875, n167);
not  g750 (n289, n59);
buf  g751 (n886, n105);
not  g752 (n716, n142);
not  g753 (n706, n178);
not  g754 (n313, n180);
buf  g755 (n725, n158);
buf  g756 (n656, n102);
not  g757 (n796, n49);
not  g758 (n787, n154);
not  g759 (n646, n177);
buf  g760 (n277, n154);
not  g761 (n508, n131);
not  g762 (n246, n143);
not  g763 (n705, n146);
not  g764 (n572, n150);
buf  g765 (n395, n130);
buf  g766 (n860, n128);
buf  g767 (n583, n69);
buf  g768 (n324, n134);
not  g769 (n667, n218);
buf  g770 (n302, n62);
not  g771 (n576, n70);
buf  g772 (n717, n101);
not  g773 (n541, n68);
buf  g774 (n281, n77);
not  g775 (n223, n81);
not  g776 (n620, n139);
not  g777 (n874, n170);
not  g778 (n507, n186);
not  g779 (n419, n216);
buf  g780 (n742, n179);
not  g781 (n862, n92);
buf  g782 (n797, n122);
not  g783 (n590, n92);
not  g784 (n615, n160);
not  g785 (n517, n153);
not  g786 (n803, n103);
buf  g787 (n846, n148);
buf  g788 (n240, n80);
not  g789 (n292, n61);
not  g790 (n312, n109);
buf  g791 (n455, n204);
buf  g792 (n866, n65);
buf  g793 (n229, n190);
not  g794 (n569, n206);
buf  g795 (n383, n193);
not  g796 (n444, n155);
buf  g797 (n679, n209);
buf  g798 (n377, n98);
buf  g799 (n752, n116);
not  g800 (n473, n121);
not  g801 (n439, n212);
buf  g802 (n587, n147);
buf  g803 (n397, n148);
not  g804 (n502, n89);
not  g805 (n394, n143);
not  g806 (n261, n67);
buf  g807 (n738, n46);
buf  g808 (n684, n78);
not  g809 (n553, n105);
buf  g810 (n571, n180);
buf  g811 (n275, n89);
buf  g812 (n255, n121);
not  g813 (n891, n91);
buf  g814 (n749, n201);
buf  g815 (n232, n102);
buf  g816 (n841, n207);
not  g817 (n628, n145);
not  g818 (n768, n139);
buf  g819 (n622, n137);
buf  g820 (n879, n106);
not  g821 (n634, n166);
buf  g822 (n673, n173);
buf  g823 (n775, n60);
not  g824 (n434, n117);
not  g825 (n876, n114);
not  g826 (n919, n108);
buf  g827 (n461, n50);
not  g828 (n529, n116);
not  g829 (n264, n195);
buf  g830 (n251, n57);
not  g831 (n843, n153);
not  g832 (n417, n135);
not  g833 (n452, n193);
buf  g834 (n542, n77);
buf  g835 (n447, n146);
buf  g836 (n369, n103);
not  g837 (n341, n204);
buf  g838 (n224, n54);
buf  g839 (n360, n183);
buf  g840 (n692, n45);
buf  g841 (n849, n196);
not  g842 (n924, n128);
not  g843 (n631, n52);
not  g844 (n350, n129);
not  g845 (n832, n142);
buf  g846 (n757, n150);
buf  g847 (n295, n218);
not  g848 (n250, n162);
not  g849 (n426, n107);
buf  g850 (n685, n184);
buf  g851 (n408, n202);
buf  g852 (n353, n110);
buf  g853 (n475, n69);
buf  g854 (n398, n111);
not  g855 (n401, n174);
buf  g856 (n868, n154);
buf  g857 (n619, n127);
buf  g858 (n682, n156);
not  g859 (n739, n137);
not  g860 (n453, n131);
buf  g861 (n392, n152);
not  g862 (n349, n88);
not  g863 (n468, n137);
buf  g864 (n436, n110);
not  g865 (n714, n211);
buf  g866 (n363, n58);
not  g867 (n272, n53);
buf  g868 (n683, n185);
buf  g869 (n767, n157);
not  g870 (n413, n124);
not  g871 (n850, n153);
not  g872 (n771, n133);
buf  g873 (n494, n211);
not  g874 (n515, n96);
not  g875 (n262, n196);
buf  g876 (n304, n218);
buf  g877 (n528, n211);
not  g878 (n339, n95);
buf  g879 (n278, n156);
xor  g880 (n931, n234, n238, n242, n221);
xnor g881 (n930, n252, n248, n249, n233);
xnor g882 (n936, n245, n234, n240, n228);
xnor g883 (n929, n227, n230, n241, n248);
nor  g884 (n938, n246, n251, n229, n244);
xor  g885 (n935, n246, n229, n231, n240);
nand g886 (n933, n232, n237, n247, n223);
and  g887 (n937, n236, n250, n252);
xnor g888 (n934, n239, n241, n245, n224);
nor  g889 (n939, n228, n236, n226, n235);
and  g890 (n940, n242, n233, n226, n247);
and  g891 (n932, n249, n243, n224, n238);
xnor g892 (n928, n243, n223, n221, n231);
and  g893 (n925, n230, n244, n222);
and  g894 (n926, n237, n225, n232, n227);
nor  g895 (n927, n235, n239, n251, n225);
not  g896 (n941, n939);
buf  g897 (n942, n940);
buf  g898 (n943, n942);
buf  g899 (n944, n942);
not  g900 (n945, n942);
not  g901 (n947, n942);
not  g902 (n950, n941);
not  g903 (n948, n941);
buf  g904 (n946, n941);
not  g905 (n949, n941);
not  g906 (n954, n944);
not  g907 (n953, n943);
buf  g908 (n955, n943);
buf  g909 (n951, n943);
not  g910 (n952, n943);
nor  g911 (n957, n944, n955, n945, n954);
nor  g912 (n956, n256, n256, n955, n255);
xnor g913 (n963, n947, n945, n953);
or   g914 (n958, n257, n945, n954, n952);
and  g915 (n959, n254, n254, n944, n952);
nor  g916 (n960, n253, n255, n944, n946);
or   g917 (n961, n953, n951, n946, n253);
nor  g918 (n962, n257, n946, n951);
not  g919 (n968, n961);
buf  g920 (n973, n963);
buf  g921 (n971, n959);
buf  g922 (n967, n956);
not  g923 (n965, n958);
not  g924 (n970, n960);
buf  g925 (n966, n962);
buf  g926 (n969, n957);
not  g927 (n964, n962);
not  g928 (n972, n963);
xnor g929 (n979, n969, n264, n276, n291);
or   g930 (n977, n296, n273, n259, n279);
nand g931 (n982, n281, n293, n270, n966);
and  g932 (n989, n971, n288, n966, n264);
nand g933 (n978, n278, n296, n275, n277);
or   g934 (n994, n290, n276, n294, n277);
xor  g935 (n976, n267, n971, n283, n299);
and  g936 (n992, n287, n269, n289, n279);
nor  g937 (n983, n295, n268, n272, n266);
and  g938 (n988, n263, n964, n274, n265);
xnor g939 (n999, n299, n967, n965);
xor  g940 (n991, n968, n259, n290, n289);
nand g941 (n975, n292, n970, n273, n964);
or   g942 (n1003, n260, n285, n965, n291);
xor  g943 (n985, n293, n292, n297, n301);
or   g944 (n1000, n262, n258, n969, n298);
xnor g945 (n998, n280, n300, n287, n970);
xor  g946 (n1002, n261, n969, n284, n274);
xnor g947 (n984, n272, n280, n966, n269);
and  g948 (n990, n278, n268, n286, n263);
or   g949 (n980, n275, n266, n260, n285);
nor  g950 (n1001, n286, n282, n967);
xnor g951 (n986, n968, n294, n964, n261);
or   g952 (n974, n265, n965, n281, n283);
xor  g953 (n997, n302, n295, n301, n297);
nor  g954 (n987, n271, n298, n968, n288);
nand g955 (n995, n965, n300, n271, n969);
nor  g956 (n996, n282, n270, n970, n966);
or   g957 (n993, n284, n258, n262, n968);
or   g958 (n981, n302, n964, n267, n970);
not  g959 (n1014, n977);
buf  g960 (n1005, n975);
not  g961 (n1012, n974);
buf  g962 (n1007, n979);
not  g963 (n1013, n981);
not  g964 (n1008, n981);
buf  g965 (n1006, n978);
not  g966 (n1015, n976);
not  g967 (n1004, n976);
not  g968 (n1010, n978);
nand g969 (n1011, n974, n979);
and  g970 (n1009, n975, n980, n977);
not  g971 (n1024, n1004);
buf  g972 (n1021, n1005);
not  g973 (n1031, n1005);
buf  g974 (n1017, n1004);
not  g975 (n1030, n1007);
buf  g976 (n1023, n1005);
buf  g977 (n1019, n1007);
buf  g978 (n1022, n1006);
buf  g979 (n1016, n1006);
not  g980 (n1028, n1004);
buf  g981 (n1025, n1004);
buf  g982 (n1029, n1007);
not  g983 (n1020, n1005);
not  g984 (n1027, n1007);
not  g985 (n1026, n1006);
not  g986 (n1018, n1006);
buf  g987 (n1033, n1016);
not  g988 (n1032, n1016);
xnor g989 (n1040, n1032, n1017, n1033);
or   g990 (n1034, n1025, n1021, n304, n1020);
xnor g991 (n1035, n1022, n1017, n1024);
or   g992 (n1039, n1019, n303, n1018, n1023);
nor  g993 (n1036, n1026, n1032, n1033, n1023);
and  g994 (n1038, n1032, n1019, n1033, n947);
xnor g995 (n1041, n303, n1032, n1021, n1025);
and  g996 (n1037, n304, n1020, n1022, n1018);
not  g997 (n1050, n982);
not  g998 (n1043, n1040);
not  g999 (n1053, n305);
not  g1000 (n1047, n973);
not  g1001 (n1049, n1034);
not  g1002 (n1045, n1041);
not  g1003 (n1044, n972);
or   g1004 (n1042, n1037, n1040, n972);
and  g1005 (n1048, n1036, n1039, n971, n1038);
xnor g1006 (n1051, n982, n972, n983, n306);
nor  g1007 (n1052, n1038, n1041, n971, n305);
nor  g1008 (n1046, n973, n1039, n1035, n972);
not  g1009 (n1066, n1048);
buf  g1010 (n1074, n1051);
buf  g1011 (n1069, n1049);
buf  g1012 (n1060, n1047);
buf  g1013 (n1063, n1049);
not  g1014 (n1081, n1047);
buf  g1015 (n1070, n1050);
not  g1016 (n1078, n1045);
not  g1017 (n1073, n1044);
not  g1018 (n1064, n1043);
not  g1019 (n1079, n1044);
buf  g1020 (n1075, n1048);
not  g1021 (n1080, n1045);
not  g1022 (n1077, n1042);
not  g1023 (n1059, n1043);
buf  g1024 (n1067, n1044);
not  g1025 (n1056, n1046);
buf  g1026 (n1072, n1050);
not  g1027 (n1054, n1046);
not  g1028 (n1062, n1051);
buf  g1029 (n1068, n1042);
buf  g1030 (n1061, n1048);
not  g1031 (n1055, n1049);
buf  g1032 (n1065, n1045);
buf  g1033 (n1057, n1046);
buf  g1034 (n1071, n1047);
buf  g1035 (n1076, n1050);
buf  g1036 (n1058, n1043);
not  g1037 (n1137, n1057);
not  g1038 (n1149, n1064);
buf  g1039 (n1127, n1074);
buf  g1040 (n1131, n1075);
not  g1041 (n1155, n1009);
not  g1042 (n1083, n1014);
not  g1043 (n1100, n1013);
not  g1044 (n1090, n1000);
buf  g1045 (n1092, n1057);
not  g1046 (n1128, n1071);
not  g1047 (n1104, n1067);
not  g1048 (n1160, n1065);
not  g1049 (n1101, n987);
buf  g1050 (n1157, n1080);
not  g1051 (n1165, n1012);
buf  g1052 (n1088, n1064);
buf  g1053 (n1141, n1075);
buf  g1054 (n1097, n1013);
buf  g1055 (n1122, n1055);
buf  g1056 (n1188, n1009);
buf  g1057 (n1171, n1079);
buf  g1058 (n1173, n1071);
not  g1059 (n1093, n1061);
not  g1060 (n1091, n1081);
buf  g1061 (n1106, n990);
not  g1062 (n1145, n1012);
not  g1063 (n1151, n1063);
buf  g1064 (n1189, n1011);
not  g1065 (n1094, n1070);
buf  g1066 (n1182, n1014);
buf  g1067 (n1191, n985);
not  g1068 (n1169, n1077);
not  g1069 (n1115, n994);
buf  g1070 (n1193, n1069);
buf  g1071 (n1132, n1080);
not  g1072 (n1111, n1054);
buf  g1073 (n1146, n991);
buf  g1074 (n1087, n1008);
not  g1075 (n1129, n1072);
not  g1076 (n1139, n1002);
not  g1077 (n1161, n1060);
not  g1078 (n1109, n1081);
buf  g1079 (n1159, n1063);
not  g1080 (n1192, n1062);
not  g1081 (n1110, n1059);
not  g1082 (n1130, n1061);
buf  g1083 (n1095, n1081);
not  g1084 (n1086, n991);
not  g1085 (n1153, n1078);
buf  g1086 (n1140, n1070);
buf  g1087 (n1150, n1062);
not  g1088 (n1098, n1055);
buf  g1089 (n1120, n1002);
not  g1090 (n1183, n1073);
buf  g1091 (n1180, n1071);
not  g1092 (n1099, n1015);
buf  g1093 (n1158, n1070);
buf  g1094 (n1112, n1057);
not  g1095 (n1166, n1067);
buf  g1096 (n1142, n1080);
buf  g1097 (n1163, n1073);
not  g1098 (n1176, n1059);
not  g1099 (n1103, n992);
buf  g1100 (n1156, n1062);
not  g1101 (n1118, n1059);
buf  g1102 (n1134, n1068);
not  g1103 (n1108, n1076);
buf  g1104 (n1154, n1008);
buf  g1105 (n1167, n1011);
buf  g1106 (n1121, n997);
not  g1107 (n1187, n1011);
buf  g1108 (n1172, n1073);
buf  g1109 (n1102, n989);
buf  g1110 (n1190, n1054);
not  g1111 (n1175, n990);
buf  g1112 (n1136, n1079);
buf  g1113 (n1089, n987);
not  g1114 (n1105, n988);
not  g1115 (n1174, n996);
buf  g1116 (n1082, n985);
not  g1117 (n1135, n1061);
buf  g1118 (n1143, n1067);
buf  g1119 (n1152, n993);
buf  g1120 (n1186, n1081);
buf  g1121 (n1147, n1078);
not  g1122 (n1144, n1056);
buf  g1123 (n1107, n1068);
not  g1124 (n1117, n1058);
not  g1125 (n1133, n988);
or   g1126 (n1177, n1064, n1066, n1001, n1071);
nand g1127 (n1168, n1065, n995, n1010, n1068);
or   g1128 (n1162, n983, n1056, n1078);
xor  g1129 (n1126, n1054, n1069, n1070, n1075);
xor  g1130 (n1164, n1013, n1079, n1010, n1000);
nor  g1131 (n1185, n1079, n1060, n1015, n1058);
and  g1132 (n1123, n1066, n1074, n1065, n1063);
or   g1133 (n1124, n1008, n989, n992, n1056);
xnor g1134 (n1116, n1014, n995, n1009, n1069);
xnor g1135 (n1170, n1077, n1060, n1054, n1008);
nor  g1136 (n1096, n1072, n1065, n1080, n1009);
xor  g1137 (n1113, n1055, n1058);
nor  g1138 (n1138, n1061, n1010, n1059, n1011);
xor  g1139 (n1178, n1062, n984, n1063);
nand g1140 (n1148, n1074, n994, n1001, n1067);
xor  g1141 (n1114, n999, n1077, n1076, n998);
xnor g1142 (n1119, n999, n996, n1060, n1077);
xor  g1143 (n1084, n1074, n998, n1073, n986);
and  g1144 (n1125, n1076, n1075, n993, n1069);
xnor g1145 (n1179, n997, n1076, n1066, n1068);
xnor g1146 (n1184, n1072, n986, n1010, n1066);
xor  g1147 (n1085, n1012, n1014, n1056, n1064);
xor  g1148 (n1181, n1072, n1012, n1057, n1013);
xor  g1149 (n1208, n623, n559, n562, n658);
nor  g1150 (n1332, n1144, n351, n695, n347);
and  g1151 (n1444, n599, n650, n1098, n364);
xnor g1152 (n1634, n1088, n556, n377, n561);
and  g1153 (n1238, n535, n625, n611, n643);
xor  g1154 (n1350, n666, n1127, n1137, n550);
nor  g1155 (n1380, n440, n568, n550, n655);
nand g1156 (n1612, n527, n630, n1146, n679);
and  g1157 (n1475, n654, n680, n1103, n595);
nor  g1158 (n1225, n431, n1165, n691, n1126);
nand g1159 (n1462, n395, n649, n583, n481);
and  g1160 (n1284, n340, n564, n523, n463);
xor  g1161 (n1546, n713, n500, n346, n1145);
nor  g1162 (n1430, n1131, n501, n651, n641);
nand g1163 (n1469, n1170, n499, n629, n1147);
and  g1164 (n1236, n306, n509, n712, n611);
xnor g1165 (n1479, n360, n644, n598, n630);
nor  g1166 (n1484, n526, n1148, n380, n1121);
and  g1167 (n1261, n609, n666, n569, n659);
xor  g1168 (n1221, n1084, n651, n459, n566);
nor  g1169 (n1386, n1175, n486, n1120, n553);
and  g1170 (n1521, n522, n397, n578, n390);
xor  g1171 (n1579, n644, n724, n693, n530);
xnor g1172 (n1533, n361, n1126, n1125, n1110);
nor  g1173 (n1200, n430, n632, n667, n564);
nor  g1174 (n1424, n607, n425, n522, n400);
xor  g1175 (n1381, n369, n680, n665, n1107);
or   g1176 (n1554, n617, n1090, n623, n535);
xnor g1177 (n1576, n528, n545, n506, n422);
xnor g1178 (n1405, n578, n683, n625, n433);
nand g1179 (n1325, n525, n515, n617, n701);
xor  g1180 (n1348, n602, n649, n1111, n546);
nor  g1181 (n1594, n396, n1186, n1161, n1136);
xnor g1182 (n1529, n578, n718, n653, n668);
xnor g1183 (n1624, n1029, n693, n457, n1171);
and  g1184 (n1467, n1137, n728, n637, n594);
xor  g1185 (n1361, n684, n570, n1158, n647);
xor  g1186 (n1440, n498, n1105, n460, n1136);
xor  g1187 (n1548, n1102, n363, n461, n343);
and  g1188 (n1447, n373, n541, n1193, n596);
xor  g1189 (n1500, n514, n538, n1112, n661);
nand g1190 (n1247, n626, n1113, n1156, n609);
and  g1191 (n1297, n540, n540, n1094, n491);
or   g1192 (n1404, n669, n585, n561, n640);
xor  g1193 (n1436, n551, n1138, n335, n1127);
and  g1194 (n1491, n485, n326, n566, n1127);
and  g1195 (n1626, n647, n1127, n648, n589);
nor  g1196 (n1274, n579, n533, n430, n322);
nand g1197 (n1555, n1145, n308, n419, n646);
nand g1198 (n1618, n603, n344, n539, n1160);
xor  g1199 (n1566, n358, n362, n502, n313);
nor  g1200 (n1291, n451, n1192, n1181, n472);
and  g1201 (n1419, n530, n644, n513, n1093);
and  g1202 (n1453, n622, n705, n670, n460);
xor  g1203 (n1542, n723, n1161, n578, n1092);
nand g1204 (n1636, n1164, n434, n1097, n1136);
nand g1205 (n1613, n481, n1188, n478, n495);
nand g1206 (n1222, n1107, n1130, n449, n532);
xor  g1207 (n1329, n1135, n649, n714, n1097);
nand g1208 (n1226, n1128, n456, n703, n608);
and  g1209 (n1206, n1189, n610, n433, n728);
nor  g1210 (n1232, n615, n630, n649, n565);
nor  g1211 (n1316, n553, n499, n331, n597);
or   g1212 (n1330, n428, n720, n1139, n608);
nand g1213 (n1421, n711, n548, n1189, n628);
or   g1214 (n1408, n1028, n720, n678, n725);
xor  g1215 (n1627, n632, n379, n375, n691);
xnor g1216 (n1456, n1123, n432, n549, n658);
xnor g1217 (n1582, n531, n1135, n501, n539);
xnor g1218 (n1287, n626, n1086, n583, n554);
nand g1219 (n1270, n528, n1157, n557, n478);
nor  g1220 (n1610, n516, n1146, n595, n669);
xnor g1221 (n1459, n1135, n1119, n1124, n1095);
or   g1222 (n1292, n614, n662, n414, n1154);
or   g1223 (n1517, n1170, n650, n681, n359);
xor  g1224 (n1464, n314, n708, n704, n657);
xnor g1225 (n1488, n1087, n319, n489, n628);
xnor g1226 (n1277, n1104, n1028, n1107, n508);
xnor g1227 (n1558, n418, n1156, n387, n495);
nor  g1228 (n1543, n1083, n556, n409, n507);
xor  g1229 (n1617, n549, n612, n1144, n575);
nand g1230 (n1468, n431, n1184, n654, n546);
nor  g1231 (n1472, n463, n661, n682, n459);
nand g1232 (n1333, n1185, n576, n1118, n1188);
or   g1233 (n1429, n332, n593, n1096, n629);
or   g1234 (n1389, n311, n675, n1156, n1153);
and  g1235 (n1514, n524, n612, n688, n510);
xor  g1236 (n1253, n568, n707, n685, n598);
or   g1237 (n1375, n718, n601, n1093, n1182);
nand g1238 (n1229, n648, n542, n646, n602);
xnor g1239 (n1283, n613, n450, n1187, n597);
or   g1240 (n1512, n1093, n468, n504, n469);
and  g1241 (n1476, n446, n385, n389, n1097);
nor  g1242 (n1262, n355, n636, n639, n562);
xor  g1243 (n1390, n1122, n692, n404, n1094);
xnor g1244 (n1377, n422, n452, n516, n1193);
nor  g1245 (n1527, n582, n333, n585, n711);
or   g1246 (n1557, n1120, n717, n328, n329);
xnor g1247 (n1489, n1145, n1144, n1142, n693);
xor  g1248 (n1511, n650, n1177, n654, n560);
or   g1249 (n1591, n1182, n310, n1151, n706);
nor  g1250 (n1535, n594, n1114, n1176, n715);
xnor g1251 (n1526, n1154, n523, n1166, n1191);
or   g1252 (n1347, n697, n712, n620, n595);
nor  g1253 (n1311, n547, n572, n670, n592);
nor  g1254 (n1205, n1176, n331, n574, n666);
xnor g1255 (n1321, n1118, n494, n624, n1115);
nand g1256 (n1379, n642, n502, n584, n456);
or   g1257 (n1231, n577, n1193, n621, n309);
nand g1258 (n1368, n1129, n585, n1112, n634);
and  g1259 (n1528, n1150, n1087, n637, n669);
xor  g1260 (n1412, n542, n546, n462, n379);
nor  g1261 (n1267, n671, n337, n548, n1162);
nor  g1262 (n1493, n443, n634, n1099, n703);
or   g1263 (n1196, n349, n448, n635, n442);
xnor g1264 (n1595, n1158, n487, n634, n382);
nand g1265 (n1217, n687, n1152, n371, n537);
and  g1266 (n1400, n558, n1110, n607, n727);
xor  g1267 (n1230, n412, n1125, n1112, n686);
nor  g1268 (n1631, n370, n678, n416, n708);
or   g1269 (n1531, n1083, n535, n582, n673);
nand g1270 (n1248, n1083, n333, n678, n1161);
xor  g1271 (n1490, n381, n1169, n643, n633);
or   g1272 (n1289, n397, n643, n616, n324);
and  g1273 (n1417, n1166, n694, n708, n1147);
or   g1274 (n1411, n590, n481, n683, n1102);
xnor g1275 (n1515, n615, n374, n707, n599);
nand g1276 (n1346, n548, n700, n668, n437);
xor  g1277 (n1265, n627, n493, n581, n694);
xor  g1278 (n1483, n536, n670, n659, n671);
nand g1279 (n1194, n525, n698, n590, n699);
nand g1280 (n1499, n1193, n678, n606, n629);
nand g1281 (n1420, n512, n601, n500, n544);
or   g1282 (n1240, n658, n1139, n1118, n312);
nor  g1283 (n1498, n365, n1108, n1164, n372);
nand g1284 (n1207, n497, n621, n1088, n567);
xnor g1285 (n1621, n538, n1168, n1092, n1091);
nand g1286 (n1245, n698, n1099, n639, n577);
and  g1287 (n1536, n502, n1103, n1152, n482);
xnor g1288 (n1427, n420, n1148, n606, n1104);
xor  g1289 (n1562, n1138, n472, n684, n378);
nor  g1290 (n1314, n672, n386, n700, n532);
xnor g1291 (n1278, n512, n1116, n718, n1155);
nand g1292 (n1598, n539, n1106, n339, n1087);
or   g1293 (n1426, n1188, n1185, n517, n1174);
nand g1294 (n1423, n1166, n1181, n1105, n690);
xnor g1295 (n1622, n487, n522, n620, n605);
xnor g1296 (n1435, n1121, n468, n1140, n656);
nor  g1297 (n1252, n537, n450, n497, n611);
and  g1298 (n1446, n1095, n528, n447, n497);
or   g1299 (n1606, n376, n435, n617, n458);
or   g1300 (n1506, n519, n645, n565, n1149);
and  g1301 (n1603, n587, n675, n464, n677);
xor  g1302 (n1549, n520, n417, n601, n663);
nor  g1303 (n1522, n567, n471, n661, n625);
nand g1304 (n1286, n361, n514, n1176, n348);
or   g1305 (n1471, n496, n1156, n582, n1119);
nand g1306 (n1224, n554, n1134, n367, n513);
nor  g1307 (n1353, n723, n413, n475, n653);
or   g1308 (n1369, n525, n1147, n715, n543);
nand g1309 (n1215, n662, n320, n574, n1175);
xor  g1310 (n1586, n1117, n543, n527, n493);
and  g1311 (n1313, n664, n338, n1139, n618);
nor  g1312 (n1349, n1092, n624, n708, n628);
or   g1313 (n1384, n480, n571, n636, n517);
or   g1314 (n1524, n1133, n489, n408, n351);
and  g1315 (n1233, n470, n695, n551, n1176);
xor  g1316 (n1373, n455, n321, n439, n383);
or   g1317 (n1338, n1189, n1110, n660, n694);
or   g1318 (n1520, n659, n727, n1126, n512);
xor  g1319 (n1320, n1094, n545, n1027, n642);
xnor g1320 (n1538, n1171, n686, n1147, n634);
xor  g1321 (n1395, n381, n660, n631, n715);
xnor g1322 (n1388, n488, n1115, n1146, n591);
and  g1323 (n1319, n663, n562, n537, n608);
nor  g1324 (n1448, n490, n707, n1167, n545);
and  g1325 (n1441, n321, n524, n562, n1186);
and  g1326 (n1590, n716, n676, n1160, n508);
or   g1327 (n1281, n596, n668, n1151, n676);
nand g1328 (n1303, n590, n1101, n1186, n551);
or   g1329 (n1326, n1086, n511, n1164, n690);
and  g1330 (n1492, n656, n587, n689, n444);
nor  g1331 (n1523, n552, n507, n633, n581);
or   g1332 (n1630, n688, n507, n445, n665);
and  g1333 (n1615, n584, n490, n696, n511);
and  g1334 (n1415, n549, n580, n1150, n457);
and  g1335 (n1561, n1129, n710, n1132);
and  g1336 (n1628, n1152, n1181, n438, n1099);
nand g1337 (n1596, n705, n336, n672, n491);
and  g1338 (n1366, n664, n543, n636, n363);
and  g1339 (n1431, n489, n684, n488, n1188);
nand g1340 (n1308, n559, n1151, n538, n467);
or   g1341 (n1547, n610, n1155, n1111, n1150);
nor  g1342 (n1530, n346, n1085, n546, n652);
or   g1343 (n1478, n645, n327, n657, n650);
or   g1344 (n1604, n1148, n670, n622, n602);
xor  g1345 (n1541, n721, n311, n685, n336);
nor  g1346 (n1195, n1029, n620, n492, n721);
nor  g1347 (n1363, n335, n1168, n576, n721);
nand g1348 (n1495, n687, n635, n591, n555);
xnor g1349 (n1199, n709, n1166, n443, n1182);
xor  g1350 (n1241, n647, n366, n499, n722);
nand g1351 (n1213, n633, n657, n1179, n526);
and  g1352 (n1422, n607, n343, n1133, n1112);
nor  g1353 (n1633, n521, n682, n719, n1142);
xor  g1354 (n1409, n1113, n699, n519, n1135);
or   g1355 (n1559, n681, n1160, n386, n675);
nand g1356 (n1306, n1180, n552, n555, n611);
xnor g1357 (n1445, n680, n586, n515, n1128);
nor  g1358 (n1545, n613, n501, n410, n1123);
nor  g1359 (n1519, n544, n1100, n683, n1111);
nand g1360 (n1357, n1159, n1091, n681, n1101);
and  g1361 (n1391, n503, n691, n606, n444);
or   g1362 (n1300, n572, n702, n1187, n696);
and  g1363 (n1525, n503, n341, n408, n620);
nor  g1364 (n1382, n672, n440, n325, n517);
and  g1365 (n1556, n585, n712, n403, n679);
and  g1366 (n1301, n446, n558, n429, n509);
and  g1367 (n1428, n1113, n552, n563, n1178);
xor  g1368 (n1312, n517, n1149, n726, n382);
or   g1369 (n1480, n536, n502, n587, n692);
or   g1370 (n1372, n498, n454, n631, n485);
nor  g1371 (n1370, n576, n557, n1192, n483);
nor  g1372 (n1583, n603, n1109, n375, n395);
xnor g1373 (n1605, n622, n514, n577, n509);
nor  g1374 (n1564, n594, n1172, n388, n610);
or   g1375 (n1454, n477, n436, n358, n313);
nand g1376 (n1601, n579, n534, n591, n326);
or   g1377 (n1451, n676, n725, n698, n1171);
xnor g1378 (n1282, n1164, n1116, n550, n1083);
nand g1379 (n1563, n526, n1142, n461, n690);
and  g1380 (n1259, n709, n1132, n642, n1109);
and  g1381 (n1641, n523, n667, n532, n322);
xnor g1382 (n1629, n614, n614, n674, n667);
xor  g1383 (n1219, n618, n398, n586, n1134);
and  g1384 (n1458, n1179, n713, n516, n501);
and  g1385 (n1510, n1178, n701, n407, n706);
xor  g1386 (n1578, n1084, n494, n1175, n448);
xor  g1387 (n1584, n309, n402, n657, n694);
or   g1388 (n1355, n1162, n581, n631, n522);
nand g1389 (n1279, n718, n402, n492, n627);
nor  g1390 (n1269, n1143, n334, n1162, n655);
nor  g1391 (n1602, n589, n647, n1030, n1089);
nand g1392 (n1587, n1133, n1173, n415, n424);
nor  g1393 (n1474, n480, n1169, n420, n510);
nand g1394 (n1477, n315, n453, n687, n1096);
and  g1395 (n1570, n324, n719, n619, n1089);
xnor g1396 (n1345, n1133, n307, n672, n717);
xor  g1397 (n1296, n371, n413, n563, n504);
nand g1398 (n1638, n1128, n583, n593, n529);
or   g1399 (n1619, n508, n474, n1098, n436);
or   g1400 (n1371, n704, n556, n1104, n690);
or   g1401 (n1273, n721, n390, n1138, n704);
nand g1402 (n1227, n1109, n612, n720, n609);
xor  g1403 (n1496, n569, n1121, n689, n638);
xor  g1404 (n1608, n445, n725, n1161, n1090);
nand g1405 (n1437, n664, n1191, n593, n588);
xor  g1406 (n1365, n505, n584, n354, n600);
or   g1407 (n1509, n477, n345, n1184, n421);
nand g1408 (n1214, n539, n705, n1168, n1167);
xnor g1409 (n1336, n411, n486, n582, n641);
xnor g1410 (n1565, n553, n682, n545, n631);
nor  g1411 (n1254, n709, n356, n704, n1170);
and  g1412 (n1414, n1167, n1138, n1122, n464);
and  g1413 (n1569, n1130, n352, n1108, n667);
or   g1414 (n1290, n1117, n619, n573, n604);
and  g1415 (n1276, n615, n1125, n503, n1178);
xor  g1416 (n1212, n373, n1100, n626, n1114);
nor  g1417 (n1518, n701, n426, n573, n466);
xor  g1418 (n1625, n613, n727, n549, n1157);
nand g1419 (n1211, n716, n1154, n1172, n434);
nand g1420 (n1374, n427, n1084, n1131, n1141);
or   g1421 (n1487, n469, n1091, n572, n646);
nor  g1422 (n1637, n599, n567, n536, n534);
or   g1423 (n1255, n394, n671, n540, n640);
nand g1424 (n1577, n607, n1177, n1149, n637);
nand g1425 (n1600, n625, n1085, n1084, n604);
or   g1426 (n1358, n534, n1184, n697, n633);
or   g1427 (n1399, n570, n362, n554, n1096);
xnor g1428 (n1235, n1105, n571, n1140, n640);
or   g1429 (n1457, n1082, n465, n368, n345);
or   g1430 (n1216, n406, n554, n673, n1174);
xnor g1431 (n1402, n1178, n711, n325, n447);
or   g1432 (n1367, n567, n317, n418, n1173);
and  g1433 (n1532, n1159, n584, n617, n1165);
nor  g1434 (n1589, n1165, n1170, n483, n510);
nor  g1435 (n1251, n334, n474, n494, n528);
nor  g1436 (n1508, n383, n316, n406, n1026);
xor  g1437 (n1202, n471, n662, n559, n616);
or   g1438 (n1197, n656, n466, n1155, n693);
or   g1439 (n1328, n425, n1141, n477, n1110);
xor  g1440 (n1237, n389, n479, n511, n421);
nand g1441 (n1317, n1180, n640, n509, n661);
xor  g1442 (n1359, n409, n599, n600, n656);
or   g1443 (n1432, n726, n566, n594, n475);
nand g1444 (n1434, n400, n1113, n329, n533);
or   g1445 (n1271, n665, n544, n641, n592);
xor  g1446 (n1580, n699, n1130, n695, n330);
xor  g1447 (n1539, n495, n1099, n586, n1119);
nand g1448 (n1481, n618, n652, n1151, n467);
and  g1449 (n1442, n1163, n458, n561, n685);
and  g1450 (n1323, n439, n591, n1082, n513);
nor  g1451 (n1360, n1140, n714, n1190, n531);
xor  g1452 (n1204, n676, n662, n529, n665);
nor  g1453 (n1397, n1173, n350, n518, n574);
xnor g1454 (n1593, n1145, n357, n1162, n511);
nand g1455 (n1620, n679, n1125, n604, n1180);
xor  g1456 (n1244, n596, n392, n573, n1184);
xnor g1457 (n1356, n560, n490, n530, n519);
nor  g1458 (n1243, n1089, n388, n580, n710);
xnor g1459 (n1567, n1153, n1093, n342, n512);
xor  g1460 (n1198, n684, n586, n653, n349);
nand g1461 (n1537, n479, n454, n1132, n608);
nor  g1462 (n1310, n486, n638, n484, n658);
xnor g1463 (n1607, n698, n1154, n527, n555);
nand g1464 (n1383, n416, n385, n515, n376);
nor  g1465 (n1497, n380, n600, n1155, n559);
and  g1466 (n1568, n573, n534, n1168, n487);
nand g1467 (n1257, n1192, n1163, n344, n587);
xor  g1468 (n1352, n523, n547, n677, n597);
nand g1469 (n1343, n1124, n374, n671, n1118);
and  g1470 (n1376, n540, n1153, n1097, n1148);
xnor g1471 (n1413, n711, n482, n551, n544);
nand g1472 (n1407, n580, n724, n553, n1136);
nand g1473 (n1473, n568, n556, n535, n1115);
nand g1474 (n1299, n340, n1122, n465, n537);
xor  g1475 (n1507, n496, n500, n410, n1124);
or   g1476 (n1298, n407, n569, n1183, n638);
xnor g1477 (n1307, n506, n705, n548, n651);
and  g1478 (n1588, n393, n1190, n716, n515);
and  g1479 (n1334, n428, n393, n1114, n347);
xor  g1480 (n1632, n1092, n1117, n720, n710);
xor  g1481 (n1396, n726, n531, n571, n1165);
and  g1482 (n1295, n629, n520, n637);
xor  g1483 (n1246, n613, n435, n1174, n526);
nor  g1484 (n1394, n600, n1134, n714, n396);
and  g1485 (n1450, n557, n417, n318, n635);
xnor g1486 (n1344, n1132, n476, n563, n498);
nand g1487 (n1364, n521, n415, n643, n648);
nand g1488 (n1597, n1121, n482, n1126, n673);
and  g1489 (n1266, n655, n1185, n1103, n713);
nand g1490 (n1339, n571, n508, n635, n524);
nor  g1491 (n1540, n404, n438, n521, n1116);
and  g1492 (n1410, n639, n697, n538, n610);
xor  g1493 (n1228, n1183, n378, n589, n1139);
nand g1494 (n1463, n1100, n619, n558, n702);
nor  g1495 (n1392, n1158, n1158, n1111, n574);
xor  g1496 (n1482, n518, n580, n646, n1119);
and  g1497 (n1293, n621, n1171, n498, n579);
or   g1498 (n1550, n419, n352, n1169, n570);
or   g1499 (n1571, n504, n348, n583, n1146);
and  g1500 (n1501, n682, n424, n604, n1157);
nand g1501 (n1264, n616, n499, n1088, n484);
or   g1502 (n1572, n308, n441, n663, n1090);
or   g1503 (n1616, n1108, n581, n598, n330);
or   g1504 (n1249, n683, n618, n727, n368);
xnor g1505 (n1552, n492, n664, n725, n480);
or   g1506 (n1513, n372, n685, n728, n561);
nand g1507 (n1354, n449, n1186, n606, n714);
xnor g1508 (n1260, n575, n1150, n1187, n654);
xor  g1509 (n1401, n565, n1177, n332, n1128);
xnor g1510 (n1439, n645, n689, n1143, n391);
xnor g1511 (n1342, n626, n615, n1142, n1143);
nand g1512 (n1560, n707, n513, n505, n1180);
xnor g1513 (n1331, n687, n1096, n1137, n524);
and  g1514 (n1351, n455, n1100, n644, n1116);
xnor g1515 (n1574, n1088, n1115, n518, n492);
nor  g1516 (n1592, n1190, n652, n603, n1173);
xor  g1517 (n1609, n666, n706, n1105, n529);
xnor g1518 (n1418, n597, n1149, n642, n541);
xor  g1519 (n1575, n310, n350, n564, n1114);
nand g1520 (n1272, n639, n560, n1191, n645);
xnor g1521 (n1452, n1102, n442, n488, n1106);
xor  g1522 (n1250, n1174, n636, n365, n533);
xnor g1523 (n1438, n485, n1122, n588, n314);
xnor g1524 (n1614, n369, n1082, n394, n353);
or   g1525 (n1466, n595, n367, n414, n312);
nor  g1526 (n1470, n723, n441, n478, n495);
xor  g1527 (n1335, n401, n1157, n1141, n652);
xor  g1528 (n1210, n719, n339, n697, n575);
xnor g1529 (n1551, n1185, n592, n1160, n1123);
and  g1530 (n1611, n623, n1085, n1130, n423);
or   g1531 (n1461, n622, n1027, n398, n1102);
or   g1532 (n1635, n483, n510, n653, n337);
and  g1533 (n1416, n533, n627, n560, n412);
xnor g1534 (n1239, n593, n342, n525, n1085);
nor  g1535 (n1503, n521, n496, n552, n1169);
nor  g1536 (n1218, n716, n547, n550, n723);
nor  g1537 (n1494, n423, n1134, n568, n590);
nand g1538 (n1465, n1190, n527, n619, n703);
or   g1539 (n1516, n366, n1098, n359, n505);
xor  g1540 (n1425, n479, n702, n491, n1087);
nor  g1541 (n1443, n387, n1103, n630, n1095);
xnor g1542 (n1304, n692, n576, n518, n566);
nor  g1543 (n1387, n403, n1129, n1090, n713);
or   g1544 (n1581, n692, n437, n726, n391);
nor  g1545 (n1340, n1179, n592, n1120, n405);
xnor g1546 (n1378, n1089, n328, n689, n695);
or   g1547 (n1327, n712, n541, n605, n1153);
xor  g1548 (n1209, n1094, n605, n532, n589);
nor  g1549 (n1302, n506, n1191, n557, n686);
xor  g1550 (n1398, n520, n1120, n1124, n703);
xor  g1551 (n1486, n1106, n688, n494, n1131);
nor  g1552 (n1406, n453, n717, n628, n1091);
or   g1553 (n1294, n505, n1144, n1181, n728);
and  g1554 (n1201, n1107, n491, n506, n1143);
or   g1555 (n1220, n1163, n696, n621, n677);
or   g1556 (n1502, n401, n356, n1172, n354);
nor  g1557 (n1449, n588, n570, n451, n688);
and  g1558 (n1256, n316, n519, n360, n674);
xnor g1559 (n1623, n632, n427, n1189, n1129);
or   g1560 (n1460, n616, n319, n719, n648);
and  g1561 (n1318, n529, n315, n691, n680);
nand g1562 (n1385, n699, n473, n558, n470);
and  g1563 (n1258, n677, n432, n596, n497);
or   g1564 (n1341, n575, n323, n669, n1029);
xnor g1565 (n1504, n476, n1123, n357, n1152);
nand g1566 (n1639, n577, n320, n627, n473);
xor  g1567 (n1485, n555, n601, n681, n503);
nand g1568 (n1403, n514, n641, n569, n452);
or   g1569 (n1534, n338, n709, n1141, n1179);
or   g1570 (n1275, n724, n572, n659, n399);
nor  g1571 (n1640, n624, n493, n1108, n663);
nor  g1572 (n1599, n1137, n588, n500, n1117);
nand g1573 (n1242, n605, n1101, n722, n531);
nor  g1574 (n1505, n660, n701, n1086, n632);
nand g1575 (n1288, n541, n1182, n1175, n565);
xnor g1576 (n1573, n651, n1159, n579, n1095);
nand g1577 (n1305, n1106, n542, n327, n496);
or   g1578 (n1544, n547, n543, n706, n493);
xnor g1579 (n1234, n724, n462, n1177, n624);
xor  g1580 (n1322, n411, n323, n1183, n384);
xor  g1581 (n1585, n614, n1140, n700, n673);
nand g1582 (n1280, n399, n700, n353, n696);
or   g1583 (n1263, n1101, n668, n484, n536);
xnor g1584 (n1268, n426, n660, n318, n702);
xor  g1585 (n1285, n686, n1104, n307, n504);
and  g1586 (n1553, n405, n598, n1172, n1192);
nand g1587 (n1315, n722, n655, n1183, n715);
and  g1588 (n1324, n364, n722, n623, n1082);
xor  g1589 (n1337, n564, n674, n638, n355);
or   g1590 (n1362, n612, n384, n317, n530);
xnor g1591 (n1203, n675, n1163, n1187, n1109);
xnor g1592 (n1223, n341, n679, n429, n563);
or   g1593 (n1309, n1098, n1131, n602, n1159);
nor  g1594 (n1433, n674, n516, n370, n609);
nand g1595 (n1393, n603, n1086, n717, n542);
or   g1596 (n1455, n507, n1167, n392, n377);
xnor g1597 (n1642, n729, n1194);
nor  g1598 (n1644, n729, n730);
nor  g1599 (n1643, n729, n1642);
not  g1600 (n1647, n1644);
buf  g1601 (n1650, n730);
buf  g1602 (n1649, n1643);
not  g1603 (n1651, n1644);
buf  g1604 (n1648, n1643);
buf  g1605 (n1646, n1643);
xor  g1606 (n1645, n1643, n1644);
not  g1607 (n1663, n731);
buf  g1608 (n1664, n1648);
not  g1609 (n1660, n736);
buf  g1610 (n1661, n738);
and  g1611 (n1656, n734, n1649, n733, n737);
xnor g1612 (n1657, n737, n732, n1647);
or   g1613 (n1652, n734, n737, n1649, n1646);
or   g1614 (n1662, n736, n738, n733, n1646);
xor  g1615 (n1654, n734, n1648, n735, n1650);
xnor g1616 (n1658, n1651, n735, n1650, n737);
nor  g1617 (n1659, n736, n1647, n732, n1645);
xnor g1618 (n1655, n733, n731, n1645, n735);
or   g1619 (n1665, n735, n731, n1651);
and  g1620 (n1653, n736, n732, n734, n733);
buf  g1621 (n1705, n738);
buf  g1622 (n1706, n1662);
not  g1623 (n1695, n1656);
buf  g1624 (n1668, n1660);
buf  g1625 (n1708, n1661);
not  g1626 (n1670, n1664);
buf  g1627 (n1678, n950);
buf  g1628 (n1674, n1661);
not  g1629 (n1721, n1655);
buf  g1630 (n1713, n948);
buf  g1631 (n1675, n1661);
not  g1632 (n1707, n949);
buf  g1633 (n1666, n1662);
buf  g1634 (n1690, n1659);
buf  g1635 (n1683, n1665);
buf  g1636 (n1704, n949);
buf  g1637 (n1720, n1652);
buf  g1638 (n1710, n1657);
not  g1639 (n1703, n1663);
not  g1640 (n1679, n1657);
not  g1641 (n1684, n950);
not  g1642 (n1716, n1664);
buf  g1643 (n1715, n1662);
not  g1644 (n1688, n1663);
not  g1645 (n1687, n1658);
not  g1646 (n1702, n1654);
buf  g1647 (n1700, n1659);
buf  g1648 (n1681, n1665);
buf  g1649 (n1669, n1657);
buf  g1650 (n1712, n1656);
buf  g1651 (n1671, n1660);
not  g1652 (n1667, n1659);
buf  g1653 (n1699, n740);
not  g1654 (n1718, n1655);
not  g1655 (n1697, n739);
buf  g1656 (n1709, n1664);
nor  g1657 (n1701, n1658, n740);
or   g1658 (n1676, n1663, n1654);
and  g1659 (n1677, n948, n1655);
nor  g1660 (n1689, n1665, n1654);
nand g1661 (n1680, n1658, n1655);
xor  g1662 (n1694, n1665, n1658);
or   g1663 (n1719, n1661, n947);
nand g1664 (n1698, n1657, n1652);
and  g1665 (n1711, n948, n1653);
xor  g1666 (n1692, n947, n1659);
nand g1667 (n1691, n739, n1656);
xor  g1668 (n1714, n948, n1654);
nand g1669 (n1693, n1656, n949);
nor  g1670 (n1686, n1664, n739);
and  g1671 (n1673, n738, n1660);
and  g1672 (n1682, n949, n1660);
buf  g1673 (n1672, n1653);
and  g1674 (n1717, n1652, n1662);
and  g1675 (n1696, n739, n1653);
xnor g1676 (n1685, n1652, n1663);
xor  g1677 (n1869, n1505, n1353, n1430, n1370);
or   g1678 (n1824, n1467, n1703, n1678, n1477);
xnor g1679 (n1755, n1461, n1448, n1293, n1236);
xor  g1680 (n1866, n1711, n1315, n1460, n1701);
xor  g1681 (n1884, n1371, n1200, n1670, n1674);
xnor g1682 (n1756, n1253, n1683, n1213, n1313);
and  g1683 (n1753, n1226, n1451, n1294, n1385);
and  g1684 (n1877, n1346, n1690, n1519, n1286);
and  g1685 (n1848, n1458, n1716, n1366, n1692);
nand g1686 (n1921, n1247, n1686, n1237, n1254);
xor  g1687 (n1777, n1506, n1429, n1680, n1426);
or   g1688 (n1727, n1509, n1515, n1490, n1326);
or   g1689 (n1782, n1271, n1523, n1485);
xnor g1690 (n1734, n1470, n1217, n1503, n1348);
nand g1691 (n1752, n1239, n1702, n1697, n1400);
xor  g1692 (n1807, n1333, n1517, n1298, n1205);
and  g1693 (n1793, n1673, n1198, n1700, n1669);
nor  g1694 (n1934, n1404, n1295, n1264, n1402);
and  g1695 (n1754, n1203, n1479, n1687, n1484);
nor  g1696 (n1938, n1272, n1335, n1443, n1332);
xnor g1697 (n1894, n1718, n1256, n1462, n1678);
nand g1698 (n1862, n1691, n1447, n1411, n1522);
nand g1699 (n1937, n1299, n1680, n1387, n1310);
nand g1700 (n1745, n1427, n1475, n1412, n1311);
xnor g1701 (n1853, n1423, n1481, n1671, n1716);
nor  g1702 (n1916, n1255, n1710, n1712, n1407);
nor  g1703 (n1943, n1418, n1291, n1357, n1227);
or   g1704 (n1933, n1344, n1715, n1201, n1666);
or   g1705 (n1942, n1452, n1509, n1683, n1669);
nand g1706 (n1809, n1472, n1365, n1478, n1720);
nand g1707 (n1749, n1273, n1238, n1359, n1484);
xnor g1708 (n1819, n1339, n1717, n1489, n1214);
or   g1709 (n1922, n1525, n1197, n1711, n1440);
xor  g1710 (n1902, n1324, n1392, n1415, n1224);
or   g1711 (n1863, n1402, n1249, n1666, n1520);
xnor g1712 (n1735, n1499, n1326, n1691, n1377);
and  g1713 (n1914, n1690, n1711, n1353, n1677);
xor  g1714 (n1924, n1414, n1694, n1222, n1667);
or   g1715 (n1932, n1398, n1268, n1475, n1306);
xnor g1716 (n1931, n1498, n1380, n1696, n1464);
xnor g1717 (n1817, n1403, n1410, n1279, n1708);
xor  g1718 (n1743, n1284, n1204, n1711, n1699);
xor  g1719 (n1887, n1294, n1252, n1208, n1695);
xnor g1720 (n1876, n1396, n1720, n1684, n1457);
nand g1721 (n1904, n1677, n1310, n1527, n1218);
nor  g1722 (n1882, n1221, n1308, n1705, n1693);
xor  g1723 (n1733, n1416, n1707, n1283, n1299);
or   g1724 (n1805, n1325, n1261, n1508, n1300);
nor  g1725 (n1913, n1694, n1721, n1376, n1290);
nand g1726 (n1917, n1258, n1674, n1447, n1325);
or   g1727 (n1796, n1221, n1675, n1211, n1695);
or   g1728 (n1927, n1235, n1454, n1522, n1521);
xnor g1729 (n1845, n1213, n1321, n1492, n1231);
nand g1730 (n1764, n1705, n1700, n1514, n1273);
nand g1731 (n1738, n1673, n1363, n1362, n1230);
nand g1732 (n1801, n1250, n1513, n1501, n1383);
or   g1733 (n1945, n1199, n1276, n1708, n1435);
nand g1734 (n1784, n1317, n1358, n1223, n1301);
xnor g1735 (n1732, n1335, n1681, n1458, n1246);
or   g1736 (n1830, n1361, n1279, n1338, n1263);
nor  g1737 (n1873, n1671, n1518, n1322, n1684);
nor  g1738 (n1911, n1449, n1212, n1375, n1333);
nor  g1739 (n1790, n1319, n1237, n1376, n1682);
and  g1740 (n1729, n1697, n1667, n1291, n1719);
xnor g1741 (n1818, n1685, n1349, n1476, n1448);
xnor g1742 (n1840, n1429, n1394, n1362, n1316);
nor  g1743 (n1905, n1503, n1679, n1491, n1410);
or   g1744 (n1821, n1331, n1255, n1283, n1232);
or   g1745 (n1891, n1675, n1220, n1420, n1365);
and  g1746 (n1815, n1378, n1479, n1707, n1675);
nor  g1747 (n1847, n1334, n1343, n1232, n1488);
and  g1748 (n1772, n1701, n1305, n1312, n1244);
xnor g1749 (n1747, n1405, n1721, n1323, n1417);
or   g1750 (n1926, n1713, n1369, n1425, n1201);
nor  g1751 (n1810, n1225, n1524, n1323, n1709);
xnor g1752 (n1901, n1674, n1408, n1340, n1409);
nand g1753 (n1737, n1216, n1496, n1408, n1694);
nor  g1754 (n1800, n1680, n1462, n1206, n1241);
nand g1755 (n1778, n1205, n1337, n1468, n1307);
or   g1756 (n1892, n1530, n1682, n1498, n1710);
and  g1757 (n1920, n1501, n1206, n1330, n1267);
xor  g1758 (n1751, n1262, n1349, n1413, n1712);
xor  g1759 (n1872, n1710, n1435, n1293, n1217);
nand g1760 (n1896, n1225, n1202, n1395, n1425);
nor  g1761 (n1730, n1352, n1691, n1233, n1274);
nand g1762 (n1803, n1668, n1342, n1382, n1302);
or   g1763 (n1785, n1690, n1396, n1679, n1714);
xnor g1764 (n1919, n1504, n1336, n1392, n1407);
or   g1765 (n1762, n1451, n1719, n1687, n1266);
xnor g1766 (n1893, n1687, n1383, n1247, n1228);
nand g1767 (n1774, n1494, n1379, n1249, n1469);
nand g1768 (n1795, n1271, n1346, n1388, n1463);
xor  g1769 (n1910, n1420, n1292, n1252, n1257);
xor  g1770 (n1741, n1482, n1713, n1441, n1275);
nand g1771 (n1832, n1384, n1197, n1678, n1214);
xor  g1772 (n1844, n1690, n1318, n1263, n1708);
nand g1773 (n1890, n1430, n1385, n1389, n1443);
xor  g1774 (n1728, n1477, n1324, n1703, n1391);
nor  g1775 (n1874, n1715, n1320, n1210, n1282);
nand g1776 (n1804, n1703, n1287, n1675, n1270);
or   g1777 (n1771, n1388, n1697, n1288, n1670);
xnor g1778 (n1744, n1504, n1269, n1245, n1207);
or   g1779 (n1767, n1523, n1281, n1461, n1386);
xnor g1780 (n1842, n1517, n1219, n1666, n1489);
or   g1781 (n1806, n1234, n1195, n1478, n1483);
xnor g1782 (n1798, n1681, n1238, n1227, n1280);
or   g1783 (n1835, n1713, n1423, n1696, n1413);
nand g1784 (n1731, n1712, n1487, n1695, n1672);
nor  g1785 (n1836, n1222, n1709, n1700, n1267);
and  g1786 (n1859, n1719, n1511, n1455, n1260);
nand g1787 (n1822, n1715, n1199, n1309, n1520);
nand g1788 (n1812, n1240, n1328, n1386, n1695);
and  g1789 (n1739, n1356, n1209, n1387, n1304);
or   g1790 (n1829, n1702, n1720, n1196, n1474);
or   g1791 (n1907, n1524, n1360, n1699, n1331);
or   g1792 (n1870, n1516, n1529, n1671, n1287);
and  g1793 (n1799, n1688, n1668, n1431, n1313);
or   g1794 (n1879, n1345, n1709, n1433, n1401);
and  g1795 (n1928, n1704, n1216, n1717, n1518);
nor  g1796 (n1871, n1218, n1681, n1483);
nor  g1797 (n1758, n1466, n1277, n1317, n1521);
nor  g1798 (n1776, n1364, n1278, n1228, n1511);
and  g1799 (n1827, n1231, n1482, n1262, n1699);
xor  g1800 (n1912, n1394, n1463, n1683, n1328);
or   g1801 (n1820, n1209, n1716, n1366, n1693);
xnor g1802 (n1779, n1347, n1710, n1230, n1411);
or   g1803 (n1857, n1258, n1241, n1330, n1676);
and  g1804 (n1823, n1371, n1688, n1424, n1373);
or   g1805 (n1723, n1373, n1672, n1685, n1698);
or   g1806 (n1944, n1459, n1309, n1400, n1372);
xnor g1807 (n1722, n1297, n1264, n1680, n1502);
and  g1808 (n1761, n1314, n1714, n1246, n1704);
and  g1809 (n1833, n1686, n1245, n1421, n1490);
xnor g1810 (n1864, n1314, n1256, n1381, n1673);
and  g1811 (n1897, n1355, n1699, n1714, n1307);
nand g1812 (n1787, n1244, n1397, n1459, n1677);
nor  g1813 (n1881, n1514, n1696, n1669, n1480);
or   g1814 (n1856, n1334, n1526, n1250, n1248);
and  g1815 (n1935, n1322, n1329, n1220, n1452);
or   g1816 (n1808, n1525, n1370, n1679);
or   g1817 (n1781, n1401, n1465, n1687, n1685);
xor  g1818 (n1865, n1327, n1670, n1254, n1442);
and  g1819 (n1736, n1445, n1682, n1471, n1357);
and  g1820 (n1825, n1395, n1487, n1194, n1364);
or   g1821 (n1861, n1686, n1721, n1708, n1409);
or   g1822 (n1794, n1692, n1706, n1721, n1368);
and  g1823 (n1826, n1278, n1354, n1456, n1368);
nand g1824 (n1757, n1689, n1464, n1688, n1332);
or   g1825 (n1852, n1450, n1393, n1242, n1471);
or   g1826 (n1918, n1265, n1692, n1374, n1486);
nand g1827 (n1834, n1689, n1704, n1718, n1340);
or   g1828 (n1929, n1426, n1693, n1207, n1422);
or   g1829 (n1750, n1363, n1428, n1678, n1285);
nand g1830 (n1791, n1688, n1236, n1285, n1269);
or   g1831 (n1868, n1441, n1251, n1668, n1442);
or   g1832 (n1802, n1507, n1350, n1212, n1701);
xnor g1833 (n1936, n1202, n1677, n1500, n1684);
and  g1834 (n1792, n1434, n1399, n1277, n1203);
nand g1835 (n1930, n1223, n1476, n1359, n1516);
nand g1836 (n1814, n1488, n1327, n1268, n1718);
xor  g1837 (n1813, n1397, n1280, n1347, n1248);
nor  g1838 (n1828, n1713, n1444, n1367, n1235);
xnor g1839 (n1766, n1446, n1412, n1390, n1707);
and  g1840 (n1850, n1515, n1261, n1449, n1434);
xnor g1841 (n1726, n1684, n1527, n1281, n1378);
xnor g1842 (n1775, n1303, n1705, n1706);
xnor g1843 (n1760, n1682, n1224, n1703, n1436);
nand g1844 (n1769, n1427, n1469, n1276, n1473);
xnor g1845 (n1858, n1676, n1374, n1667, n1508);
nor  g1846 (n1789, n1671, n1337, n1338, n1305);
or   g1847 (n1746, n1672, n1432, n1265, n1718);
xnor g1848 (n1878, n1272, n1382, n1714, n1303);
xor  g1849 (n1940, n1361, n1473, n1666, n1715);
xnor g1850 (n1788, n1355, n1507, n1226, n1505);
and  g1851 (n1851, n1502, n1513, n1494, n1219);
nor  g1852 (n1880, n1351, n1510, n1512, n1290);
and  g1853 (n1909, n1438, n1707, n1360, n1210);
nor  g1854 (n1843, n1312, n1422, n1344, n1297);
nand g1855 (n1816, n1686, n1369, n1416, n1234);
and  g1856 (n1923, n1289, n1381, n1419, n1698);
nand g1857 (n1875, n1345, n1233, n1251, n1295);
and  g1858 (n1831, n1292, n1689, n1698, n1493);
and  g1859 (n1860, n1491, n1379, n1445, n1384);
xnor g1860 (n1765, n1354, n1242, n1717, n1352);
nor  g1861 (n1786, n1480, n1367, n1301, n1428);
nand g1862 (n1724, n1495, n1404, n1437, n1351);
nor  g1863 (n1841, n1702, n1691, n1257, n1418);
and  g1864 (n1759, n1296, n1393, n1302, n1284);
and  g1865 (n1903, n1709, n1319, n1424, n1229);
or   g1866 (n1886, n1700, n1467, n1372, n1380);
or   g1867 (n1838, n1415, n1685, n1497, n1229);
xor  g1868 (n1925, n1282, n1667, n1315, n1274);
nor  g1869 (n1908, n1198, n1674, n1286, n1196);
xor  g1870 (n1895, n1453, n1243, n1239, n1676);
or   g1871 (n1883, n1253, n1712, n1270, n1719);
and  g1872 (n1742, n1195, n1474, n1702, n1243);
xor  g1873 (n1939, n1720, n1529, n1500, n1439);
xnor g1874 (n1740, n1512, n1468, n1215, n1266);
and  g1875 (n1837, n1336, n1438, n1358, n1298);
xnor g1876 (n1725, n1389, n1275, n1470, n1704);
or   g1877 (n1768, n1453, n1436, n1676, n1454);
or   g1878 (n1900, n1433, n1450, n1697, n1444);
nand g1879 (n1888, n1701, n1446, n1432, n1495);
and  g1880 (n1846, n1717, n1406, n1403, n1670);
nor  g1881 (n1811, n1304, n1350, n1716, n1672);
and  g1882 (n1855, n1497, n1506, n1668, n1419);
nor  g1883 (n1889, n1320, n1405, n1316, n1492);
or   g1884 (n1780, n1431, n1694, n1215, n1342);
xor  g1885 (n1899, n1705, n1200, n1706, n1692);
xnor g1886 (n1915, n1375, n1204, n1414, n1499);
nor  g1887 (n1783, n1465, n1683, n1437, n1208);
nor  g1888 (n1839, n1439, n1339, n1308, n1460);
xnor g1889 (n1773, n1288, n1696, n1417, n1348);
nand g1890 (n1770, n1456, n1457, n1289, n1698);
and  g1891 (n1867, n1496, n1486, n1669, n1329);
or   g1892 (n1898, n1455, n1528, n1240, n1391);
nor  g1893 (n1763, n1211, n1472, n1406, n1341);
and  g1894 (n1906, n1440, n1318, n1399, n1311);
nor  g1895 (n1885, n1356, n1673, n1259, n1321);
nor  g1896 (n1941, n1300, n1466, n1306, n1526);
or   g1897 (n1748, n1343, n1296, n1260, n1481);
nor  g1898 (n1849, n1519, n1341, n1259, n1377);
xnor g1899 (n1797, n1390, n1528, n1493, n1421);
or   g1900 (n1854, n1693, n1689, n1510, n1398);
xor  g1901 (n2077, n743, n866, n1936, n1843);
and  g1902 (n2159, n744, n895, n1544, n1883);
nand g1903 (n2071, n1875, n1585, n766, n922);
xor  g1904 (n2243, n1597, n1766, n1885, n1769);
or   g1905 (n1974, n819, n1614, n1926, n1930);
or   g1906 (n2078, n1820, n813, n784, n1726);
xnor g1907 (n2124, n1736, n892, n1551, n820);
nor  g1908 (n1961, n791, n753, n1933, n1547);
nor  g1909 (n2001, n1909, n808, n1908, n1934);
nand g1910 (n2149, n1930, n877, n1887, n774);
nor  g1911 (n2235, n1912, n1741, n1586, n1605);
nand g1912 (n2215, n853, n781, n907, n1586);
nand g1913 (n2041, n875, n1866, n1589, n1582);
xnor g1914 (n2157, n751, n910, n1913, n877);
nor  g1915 (n2282, n1621, n794, n782, n888);
xnor g1916 (n2017, n1830, n741, n921, n1557);
nor  g1917 (n2137, n812, n1850, n867, n852);
nor  g1918 (n2161, n908, n1862, n817, n1608);
and  g1919 (n2257, n1943, n1560, n863, n1740);
and  g1920 (n2117, n770, n1562, n846, n915);
and  g1921 (n2092, n1878, n1901, n900, n889);
or   g1922 (n2125, n817, n1724, n1592, n783);
xor  g1923 (n2059, n1536, n744, n899, n752);
or   g1924 (n1975, n754, n749, n862, n1542);
nor  g1925 (n2290, n1536, n1945, n807, n848);
nand g1926 (n2070, n1728, n872, n800, n754);
nor  g1927 (n1956, n920, n1753, n800, n888);
and  g1928 (n2134, n795, n769, n747, n1912);
nand g1929 (n1976, n823, n1895, n841, n1605);
and  g1930 (n2160, n1577, n875, n1612, n916);
and  g1931 (n2111, n915, n824, n762, n1792);
or   g1932 (n2042, n846, n1593, n1576, n1778);
nand g1933 (n2130, n864, n1794, n904, n1833);
nor  g1934 (n2270, n1797, n756, n837, n1844);
nor  g1935 (n2007, n844, n872, n868, n1600);
nor  g1936 (n2062, n862, n1889, n1798, n1845);
and  g1937 (n2028, n1740, n911, n1801, n1874);
and  g1938 (n2139, n1903, n898, n904, n1623);
nand g1939 (n1977, n1825, n749, n875, n870);
and  g1940 (n1972, n1921, n1756, n1749, n1869);
xor  g1941 (n1953, n1839, n757, n1817, n1750);
and  g1942 (n2067, n833, n1739, n838, n879);
xor  g1943 (n2133, n1544, n760, n1823, n878);
nor  g1944 (n2024, n1915, n881, n772, n1790);
nand g1945 (n2250, n815, n1754, n823, n1766);
and  g1946 (n1990, n883, n1942, n847, n803);
nand g1947 (n2231, n806, n883, n775, n1613);
or   g1948 (n2104, n787, n760, n1770, n1747);
nand g1949 (n2262, n881, n843, n923, n1602);
xor  g1950 (n2255, n919, n1783, n1599, n898);
nand g1951 (n2198, n755, n816, n799, n1920);
xnor g1952 (n2277, n1816, n855, n890, n869);
nor  g1953 (n2034, n780, n772, n1537, n774);
xor  g1954 (n1991, n1893, n1589, n837, n1842);
xor  g1955 (n2239, n786, n741, n1848, n828);
nor  g1956 (n2109, n1533, n856, n825, n1762);
nand g1957 (n2146, n751, n1836, n1577, n820);
and  g1958 (n2002, n1920, n1615, n748, n744);
or   g1959 (n1963, n1882, n1768, n783, n873);
or   g1960 (n2174, n1541, n835, n1889, n747);
xor  g1961 (n2088, n1780, n884, n1558);
and  g1962 (n2266, n822, n794, n1863, n782);
and  g1963 (n2199, n1563, n917, n1798, n1590);
xor  g1964 (n1964, n831, n1917, n905, n906);
or   g1965 (n2195, n1869, n769, n1781, n1550);
nand g1966 (n2275, n757, n1729, n853, n1880);
or   g1967 (n2165, n1610, n1744, n1893, n1859);
xnor g1968 (n2208, n778, n1545, n1738, n1799);
or   g1969 (n2203, n913, n870, n1574, n920);
xor  g1970 (n2144, n766, n906, n1882, n851);
xnor g1971 (n2248, n878, n1885, n806, n748);
nand g1972 (n2283, n901, n1779, n858, n771);
xor  g1973 (n2219, n1813, n1905, n1846, n1726);
nor  g1974 (n2022, n809, n902, n1552, n1918);
or   g1975 (n2057, n1732, n912, n1932, n914);
or   g1976 (n1994, n1813, n814, n1823, n1572);
nor  g1977 (n2206, n758, n747, n1853, n831);
nand g1978 (n1989, n1620, n1533, n833, n791);
or   g1979 (n1960, n810, n825, n771, n767);
nor  g1980 (n2014, n758, n1617, n845, n1734);
nand g1981 (n2269, n740, n1750, n1561, n1731);
or   g1982 (n1987, n1548, n755, n858, n786);
nand g1983 (n2260, n1864, n853, n1830, n1600);
xor  g1984 (n2240, n900, n1617, n1723, n914);
xor  g1985 (n2251, n804, n885, n857, n746);
nor  g1986 (n2006, n850, n1582, n788, n832);
nand g1987 (n2263, n1770, n1847, n797, n908);
xor  g1988 (n2136, n792, n1795, n886, n862);
xor  g1989 (n2214, n1767, n849, n776, n1596);
nand g1990 (n2020, n790, n879, n893, n832);
and  g1991 (n2032, n1923, n1916, n1572, n1551);
xor  g1992 (n2023, n1738, n1865, n1858, n909);
or   g1993 (n2035, n1879, n1924, n889, n1538);
and  g1994 (n2181, n779, n1918, n836, n1751);
and  g1995 (n2221, n784, n1532, n1744, n1768);
xor  g1996 (n2210, n859, n1809, n811, n801);
nor  g1997 (n2039, n1587, n1545, n761, n919);
or   g1998 (n2220, n1769, n923, n1877, n1802);
and  g1999 (n2018, n762, n763, n798, n760);
and  g2000 (n2000, n847, n1794, n1530, n1616);
nor  g2001 (n1978, n840, n904, n1786, n1821);
nor  g2002 (n2213, n810, n1896, n892, n798);
nand g2003 (n2202, n886, n815, n1914, n1888);
nand g2004 (n2033, n1575, n1917, n803, n780);
or   g2005 (n2253, n791, n797, n1759, n1902);
or   g2006 (n2147, n805, n920, n1729, n1868);
nand g2007 (n2140, n1618, n887, n1776, n1570);
nand g2008 (n1970, n1598, n1611, n755, n861);
nand g2009 (n1997, n758, n909, n776, n767);
or   g2010 (n2279, n918, n1807, n783, n830);
xor  g2011 (n2172, n841, n911, n1585, n1827);
nor  g2012 (n2040, n924, n1584, n776, n1751);
xor  g2013 (n2212, n808, n1833, n822, n1540);
xor  g2014 (n2112, n1815, n1852, n850, n801);
and  g2015 (n1955, n1847, n1787, n852, n779);
nor  g2016 (n2191, n759, n1797, n830, n1782);
xor  g2017 (n1966, n797, n833, n754, n1940);
nand g2018 (n2064, n1932, n917, n773, n841);
xnor g2019 (n2110, n1836, n824, n1607, n1808);
nand g2020 (n2065, n835, n1939, n762, n1725);
or   g2021 (n2265, n892, n824, n760, n786);
nand g2022 (n2060, n802, n857, n1848, n1878);
xor  g2023 (n2115, n1810, n761, n874, n1743);
xor  g2024 (n2089, n918, n1565, n1929, n1619);
nor  g2025 (n1951, n1834, n912, n1831, n893);
and  g2026 (n2222, n740, n890, n822, n1552);
and  g2027 (n2171, n1888, n1565, n859, n1887);
or   g2028 (n2236, n1567, n865, n792, n1737);
xnor g2029 (n2047, n863, n1602, n1825, n1730);
and  g2030 (n2186, n826, n773, n818, n1872);
nor  g2031 (n2087, n795, n1614, n861, n1884);
nand g2032 (n2197, n770, n821, n843, n757);
nand g2033 (n2167, n1616, n1627, n801, n887);
nor  g2034 (n2106, n1580, n1904, n818, n855);
and  g2035 (n1949, n832, n777, n834, n752);
xor  g2036 (n2114, n771, n767, n1790, n754);
and  g2037 (n2247, n1553, n1782, n766, n1804);
xnor g2038 (n2019, n1838, n751, n898, n883);
xor  g2039 (n2141, n822, n889, n1784, n1774);
nor  g2040 (n2154, n1815, n1806, n1743, n1626);
and  g2041 (n2216, n769, n842, n1849, n1880);
xnor g2042 (n2101, n1858, n749, n829, n899);
or   g2043 (n1995, n823, n849, n782, n799);
xnor g2044 (n1983, n804, n1931, n1570, n1554);
nand g2045 (n2152, n1856, n845, n1754, n813);
nor  g2046 (n2090, n905, n1891, n781, n1560);
nand g2047 (n1959, n874, n1745, n1550, n1876);
xor  g2048 (n2038, n859, n1890, n1580, n1826);
xnor g2049 (n2280, n787, n781, n819, n1911);
nand g2050 (n2268, n916, n911, n838, n819);
xnor g2051 (n2234, n1817, n795, n877, n1566);
or   g2052 (n1986, n1573, n814, n857, n750);
and  g2053 (n2063, n833, n1837, n887, n879);
nor  g2054 (n2244, n1569, n1827, n1757, n877);
nor  g2055 (n2192, n775, n1892, n747, n869);
xnor g2056 (n2180, n913, n1855, n921, n860);
nand g2057 (n2122, n852, n897, n1819, n888);
and  g2058 (n2272, n1832, n869, n1741, n1591);
and  g2059 (n2100, n815, n826, n1787, n775);
nand g2060 (n2037, n840, n1844, n880, n895);
nor  g2061 (n2026, n1622, n1764, n867, n756);
xnor g2062 (n1980, n874, n1875, n1546, n1922);
and  g2063 (n2223, n1615, n1800, n922, n1891);
or   g2064 (n2278, n882, n758, n1724, n893);
and  g2065 (n2211, n1543, n1538, n1804, n882);
or   g2066 (n2098, n1780, n886, n1599, n1596);
xnor g2067 (n2209, n821, n742, n830, n1877);
nand g2068 (n2031, n798, n839, n1543, n1742);
xnor g2069 (n2258, n1808, n766, n1755, n897);
nor  g2070 (n1993, n1776, n1913, n768, n894);
or   g2071 (n1981, n1775, n787, n1559, n1537);
nand g2072 (n2185, n894, n1857, n844, n1826);
and  g2073 (n2103, n801, n780, n1862, n1564);
nand g2074 (n2113, n1777, n891, n1748, n903);
nand g2075 (n2175, n1608, n1828, n905, n844);
xor  g2076 (n2121, n896, n880, n838, n1627);
nand g2077 (n2230, n742, n880, n1837, n834);
and  g2078 (n1982, n1802, n764, n809, n897);
and  g2079 (n2027, n1843, n1890, n1898, n815);
and  g2080 (n2120, n1789, n834, n788, n1900);
nor  g2081 (n1984, n1871, n1783, n746, n1779);
nand g2082 (n1988, n789, n1730, n1903, n851);
nand g2083 (n1992, n867, n799, n1884, n1806);
xnor g2084 (n2158, n780, n768, n827, n1597);
nor  g2085 (n2075, n1535, n890, n1727, n1777);
nor  g2086 (n2004, n835, n868, n809, n1811);
and  g2087 (n2123, n828, n914, n1910, n1938);
xnor g2088 (n2178, n1935, n800, n861, n864);
nand g2089 (n2030, n764, n1540, n1534, n1816);
xor  g2090 (n2094, n804, n813, n884, n881);
nand g2091 (n2205, n844, n871, n1886, n916);
nor  g2092 (n2054, n790, n1814, n1619, n828);
nor  g2093 (n1948, n1745, n1943, n1941, n854);
nand g2094 (n2058, n753, n773, n1598, n891);
xnor g2095 (n2238, n1581, n785, n778, n869);
and  g2096 (n2008, n856, n899, n1865, n765);
xor  g2097 (n1952, n1872, n882, n746, n890);
or   g2098 (n2189, n806, n853, n860, n907);
xnor g2099 (n2015, n745, n854, n866, n1611);
or   g2100 (n2029, n1557, n1934, n1625, n1841);
and  g2101 (n2095, n1732, n1840, n1773);
nor  g2102 (n1998, n1805, n1924, n1907, n1739);
xnor g2103 (n1958, n894, n746, n817, n1603);
or   g2104 (n1996, n1854, n793, n1612, n1556);
or   g2105 (n2153, n842, n1906, n892, n912);
nand g2106 (n2048, n871, n763, n897, n789);
xnor g2107 (n2036, n1727, n881, n870, n834);
nand g2108 (n2273, n891, n1756, n1748, n1735);
xor  g2109 (n2150, n827, n1881, n787, n814);
and  g2110 (n2091, n1548, n1927, n850, n808);
and  g2111 (n2143, n868, n768, n1623, n788);
or   g2112 (n2256, n1831, n761, n785, n860);
or   g2113 (n2188, n1764, n1860, n1583, n866);
nor  g2114 (n2267, n1935, n1604, n774, n1921);
or   g2115 (n2055, n755, n1838, n902, n1938);
or   g2116 (n2142, n1583, n1563, n782, n1807);
and  g2117 (n2050, n1576, n1723, n820, n793);
xor  g2118 (n2162, n846, n916, n854, n796);
xor  g2119 (n2168, n880, n829, n868, n792);
nand g2120 (n2099, n1531, n784, n1933, n878);
xor  g2121 (n2176, n829, n896, n1594, n1892);
xor  g2122 (n1947, n808, n1579, n1899, n763);
nand g2123 (n2288, n1568, n839, n770, n818);
nand g2124 (n1968, n1812, n745, n895, n807);
nor  g2125 (n1950, n1568, n1795, n1812, n792);
and  g2126 (n1973, n804, n875, n873, n866);
or   g2127 (n2184, n1799, n810, n913, n1822);
nor  g2128 (n2228, n1791, n1604, n1542, n1603);
xnor g2129 (n2045, n1532, n789, n921);
nor  g2130 (n2066, n858, n816, n1626, n843);
or   g2131 (n2164, n812, n796, n1575, n745);
or   g2132 (n2190, n863, n1855, n748, n864);
nor  g2133 (n2148, n1607, n888, n785, n903);
or   g2134 (n2177, n1925, n1854, n1909, n1868);
nor  g2135 (n2227, n914, n777, n1555, n825);
xnor g2136 (n1971, n1852, n743, n1584, n1722);
or   g2137 (n2056, n950, n1870, n1796, n1820);
or   g2138 (n2271, n1883, n906, n1939, n1749);
and  g2139 (n2052, n744, n1851, n745, n1845);
and  g2140 (n2009, n759, n803, n1613, n1767);
and  g2141 (n1967, n827, n1898, n922, n899);
and  g2142 (n2131, n774, n1905, n839, n764);
or   g2143 (n2108, n1937, n873, n903, n752);
xnor g2144 (n2082, n765, n847, n1900, n887);
or   g2145 (n2201, n1765, n922, n865, n1574);
nand g2146 (n2252, n885, n797, n1809, n828);
nand g2147 (n1979, n1904, n786, n803, n1871);
xnor g2148 (n2207, n920, n1908, n847, n1587);
nor  g2149 (n2072, n1906, n865, n1914, n902);
nand g2150 (n2170, n1731, n1910, n1879, n743);
xnor g2151 (n2119, n849, n912, n1911, n840);
xnor g2152 (n2237, n873, n1829, n1774, n1772);
and  g2153 (n2053, n1942, n1788, n1725, n1571);
xnor g2154 (n1999, n891, n1566, n818, n1927);
or   g2155 (n2232, n783, n1592, n852, n743);
xor  g2156 (n2285, n759, n902, n1894, n1558);
or   g2157 (n2126, n751, n1819, n805, n1553);
xnor g2158 (n2005, n1606, n841, n769, n1864);
and  g2159 (n2138, n1781, n848, n753, n872);
nand g2160 (n2196, n790, n900, n796, n845);
xnor g2161 (n2274, n1853, n832, n1734, n1578);
nor  g2162 (n2127, n768, n842, n1928, n1922);
or   g2163 (n2097, n1610, n772, n809, n1896);
xor  g2164 (n2093, n1945, n827, n1840, n1867);
nand g2165 (n2051, n1841, n1801, n1578, n1554);
xnor g2166 (n2151, n855, n856, n846, n1941);
nor  g2167 (n2261, n923, n896, n838, n876);
and  g2168 (n2204, n826, n773, n1539, n1549);
nor  g2169 (n2069, n850, n1534, n884, n793);
nand g2170 (n2128, n756, n811, n918, n1863);
nand g2171 (n2074, n1539, n1728, n1785, n1561);
xor  g2172 (n2102, n872, n816, n1755, n1894);
and  g2173 (n1946, n876, n1609, n1861, n1873);
xor  g2174 (n2179, n917, n807, n860, n1936);
or   g2175 (n2135, n795, n1834, n1793, n779);
xor  g2176 (n2013, n910, n859, n921, n1842);
nor  g2177 (n1985, n1556, n1733, n1788, n830);
xor  g2178 (n2118, n805, n910, n1818, n915);
nor  g2179 (n2046, n790, n905, n1784, n1861);
nor  g2180 (n2200, n1822, n1549, n1796, n1928);
nor  g2181 (n2011, n919, n1588, n867, n901);
nand g2182 (n2281, n1814, n1874, n1899, n1897);
and  g2183 (n1962, n1569, n1824, n864, n1907);
and  g2184 (n2049, n855, n840, n1886, n919);
xor  g2185 (n2025, n767, n904, n1546, n907);
nor  g2186 (n1957, n741, n896, n885, n1803);
xnor g2187 (n2264, n1791, n1916, n1860, n759);
or   g2188 (n2079, n862, n842, n806, n765);
or   g2189 (n2083, n826, n1763, n820, n1606);
nor  g2190 (n2218, n1919, n1562, n794, n908);
and  g2191 (n2012, n1761, n1573, n1747, n1785);
xor  g2192 (n2068, n1759, n1805, n1594, n849);
and  g2193 (n2194, n742, n781, n1940, n1601);
or   g2194 (n2016, n788, n913, n810, n1824);
xnor g2195 (n2245, n791, n777, n1620, n1775);
and  g2196 (n2129, n814, n771, n1800, n1593);
nand g2197 (n2073, n1762, n753, n908, n909);
and  g2198 (n2187, n1625, n1609, n879, n1761);
or   g2199 (n2156, n1870, n1763, n1867, n807);
and  g2200 (n2193, n1579, n1624, n901, n1595);
and  g2201 (n2010, n1902, n1931, n798, n898);
nor  g2202 (n2076, n848, n817, n1590, n1859);
nand g2203 (n2086, n915, n750, n851, n1835);
xor  g2204 (n2224, n845, n1628, n856, n799);
nor  g2205 (n2105, n1771, n1722, n876, n835);
xor  g2206 (n2155, n883, n1772, n813, n1757);
nand g2207 (n1954, n750, n1588, n1765, n901);
nor  g2208 (n2287, n1601, n1559, n874, n821);
xnor g2209 (n2084, n1535, n836, n851, n1915);
or   g2210 (n1965, n1944, n894, n1778, n843);
nand g2211 (n2166, n750, n765, n824, n1857);
xor  g2212 (n2173, n785, n777, n1850, n906);
and  g2213 (n2116, n778, n1846, n1752, n857);
and  g2214 (n2043, n865, n1866, n1829, n1839);
xor  g2215 (n2217, n1786, n1789, n742, n831);
xnor g2216 (n2021, n1760, n882, n1737, n900);
and  g2217 (n2145, n1925, n1923, n1771, n819);
xor  g2218 (n2254, n1929, n1746, n1881, n870);
xor  g2219 (n2276, n917, n909, n1876, n1733);
or   g2220 (n2226, n761, n871, n764, n1618);
nand g2221 (n2061, n1555, n1792, n839, n889);
xnor g2222 (n2163, n1818, n794, n907, n836);
nand g2223 (n2225, n812, n816, n903, n1811);
xnor g2224 (n2259, n779, n885, n770, n1581);
and  g2225 (n2183, n772, n811, n749, n1897);
xor  g2226 (n2246, n836, n1531, n1919, n1926);
or   g2227 (n2085, n776, n1567, n831, n1803);
and  g2228 (n1969, n878, n821, n1828, n1760);
nor  g2229 (n2242, n811, n858, n1752, n741);
xor  g2230 (n2289, n911, n748, n1746, n886);
nor  g2231 (n2241, n1541, n800, n1735, n1753);
nor  g2232 (n2286, n1742, n1851, n793, n1564);
nand g2233 (n2107, n1571, n895, n1622, n829);
xor  g2234 (n2080, n756, n802, n876, n1849);
or   g2235 (n2249, n805, n1835, n812, n752);
xor  g2236 (n2229, n923, n837, n861, n784);
nor  g2237 (n2284, n837, n796, n1901, n918);
xnor g2238 (n2003, n1595, n1758, n757, n1621);
nor  g2239 (n2169, n1810, n1736, n825, n762);
and  g2240 (n2132, n823, n775, n863, n1937);
xor  g2241 (n2044, n778, n854, n1873, n802);
and  g2242 (n2081, n1832, n1758, n763, n1856);
xnor g2243 (n2096, n910, n1591, n1944, n848);
xor  g2244 (n2182, n1547, n1895, n871, n1821);
nand g2245 (n2233, n1793, n802, n893, n1624);
xor  g2246 (n2307, n2094, n1956, n2081, n2175);
nor  g2247 (n2301, n2034, n1951, n2189, n2155);
nor  g2248 (n2379, n2236, n1985, n2017, n2158);
nor  g2249 (n2341, n1996, n2254, n2154, n2073);
or   g2250 (n2387, n1990, n2184, n2009, n2064);
nor  g2251 (n2365, n2083, n1983, n2260, n2008);
xor  g2252 (n2380, n1984, n2010, n2071, n2230);
nor  g2253 (n2393, n2139, n2178, n1975, n2179);
nor  g2254 (n2423, n2176, n2046, n1962, n2134);
or   g2255 (n2319, n1949, n2164, n2225, n2018);
nor  g2256 (n2364, n2002, n2028, n2070, n2029);
nand g2257 (n2315, n2152, n2115, n2058, n1982);
nand g2258 (n2360, n2077, n2204, n2145, n1961);
xor  g2259 (n2349, n1993, n1982, n1963, n2197);
nand g2260 (n2442, n2257, n2109, n2019, n2006);
nor  g2261 (n2425, n2160, n2198, n2255, n2171);
xor  g2262 (n2424, n1967, n1979, n2126, n2233);
nand g2263 (n2297, n2234, n2224, n2129, n2112);
xor  g2264 (n2299, n1952, n2111, n2050, n2216);
xor  g2265 (n2416, n1966, n2227, n2027, n2246);
and  g2266 (n2399, n2269, n2059, n2214, n2154);
xnor g2267 (n2342, n2200, n1965, n1983, n2078);
xor  g2268 (n2436, n1999, n2016, n2048, n1948);
xor  g2269 (n2439, n2190, n2036, n1997, n2197);
or   g2270 (n2396, n2148, n2003, n2121, n2267);
and  g2271 (n2420, n2006, n2260, n2156, n1970);
nor  g2272 (n2303, n2001, n2052, n2069, n2034);
xor  g2273 (n2384, n2259, n2139, n2090, n2255);
nand g2274 (n2441, n2016, n2040, n1989, n2194);
or   g2275 (n2382, n2012, n2207, n2246, n2212);
nor  g2276 (n2337, n2211, n1964, n2262, n2159);
nand g2277 (n2421, n2076, n2052, n2110, n1995);
xnor g2278 (n2359, n2053, n2241, n2103, n2151);
xor  g2279 (n2386, n2089, n2126, n2230, n2263);
nand g2280 (n2374, n2263, n2147, n2184, n2210);
xnor g2281 (n2409, n2042, n2183, n2082, n1976);
nand g2282 (n2317, n2026, n2108, n2058, n2014);
nand g2283 (n2357, n2086, n2025, n1977, n2217);
xor  g2284 (n2348, n2186, n2047, n1947, n2232);
nor  g2285 (n2391, n2161, n2000, n2075, n2209);
xnor g2286 (n2309, n1969, n2131, n2024, n2037);
xnor g2287 (n2346, n2007, n2211, n2118, n2251);
xor  g2288 (n2328, n2187, n2178, n2203, n2256);
nor  g2289 (n2339, n2202, n2103, n1999, n2113);
xor  g2290 (n2397, n2258, n1985, n2125, n2001);
nand g2291 (n2295, n2169, n2079, n2193, n1972);
and  g2292 (n2310, n1960, n2195, n2250, n2168);
xnor g2293 (n2318, n2023, n2152, n2074, n2142);
nand g2294 (n2389, n2020, n2060, n2043, n2192);
and  g2295 (n2340, n2065, n2241, n2170, n1965);
nor  g2296 (n2408, n2240, n2079, n2203, n2251);
or   g2297 (n2437, n2244, n2173, n2132, n1991);
or   g2298 (n2324, n2123, n2008, n2149, n2143);
nor  g2299 (n2358, n2031, n2088, n2141, n2242);
or   g2300 (n2417, n1992, n2061, n1980, n2073);
xnor g2301 (n2450, n2035, n1946, n2122, n2096);
and  g2302 (n2445, n1958, n2084, n2082, n2261);
nor  g2303 (n2291, n2237, n2117, n1949, n2156);
or   g2304 (n2313, n2031, n2224, n1956, n1957);
or   g2305 (n2347, n2049, n2261, n2015, n1959);
and  g2306 (n2452, n2011, n2166, n1970, n2124);
and  g2307 (n2363, n2225, n2022, n1973, n1977);
xnor g2308 (n2395, n2028, n2032, n2071, n2080);
or   g2309 (n2333, n2039, n2041, n2004, n2248);
nor  g2310 (n2376, n2259, n2022, n2137, n2056);
xor  g2311 (n2311, n2145, n2165, n2213, n2134);
xor  g2312 (n2398, n2219, n2209, n2256, n2228);
and  g2313 (n2426, n2097, n2170, n2137, n2038);
xnor g2314 (n2418, n2242, n2207, n1987, n2039);
xnor g2315 (n2413, n2101, n2267, n2102, n2062);
and  g2316 (n2381, n2151, n2176, n2217, n2102);
and  g2317 (n2373, n2243, n1974, n1990, n2168);
xnor g2318 (n2448, n2252, n2253, n2005, n2074);
xnor g2319 (n2296, n2220, n2061, n2188, n2021);
xor  g2320 (n2435, n1946, n2192, n2144, n2147);
and  g2321 (n2407, n2113, n2063, n2269, n2081);
nand g2322 (n2321, n1963, n1979, n2215, n2221);
nor  g2323 (n2371, n2012, n2153, n2140, n1998);
and  g2324 (n2343, n2245, n2062, n1976, n2116);
nand g2325 (n2306, n2084, n2050, n2185, n1988);
or   g2326 (n2332, n2229, n2040, n2112, n2171);
nor  g2327 (n2304, n2085, n2138, n2066, n1989);
and  g2328 (n2327, n2086, n2208, n2244, n2093);
nand g2329 (n2316, n2146, n2108, n2070, n2055);
xnor g2330 (n2350, n2106, n1968, n2268, n1957);
or   g2331 (n2404, n2198, n2033, n2193, n2010);
nor  g2332 (n2427, n1958, n2100, n2181, n1967);
and  g2333 (n2394, n1948, n2130, n2098, n2090);
xor  g2334 (n2366, n2142, n2257, n2076, n2120);
xor  g2335 (n2434, n2119, n2000, n2166, n2191);
and  g2336 (n2432, n2132, n2054, n2239, n2165);
xnor g2337 (n2293, n1955, n2115, n2180, n2107);
xor  g2338 (n2429, n2240, n2023, n2232, n2049);
nand g2339 (n2403, n2199, n2186, n2128, n2140);
and  g2340 (n2338, n2179, n2053, n2215, n2045);
xnor g2341 (n2402, n2177, n2136, n2247, n1997);
nand g2342 (n2353, n2092, n2222, n2221, n2105);
and  g2343 (n2430, n2169, n2119, n2109, n2057);
xnor g2344 (n2300, n2174, n2167, n2072, n2021);
nor  g2345 (n2362, n2048, n2149, n2249, n2030);
xor  g2346 (n2370, n2219, n1984, n1978, n1952);
and  g2347 (n2344, n2264, n1998, n1954, n2127);
and  g2348 (n2361, n2226, n2044, n2206, n2135);
xnor g2349 (n2329, n2223, n2265, n2172, n2235);
nor  g2350 (n2411, n2133, n2067, n2174, n2041);
nand g2351 (n2314, n2208, n2004, n2005, n2007);
and  g2352 (n2447, n1951, n2087, n2243, n1955);
xor  g2353 (n2449, n2032, n1994, n2066, n2051);
nor  g2354 (n2400, n2124, n2180, n1971, n2143);
xor  g2355 (n2330, n2069, n2185, n2253, n2254);
and  g2356 (n2312, n1974, n2104, n2116, n2059);
or   g2357 (n2444, n1973, n2068, n2250, n1960);
nand g2358 (n2438, n2196, n2128, n1950, n2056);
nand g2359 (n2331, n2064, n2033, n2155, n2196);
nand g2360 (n2345, n2172, n2054, n2017, n2099);
nand g2361 (n2415, n2191, n1972, n2089, n2194);
and  g2362 (n2336, n1966, n2121, n2038, n2092);
and  g2363 (n2355, n1978, n2051, n2200, n2248);
and  g2364 (n2428, n2160, n2262, n1975, n2015);
xnor g2365 (n2368, n2047, n2019, n2105, n2159);
and  g2366 (n2405, n2231, n1962, n2029, n1953);
nor  g2367 (n2372, n1947, n2236, n2216, n2043);
nand g2368 (n2326, n2104, n2150, n1991, n2144);
and  g2369 (n2422, n2229, n2205, n2201, n2037);
nor  g2370 (n2378, n1953, n2264, n2163, n2093);
nand g2371 (n2302, n2057, n2183, n2018, n2095);
or   g2372 (n2305, n1954, n2003, n2223, n2222);
xor  g2373 (n2375, n2233, n2227, n2158, n2096);
nand g2374 (n2352, n2148, n2114, n2098, n2266);
or   g2375 (n2412, n2212, n2122, n2065, n2060);
xnor g2376 (n2351, n2157, n2234, n1986, n1988);
nor  g2377 (n2385, n2107, n2091, n2228, n2100);
or   g2378 (n2410, n2177, n2097, n2009, n2175);
nand g2379 (n2388, n2011, n2077, n2235, n2123);
and  g2380 (n2356, n2120, n2091, n2106, n2266);
and  g2381 (n2451, n2036, n1992, n2020, n2075);
nand g2382 (n2390, n2117, n2182, n1959, n2094);
nand g2383 (n2325, n2201, n2173, n2249, n2218);
xnor g2384 (n2446, n2099, n2162, n2042, n1995);
nor  g2385 (n2320, n2252, n2210, n2068, n1987);
nand g2386 (n2406, n2202, n2214, n2161, n2181);
and  g2387 (n2414, n2055, n1950, n2182, n2220);
xnor g2388 (n2322, n1981, n2125, n2027, n2014);
xnor g2389 (n2431, n2111, n2044, n2085, n2226);
and  g2390 (n2308, n1994, n2231, n2204, n1986);
nor  g2391 (n2367, n2218, n2135, n2045, n2153);
nand g2392 (n2443, n2035, n2187, n2206, n2088);
nor  g2393 (n2392, n2188, n2080, n2245, n2129);
xnor g2394 (n2440, n2025, n2026, n1969, n2114);
and  g2395 (n2292, n1964, n1971, n2133, n2213);
and  g2396 (n2323, n2013, n2127, n2237, n2072);
and  g2397 (n2369, n2238, n2195, n1996, n2118);
and  g2398 (n2377, n1961, n2002, n2138, n2205);
xor  g2399 (n2298, n2164, n2078, n2162, n2046);
xnor g2400 (n2433, n2268, n2136, n2146, n2238);
xnor g2401 (n2383, n2101, n2199, n2258, n1993);
nor  g2402 (n2294, n2150, n1980, n2190, n2013);
and  g2403 (n2354, n2130, n2095, n2131, n2265);
and  g2404 (n2419, n2083, n2087, n2067, n2239);
xor  g2405 (n2334, n2247, n2189, n2157, n2167);
xnor g2406 (n2335, n2163, n2110, n1981, n2063);
xnor g2407 (n2401, n2024, n1968, n2030, n2141);
xnor g2408 (n2457, n2294, n2303, n2302, n2293);
and  g2409 (n2454, n2304, n2299, n2291, n2307);
nor  g2410 (n2455, n2295, n2309, n2298, n2310);
nor  g2411 (n2453, n2297, n2305, n2300, n2296);
xnor g2412 (n2456, n2306, n2292, n2301, n2308);
not  g2413 (n2458, n2457);
buf  g2414 (n2461, n2455);
not  g2415 (n2460, n2454);
not  g2416 (n2459, n2456);
buf  g2417 (n2462, n2458);
not  g2418 (n2463, n2458);
buf  g2419 (n2464, n2463);
not  g2420 (n2466, n1030);
xor  g2421 (n2467, n2463, n2270, n1031, n2311);
nand g2422 (n2465, n1030, n2270, n2462);
xor  g2423 (n2470, n2317, n2314, n2465);
nor  g2424 (n2469, n2315, n2316, n2318);
xor  g2425 (n2468, n2312, n2464, n2313);
nand g2426 (n2478, n2319, n2339, n2345, n2468);
nor  g2427 (n2477, n2341, n2468, n2338);
and  g2428 (n2474, n2334, n2324, n2469);
nor  g2429 (n2473, n2331, n2470, n2335, n2329);
or   g2430 (n2472, n2470, n2320, n2343, n2322);
xor  g2431 (n2476, n2340, n2337, n2469, n2328);
xor  g2432 (n2479, n2327, n2325, n2333, n2336);
or   g2433 (n2475, n2326, n2344, n2321, n2342);
xor  g2434 (n2471, n2470, n2323, n2330, n2332);
nand g2435 (n2484, n2358, n2346, n2357, n2474);
or   g2436 (n2480, n2352, n2359, n2356, n2350);
or   g2437 (n2482, n2354, n2472, n2473, n2360);
or   g2438 (n2481, n2347, n2348, n2475, n2349);
nor  g2439 (n2483, n2351, n2471, n2355, n2353);
nand g2440 (n2486, n2364, n2372, n2369, n2363);
nand g2441 (n2488, n2365, n2484, n2361, n2362);
nor  g2442 (n2485, n2481, n2366, n2371, n2368);
xor  g2443 (n2487, n2367, n2483, n2482, n2370);
xor  g2444 (n2500, n1633, n2458, n2459, n2486);
nand g2445 (n2499, n2467, n2488, n2485, n2460);
nand g2446 (n2493, n2373, n2461, n2459);
nor  g2447 (n2490, n1631, n2486, n2487);
or   g2448 (n2489, n2458, n1640, n2460, n1628);
xnor g2449 (n2491, n1634, n2485, n2486, n1639);
xor  g2450 (n2497, n1634, n2485, n2461);
xor  g2451 (n2503, n1641, n2461, n2465, n1637);
or   g2452 (n2504, n2487, n2488, n1638, n2466);
xnor g2453 (n2501, n2466, n2485, n1630, n1629);
nand g2454 (n2502, n1640, n1636, n1630, n1641);
nand g2455 (n2498, n2487, n2488, n1632, n1031);
and  g2456 (n2494, n2460, n1631, n1638, n2374);
xor  g2457 (n2496, n2460, n2487, n1636, n1639);
xnor g2458 (n2495, n2488, n1635, n1633, n2459);
xnor g2459 (n2492, n1632, n1635, n1629, n1637);
and  g2460 (n2517, n2496, n2500, n1003, n2377);
or   g2461 (n2508, n2499, n2497, n2491, n2496);
nor  g2462 (n2516, n2495, n2381, n2501, n950);
and  g2463 (n2511, n2498, n2492, n2490, n2495);
xnor g2464 (n2510, n2491, n2504, n2500);
nand g2465 (n2506, n2494, n2378, n2492, n2376);
xor  g2466 (n2512, n2382, n2498, n2500, n2467);
xor  g2467 (n2513, n2502, n2499, n2489, n2380);
or   g2468 (n2519, n2500, n2497, n2501);
and  g2469 (n2518, n2497, n2503, n2498, n2504);
or   g2470 (n2514, n2494, n2499, n2501);
and  g2471 (n2507, n2490, n2502, n2504, n2493);
nand g2472 (n2509, n2375, n1003, n2503);
nor  g2473 (n2505, n2379, n2497, n2489, n2502);
nor  g2474 (n2515, n2502, n2503, n2498, n2493);
nor  g2475 (n2524, n2516, n2508, n2510, n2505);
or   g2476 (n2521, n2513, n2515, n2506, n2517);
nor  g2477 (n2522, n2518, n2511, n2512, n2515);
xnor g2478 (n2520, n2510, n2509, n2514, n2508);
xnor g2479 (n2526, n2512, n2505, n2507, n2509);
xor  g2480 (n2523, n2507, n2513, n2518, n2516);
and  g2481 (n2525, n2514, n2517, n2511, n2506);
nand g2482 (n2527, n2384, n2387, n2526, n2386);
and  g2483 (n2528, n2388, n2525, n2385, n2383);
nor  g2484 (n2532, n2527, n2528, n1052, n2477);
nor  g2485 (n2534, n2519, n2527, n2478, n2391);
nand g2486 (n2531, n2528, n1053, n2390);
nand g2487 (n2530, n2528, n1015, n2527, n2479);
nand g2488 (n2533, n2527, n2528, n2389, n2479);
xor  g2489 (n2529, n2476, n1015, n924, n1644);
nand g2490 (n2536, n1031, n1052, n1051);
and  g2491 (n2535, n1053, n924, n2519);
nor  g2492 (n2544, n2529, n2284, n2282, n2277);
or   g2493 (n2537, n2536, n2286, n973, n2280);
nor  g2494 (n2549, n2272, n2290, n2533, n2273);
nand g2495 (n2543, n2286, n2283, n2287, n2532);
xnor g2496 (n2552, n2394, n2281, n2397, n2534);
or   g2497 (n2547, n2275, n2278, n2289, n2271);
nor  g2498 (n2538, n2279, n2288, n2393, n2532);
xnor g2499 (n2539, n2281, n2276, n2535);
xnor g2500 (n2551, n2279, n2277, n973, n2534);
or   g2501 (n2540, n2282, n2536, n2392, n2531);
xor  g2502 (n2548, n2290, n2274, n2272, n2531);
or   g2503 (n2546, n2284, n2396, n2280, n2530);
nor  g2504 (n2542, n2289, n2288, n2395, n2287);
nand g2505 (n2541, n2285, n2529, n2273, n2274);
nor  g2506 (n2545, n2285, n2271, n2275, n2278);
nor  g2507 (n2550, n2530, n2533, n2283, n2535);
xor  g2508 (n2576, n2446, n2540, n2544, n2452);
xnor g2509 (n2562, n2551, n2428, n2430, n2548);
and  g2510 (n2573, n2418, n2444, n2542, n2420);
xor  g2511 (n2559, n2539, n2404, n2552, n2448);
and  g2512 (n2564, n2405, n2542, n2440, n2452);
xor  g2513 (n2565, n2444, n2436, n2417, n2410);
xnor g2514 (n2556, n2451, n2412, n2422, n2450);
xnor g2515 (n2572, n2449, n2428, n2437, n2540);
nor  g2516 (n2577, n2547, n2543, n2439, n2415);
and  g2517 (n2580, n2401, n2430, n2431, n2451);
nand g2518 (n2583, n2445, n2550, n2426, n2425);
or   g2519 (n2568, n2441, n2538, n2424, n2413);
xnor g2520 (n2579, n2450, n2408, n2411, n2399);
and  g2521 (n2563, n2543, n2435, n2551, n2446);
nor  g2522 (n2558, n2549, n2443, n2437, n2422);
xnor g2523 (n2554, n2416, n2546, n2442, n2420);
and  g2524 (n2578, n2429, n2545, n2447, n2441);
xnor g2525 (n2553, n2439, n2541, n2539, n2424);
or   g2526 (n2574, n2414, n2415, n2541, n2421);
or   g2527 (n2582, n2445, n2426, n2416, n2425);
and  g2528 (n2571, n2547, n2545, n2438, n2419);
xor  g2529 (n2584, n2537, n2447, n2433, n2436);
nand g2530 (n2561, n2449, n2412, n2423, n2442);
xnor g2531 (n2581, n2548, n2431, n2413, n2427);
nor  g2532 (n2566, n2421, n2432, n2418, n2414);
xor  g2533 (n2567, n2538, n2409, n2448, n2433);
nor  g2534 (n2560, n2423, n2427, n2440, n2398);
xnor g2535 (n2575, n2403, n2406, n2550, n2435);
and  g2536 (n2557, n2419, n2549, n2546, n2417);
xnor g2537 (n2570, n2432, n2438, n2402, n2434);
xnor g2538 (n2569, n2434, n2544, n2552, n2537);
and  g2539 (n2555, n2429, n2400, n2407, n2443);
endmodule
