// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_436 written by SynthGen on 2021/04/05 11:24:27
module Stat_3000_436( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n2746, n2898, n2901, n2902, n2897, n2911, n2910, n2914,
 n2917, n2979, n2992, n2988, n2997, n2993, n2999, n3000,
 n3004, n2998, n3001, n3003, n3022, n3027, n3024, n3032,
 n3029, n3030, n3023, n3025, n3021, n3031, n3028, n3026);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n2746, n2898, n2901, n2902, n2897, n2911, n2910, n2914,
 n2917, n2979, n2992, n2988, n2997, n2993, n2999, n3000,
 n3004, n2998, n3001, n3003, n3022, n3027, n3024, n3032,
 n3029, n3030, n3023, n3025, n3021, n3031, n3028, n3026;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
 n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
 n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
 n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
 n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
 n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
 n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
 n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
 n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
 n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
 n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
 n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
 n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
 n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
 n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
 n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
 n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
 n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
 n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
 n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
 n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
 n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
 n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
 n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
 n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
 n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
 n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
 n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
 n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
 n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
 n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
 n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
 n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
 n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
 n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
 n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
 n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
 n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
 n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
 n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
 n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
 n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
 n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
 n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
 n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
 n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
 n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
 n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
 n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
 n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
 n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
 n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
 n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
 n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
 n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
 n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
 n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
 n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
 n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
 n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
 n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
 n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
 n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
 n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
 n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
 n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
 n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
 n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
 n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
 n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
 n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
 n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
 n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
 n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
 n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
 n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
 n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
 n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
 n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
 n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
 n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
 n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
 n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
 n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
 n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
 n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
 n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
 n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
 n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
 n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
 n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
 n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
 n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
 n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
 n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
 n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
 n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
 n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
 n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
 n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
 n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
 n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
 n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
 n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
 n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
 n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
 n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
 n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
 n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
 n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
 n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
 n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
 n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
 n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
 n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
 n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
 n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
 n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
 n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
 n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
 n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
 n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
 n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
 n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
 n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
 n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
 n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
 n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
 n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
 n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
 n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
 n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
 n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
 n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
 n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
 n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
 n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
 n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
 n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
 n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
 n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
 n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
 n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
 n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
 n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
 n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
 n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
 n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
 n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
 n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
 n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
 n2745, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
 n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
 n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
 n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
 n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
 n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
 n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
 n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
 n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
 n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
 n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
 n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
 n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
 n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
 n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
 n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
 n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
 n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
 n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2899,
 n2900, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
 n2912, n2913, n2915, n2916, n2918, n2919, n2920, n2921,
 n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
 n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
 n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
 n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
 n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
 n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
 n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
 n2978, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
 n2987, n2989, n2990, n2991, n2994, n2995, n2996, n3002,
 n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
 n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020;

not  g0 (n140, n19);
buf  g1 (n117, n6);
buf  g2 (n100, n7);
buf  g3 (n111, n1);
not  g4 (n128, n11);
not  g5 (n132, n23);
buf  g6 (n41, n4);
not  g7 (n88, n20);
buf  g8 (n83, n17);
buf  g9 (n42, n14);
not  g10 (n110, n13);
buf  g11 (n102, n12);
not  g12 (n82, n16);
not  g13 (n142, n24);
buf  g14 (n54, n6);
not  g15 (n46, n17);
not  g16 (n47, n9);
not  g17 (n92, n13);
buf  g18 (n121, n25);
buf  g19 (n67, n32);
buf  g20 (n149, n11);
buf  g21 (n130, n19);
not  g22 (n72, n13);
not  g23 (n33, n29);
not  g24 (n157, n5);
not  g25 (n153, n16);
buf  g26 (n56, n23);
buf  g27 (n65, n19);
buf  g28 (n76, n3);
not  g29 (n40, n20);
buf  g30 (n118, n30);
buf  g31 (n91, n28);
buf  g32 (n107, n2);
buf  g33 (n95, n10);
not  g34 (n68, n15);
buf  g35 (n146, n16);
not  g36 (n66, n24);
not  g37 (n115, n30);
not  g38 (n77, n9);
not  g39 (n71, n26);
not  g40 (n138, n9);
not  g41 (n135, n5);
buf  g42 (n127, n8);
buf  g43 (n120, n28);
not  g44 (n155, n31);
not  g45 (n55, n28);
buf  g46 (n160, n32);
buf  g47 (n53, n31);
not  g48 (n38, n6);
not  g49 (n87, n20);
not  g50 (n35, n22);
buf  g51 (n106, n4);
buf  g52 (n80, n26);
not  g53 (n36, n8);
not  g54 (n156, n31);
buf  g55 (n133, n23);
buf  g56 (n109, n29);
buf  g57 (n62, n27);
buf  g58 (n86, n12);
buf  g59 (n113, n2);
not  g60 (n43, n2);
buf  g61 (n51, n10);
buf  g62 (n48, n3);
not  g63 (n143, n27);
not  g64 (n85, n18);
not  g65 (n134, n7);
buf  g66 (n159, n8);
not  g67 (n58, n6);
not  g68 (n94, n15);
not  g69 (n126, n17);
buf  g70 (n37, n18);
not  g71 (n57, n14);
not  g72 (n59, n32);
not  g73 (n108, n22);
buf  g74 (n103, n29);
buf  g75 (n63, n30);
buf  g76 (n70, n3);
buf  g77 (n52, n26);
buf  g78 (n122, n21);
not  g79 (n81, n3);
buf  g80 (n116, n17);
buf  g81 (n61, n1);
not  g82 (n124, n21);
not  g83 (n50, n32);
buf  g84 (n154, n22);
buf  g85 (n90, n22);
not  g86 (n98, n25);
buf  g87 (n69, n31);
buf  g88 (n125, n5);
not  g89 (n60, n11);
buf  g90 (n73, n21);
not  g91 (n151, n28);
not  g92 (n93, n26);
buf  g93 (n139, n7);
buf  g94 (n44, n2);
not  g95 (n64, n15);
not  g96 (n45, n24);
not  g97 (n39, n19);
not  g98 (n99, n1);
not  g99 (n97, n20);
not  g100 (n148, n1);
not  g101 (n129, n15);
buf  g102 (n101, n4);
buf  g103 (n96, n10);
not  g104 (n145, n16);
not  g105 (n150, n14);
buf  g106 (n89, n18);
buf  g107 (n105, n27);
not  g108 (n158, n9);
buf  g109 (n34, n14);
buf  g110 (n74, n23);
not  g111 (n136, n4);
buf  g112 (n147, n7);
buf  g113 (n137, n21);
buf  g114 (n79, n30);
buf  g115 (n119, n18);
not  g116 (n104, n12);
buf  g117 (n131, n24);
not  g118 (n152, n5);
not  g119 (n78, n12);
not  g120 (n112, n29);
not  g121 (n84, n8);
buf  g122 (n49, n25);
not  g123 (n114, n13);
not  g124 (n123, n25);
not  g125 (n144, n11);
buf  g126 (n75, n27);
not  g127 (n141, n10);
buf  g128 (n324, n89);
not  g129 (n350, n38);
buf  g130 (n222, n70);
buf  g131 (n413, n71);
buf  g132 (n617, n152);
buf  g133 (n548, n98);
buf  g134 (n655, n60);
not  g135 (n373, n153);
not  g136 (n492, n37);
not  g137 (n487, n82);
buf  g138 (n543, n66);
buf  g139 (n612, n55);
buf  g140 (n211, n68);
buf  g141 (n604, n88);
not  g142 (n316, n43);
not  g143 (n601, n148);
not  g144 (n508, n102);
buf  g145 (n255, n91);
not  g146 (n183, n142);
not  g147 (n459, n154);
buf  g148 (n639, n47);
not  g149 (n611, n147);
buf  g150 (n591, n79);
buf  g151 (n454, n126);
not  g152 (n257, n96);
not  g153 (n224, n111);
not  g154 (n565, n41);
buf  g155 (n615, n113);
not  g156 (n248, n96);
buf  g157 (n504, n140);
buf  g158 (n312, n57);
not  g159 (n481, n144);
not  g160 (n215, n68);
not  g161 (n243, n35);
not  g162 (n587, n155);
buf  g163 (n297, n136);
not  g164 (n456, n54);
not  g165 (n357, n52);
buf  g166 (n666, n41);
not  g167 (n621, n55);
buf  g168 (n438, n46);
not  g169 (n370, n125);
not  g170 (n506, n112);
buf  g171 (n630, n151);
not  g172 (n545, n127);
buf  g173 (n218, n124);
buf  g174 (n187, n54);
buf  g175 (n217, n135);
not  g176 (n397, n112);
buf  g177 (n237, n70);
buf  g178 (n606, n39);
not  g179 (n480, n123);
buf  g180 (n175, n123);
not  g181 (n529, n62);
not  g182 (n346, n109);
not  g183 (n194, n51);
not  g184 (n616, n116);
buf  g185 (n193, n83);
not  g186 (n245, n142);
buf  g187 (n633, n43);
buf  g188 (n625, n55);
not  g189 (n602, n134);
not  g190 (n582, n138);
not  g191 (n343, n93);
not  g192 (n528, n140);
buf  g193 (n323, n45);
buf  g194 (n540, n150);
buf  g195 (n605, n123);
not  g196 (n414, n80);
not  g197 (n272, n65);
buf  g198 (n399, n72);
buf  g199 (n198, n105);
not  g200 (n180, n59);
buf  g201 (n286, n118);
not  g202 (n599, n135);
not  g203 (n330, n83);
not  g204 (n433, n80);
buf  g205 (n518, n117);
buf  g206 (n573, n105);
not  g207 (n522, n81);
not  g208 (n331, n49);
buf  g209 (n184, n113);
not  g210 (n500, n35);
buf  g211 (n279, n53);
buf  g212 (n449, n59);
not  g213 (n620, n112);
buf  g214 (n539, n145);
buf  g215 (n364, n122);
not  g216 (n436, n82);
buf  g217 (n496, n102);
not  g218 (n319, n37);
buf  g219 (n420, n117);
buf  g220 (n260, n147);
buf  g221 (n670, n92);
buf  g222 (n253, n35);
buf  g223 (n483, n62);
not  g224 (n242, n146);
not  g225 (n661, n155);
buf  g226 (n585, n116);
not  g227 (n204, n44);
buf  g228 (n179, n158);
not  g229 (n645, n42);
buf  g230 (n419, n132);
not  g231 (n552, n128);
not  g232 (n473, n124);
buf  g233 (n344, n150);
buf  g234 (n556, n75);
not  g235 (n572, n105);
not  g236 (n246, n52);
not  g237 (n202, n130);
not  g238 (n327, n129);
buf  g239 (n287, n97);
not  g240 (n482, n146);
not  g241 (n486, n45);
buf  g242 (n668, n108);
not  g243 (n403, n56);
buf  g244 (n369, n58);
not  g245 (n443, n40);
buf  g246 (n186, n102);
not  g247 (n283, n94);
buf  g248 (n335, n86);
buf  g249 (n466, n128);
not  g250 (n295, n34);
not  g251 (n610, n99);
buf  g252 (n355, n155);
not  g253 (n376, n149);
buf  g254 (n244, n119);
not  g255 (n407, n41);
buf  g256 (n643, n71);
not  g257 (n538, n79);
not  g258 (n626, n125);
not  g259 (n411, n151);
buf  g260 (n226, n58);
buf  g261 (n519, n39);
buf  g262 (n447, n160);
not  g263 (n307, n158);
buf  g264 (n589, n54);
buf  g265 (n444, n34);
not  g266 (n448, n71);
buf  g267 (n329, n95);
not  g268 (n209, n131);
not  g269 (n471, n94);
not  g270 (n468, n118);
not  g271 (n490, n124);
buf  g272 (n195, n97);
buf  g273 (n306, n111);
not  g274 (n258, n109);
not  g275 (n635, n110);
not  g276 (n450, n153);
buf  g277 (n631, n59);
buf  g278 (n298, n100);
not  g279 (n168, n78);
buf  g280 (n304, n141);
buf  g281 (n374, n49);
not  g282 (n584, n79);
not  g283 (n446, n68);
not  g284 (n542, n47);
buf  g285 (n395, n43);
not  g286 (n555, n99);
not  g287 (n417, n84);
buf  g288 (n649, n40);
not  g289 (n416, n54);
buf  g290 (n356, n40);
not  g291 (n614, n33);
buf  g292 (n600, n117);
not  g293 (n619, n157);
buf  g294 (n234, n150);
not  g295 (n402, n56);
not  g296 (n644, n35);
not  g297 (n240, n66);
buf  g298 (n659, n63);
buf  g299 (n618, n72);
not  g300 (n557, n121);
buf  g301 (n284, n130);
not  g302 (n231, n46);
buf  g303 (n477, n43);
buf  g304 (n535, n85);
not  g305 (n568, n77);
buf  g306 (n465, n132);
buf  g307 (n185, n73);
not  g308 (n321, n70);
not  g309 (n250, n81);
buf  g310 (n200, n78);
buf  g311 (n230, n71);
buf  g312 (n415, n109);
buf  g313 (n391, n115);
not  g314 (n206, n57);
buf  g315 (n377, n66);
buf  g316 (n334, n131);
not  g317 (n652, n89);
buf  g318 (n362, n101);
not  g319 (n276, n152);
buf  g320 (n269, n84);
buf  g321 (n261, n73);
not  g322 (n654, n110);
not  g323 (n164, n136);
buf  g324 (n424, n38);
not  g325 (n282, n85);
not  g326 (n271, n108);
buf  g327 (n603, n135);
not  g328 (n241, n144);
buf  g329 (n384, n38);
buf  g330 (n262, n101);
buf  g331 (n278, n93);
not  g332 (n342, n49);
not  g333 (n580, n127);
buf  g334 (n537, n36);
not  g335 (n463, n77);
buf  g336 (n515, n84);
not  g337 (n317, n133);
buf  g338 (n340, n73);
buf  g339 (n484, n90);
buf  g340 (n190, n125);
buf  g341 (n267, n159);
buf  g342 (n623, n36);
buf  g343 (n351, n101);
not  g344 (n440, n87);
buf  g345 (n534, n145);
buf  g346 (n469, n95);
not  g347 (n553, n111);
buf  g348 (n220, n156);
not  g349 (n656, n130);
buf  g350 (n562, n120);
buf  g351 (n390, n58);
buf  g352 (n550, n99);
buf  g353 (n453, n134);
not  g354 (n434, n67);
buf  g355 (n285, n122);
buf  g356 (n409, n157);
not  g357 (n594, n37);
not  g358 (n396, n90);
not  g359 (n478, n73);
not  g360 (n634, n107);
not  g361 (n520, n92);
buf  g362 (n169, n45);
buf  g363 (n461, n158);
not  g364 (n646, n44);
not  g365 (n502, n90);
not  g366 (n341, n145);
not  g367 (n641, n64);
buf  g368 (n592, n131);
not  g369 (n583, n144);
not  g370 (n665, n128);
not  g371 (n406, n148);
buf  g372 (n642, n136);
buf  g373 (n208, n68);
buf  g374 (n577, n127);
buf  g375 (n299, n50);
not  g376 (n308, n139);
not  g377 (n638, n97);
not  g378 (n554, n46);
buf  g379 (n628, n132);
buf  g380 (n173, n87);
buf  g381 (n410, n57);
buf  g382 (n336, n159);
not  g383 (n613, n154);
not  g384 (n517, n46);
buf  g385 (n511, n84);
buf  g386 (n233, n38);
buf  g387 (n509, n129);
buf  g388 (n338, n50);
buf  g389 (n358, n155);
not  g390 (n445, n47);
not  g391 (n647, n156);
buf  g392 (n265, n107);
buf  g393 (n576, n76);
buf  g394 (n216, n101);
not  g395 (n212, n36);
not  g396 (n273, n138);
buf  g397 (n177, n91);
buf  g398 (n361, n115);
not  g399 (n266, n139);
not  g400 (n629, n81);
not  g401 (n162, n69);
buf  g402 (n219, n94);
buf  g403 (n203, n62);
buf  g404 (n228, n112);
buf  g405 (n663, n151);
not  g406 (n315, n102);
buf  g407 (n236, n131);
not  g408 (n525, n92);
buf  g409 (n401, n144);
buf  g410 (n232, n51);
buf  g411 (n288, n95);
not  g412 (n653, n143);
buf  g413 (n264, n122);
not  g414 (n326, n64);
not  g415 (n263, n78);
not  g416 (n404, n42);
not  g417 (n239, n134);
buf  g418 (n280, n48);
buf  g419 (n514, n139);
buf  g420 (n593, n119);
buf  g421 (n451, n61);
buf  g422 (n191, n44);
buf  g423 (n325, n88);
buf  g424 (n313, n110);
buf  g425 (n394, n85);
buf  g426 (n464, n119);
buf  g427 (n385, n69);
not  g428 (n167, n52);
buf  g429 (n381, n44);
not  g430 (n353, n140);
buf  g431 (n210, n141);
not  g432 (n598, n91);
not  g433 (n229, n50);
not  g434 (n435, n93);
buf  g435 (n339, n129);
buf  g436 (n165, n133);
buf  g437 (n441, n74);
not  g438 (n178, n148);
buf  g439 (n664, n42);
not  g440 (n170, n108);
buf  g441 (n268, n48);
buf  g442 (n379, n117);
not  g443 (n201, n119);
buf  g444 (n521, n67);
not  g445 (n457, n107);
buf  g446 (n491, n137);
buf  g447 (n328, n82);
buf  g448 (n259, n74);
buf  g449 (n371, n128);
buf  g450 (n530, n52);
buf  g451 (n305, n104);
buf  g452 (n505, n57);
buf  g453 (n488, n51);
not  g454 (n387, n45);
buf  g455 (n289, n72);
buf  g456 (n512, n116);
not  g457 (n181, n157);
not  g458 (n581, n114);
buf  g459 (n311, n85);
not  g460 (n662, n113);
not  g461 (n531, n124);
not  g462 (n254, n76);
buf  g463 (n205, n86);
buf  g464 (n588, n115);
not  g465 (n474, n121);
not  g466 (n207, n78);
buf  g467 (n393, n107);
buf  g468 (n274, n62);
buf  g469 (n561, n157);
buf  g470 (n493, n56);
buf  g471 (n418, n145);
buf  g472 (n345, n115);
buf  g473 (n475, n130);
buf  g474 (n526, n141);
buf  g475 (n292, n121);
not  g476 (n523, n63);
buf  g477 (n412, n126);
not  g478 (n536, n137);
not  g479 (n290, n103);
not  g480 (n388, n146);
buf  g481 (n349, n75);
buf  g482 (n546, n103);
buf  g483 (n503, n63);
buf  g484 (n174, n61);
not  g485 (n559, n122);
not  g486 (n352, n132);
not  g487 (n609, n59);
buf  g488 (n510, n123);
buf  g489 (n363, n106);
not  g490 (n197, n139);
not  g491 (n476, n120);
buf  g492 (n368, n99);
buf  g493 (n527, n153);
buf  g494 (n366, n90);
buf  g495 (n636, n74);
buf  g496 (n648, n51);
not  g497 (n354, n152);
buf  g498 (n541, n49);
buf  g499 (n651, n75);
buf  g500 (n564, n37);
not  g501 (n382, n135);
buf  g502 (n252, n113);
not  g503 (n558, n47);
not  g504 (n516, n104);
buf  g505 (n494, n118);
buf  g506 (n221, n69);
buf  g507 (n650, n149);
buf  g508 (n579, n147);
buf  g509 (n563, n76);
not  g510 (n256, n126);
not  g511 (n507, n156);
buf  g512 (n188, n88);
not  g513 (n189, n96);
buf  g514 (n172, n100);
not  g515 (n426, n118);
buf  g516 (n575, n105);
buf  g517 (n367, n98);
not  g518 (n199, n40);
buf  g519 (n551, n61);
not  g520 (n428, n156);
buf  g521 (n360, n100);
not  g522 (n405, n41);
not  g523 (n275, n138);
buf  g524 (n501, n114);
buf  g525 (n163, n42);
not  g526 (n247, n66);
not  g527 (n658, n120);
not  g528 (n607, n152);
not  g529 (n432, n53);
buf  g530 (n270, n143);
not  g531 (n337, n153);
not  g532 (n590, n106);
not  g533 (n608, n80);
not  g534 (n570, n91);
buf  g535 (n171, n56);
not  g536 (n458, n116);
buf  g537 (n431, n34);
not  g538 (n303, n79);
buf  g539 (n467, n65);
not  g540 (n348, n154);
not  g541 (n359, n106);
not  g542 (n567, n137);
not  g543 (n251, n76);
buf  g544 (n166, n158);
not  g545 (n657, n89);
not  g546 (n161, n74);
not  g547 (n301, n148);
buf  g548 (n566, n36);
not  g549 (n586, n97);
buf  g550 (n425, n109);
buf  g551 (n660, n98);
not  g552 (n322, n80);
not  g553 (n430, n100);
not  g554 (n495, n146);
buf  g555 (n227, n93);
not  g556 (n627, n114);
not  g557 (n365, n77);
buf  g558 (n213, n104);
buf  g559 (n533, n159);
not  g560 (n223, n149);
buf  g561 (n293, n39);
buf  g562 (n460, n82);
buf  g563 (n392, n147);
not  g564 (n439, n120);
buf  g565 (n225, n129);
buf  g566 (n176, n86);
not  g567 (n310, n55);
buf  g568 (n524, n142);
buf  g569 (n291, n111);
buf  g570 (n578, n60);
buf  g571 (n452, n87);
not  g572 (n571, n127);
buf  g573 (n235, n58);
buf  g574 (n442, n67);
not  g575 (n632, n141);
not  g576 (n498, n121);
buf  g577 (n302, n134);
buf  g578 (n427, n136);
not  g579 (n281, n48);
buf  g580 (n277, n140);
not  g581 (n637, n67);
buf  g582 (n622, n143);
buf  g583 (n596, n104);
not  g584 (n249, n126);
buf  g585 (n320, n72);
not  g586 (n408, n133);
not  g587 (n472, n86);
buf  g588 (n294, n103);
not  g589 (n489, n150);
not  g590 (n544, n87);
buf  g591 (n640, n64);
not  g592 (n375, n53);
buf  g593 (n574, n70);
not  g594 (n383, n88);
buf  g595 (n497, n50);
not  g596 (n547, n154);
buf  g597 (n455, n149);
not  g598 (n398, n77);
not  g599 (n479, n63);
not  g600 (n423, n81);
buf  g601 (n380, n65);
buf  g602 (n378, n114);
buf  g603 (n182, n106);
buf  g604 (n499, n33);
not  g605 (n196, n96);
buf  g606 (n192, n34);
not  g607 (n347, n159);
not  g608 (n624, n75);
not  g609 (n549, n83);
buf  g610 (n595, n64);
not  g611 (n296, n61);
not  g612 (n470, n133);
buf  g613 (n389, n98);
not  g614 (n214, n89);
buf  g615 (n667, n95);
not  g616 (n560, n137);
buf  g617 (n437, n39);
buf  g618 (n485, n103);
not  g619 (n462, n83);
not  g620 (n532, n110);
buf  g621 (n669, n160);
buf  g622 (n372, n151);
not  g623 (n400, n60);
not  g624 (n569, n33);
buf  g625 (n513, n60);
not  g626 (n386, n92);
not  g627 (n238, n69);
buf  g628 (n429, n138);
buf  g629 (n422, n143);
buf  g630 (n318, n142);
buf  g631 (n309, n94);
not  g632 (n314, n53);
not  g633 (n300, n48);
buf  g634 (n333, n125);
not  g635 (n597, n33);
not  g636 (n421, n65);
buf  g637 (n332, n108);
not  g638 (n1685, n489);
buf  g639 (n1613, n504);
buf  g640 (n868, n598);
not  g641 (n1854, n347);
not  g642 (n906, n447);
not  g643 (n2034, n599);
not  g644 (n845, n282);
buf  g645 (n770, n378);
not  g646 (n772, n394);
not  g647 (n2003, n355);
not  g648 (n1479, n489);
buf  g649 (n1572, n238);
buf  g650 (n1413, n584);
not  g651 (n1268, n665);
buf  g652 (n920, n243);
buf  g653 (n865, n402);
buf  g654 (n1954, n368);
buf  g655 (n1238, n175);
not  g656 (n690, n496);
buf  g657 (n1064, n628);
not  g658 (n1197, n349);
not  g659 (n1768, n312);
buf  g660 (n1510, n166);
not  g661 (n1323, n662);
buf  g662 (n1111, n460);
not  g663 (n2022, n481);
buf  g664 (n740, n589);
not  g665 (n981, n462);
not  g666 (n1467, n515);
not  g667 (n1407, n162);
not  g668 (n1624, n593);
buf  g669 (n1418, n456);
not  g670 (n1408, n306);
not  g671 (n753, n594);
not  g672 (n1899, n283);
not  g673 (n673, n181);
buf  g674 (n1020, n484);
not  g675 (n1426, n623);
buf  g676 (n875, n561);
buf  g677 (n998, n272);
buf  g678 (n1061, n576);
buf  g679 (n1599, n464);
buf  g680 (n1770, n619);
buf  g681 (n1511, n424);
not  g682 (n1481, n241);
not  g683 (n798, n447);
buf  g684 (n1777, n301);
buf  g685 (n688, n475);
buf  g686 (n1112, n341);
not  g687 (n1300, n440);
buf  g688 (n718, n614);
not  g689 (n1900, n248);
buf  g690 (n2056, n233);
not  g691 (n2057, n357);
buf  g692 (n1218, n221);
buf  g693 (n1556, n598);
not  g694 (n1366, n229);
not  g695 (n1384, n163);
buf  g696 (n1139, n171);
not  g697 (n1412, n459);
not  g698 (n1494, n570);
not  g699 (n1187, n250);
buf  g700 (n788, n404);
buf  g701 (n1944, n478);
not  g702 (n1231, n447);
not  g703 (n1387, n473);
not  g704 (n1049, n555);
buf  g705 (n2068, n551);
buf  g706 (n1847, n428);
not  g707 (n1441, n182);
not  g708 (n1639, n345);
not  g709 (n1918, n467);
not  g710 (n1881, n380);
buf  g711 (n1215, n161);
not  g712 (n1278, n235);
buf  g713 (n877, n565);
not  g714 (n1023, n511);
not  g715 (n1969, n355);
buf  g716 (n914, n465);
not  g717 (n844, n406);
not  g718 (n1839, n658);
buf  g719 (n1791, n437);
buf  g720 (n856, n488);
buf  g721 (n1836, n210);
buf  g722 (n803, n240);
buf  g723 (n1217, n222);
buf  g724 (n1505, n253);
not  g725 (n1739, n573);
not  g726 (n1107, n232);
buf  g727 (n1496, n644);
not  g728 (n1805, n266);
not  g729 (n797, n471);
not  g730 (n1234, n539);
buf  g731 (n1794, n616);
not  g732 (n2075, n218);
not  g733 (n1977, n230);
buf  g734 (n1228, n559);
not  g735 (n1573, n489);
not  g736 (n967, n237);
not  g737 (n1726, n554);
not  g738 (n702, n520);
not  g739 (n742, n555);
not  g740 (n1593, n469);
not  g741 (n1831, n285);
not  g742 (n1731, n548);
not  g743 (n1483, n282);
not  g744 (n1933, n402);
buf  g745 (n1178, n530);
buf  g746 (n1760, n589);
not  g747 (n795, n479);
not  g748 (n1611, n220);
buf  g749 (n1216, n439);
buf  g750 (n1955, n603);
buf  g751 (n961, n201);
buf  g752 (n1358, n220);
buf  g753 (n1751, n362);
not  g754 (n1406, n430);
not  g755 (n995, n662);
not  g756 (n1236, n486);
not  g757 (n1584, n610);
buf  g758 (n2058, n247);
buf  g759 (n1008, n496);
not  g760 (n1750, n544);
not  g761 (n1331, n512);
buf  g762 (n2074, n538);
not  g763 (n999, n555);
buf  g764 (n1605, n319);
not  g765 (n1273, n250);
buf  g766 (n1558, n499);
not  g767 (n942, n264);
not  g768 (n1834, n533);
buf  g769 (n983, n443);
not  g770 (n1263, n381);
not  g771 (n872, n252);
not  g772 (n769, n207);
not  g773 (n889, n185);
not  g774 (n1783, n389);
not  g775 (n1184, n312);
buf  g776 (n1206, n414);
not  g777 (n1676, n333);
not  g778 (n1893, n471);
buf  g779 (n1198, n214);
not  g780 (n1142, n586);
buf  g781 (n1655, n374);
buf  g782 (n1269, n634);
not  g783 (n1041, n176);
buf  g784 (n963, n351);
buf  g785 (n2044, n581);
buf  g786 (n1801, n344);
not  g787 (n1080, n339);
not  g788 (n1724, n509);
buf  g789 (n902, n452);
not  g790 (n1083, n392);
not  g791 (n1381, n283);
buf  g792 (n750, n274);
buf  g793 (n1361, n480);
buf  g794 (n1934, n525);
buf  g795 (n804, n213);
not  g796 (n2048, n451);
buf  g797 (n1473, n405);
buf  g798 (n760, n566);
not  g799 (n1488, n556);
buf  g800 (n2039, n272);
not  g801 (n1594, n171);
not  g802 (n1745, n408);
buf  g803 (n1811, n232);
not  g804 (n956, n625);
not  g805 (n775, n586);
not  g806 (n1424, n291);
not  g807 (n2077, n393);
not  g808 (n1249, n476);
not  g809 (n1815, n343);
buf  g810 (n764, n590);
not  g811 (n936, n612);
buf  g812 (n930, n596);
not  g813 (n1964, n499);
buf  g814 (n1932, n635);
not  g815 (n1749, n167);
buf  g816 (n1545, n177);
not  g817 (n1043, n398);
not  g818 (n1019, n195);
not  g819 (n1290, n251);
buf  g820 (n1714, n412);
buf  g821 (n1247, n445);
not  g822 (n1264, n307);
not  g823 (n1525, n382);
not  g824 (n900, n563);
not  g825 (n736, n334);
buf  g826 (n1260, n231);
buf  g827 (n1705, n595);
buf  g828 (n1501, n354);
not  g829 (n1179, n591);
buf  g830 (n689, n462);
not  g831 (n825, n238);
not  g832 (n782, n446);
buf  g833 (n1856, n388);
buf  g834 (n1255, n445);
buf  g835 (n1102, n547);
not  g836 (n1118, n602);
buf  g837 (n980, n227);
not  g838 (n1324, n646);
buf  g839 (n1938, n216);
buf  g840 (n1988, n437);
buf  g841 (n1096, n579);
not  g842 (n705, n554);
buf  g843 (n1258, n517);
not  g844 (n1981, n254);
buf  g845 (n1844, n359);
not  g846 (n1671, n434);
buf  g847 (n1892, n317);
not  g848 (n784, n567);
not  g849 (n1972, n592);
not  g850 (n1310, n400);
not  g851 (n982, n192);
buf  g852 (n977, n646);
not  g853 (n1493, n650);
buf  g854 (n1338, n433);
buf  g855 (n1031, n336);
buf  g856 (n1209, n426);
buf  g857 (n916, n607);
buf  g858 (n1992, n282);
not  g859 (n717, n299);
buf  g860 (n1151, n411);
buf  g861 (n1070, n593);
not  g862 (n974, n269);
buf  g863 (n1207, n333);
buf  g864 (n2011, n585);
not  g865 (n1033, n416);
not  g866 (n1549, n197);
not  g867 (n1298, n308);
buf  g868 (n1194, n321);
not  g869 (n1251, n628);
not  g870 (n996, n333);
not  g871 (n852, n639);
not  g872 (n1502, n275);
not  g873 (n1073, n626);
buf  g874 (n1636, n574);
buf  g875 (n1653, n466);
not  g876 (n976, n253);
buf  g877 (n2019, n206);
not  g878 (n1528, n281);
buf  g879 (n1245, n491);
buf  g880 (n921, n633);
not  g881 (n1451, n393);
buf  g882 (n1474, n399);
buf  g883 (n1166, n382);
not  g884 (n683, n479);
buf  g885 (n1414, n434);
buf  g886 (n1617, n423);
not  g887 (n1641, n381);
buf  g888 (n1845, n581);
buf  g889 (n732, n262);
buf  g890 (n824, n474);
not  g891 (n722, n441);
buf  g892 (n1240, n420);
buf  g893 (n932, n556);
not  g894 (n789, n403);
buf  g895 (n1926, n594);
buf  g896 (n1094, n261);
buf  g897 (n1442, n431);
buf  g898 (n1165, n242);
not  g899 (n1663, n664);
buf  g900 (n846, n470);
not  g901 (n1156, n173);
buf  g902 (n878, n329);
not  g903 (n1660, n299);
not  g904 (n978, n548);
not  g905 (n1335, n532);
buf  g906 (n1861, n419);
buf  g907 (n1914, n260);
not  g908 (n1349, n601);
not  g909 (n1767, n226);
buf  g910 (n699, n593);
buf  g911 (n2067, n324);
not  g912 (n1723, n331);
buf  g913 (n1769, n369);
buf  g914 (n1512, n233);
buf  g915 (n1293, n583);
buf  g916 (n1065, n247);
not  g917 (n909, n347);
buf  g918 (n1633, n270);
not  g919 (n1984, n466);
buf  g920 (n1646, n272);
not  g921 (n1321, n513);
not  g922 (n1146, n613);
buf  g923 (n2055, n528);
not  g924 (n1021, n662);
buf  g925 (n1476, n348);
buf  g926 (n1687, n306);
not  g927 (n1145, n374);
buf  g928 (n1703, n402);
buf  g929 (n1379, n477);
not  g930 (n1725, n278);
buf  g931 (n1202, n433);
buf  g932 (n1686, n652);
not  g933 (n1138, n169);
not  g934 (n1508, n564);
buf  g935 (n919, n429);
buf  g936 (n743, n498);
buf  g937 (n1322, n247);
not  g938 (n1105, n501);
not  g939 (n1224, n418);
not  g940 (n1009, n562);
buf  g941 (n1109, n511);
not  g942 (n1896, n197);
not  g943 (n1911, n164);
buf  g944 (n1532, n283);
not  g945 (n678, n496);
buf  g946 (n1128, n194);
not  g947 (n870, n541);
buf  g948 (n1882, n624);
buf  g949 (n2043, n628);
not  g950 (n1889, n425);
not  g951 (n1339, n576);
buf  g952 (n1588, n600);
buf  g953 (n1318, n194);
buf  g954 (n1223, n476);
buf  g955 (n1312, n414);
buf  g956 (n1905, n525);
buf  g957 (n1658, n403);
buf  g958 (n783, n590);
buf  g959 (n1484, n503);
not  g960 (n858, n493);
not  g961 (n1780, n548);
not  g962 (n1086, n398);
not  g963 (n693, n529);
buf  g964 (n2047, n580);
not  g965 (n1566, n343);
buf  g966 (n968, n444);
buf  g967 (n1272, n311);
not  g968 (n1662, n523);
buf  g969 (n1182, n359);
not  g970 (n1776, n329);
not  g971 (n1454, n259);
buf  g972 (n1652, n457);
buf  g973 (n1014, n394);
not  g974 (n1855, n415);
buf  g975 (n720, n356);
not  g976 (n1159, n582);
buf  g977 (n1849, n538);
not  g978 (n757, n336);
not  g979 (n1059, n567);
not  g980 (n1616, n296);
buf  g981 (n786, n457);
not  g982 (n1922, n174);
not  g983 (n1325, n551);
not  g984 (n1468, n215);
buf  g985 (n1066, n186);
buf  g986 (n1492, n420);
not  g987 (n1553, n586);
not  g988 (n954, n626);
not  g989 (n989, n216);
not  g990 (n1623, n351);
buf  g991 (n990, n405);
not  g992 (n1005, n506);
not  g993 (n1125, n435);
not  g994 (n1087, n516);
buf  g995 (n840, n595);
not  g996 (n927, n360);
buf  g997 (n1656, n621);
not  g998 (n946, n240);
buf  g999 (n1742, n386);
buf  g1000 (n2009, n553);
not  g1001 (n1910, n415);
buf  g1002 (n2021, n369);
not  g1003 (n1256, n303);
buf  g1004 (n2030, n307);
buf  g1005 (n1574, n445);
buf  g1006 (n1500, n330);
buf  g1007 (n1946, n619);
buf  g1008 (n2020, n665);
buf  g1009 (n1542, n474);
buf  g1010 (n1482, n484);
buf  g1011 (n1036, n423);
buf  g1012 (n787, n239);
buf  g1013 (n1581, n334);
not  g1014 (n1945, n261);
not  g1015 (n1632, n178);
buf  g1016 (n1504, n399);
not  g1017 (n1174, n191);
not  g1018 (n1190, n603);
buf  g1019 (n1894, n563);
not  g1020 (n894, n224);
not  g1021 (n1610, n282);
not  g1022 (n895, n512);
not  g1023 (n2005, n520);
not  g1024 (n1060, n305);
not  g1025 (n2051, n372);
buf  g1026 (n2061, n376);
buf  g1027 (n1679, n385);
buf  g1028 (n1093, n186);
buf  g1029 (n1962, n449);
not  g1030 (n1943, n638);
buf  g1031 (n1620, n590);
not  g1032 (n765, n256);
not  g1033 (n1316, n550);
buf  g1034 (n1498, n243);
not  g1035 (n1003, n667);
not  g1036 (n1051, n221);
not  g1037 (n1092, n163);
not  g1038 (n1570, n310);
not  g1039 (n721, n229);
buf  g1040 (n1434, n370);
not  g1041 (n1692, n205);
not  g1042 (n1503, n510);
not  g1043 (n1852, n513);
not  g1044 (n1044, n413);
buf  g1045 (n1579, n450);
buf  g1046 (n1600, n277);
buf  g1047 (n2013, n427);
not  g1048 (n1898, n175);
not  g1049 (n1078, n308);
not  g1050 (n1615, n270);
not  g1051 (n1459, n170);
buf  g1052 (n1718, n371);
not  g1053 (n973, n479);
buf  g1054 (n869, n390);
buf  g1055 (n848, n241);
buf  g1056 (n1773, n410);
not  g1057 (n1432, n536);
buf  g1058 (n1763, n584);
not  g1059 (n1651, n530);
not  g1060 (n965, n493);
not  g1061 (n1698, n508);
not  g1062 (n1930, n234);
buf  g1063 (n1239, n214);
buf  g1064 (n1333, n435);
not  g1065 (n1784, n459);
not  g1066 (n1526, n300);
buf  g1067 (n1114, n209);
not  g1068 (n859, n552);
buf  g1069 (n1229, n489);
buf  g1070 (n2018, n407);
not  g1071 (n1989, n180);
not  g1072 (n1135, n485);
not  g1073 (n862, n579);
not  g1074 (n821, n423);
not  g1075 (n679, n548);
buf  g1076 (n1567, n636);
not  g1077 (n1495, n330);
buf  g1078 (n1666, n656);
not  g1079 (n1004, n350);
not  g1080 (n843, n497);
not  g1081 (n1365, n645);
buf  g1082 (n1439, n213);
buf  g1083 (n1822, n388);
not  g1084 (n1226, n604);
not  g1085 (n1524, n256);
not  g1086 (n2006, n373);
buf  g1087 (n2014, n355);
not  g1088 (n1916, n569);
buf  g1089 (n1039, n369);
buf  g1090 (n1643, n366);
buf  g1091 (n1865, n311);
not  g1092 (n794, n516);
buf  g1093 (n1927, n200);
buf  g1094 (n1377, n503);
not  g1095 (n1735, n524);
buf  g1096 (n1035, n467);
not  g1097 (n1765, n609);
buf  g1098 (n1047, n448);
buf  g1099 (n1193, n430);
buf  g1100 (n1688, n531);
buf  g1101 (n880, n579);
not  g1102 (n1411, n421);
not  g1103 (n1848, n421);
buf  g1104 (n767, n577);
not  g1105 (n1609, n640);
not  g1106 (n1562, n305);
buf  g1107 (n1967, n434);
buf  g1108 (n1995, n235);
buf  g1109 (n807, n370);
not  g1110 (n922, n389);
not  g1111 (n1888, n276);
buf  g1112 (n1982, n398);
not  g1113 (n1824, n635);
buf  g1114 (n1704, n190);
buf  g1115 (n1909, n249);
buf  g1116 (n749, n398);
buf  g1117 (n1436, n234);
not  g1118 (n1957, n316);
buf  g1119 (n1953, n325);
not  g1120 (n1397, n582);
buf  g1121 (n1211, n577);
not  g1122 (n1912, n622);
buf  g1123 (n1798, n234);
buf  g1124 (n992, n557);
not  g1125 (n1961, n386);
not  g1126 (n2002, n361);
not  g1127 (n1531, n166);
buf  g1128 (n759, n410);
not  g1129 (n1160, n339);
not  g1130 (n1376, n309);
not  g1131 (n1947, n664);
not  g1132 (n1552, n396);
not  g1133 (n836, n570);
not  g1134 (n882, n631);
buf  g1135 (n1425, n358);
not  g1136 (n1752, n375);
buf  g1137 (n704, n404);
buf  g1138 (n1359, n582);
buf  g1139 (n984, n257);
buf  g1140 (n827, n337);
buf  g1141 (n898, n553);
buf  g1142 (n1604, n655);
not  g1143 (n680, n224);
not  g1144 (n1877, n241);
buf  g1145 (n1821, n433);
buf  g1146 (n1172, n345);
buf  g1147 (n1429, n244);
not  g1148 (n1176, n442);
buf  g1149 (n993, n556);
not  g1150 (n1121, n558);
buf  g1151 (n1627, n350);
buf  g1152 (n1998, n560);
buf  g1153 (n1281, n254);
buf  g1154 (n1991, n163);
buf  g1155 (n913, n338);
not  g1156 (n896, n522);
buf  g1157 (n1191, n618);
buf  g1158 (n1748, n268);
buf  g1159 (n1431, n363);
buf  g1160 (n1097, n606);
buf  g1161 (n1284, n180);
buf  g1162 (n1013, n335);
buf  g1163 (n711, n435);
not  g1164 (n708, n180);
not  g1165 (n1607, n395);
buf  g1166 (n1419, n416);
buf  g1167 (n1591, n376);
buf  g1168 (n1219, n552);
not  g1169 (n1979, n565);
not  g1170 (n957, n647);
buf  g1171 (n1903, n342);
not  g1172 (n1618, n294);
buf  g1173 (n1410, n275);
not  g1174 (n793, n191);
buf  g1175 (n1010, n526);
not  g1176 (n861, n209);
not  g1177 (n1313, n320);
not  g1178 (n1997, n255);
not  g1179 (n1277, n285);
buf  g1180 (n1443, n165);
not  g1181 (n1522, n601);
not  g1182 (n1650, n309);
not  g1183 (n1106, n594);
buf  g1184 (n805, n301);
not  g1185 (n1022, n611);
not  g1186 (n2023, n292);
not  g1187 (n731, n379);
buf  g1188 (n1818, n325);
not  g1189 (n1129, n512);
buf  g1190 (n1983, n615);
not  g1191 (n785, n267);
not  g1192 (n1056, n390);
not  g1193 (n1233, n485);
not  g1194 (n1832, n173);
buf  g1195 (n1067, n213);
not  g1196 (n812, n387);
not  g1197 (n1843, n260);
not  g1198 (n2073, n420);
buf  g1199 (n1416, n177);
buf  g1200 (n1630, n337);
not  g1201 (n1344, n296);
not  g1202 (n745, n626);
not  g1203 (n1544, n167);
buf  g1204 (n796, n353);
buf  g1205 (n2008, n472);
not  g1206 (n1555, n492);
not  g1207 (n1052, n176);
buf  g1208 (n1948, n171);
buf  g1209 (n908, n556);
buf  g1210 (n1779, n561);
not  g1211 (n1701, n265);
not  g1212 (n1375, n235);
not  g1213 (n747, n318);
buf  g1214 (n1354, n490);
buf  g1215 (n1405, n280);
buf  g1216 (n1450, n550);
buf  g1217 (n1634, n372);
not  g1218 (n1876, n374);
buf  g1219 (n737, n226);
buf  g1220 (n1587, n166);
not  g1221 (n867, n383);
buf  g1222 (n1833, n524);
not  g1223 (n1485, n189);
not  g1224 (n1668, n452);
not  g1225 (n1864, n401);
not  g1226 (n864, n181);
not  g1227 (n776, n455);
not  g1228 (n1382, n499);
buf  g1229 (n1858, n440);
buf  g1230 (n1458, n587);
buf  g1231 (n1314, n334);
buf  g1232 (n1385, n278);
buf  g1233 (n1140, n634);
buf  g1234 (n1472, n271);
buf  g1235 (n1243, n421);
buf  g1236 (n1422, n376);
not  g1237 (n1355, n174);
not  g1238 (n1951, n637);
buf  g1239 (n1559, n555);
buf  g1240 (n1601, n248);
not  g1241 (n1068, n474);
not  g1242 (n1744, n274);
buf  g1243 (n873, n510);
not  g1244 (n1551, n592);
buf  g1245 (n2050, n335);
buf  g1246 (n1994, n558);
buf  g1247 (n1754, n185);
buf  g1248 (n1654, n656);
not  g1249 (n1402, n390);
buf  g1250 (n710, n190);
buf  g1251 (n2041, n632);
not  g1252 (n1799, n661);
not  g1253 (n685, n400);
buf  g1254 (n1282, n515);
not  g1255 (n834, n202);
buf  g1256 (n815, n457);
buf  g1257 (n1444, n389);
buf  g1258 (n910, n468);
not  g1259 (n1115, n449);
buf  g1260 (n881, n589);
not  g1261 (n1840, n259);
not  g1262 (n1965, n610);
buf  g1263 (n818, n338);
not  g1264 (n1403, n575);
not  g1265 (n1716, n647);
buf  g1266 (n1842, n600);
buf  g1267 (n726, n592);
not  g1268 (n929, n225);
not  g1269 (n768, n193);
buf  g1270 (n1734, n232);
not  g1271 (n888, n200);
not  g1272 (n1262, n219);
not  g1273 (n819, n627);
buf  g1274 (n1200, n474);
not  g1275 (n1225, n487);
buf  g1276 (n1347, n498);
not  g1277 (n1210, n514);
not  g1278 (n814, n289);
not  g1279 (n1756, n230);
buf  g1280 (n1732, n207);
not  g1281 (n780, n239);
not  g1282 (n1917, n161);
buf  g1283 (n1571, n616);
buf  g1284 (n1875, n667);
buf  g1285 (n1682, n294);
not  g1286 (n2004, n252);
buf  g1287 (n1259, n580);
buf  g1288 (n951, n549);
buf  g1289 (n1672, n315);
buf  g1290 (n1328, n317);
not  g1291 (n1370, n184);
buf  g1292 (n700, n524);
not  g1293 (n1058, n409);
not  g1294 (n1857, n463);
buf  g1295 (n1885, n464);
buf  g1296 (n1072, n306);
not  g1297 (n1133, n572);
not  g1298 (n917, n467);
buf  g1299 (n972, n466);
not  g1300 (n701, n417);
buf  g1301 (n1006, n462);
not  g1302 (n2012, n495);
not  g1303 (n950, n628);
buf  g1304 (n1235, n254);
not  g1305 (n730, n186);
buf  g1306 (n692, n379);
buf  g1307 (n1890, n539);
not  g1308 (n1490, n236);
buf  g1309 (n1212, n193);
not  g1310 (n1862, n553);
not  g1311 (n1527, n167);
not  g1312 (n1960, n363);
not  g1313 (n733, n179);
not  g1314 (n1790, n446);
not  g1315 (n2025, n544);
buf  g1316 (n1012, n414);
not  g1317 (n1461, n368);
not  g1318 (n1936, n395);
buf  g1319 (n1608, n395);
buf  g1320 (n1149, n273);
not  g1321 (n1395, n216);
buf  g1322 (n2060, n210);
not  g1323 (n1188, n416);
buf  g1324 (n1635, n242);
buf  g1325 (n1986, n203);
buf  g1326 (n1283, n173);
buf  g1327 (n903, n441);
not  g1328 (n1901, n592);
not  g1329 (n1887, n186);
not  g1330 (n2080, n259);
not  g1331 (n1099, n448);
buf  g1332 (n863, n521);
buf  g1333 (n2071, n408);
not  g1334 (n1778, n586);
buf  g1335 (n1812, n320);
not  g1336 (n817, n422);
not  g1337 (n1167, n162);
buf  g1338 (n1536, n244);
buf  g1339 (n1781, n287);
buf  g1340 (n1683, n531);
buf  g1341 (n1017, n179);
not  g1342 (n766, n289);
not  g1343 (n727, n647);
not  g1344 (n949, n293);
buf  g1345 (n801, n534);
not  g1346 (n1680, n274);
not  g1347 (n728, n477);
not  g1348 (n891, n570);
buf  g1349 (n2033, n524);
not  g1350 (n1122, n599);
not  g1351 (n1437, n343);
buf  g1352 (n744, n311);
not  g1353 (n1809, n482);
buf  g1354 (n970, n281);
not  g1355 (n1457, n296);
buf  g1356 (n1180, n302);
not  g1357 (n1759, n388);
not  g1358 (n1372, n215);
buf  g1359 (n833, n618);
buf  g1360 (n1192, n620);
not  g1361 (n991, n490);
buf  g1362 (n1973, n315);
buf  g1363 (n1048, n507);
not  g1364 (n1806, n615);
buf  g1365 (n735, n533);
buf  g1366 (n1557, n249);
not  g1367 (n1817, n331);
buf  g1368 (n1203, n607);
buf  g1369 (n707, n472);
buf  g1370 (n1730, n469);
not  g1371 (n1913, n545);
not  g1372 (n1694, n535);
buf  g1373 (n773, n211);
buf  g1374 (n1874, n561);
buf  g1375 (n1038, n375);
not  g1376 (n1647, n657);
not  g1377 (n1221, n660);
not  g1378 (n1378, n320);
not  g1379 (n781, n624);
buf  g1380 (n1371, n530);
not  g1381 (n966, n597);
buf  g1382 (n1100, n652);
not  g1383 (n1438, n629);
not  g1384 (n1626, n417);
buf  g1385 (n2049, n242);
not  g1386 (n1137, n228);
not  g1387 (n676, n478);
buf  g1388 (n1007, n173);
not  g1389 (n1873, n204);
buf  g1390 (n1353, n588);
not  g1391 (n1449, n318);
not  g1392 (n1155, n529);
not  g1393 (n854, n608);
not  g1394 (n1808, n616);
buf  g1395 (n1391, n564);
buf  g1396 (n987, n476);
buf  g1397 (n897, n323);
buf  g1398 (n1923, n166);
buf  g1399 (n1356, n559);
not  g1400 (n1119, n432);
not  g1401 (n1028, n461);
buf  g1402 (n811, n515);
not  g1403 (n1315, n507);
not  g1404 (n850, n640);
not  g1405 (n1537, n455);
buf  g1406 (n1404, n367);
buf  g1407 (n1090, n401);
not  g1408 (n1538, n324);
not  g1409 (n1421, n470);
not  g1410 (n1880, n165);
buf  g1411 (n1351, n505);
buf  g1412 (n1000, n578);
buf  g1413 (n1002, n554);
not  g1414 (n1669, n618);
not  g1415 (n841, n385);
buf  g1416 (n986, n617);
not  g1417 (n1563, n450);
buf  g1418 (n694, n645);
buf  g1419 (n1838, n381);
not  g1420 (n1295, n208);
buf  g1421 (n1810, n613);
not  g1422 (n1860, n483);
not  g1423 (n1026, n529);
buf  g1424 (n1175, n578);
buf  g1425 (n2029, n229);
buf  g1426 (n779, n325);
buf  g1427 (n1925, n311);
not  g1428 (n1303, n514);
not  g1429 (n1539, n483);
buf  g1430 (n1173, n350);
not  g1431 (n1758, n400);
buf  g1432 (n1398, n268);
buf  g1433 (n696, n304);
not  g1434 (n1866, n542);
not  g1435 (n1564, n610);
not  g1436 (n1161, n588);
not  g1437 (n1879, n604);
not  g1438 (n1774, n452);
not  g1439 (n1241, n364);
buf  g1440 (n1183, n503);
not  g1441 (n1132, n292);
buf  g1442 (n1389, n636);
not  g1443 (n1786, n578);
not  g1444 (n1428, n207);
buf  g1445 (n2079, n596);
buf  g1446 (n1050, n632);
buf  g1447 (n1867, n290);
not  g1448 (n876, n345);
not  g1449 (n1025, n643);
not  g1450 (n1162, n503);
buf  g1451 (n1757, n492);
not  g1452 (n738, n651);
not  g1453 (n1738, n319);
not  g1454 (n1851, n559);
not  g1455 (n1795, n487);
buf  g1456 (n923, n621);
buf  g1457 (n1469, n225);
buf  g1458 (n762, n304);
buf  g1459 (n945, n169);
buf  g1460 (n1733, n428);
buf  g1461 (n802, n453);
buf  g1462 (n1939, n494);
buf  g1463 (n1996, n368);
buf  g1464 (n1814, n570);
not  g1465 (n1603, n336);
buf  g1466 (n1069, n189);
buf  g1467 (n1782, n638);
buf  g1468 (n800, n338);
not  g1469 (n2028, n546);
buf  g1470 (n1227, n625);
not  g1471 (n1045, n636);
buf  g1472 (n1276, n196);
not  g1473 (n1362, n554);
buf  g1474 (n1707, n514);
buf  g1475 (n1924, n501);
not  g1476 (n1576, n568);
not  g1477 (n1301, n273);
buf  g1478 (n1435, n540);
buf  g1479 (n1829, n406);
buf  g1480 (n1163, n528);
not  g1481 (n890, n364);
buf  g1482 (n697, n203);
not  g1483 (n1706, n493);
buf  g1484 (n1237, n492);
not  g1485 (n1506, n438);
not  g1486 (n1124, n426);
buf  g1487 (n1150, n647);
not  g1488 (n1329, n409);
buf  g1489 (n1642, n178);
not  g1490 (n1091, n310);
buf  g1491 (n1736, n223);
buf  g1492 (n1185, n284);
not  g1493 (n1596, n536);
not  g1494 (n1001, n526);
not  g1495 (n1702, n225);
buf  g1496 (n962, n563);
buf  g1497 (n1959, n660);
not  g1498 (n2031, n509);
buf  g1499 (n1569, n597);
not  g1500 (n1602, n418);
not  g1501 (n1326, n425);
not  g1502 (n1648, n552);
buf  g1503 (n1775, n477);
buf  g1504 (n810, n574);
not  g1505 (n758, n522);
buf  g1506 (n1720, n559);
not  g1507 (n1835, n543);
buf  g1508 (n1568, n384);
buf  g1509 (n2076, n468);
buf  g1510 (n791, n256);
not  g1511 (n1394, n227);
not  g1512 (n1684, n342);
not  g1513 (n925, n382);
not  g1514 (n1327, n380);
not  g1515 (n935, n436);
not  g1516 (n682, n293);
buf  g1517 (n1015, n277);
not  g1518 (n1016, n490);
buf  g1519 (n1690, n275);
not  g1520 (n1621, n660);
not  g1521 (n1561, n191);
buf  g1522 (n837, n298);
not  g1523 (n1116, n309);
buf  g1524 (n1158, n415);
not  g1525 (n755, n377);
not  g1526 (n1027, n392);
buf  g1527 (n1089, n641);
buf  g1528 (n1740, n609);
buf  g1529 (n964, n506);
buf  g1530 (n2064, n433);
buf  g1531 (n1470, n446);
buf  g1532 (n1540, n659);
not  g1533 (n1638, n529);
buf  g1534 (n774, n360);
not  g1535 (n1940, n294);
buf  g1536 (n1334, n228);
buf  g1537 (n1677, n313);
not  g1538 (n1393, n659);
buf  g1539 (n1606, n204);
buf  g1540 (n1071, n422);
buf  g1541 (n1440, n356);
not  g1542 (n1110, n396);
not  g1543 (n1053, n346);
buf  g1544 (n911, n290);
not  g1545 (n1336, n567);
not  g1546 (n1074, n312);
buf  g1547 (n958, n587);
buf  g1548 (n1637, n589);
buf  g1549 (n1796, n520);
not  g1550 (n1816, n665);
not  g1551 (n1085, n536);
not  g1552 (n1287, n238);
buf  g1553 (n1550, n546);
not  g1554 (n1950, n252);
not  g1555 (n887, n611);
not  g1556 (n1521, n653);
not  g1557 (n1827, n162);
buf  g1558 (n835, n450);
buf  g1559 (n1120, n361);
not  g1560 (n1266, n257);
not  g1561 (n1063, n284);
buf  g1562 (n1034, n208);
not  g1563 (n1659, n622);
not  g1564 (n1299, n291);
not  g1565 (n1374, n491);
not  g1566 (n893, n461);
not  g1567 (n1583, n170);
buf  g1568 (n1456, n513);
not  g1569 (n1380, n533);
buf  g1570 (n1697, n516);
not  g1571 (n1657, n393);
buf  g1572 (n1722, n432);
buf  g1573 (n1915, n654);
not  g1574 (n672, n206);
not  g1575 (n1878, n608);
buf  g1576 (n1352, n631);
buf  g1577 (n741, n624);
buf  g1578 (n1471, n169);
not  g1579 (n1148, n188);
not  g1580 (n1220, n643);
buf  g1581 (n1895, n521);
not  g1582 (n1076, n517);
not  g1583 (n1970, n572);
buf  g1584 (n1291, n217);
not  g1585 (n871, n223);
buf  g1586 (n1465, n530);
not  g1587 (n1153, n397);
buf  g1588 (n1242, n168);
buf  g1589 (n1168, n567);
buf  g1590 (n1622, n593);
not  g1591 (n2063, n537);
not  g1592 (n1800, n377);
not  g1593 (n687, n300);
buf  g1594 (n2035, n342);
buf  g1595 (n1535, n517);
not  g1596 (n1279, n324);
not  g1597 (n828, n631);
not  g1598 (n1755, n341);
buf  g1599 (n754, n657);
not  g1600 (n1708, n490);
buf  g1601 (n1304, n581);
buf  g1602 (n1075, n499);
buf  g1603 (n763, n418);
not  g1604 (n1307, n526);
not  g1605 (n790, n557);
not  g1606 (n886, n537);
buf  g1607 (n1595, n505);
not  g1608 (n831, n480);
buf  g1609 (n2066, n473);
buf  g1610 (n1937, n203);
not  g1611 (n1828, n346);
not  g1612 (n1244, n557);
buf  g1613 (n1853, n437);
not  g1614 (n1369, n436);
not  g1615 (n809, n353);
buf  g1616 (n1871, n502);
not  g1617 (n2024, n179);
not  g1618 (n1024, n215);
not  g1619 (n1213, n243);
not  g1620 (n874, n417);
not  g1621 (n1409, n336);
not  g1622 (n1364, n365);
not  g1623 (n1143, n510);
buf  g1624 (n847, n477);
not  g1625 (n1448, n223);
not  g1626 (n2001, n376);
buf  g1627 (n905, n488);
not  g1628 (n813, n604);
not  g1629 (n725, n361);
not  g1630 (n1181, n302);
not  g1631 (n778, n303);
not  g1632 (n684, n651);
not  g1633 (n988, n480);
not  g1634 (n1113, n357);
buf  g1635 (n1518, n194);
not  g1636 (n1079, n378);
buf  g1637 (n1383, n206);
not  g1638 (n1747, n369);
buf  g1639 (n1597, n285);
not  g1640 (n1098, n179);
not  g1641 (n1399, n224);
buf  g1642 (n1330, n233);
buf  g1643 (n960, n643);
buf  g1644 (n1921, n663);
not  g1645 (n1396, n448);
not  g1646 (n729, n268);
not  g1647 (n947, n347);
not  g1648 (n1392, n373);
not  g1649 (n1590, n412);
buf  g1650 (n1761, n591);
buf  g1651 (n751, n367);
not  g1652 (n2053, n637);
buf  g1653 (n1308, n200);
not  g1654 (n1515, n469);
buf  g1655 (n2038, n578);
buf  g1656 (n934, n332);
not  g1657 (n716, n551);
buf  g1658 (n1802, n472);
not  g1659 (n1386, n168);
buf  g1660 (n1337, n431);
buf  g1661 (n855, n549);
buf  g1662 (n1040, n621);
not  g1663 (n2000, n211);
not  g1664 (n2016, n658);
buf  g1665 (n1088, n407);
buf  g1666 (n1103, n238);
buf  g1667 (n1753, n381);
buf  g1668 (n1147, n359);
not  g1669 (n1292, n607);
not  g1670 (n1057, n188);
buf  g1671 (n1614, n445);
not  g1672 (n1199, n240);
buf  g1673 (n2017, n276);
buf  g1674 (n1541, n383);
buf  g1675 (n1743, n329);
not  g1676 (n746, n599);
not  g1677 (n1598, n612);
buf  g1678 (n1578, n367);
not  g1679 (n1489, n230);
not  g1680 (n1030, n512);
not  g1681 (n1130, n412);
buf  g1682 (n1987, n175);
not  g1683 (n1340, n290);
not  g1684 (n860, n202);
not  g1685 (n1257, n346);
buf  g1686 (n1529, n429);
not  g1687 (n839, n564);
not  g1688 (n2032, n216);
not  g1689 (n940, n161);
buf  g1690 (n1445, n576);
buf  g1691 (n915, n174);
not  g1692 (n1830, n269);
not  g1693 (n1497, n654);
buf  g1694 (n1968, n288);
not  g1695 (n838, n270);
not  g1696 (n1908, n640);
not  g1697 (n1157, n392);
not  g1698 (n1993, n411);
not  g1699 (n1433, n323);
buf  g1700 (n1123, n574);
not  g1701 (n1363, n231);
not  g1702 (n1543, n306);
buf  g1703 (n703, n629);
not  g1704 (n1920, n313);
buf  g1705 (n723, n596);
buf  g1706 (n1230, n341);
buf  g1707 (n997, n506);
not  g1708 (n1891, n345);
not  g1709 (n1667, n440);
buf  g1710 (n1294, n251);
not  g1711 (n975, n527);
not  g1712 (n1746, n386);
not  g1713 (n1169, n518);
buf  g1714 (n1117, n274);
not  g1715 (n1737, n500);
not  g1716 (n1919, n534);
buf  g1717 (n1519, n664);
not  g1718 (n1154, n508);
not  g1719 (n1649, n419);
buf  g1720 (n1813, n412);
buf  g1721 (n1367, n263);
not  g1722 (n1275, n606);
buf  g1723 (n709, n638);
buf  g1724 (n1904, n363);
buf  g1725 (n892, n316);
buf  g1726 (n1719, n317);
not  g1727 (n1693, n340);
not  g1728 (n1475, n666);
buf  g1729 (n1530, n460);
not  g1730 (n1547, n547);
not  g1731 (n1713, n645);
not  g1732 (n724, n295);
buf  g1733 (n1317, n603);
not  g1734 (n1582, n291);
buf  g1735 (n1952, n175);
not  g1736 (n1711, n590);
buf  g1737 (n792, n401);
buf  g1738 (n2026, n366);
buf  g1739 (n1082, n568);
not  g1740 (n1400, n301);
not  g1741 (n1787, n234);
not  g1742 (n1665, n549);
buf  g1743 (n1491, n226);
buf  g1744 (n1797, n527);
buf  g1745 (n1764, n642);
buf  g1746 (n1523, n545);
not  g1747 (n1897, n446);
not  g1748 (n1546, n407);
buf  g1749 (n899, n435);
buf  g1750 (n1661, n486);
not  g1751 (n1619, n371);
not  g1752 (n808, n276);
not  g1753 (n1534, n305);
buf  g1754 (n1288, n299);
not  g1755 (n1297, n177);
not  g1756 (n931, n439);
buf  g1757 (n1678, n459);
not  g1758 (n1820, n410);
not  g1759 (n1453, n649);
buf  g1760 (n816, n544);
buf  g1761 (n1664, n485);
buf  g1762 (n1792, n349);
buf  g1763 (n1673, n641);
not  g1764 (n1640, n408);
buf  g1765 (n994, n424);
not  g1766 (n2046, n585);
buf  g1767 (n1990, n196);
not  g1768 (n1095, n261);
not  g1769 (n1101, n509);
buf  g1770 (n1208, n246);
not  g1771 (n1134, n481);
buf  g1772 (n2081, n634);
buf  g1773 (n1346, n340);
buf  g1774 (n1906, n348);
buf  g1775 (n933, n496);
not  g1776 (n1289, n305);
buf  g1777 (n1104, n448);
not  g1778 (n884, n373);
not  g1779 (n748, n611);
not  g1780 (n959, n220);
buf  g1781 (n1629, n237);
buf  g1782 (n1586, n515);
buf  g1783 (n1533, n520);
not  g1784 (n1108, n463);
not  g1785 (n1046, n199);
not  g1786 (n937, n189);
not  g1787 (n1390, n646);
not  g1788 (n1499, n184);
not  g1789 (n1084, n190);
buf  g1790 (n771, n507);
not  g1791 (n2040, n212);
buf  g1792 (n2072, n321);
buf  g1793 (n1348, n656);
buf  g1794 (n907, n537);
not  g1795 (n1825, n217);
not  g1796 (n1285, n494);
not  g1797 (n1807, n302);
buf  g1798 (n866, n288);
buf  g1799 (n1401, n278);
not  g1800 (n1729, n182);
buf  g1801 (n1712, n655);
buf  g1802 (n677, n170);
not  g1803 (n1514, n634);
buf  g1804 (n777, n181);
buf  g1805 (n912, n460);
not  g1806 (n2037, n462);
not  g1807 (n1645, n525);
buf  g1808 (n939, n341);
buf  g1809 (n1717, n605);
buf  g1810 (n1011, n380);
not  g1811 (n1585, n322);
buf  g1812 (n1804, n382);
not  g1813 (n952, n492);
not  g1814 (n822, n617);
buf  g1815 (n1980, n657);
buf  g1816 (n1274, n424);
buf  g1817 (n1319, n397);
not  g1818 (n944, n425);
buf  g1819 (n943, n452);
not  g1820 (n1343, n479);
not  g1821 (n1018, n183);
not  g1822 (n1565, n193);
not  g1823 (n969, n361);
buf  g1824 (n2054, n478);
not  g1825 (n842, n271);
buf  g1826 (n1232, n352);
buf  g1827 (n1480, n623);
not  g1828 (n1949, n500);
buf  g1829 (n1974, n526);
not  g1830 (n2070, n487);
buf  g1831 (n1252, n585);
buf  g1832 (n734, n349);
buf  g1833 (n1696, n660);
buf  g1834 (n1466, n231);
buf  g1835 (n695, n219);
buf  g1836 (n1884, n294);
buf  g1837 (n1863, n187);
buf  g1838 (n2015, n501);
not  g1839 (n1868, n664);
buf  g1840 (n2052, n523);
buf  g1841 (n1171, n298);
not  g1842 (n1462, n264);
nand g1843 (n849, n456, n300);
nand g1844 (n879, n316, n471, n214, n326);
xor  g1845 (n1486, n659, n335, n403, n576);
or   g1846 (n1999, n616, n297, n440, n164);
xnor g1847 (n1935, n650, n205, n304, n254);
nand g1848 (n1691, n245, n517, n161, n270);
nand g1849 (n1177, n273, n187, n575, n379);
and  g1850 (n713, n210, n222, n340, n366);
nor  g1851 (n1270, n191, n614, n287, n245);
xnor g1852 (n1513, n411, n189, n428, n552);
xor  g1853 (n1789, n383, n330, n283, n249);
or   g1854 (n826, n500, n413, n293, n192);
or   g1855 (n857, n321, n404, n535, n456);
and  g1856 (n1577, n571, n543, n198, n397);
and  g1857 (n1248, n476, n269, n302, n600);
nand g1858 (n1728, n441, n344, n394, n201);
nor  g1859 (n1309, n663, n444, n200);
nor  g1860 (n1214, n183, n623, n641, n614);
xnor g1861 (n1311, n372, n373, n182, n196);
xor  g1862 (n1699, n277, n265, n667, n466);
and  g1863 (n955, n454, n371, n328, n264);
nor  g1864 (n2007, n300, n635, n308, n207);
xor  g1865 (n1420, n309, n574, n169, n542);
xnor g1866 (n820, n394, n607, n516, n233);
or   g1867 (n1265, n650, n495, n493, n258);
and  g1868 (n1464, n539, n415, n501, n326);
xnor g1869 (n1727, n439, n346, n188, n278);
xnor g1870 (n674, n595, n275, n622, n405);
nand g1871 (n901, n277, n521, n504, n399);
xnor g1872 (n1460, n591, n473, n550, n214);
nor  g1873 (n1254, n541, n458, n352, n286);
nor  g1874 (n1368, n498, n482, n255, n528);
xor  g1875 (n1204, n165, n432, n642, n409);
or   g1876 (n1126, n245, n344, n180, n562);
xor  g1877 (n1341, n227, n507, n279, n172);
or   g1878 (n1592, n387, n454, n314, n212);
xor  g1879 (n938, n182, n495, n243, n658);
xnor g1880 (n1788, n327, n502, n653, n241);
nand g1881 (n1872, n314, n264, n522, n488);
or   g1882 (n1850, n333, n475, n330, n349);
xor  g1883 (n1628, n612, n184, n318, n201);
nor  g1884 (n1520, n223, n348, n560, n416);
xnor g1885 (n1430, n523, n598, n359, n314);
xor  g1886 (n1517, n308, n627, n249, n348);
nand g1887 (n1246, n615, n463, n577, n450);
or   g1888 (n1195, n331, n624, n310, n528);
xnor g1889 (n1373, n410, n281, n253, n627);
nor  g1890 (n1280, n505, n569, n465, n638);
and  g1891 (n853, n648, n194, n271, n587);
nand g1892 (n1127, n577, n313, n579, n427);
xnor g1893 (n1345, n307, n458, n632, n441);
xnor g1894 (n671, n332, n409, n237, n315);
and  g1895 (n1823, n222, n379, n250, n429);
xor  g1896 (n1360, n263, n508, n532, n210);
and  g1897 (n1985, n203, n620, n451, n375);
xor  g1898 (n1261, n286, n510, n486, n344);
and  g1899 (n1144, n594, n263, n257, n236);
or   g1900 (n953, n597, n168, n419, n202);
xor  g1901 (n1189, n500, n655, n413, n546);
nor  g1902 (n1487, n511, n425, n429, n209);
xor  g1903 (n1196, n273, n427, n615, n597);
or   g1904 (n1516, n258, n658, n188, n402);
and  g1905 (n1388, n543, n322, n625, n265);
and  g1906 (n1976, n649, n666, n437, n217);
xnor g1907 (n1575, n199, n483, n583, n350);
xor  g1908 (n1455, n571, n183, n643, n637);
xnor g1909 (n739, n531, n247, n536, n443);
nor  g1910 (n1350, n484, n334, n626, n573);
nor  g1911 (n1966, n478, n244, n506, n231);
xnor g1912 (n885, n354, n644, n195, n295);
xor  g1913 (n1762, n431, n229, n285, n276);
nor  g1914 (n1417, n218, n357, n569, n352);
nand g1915 (n1837, n591, n614, n497, n442);
and  g1916 (n2036, n205, n604, n487, n599);
nor  g1917 (n1332, n488, n251, n451, n547);
or   g1918 (n1721, n562, n370, n176, n618);
xor  g1919 (n928, n561, n321, n347, n396);
xnor g1920 (n1975, n545, n286, n442, n642);
or   g1921 (n1306, n438, n542, n198, n424);
or   g1922 (n1631, n298, n632, n661, n198);
nand g1923 (n686, n197, n541, n213, n371);
nor  g1924 (n1342, n315, n654, n370, n386);
xnor g1925 (n1709, n292, n545, n641, n580);
nor  g1926 (n1846, n212, n471, n280, n560);
xor  g1927 (n823, n406, n653, n248, n582);
nor  g1928 (n1819, n199, n475, n293, n328);
xnor g1929 (n1978, n502, n399, n217, n314);
xor  g1930 (n1886, n289, n396, n324, n280);
or   g1931 (n1963, n177, n436, n622, n389);
and  g1932 (n1452, n571, n183, n262, n625);
nand g1933 (n1136, n328, n656, n573, n449);
xnor g1934 (n1907, n375, n261, n222, n483);
nor  g1935 (n1674, n193, n584, n316, n609);
xnor g1936 (n1741, n303, n584, n271, n428);
and  g1937 (n1170, n620, n519, n289, n307);
or   g1938 (n948, n583, n176, n202, n527);
xnor g1939 (n1689, n170, n465, n558, n531);
xor  g1940 (n1772, n246, n363, n423, n498);
xnor g1941 (n985, n442, n280, n580, n317);
and  g1942 (n1958, n627, n272, n565, n482);
nand g1943 (n1131, n230, n532, n453, n620);
nand g1944 (n904, n310, n648, n587, n364);
or   g1945 (n706, n665, n245, n184, n357);
xor  g1946 (n1869, n605, n606, n253, n226);
xnor g1947 (n1560, n260, n391, n610, n256);
nand g1948 (n924, n219, n661, n568, n251);
xnor g1949 (n2062, n391, n236, n421, n267);
nor  g1950 (n1205, n400, n533, n644, n621);
xor  g1951 (n918, n258, n649, n553, n572);
nand g1952 (n1700, n473, n434, n513, n666);
or   g1953 (n1941, n613, n287, n299, n605);
xnor g1954 (n712, n318, n329, n246, n407);
and  g1955 (n1164, n246, n566, n419);
and  g1956 (n1931, n232, n588, n602, n395);
xnor g1957 (n1267, n351, n438, n342, n666);
nor  g1958 (n1478, n228, n662, n390, n239);
xnor g1959 (n926, n298, n353, n444, n461);
nand g1960 (n761, n358, n630, n312, n185);
nand g1961 (n1612, n560, n648, n659, n454);
and  g1962 (n1928, n595, n447, n366, n313);
xnor g1963 (n883, n239, n392, n633, n164);
nand g1964 (n1771, n600, n326, n295, n413);
nor  g1965 (n1929, n541, n319, n220, n509);
nor  g1966 (n681, n327, n514, n542, n255);
and  g1967 (n1826, n460, n562, n290, n568);
nand g1968 (n675, n451, n564, n436, n225);
and  g1969 (n2027, n168, n354, n455, n640);
xnor g1970 (n1253, n288, n340, n426, n468);
nor  g1971 (n851, n557, n464, n540, n215);
nand g1972 (n1675, n360, n519, n358, n172);
and  g1973 (n1463, n457, n257, n262, n384);
and  g1974 (n1956, n192, n538, n326, n208);
and  g1975 (n1062, n228, n418, n630, n420);
or   g1976 (n1625, n619, n449, n378, n258);
xor  g1977 (n698, n368, n185, n636, n504);
and  g1978 (n1785, n204, n608, n265, n588);
xor  g1979 (n1870, n323, n494, n212, n563);
nor  g1980 (n1793, n263, n292, n266, n388);
or   g1981 (n1055, n364, n443, n518, n521);
nand g1982 (n1357, n380, n221, n351, n165);
xor  g1983 (n1042, n649, n393, n601, n178);
xnor g1984 (n1152, n387, n332, n269, n171);
or   g1985 (n1644, n195, n495, n167, n252);
nand g1986 (n1841, n281, n467, n633, n297);
nand g1987 (n1710, n633, n199, n537, n644);
xnor g1988 (n1507, n569, n335, n405, n511);
xor  g1989 (n2078, n566, n206, n403, n365);
xor  g1990 (n1296, n494, n337, n301, n224);
or   g1991 (n2059, n532, n550, n320, n244);
nor  g1992 (n1029, n211, n538, n353, n385);
nor  g1993 (n1446, n367, n654, n655, n565);
and  g1994 (n719, n585, n547, n653, n259);
xnor g1995 (n1415, n374, n372, n411, n571);
xnor g1996 (n1681, n408, n485, n331, n486);
xnor g1997 (n941, n535, n205, n260, n458);
and  g1998 (n1695, n401, n602, n443, n187);
or   g1999 (n1305, n322, n491, n609, n352);
and  g2000 (n2045, n639, n540, n181, n266);
and  g2001 (n1580, n651, n192, n284, n432);
nor  g2002 (n714, n297, n284, n325, n387);
nand g2003 (n1803, n661, n404, n518, n221);
nand g2004 (n1589, n575, n430, n358, n304);
nor  g2005 (n1054, n378, n581, n534, n603);
xnor g2006 (n1037, n356, n218, n172, n240);
nand g2007 (n2010, n355, n297, n522, n362);
xor  g2008 (n1883, n287, n187, n174, n328);
xor  g2009 (n1320, n465, n219, n648, n172);
and  g2010 (n1554, n534, n303, n481, n463);
or   g2011 (n756, n365, n267, n385, n470);
nand g2012 (n1548, n422, n236, n431, n438);
nand g2013 (n1715, n539, n630, n391, n250);
nor  g2014 (n2065, n469, n623, n338, n518);
or   g2015 (n1859, n197, n455, n332, n327);
or   g2016 (n1201, n343, n646, n502, n384);
xor  g2017 (n829, n505, n208, n608, n663);
and  g2018 (n1077, n196, n218, n601, n573);
or   g2019 (n1971, n540, n211, n598, n248);
xor  g2020 (n1477, n163, n484, n198, n383);
or   g2021 (n1222, n650, n162, n266, n337);
nand g2022 (n832, n235, n397, n267, n262);
nor  g2023 (n1250, n453, n190, n619, n606);
nor  g2024 (n1427, n327, n453, n201, n365);
xnor g2025 (n1081, n523, n525, n639, n414);
and  g2026 (n979, n657, n458, n242, n164);
nor  g2027 (n2069, n551, n549, n575, n472);
xnor g2028 (n1286, n422, n291, n360, n279);
and  g2029 (n1423, n362, n527, n663, n596);
xnor g2030 (n806, n286, n279, n519, n339);
or   g2031 (n1509, n339, n572, n322, n178);
xor  g2032 (n715, n480, n617, n546, n295);
nor  g2033 (n691, n481, n255, n377, n631);
and  g2034 (n971, n519, n377, n204, n279);
xor  g2035 (n1670, n464, n611, n237, n227);
nand g2036 (n1271, n635, n209, n268, n456);
nand g2037 (n1902, n543, n602, n617, n652);
nand g2038 (n1032, n629, n417, n639, n391);
or   g2039 (n1447, n427, n651, n384, n504);
or   g2040 (n799, n544, n637, n613, n461);
and  g2041 (n1302, n426, n288, n630, n642);
nand g2042 (n2042, n535, n629, n482, n497);
and  g2043 (n1942, n497, n296, n508, n454);
nand g2044 (n1186, n354, n319, n645, n430);
or   g2045 (n830, n491, n195, n459, n356);
xor  g2046 (n1766, n362, n583, n323, n406);
xor  g2047 (n752, n652, n475, n439, n468);
nand g2048 (n1141, n612, n558, n470, n605);
xnor g2049 (n2515, n689, n1478, n1127, n1197);
xor  g2050 (n2187, n1224, n1161, n1883, n2014);
xor  g2051 (n2348, n1815, n773, n1676, n1074);
nor  g2052 (n2379, n1955, n1730, n1474, n1963);
and  g2053 (n2717, n1293, n1025, n2058, n1257);
nor  g2054 (n2646, n1427, n1112, n1199, n811);
and  g2055 (n2296, n1267, n717, n1017, n1741);
nand g2056 (n2321, n1688, n1756, n862, n1147);
nor  g2057 (n2237, n1507, n1886, n1137, n1506);
and  g2058 (n2532, n1739, n1233, n1248, n1287);
nand g2059 (n2432, n2019, n995, n678, n2068);
nor  g2060 (n2500, n1207, n1729, n1572, n1832);
xor  g2061 (n2558, n1111, n1610, n2003, n1941);
and  g2062 (n2622, n1435, n1657, n1927, n1388);
and  g2063 (n2122, n1936, n1202, n1740, n2052);
xnor g2064 (n2093, n2037, n1462, n1437, n1651);
xor  g2065 (n2088, n1685, n2028, n2023, n1180);
nand g2066 (n2227, n1326, n1973, n1397, n1242);
and  g2067 (n2120, n1675, n1470, n1588, n1347);
nor  g2068 (n2360, n1640, n1726, n1624, n1626);
nor  g2069 (n2513, n2015, n1645, n1580, n1779);
or   g2070 (n2493, n1972, n1811, n1232, n1909);
nand g2071 (n2281, n1886, n1576, n1940, n1951);
and  g2072 (n2262, n2046, n852, n1613, n1346);
nand g2073 (n2346, n1527, n1598, n1312, n801);
and  g2074 (n2685, n1919, n1990, n1737, n939);
nand g2075 (n2479, n1009, n1279, n1389, n2024);
xor  g2076 (n2620, n2061, n1683, n769, n1080);
nor  g2077 (n2437, n2003, n1289, n1998, n753);
or   g2078 (n2619, n1273, n1570, n1685, n1543);
xnor g2079 (n2430, n1867, n894, n2002, n951);
or   g2080 (n2245, n1767, n1744, n1300, n1317);
nand g2081 (n2171, n1271, n2055, n694, n1502);
xnor g2082 (n2089, n1309, n1689, n1242, n1836);
and  g2083 (n2687, n1286, n899, n1923, n1033);
xor  g2084 (n2494, n1496, n1991, n874, n1368);
nand g2085 (n2714, n1596, n2043, n1937, n1348);
nand g2086 (n2635, n1282, n1366, n982, n1479);
xor  g2087 (n2453, n1543, n1765, n1217, n1310);
nor  g2088 (n2092, n1517, n1480, n864, n1597);
or   g2089 (n2114, n1363, n1793, n2059, n1937);
xor  g2090 (n2216, n1932, n1410, n766, n1577);
xnor g2091 (n2234, n1773, n1485, n1591, n983);
nor  g2092 (n2675, n1233, n1815, n1345, n1937);
or   g2093 (n2428, n1844, n1934, n1483, n680);
nor  g2094 (n2385, n2054, n1275, n1133, n1601);
nand g2095 (n2424, n1184, n1817, n1200, n1646);
and  g2096 (n2490, n2050, n1569, n2037, n696);
nand g2097 (n2365, n1981, n1217, n806, n1916);
nand g2098 (n2377, n1160, n1380, n1759, n1584);
xnor g2099 (n2690, n1991, n2012, n1833, n963);
xnor g2100 (n2603, n1514, n879, n1515, n1304);
or   g2101 (n2408, n1382, n1995, n2053, n2040);
xor  g2102 (n2295, n731, n2003, n2030, n2062);
nor  g2103 (n2459, n1644, n1297, n1637, n1324);
nand g2104 (n2366, n1884, n1655, n1633, n1982);
or   g2105 (n2284, n1809, n1675, n2017, n2012);
xnor g2106 (n2465, n1669, n1504, n1575, n1421);
xor  g2107 (n2306, n1077, n2023, n1941, n1852);
nor  g2108 (n2156, n1966, n1358, n1474, n1457);
nor  g2109 (n2436, n940, n1686, n1176, n781);
and  g2110 (n2421, n1510, n2004, n1952, n1064);
xnor g2111 (n2451, n2045, n1913, n1013, n1937);
or   g2112 (n2405, n1827, n1290, n1385, n1894);
and  g2113 (n2688, n1220, n1835, n1621, n954);
nor  g2114 (n2559, n1436, n887, n1711, n1702);
xnor g2115 (n2653, n2026, n2027, n722, n1598);
nand g2116 (n2501, n1857, n1893, n1602, n1205);
and  g2117 (n2575, n992, n1691, n1896, n2024);
or   g2118 (n2581, n1535, n1463, n1483, n1987);
xnor g2119 (n2695, n1881, n821, n1395, n1563);
xnor g2120 (n2669, n1278, n2071, n1947, n1892);
and  g2121 (n2384, n1120, n1679, n1335, n990);
xnor g2122 (n2201, n863, n1957, n1413, n1073);
xor  g2123 (n2108, n1861, n1476, n1988, n1043);
or   g2124 (n2204, n1404, n1997, n1645, n1314);
and  g2125 (n2246, n1673, n1311, n2066, n1681);
and  g2126 (n2457, n1215, n1353, n1705, n2000);
xnor g2127 (n2263, n1254, n777, n1191, n1650);
xor  g2128 (n2336, n798, n1453, n1799, n1864);
nand g2129 (n2252, n1490, n1579, n2068, n795);
xnor g2130 (n2241, n1244, n1684, n1811, n2029);
nand g2131 (n2645, n1540, n2012, n1783, n1394);
nand g2132 (n2648, n1926, n2053, n1366, n786);
or   g2133 (n2231, n1634, n1647, n896, n2034);
nor  g2134 (n2576, n1871, n1325, n1236, n1589);
or   g2135 (n2115, n2060, n1139, n1704, n1891);
xor  g2136 (n2264, n1883, n1461, n2065, n1041);
xor  g2137 (n2309, n1845, n914, n2018, n743);
xor  g2138 (n2388, n1274, n1944, n2004, n1525);
or   g2139 (n2090, n2016, n2004, n698, n733);
xnor g2140 (n2086, n1694, n1967, n986, n1438);
xnor g2141 (n2352, n1625, n1954, n1557, n1599);
nor  g2142 (n2621, n927, n2065, n1424, n2006);
xnor g2143 (n2461, n757, n1944, n1364, n1877);
or   g2144 (n2539, n1361, n1415, n1550, n816);
xor  g2145 (n2151, n759, n2067, n1652, n1068);
nor  g2146 (n2696, n2051, n701, n1556, n1528);
and  g2147 (n2323, n1416, n809, n1393, n935);
xnor g2148 (n2111, n888, n1089, n1967, n1969);
xor  g2149 (n2382, n1873, n1611, n1868, n1051);
and  g2150 (n2230, n1976, n857, n1435, n1676);
xor  g2151 (n2105, n2049, n1984, n1440, n761);
nand g2152 (n2652, n1952, n1596, n1315, n1509);
and  g2153 (n2103, n1425, n2027, n2039, n1333);
xnor g2154 (n2137, n1249, n909, n1559, n1239);
xor  g2155 (n2387, n671, n1665, n2000, n1880);
xnor g2156 (n2126, n1602, n868, n1151, n1982);
nand g2157 (n2391, n1824, n1644, n2019, n1530);
or   g2158 (n2691, n762, n1630, n1692, n1648);
xnor g2159 (n2507, n1528, n730, n1228, n1305);
or   g2160 (n2270, n1460, n1004, n1315, n1439);
nand g2161 (n2362, n1130, n1728, n1712, n1729);
and  g2162 (n2598, n1072, n2041, n1639, n1114);
nand g2163 (n2613, n1553, n1206, n1951, n674);
xnor g2164 (n2184, n772, n1930, n1812, n1451);
nand g2165 (n2261, n1499, n2055, n1783, n1475);
nand g2166 (n2670, n1516, n1623, n1968, n1375);
nand g2167 (n2460, n2001, n1103, n890, n1225);
or   g2168 (n2548, n1251, n2019, n1323, n1997);
xnor g2169 (n2179, n1774, n1219, n1803, n1865);
or   g2170 (n2302, n2025, n1510, n1480, n1558);
and  g2171 (n2700, n1848, n1974, n1915, n2046);
xnor g2172 (n2213, n1849, n1595, n713, n1036);
xor  g2173 (n2701, n1422, n1548, n1973, n1875);
and  g2174 (n2510, n1760, n1948, n1622, n1840);
xor  g2175 (n2486, n1307, n1037, n1938, n1915);
nand g2176 (n2316, n1903, n1305, n1720, n2070);
xnor g2177 (n2340, n2009, n1971, n922, n1861);
xor  g2178 (n2170, n1971, n1954, n1988, n1749);
nand g2179 (n2466, n1326, n1355, n1990, n2021);
xnor g2180 (n2149, n1332, n1471, n1810, n1210);
or   g2181 (n2305, n1671, n1341, n897, n1777);
and  g2182 (n2516, n1030, n692, n1559, n1373);
or   g2183 (n2692, n1313, n1420, n1962, n1668);
or   g2184 (n2596, n1869, n1466, n1283, n1995);
nor  g2185 (n2469, n1563, n2002, n1722, n2015);
xor  g2186 (n2628, n1680, n1986, n1391, n985);
nor  g2187 (n2359, n1342, n2050, n972, n1946);
or   g2188 (n2082, n910, n2007, n2024, n1338);
or   g2189 (n2523, n1354, n1015, n1957, n1042);
and  g2190 (n2608, n1640, n1658, n1919, n1251);
xor  g2191 (n2444, n1858, n1261, n1411, n1443);
nor  g2192 (n2221, n2064, n690, n881, n1847);
or   g2193 (n2591, n1336, n797, n1473, n1620);
xor  g2194 (n2297, n2007, n1029, n1993, n1952);
or   g2195 (n2313, n2051, n1402, n1723, n1986);
and  g2196 (n2588, n1878, n1971, n1715, n1555);
nor  g2197 (n2565, n794, n1345, n1953, n2010);
nand g2198 (n2595, n1661, n1472, n1955, n1974);
or   g2199 (n2491, n1698, n1784, n1950, n1395);
xor  g2200 (n2573, n810, n1205, n1222, n1735);
xnor g2201 (n2146, n1243, n1673, n2066, n1451);
nor  g2202 (n2206, n1819, n1405, n1248, n1948);
nand g2203 (n2238, n2058, n867, n1503, n1822);
and  g2204 (n2470, n1960, n1898, n1132, n2009);
xnor g2205 (n2311, n1203, n2044, n1863, n1350);
xor  g2206 (n2478, n1520, n2059, n699, n980);
xnor g2207 (n2123, n728, n1939, n1859, n1319);
xor  g2208 (n2683, n1287, n1351, n1519, n755);
and  g2209 (n2593, n1316, n903, n827, n1929);
nor  g2210 (n2177, n1974, n1470, n1523, n947);
xnor g2211 (n2441, n1921, n1982, n1479, n949);
or   g2212 (n2662, n1034, n1376, n902, n1810);
nand g2213 (n2096, n2046, n1478, n2032, n2018);
and  g2214 (n2618, n1275, n1756, n2054, n1933);
xor  g2215 (n2383, n2025, n1447, n1212, n1752);
nor  g2216 (n2564, n1376, n2010, n1984, n1213);
xnor g2217 (n2167, n1235, n1956, n726, n792);
or   g2218 (n2401, n1551, n1833, n1925, n2000);
or   g2219 (n2275, n1079, n1658, n1362, n2022);
xor  g2220 (n2592, n1095, n2038, n1381, n1765);
and  g2221 (n2549, n1562, n1989, n1840, n1776);
and  g2222 (n2338, n2000, n1399, n962, n1727);
or   g2223 (n2176, n1101, n1467, n1583, n1401);
or   g2224 (n2205, n929, n978, n1799, n2031);
nand g2225 (n2250, n1800, n1962, n1674, n1784);
or   g2226 (n2310, n1016, n931, n1888, n1582);
and  g2227 (n2172, n1956, n1196, n1947, n1539);
nor  g2228 (n2681, n2038, n1457, n1335, n930);
and  g2229 (n2659, n851, n1481, n2070, n886);
xnor g2230 (n2135, n1003, n1740, n1048, n1935);
xor  g2231 (n2518, n1750, n1142, n1996, n1947);
or   g2232 (n2403, n1996, n1935, n928, n1485);
or   g2233 (n2290, n1524, n1339, n1134, n1614);
or   g2234 (n2254, n2042, n1710, n1969, n1961);
nor  g2235 (n2267, n1901, n1276, n1804, n2028);
nor  g2236 (n2330, n1999, n2009, n1738, n1945);
xnor g2237 (n2188, n2008, n1863, n1662, n1994);
and  g2238 (n2474, n1899, n1731, n1959, n2009);
nand g2239 (n2508, n1417, n1618, n1738, n1690);
and  g2240 (n2439, n1442, n1352, n2008, n2063);
xnor g2241 (n2433, n1115, n1788, n1230, n1428);
nor  g2242 (n2654, n1297, n1772, n1131, n1992);
or   g2243 (n2106, n744, n1672, n1271, n941);
xnor g2244 (n2130, n1865, n725, n2024, n1378);
xor  g2245 (n2580, n1980, n2023, n1821, n1616);
nand g2246 (n2398, n774, n1874, n735, n1413);
xor  g2247 (n2600, n758, n738, n1493, n1220);
or   g2248 (n2489, n1019, n1897, n1934, n1781);
nand g2249 (n2393, n1231, n1562, n1329, n1207);
xor  g2250 (n2158, n1223, n1396, n703, n1625);
xor  g2251 (n2319, n2039, n1818, n1464, n1928);
and  g2252 (n2165, n1953, n1965, n1285, n1542);
xor  g2253 (n2540, n1763, n1869, n943, n876);
or   g2254 (n2535, n1923, n1477, n2013, n975);
xnor g2255 (n2226, n1917, n2053, n1629, n1981);
or   g2256 (n2425, n1850, n1653, n1238, n1302);
and  g2257 (n2657, n1195, n1925, n1699, n1397);
nand g2258 (n2095, n1734, n1402, n843, n1560);
xor  g2259 (n2322, n2022, n1371, n1511, n1549);
and  g2260 (n2299, n1682, n1194, n1211, n1940);
and  g2261 (n2314, n1182, n1870, n1301, n752);
or   g2262 (n2222, n1239, n1978, n837, n1594);
nor  g2263 (n2449, n1642, n1136, n1960, n1826);
or   g2264 (n2361, n1804, n1980, n1081, n1905);
nand g2265 (n2697, n1938, n2060, n1964, n1660);
nand g2266 (n2202, n1578, n1178, n1764, n1854);
and  g2267 (n2715, n1463, n1950, n1767, n1722);
xnor g2268 (n2423, n988, n1827, n2047, n1360);
or   g2269 (n2185, n1444, n2007, n926, n2011);
nand g2270 (n2148, n1407, n1405, n1247, n875);
xor  g2271 (n2467, n1949, n2025, n1467, n977);
xnor g2272 (n2364, n1618, n1476, n1503, n853);
xnor g2273 (n2193, n1766, n1020, n1281, n1449);
nand g2274 (n2370, n1152, n2063, n1619, n1716);
and  g2275 (n2434, n1304, n1632, n1206, n1721);
xnor g2276 (n2209, n771, n1018, n1124, n1825);
and  g2277 (n2571, n1146, n1442, n1513, n685);
xnor g2278 (n2527, n2050, n1038, n1446, n2022);
or   g2279 (n2496, n1961, n1968, n1590, n1979);
and  g2280 (n2661, n765, n1724, n1953, n2036);
nand g2281 (n2504, n1600, n1778, n2033, n1951);
nor  g2282 (n2286, n1216, n1552, n1585, n1404);
nor  g2283 (n2235, n1403, n1277, n1213, n1841);
xnor g2284 (n2534, n720, n760, n1568, n2063);
nand g2285 (n2390, n1858, n1374, n1968, n848);
or   g2286 (n2686, n936, n2045, n1560, n1456);
xor  g2287 (n2712, n1193, n2050, n1791, n1949);
xor  g2288 (n2304, n957, n1994, n1262, n1963);
xor  g2289 (n2506, n1889, n1697, n1426, n1450);
nand g2290 (n2271, n1257, n1339, n1392, n2036);
nor  g2291 (n2112, n1422, n1761, n1862, n2001);
nor  g2292 (n2498, n1978, n849, n1608, n1902);
xor  g2293 (n2519, n1661, n1825, n2011, n1356);
xnor g2294 (n2169, n895, n1628, n2059, n1670);
nand g2295 (n2144, n1505, n2027, n1592, n687);
xnor g2296 (n2233, n1306, n1964, n1309, n1501);
or   g2297 (n2509, n1972, n684, n1795, n1065);
nand g2298 (n2589, n1155, n855, n1377, n1340);
and  g2299 (n2577, n1983, n1839, n712, n1002);
and  g2300 (n2339, n1747, n1230, n1331, n790);
xnor g2301 (n2279, n707, n1960, n2020, n1859);
or   g2302 (n2468, n1502, n1890, n1763, n1747);
xor  g2303 (n2642, n1224, n2023, n846, n1603);
or   g2304 (n2607, n1940, n1214, n1550, n1225);
xnor g2305 (n2255, n1914, n1683, n1188, n1360);
or   g2306 (n2312, n1942, n1236, n1484, n920);
xnor g2307 (n2599, n1914, n1508, n783, n1656);
xor  g2308 (n2409, n1145, n1209, n1986, n1511);
and  g2309 (n2578, n2025, n1379, n2048, n742);
and  g2310 (n2693, n877, n1497, n1965, n835);
xnor g2311 (n2522, n1040, n824, n856, n1584);
nand g2312 (n2372, n1617, n1637, n1157, n945);
nor  g2313 (n2650, n1604, n1448, n2070, n2056);
and  g2314 (n2288, n1876, n2057, n693, n1778);
or   g2315 (n2435, n1096, n1447, n1970, n1234);
and  g2316 (n2638, n1989, n1229, n1278, n1186);
or   g2317 (n2097, n1718, n1868, n1580, n2058);
or   g2318 (n2601, n2029, n1624, n1338, n1643);
xnor g2319 (n2634, n1121, n750, n1325, n2056);
and  g2320 (n2411, n1529, n912, n1344, n2068);
nand g2321 (n2400, n1978, n1986, n2040, n1622);
xnor g2322 (n2649, n1769, n2047, n1313, n1786);
nor  g2323 (n2538, n1258, n1630, n1319, n1499);
xor  g2324 (n2154, n1629, n1337, n2042, n1979);
nor  g2325 (n2369, n1807, n1218, n1331, n1587);
xnor g2326 (n2157, n2032, n1757, n1296, n1808);
xor  g2327 (n2197, n1520, n2002, n1250, n1035);
or   g2328 (n2716, n1280, n1605, n1210, n1334);
and  g2329 (n2667, n1090, n711, n1906, n1911);
xor  g2330 (n2525, n924, n1987, n1054, n1378);
or   g2331 (n2168, n1918, n1084, n2001, n1253);
xor  g2332 (n2568, n1464, n682, n866, n1736);
and  g2333 (n2673, n1110, n1455, n1775, n1332);
nand g2334 (n2194, n1249, n2004, n815, n1564);
xor  g2335 (n2182, n702, n1458, n1255, n803);
or   g2336 (n2229, n904, n1579, n1168, n2062);
xnor g2337 (n2265, n1597, n1717, n1636, n1943);
xnor g2338 (n2570, n1519, n1649, n1982, n1491);
nor  g2339 (n2429, n1533, n1327, n1489, n1443);
nor  g2340 (n2455, n1379, n1383, n1938, n1714);
nor  g2341 (n2085, n1642, n2049, n1659, n1888);
and  g2342 (n2129, n1264, n2020, n1546, n2028);
and  g2343 (n2274, n1650, n1704, n1429, n1367);
nor  g2344 (n2658, n1771, n1406, n1569, n1302);
or   g2345 (n2303, n1570, n1939, n1414, n1958);
nor  g2346 (n2629, n2065, n1837, n1329, n813);
nor  g2347 (n2684, n2044, n1055, n1259, n2005);
or   g2348 (n2394, n1920, n745, n1968, n2031);
or   g2349 (n2217, n1999, n1431, n1751, n1226);
or   g2350 (n2414, n1709, n793, n1386, n1785);
or   g2351 (n2412, n2057, n956, n1238, n1284);
or   g2352 (n2207, n1286, n1983, n1599, n1855);
xor  g2353 (n2614, n2005, n1860, n1979, n1250);
nand g2354 (n2416, n775, n2017, n1341, n1177);
and  g2355 (n2219, n1192, n1682, n1719, n1932);
nand g2356 (n2438, n1308, n1718, n817, n1211);
and  g2357 (n2107, n2057, n741, n1857, n2030);
nor  g2358 (n2679, n1212, n2020, n1295, n2021);
and  g2359 (n2277, n718, n1495, n1851, n2015);
or   g2360 (n2109, n1653, n1416, n847, n1684);
and  g2361 (n2672, n2043, n1299, n1291, n1056);
or   g2362 (n2402, n2010, n1289, n1936, n1246);
nand g2363 (n2463, n2041, n802, n1733, n932);
and  g2364 (n2554, n2071, n1705, n1383, n796);
xnor g2365 (n2511, n1544, n2035, n1027, n1348);
nand g2366 (n2707, n1265, n1143, n1998, n788);
xnor g2367 (n2533, n1696, n901, n1012, n1792);
and  g2368 (n2102, n1911, n1573, n1727, n1228);
xor  g2369 (n2475, n1581, n1369, n1088, n1488);
and  g2370 (n2143, n1711, n1723, n1616, n2037);
and  g2371 (n2702, n677, n2034, n1904, n2035);
nand g2372 (n2214, n1518, n1774, n916, n1730);
nand g2373 (n2483, n1945, n1589, n734, n1977);
nor  g2374 (n2442, n1805, n746, n688, n1943);
nand g2375 (n2550, n754, n1581, n1881, n1988);
and  g2376 (n2563, n1587, n1380, n1166, n1969);
or   g2377 (n2450, n1994, n1615, n1288, n2017);
nand g2378 (n2627, n1181, n1921, n1517, n1389);
xor  g2379 (n2333, n1534, n1762, n1409, n1237);
xor  g2380 (n2448, n1850, n1234, n1010, n1962);
or   g2381 (n2632, n1227, n1939, n1828, n1816);
nor  g2382 (n2704, n2049, n814, n1266, n2044);
or   g2383 (n2292, n1764, n1267, n1998, n1535);
xor  g2384 (n2236, n1743, n1766, n1449, n697);
or   g2385 (n2574, n1654, n1431, n1135, n1972);
nand g2386 (n2223, n1365, n2010, n1551, n1739);
nand g2387 (n2711, n1368, n1189, n1382, n1428);
xor  g2388 (n2396, n1609, n1958, n1907, n1554);
or   g2389 (n2117, n854, n1836, n1797, n1666);
nor  g2390 (n2445, n1272, n2016, n768, n1970);
xnor g2391 (n2514, n2037, n732, n826, n1761);
nor  g2392 (n2395, n1912, n1525, n1561, n1459);
and  g2393 (n2371, n2047, n998, n1357, n1880);
or   g2394 (n2505, n1586, n1601, n1566, n2042);
and  g2395 (n2488, n1482, n1610, n1058, n1743);
nand g2396 (n2272, n1634, n2044, n1429, n1349);
nand g2397 (n2347, n1948, n1977, n1262, n1487);
nor  g2398 (n2587, n1172, n1996, n1892, n1561);
and  g2399 (n2373, n1069, n946, n2056, n719);
nor  g2400 (n2368, n959, n1809, n1990, n1537);
or   g2401 (n2155, n1910, n1097, n865, n1752);
xnor g2402 (n2555, n1745, n1605, n1290, n1655);
xnor g2403 (n2259, n1820, n1594, n1979, n1209);
nand g2404 (n2497, n1214, n1686, n2013, n1994);
nor  g2405 (n2228, n1536, n1468, n1512, n1311);
xor  g2406 (n2584, n1390, n1781, n1022, n1667);
nand g2407 (n2285, n1999, n1252, n2033, n961);
or   g2408 (n2166, n705, n1515, n1350, n2007);
nor  g2409 (n2243, n1269, n1818, n1631, n1769);
nand g2410 (n2183, n1344, n1606, n1750, n1735);
or   g2411 (n2367, n906, n1997, n1167, n1045);
or   g2412 (n2651, n1678, n1123, n1942, n1949);
and  g2413 (n2195, n1794, n2031, n1714, n1495);
and  g2414 (n2127, n873, n1903, n1492, n1814);
nor  g2415 (n2623, n1159, n1600, n1403, n1835);
nand g2416 (n2175, n1895, n1973, n1384, n1924);
or   g2417 (n2358, n2049, n1953, n1975, n1548);
xnor g2418 (n2139, n1837, n1950, n1664, n2064);
nor  g2419 (n2191, n913, n1853, n1316, n1241);
and  g2420 (n2647, n1455, n1700, n1951, n1306);
nor  g2421 (n2280, n1977, n1523, n1963, n1990);
nor  g2422 (n2606, n1509, n1462, n1489, n1169);
and  g2423 (n2328, n1340, n1093, n1993, n1877);
xnor g2424 (n2212, n1713, n1945, n1343, n1843);
xor  g2425 (n2521, n1076, n1534, n1050, n1526);
or   g2426 (n2150, n1957, n1328, n710, n1218);
and  g2427 (n2590, n1541, n1963, n1882, n1418);
nor  g2428 (n2345, n1314, n1407, n1521, n1494);
and  g2429 (n2529, n1237, n1606, n1999, n1202);
and  g2430 (n2583, n965, n1240, n1959, n950);
nand g2431 (n2705, n1370, n2001, n1847, n1298);
or   g2432 (n2335, n1633, n1894, n1802, n1039);
nor  g2433 (n2477, n1393, n1500, n1370, n1272);
xnor g2434 (n2553, n1417, n1668, n1762, n708);
or   g2435 (n2342, n1179, n1285, n1697, n1641);
xor  g2436 (n2476, n1109, n1666, n1001, n1558);
or   g2437 (n2616, n1940, n917, n1162, n1952);
xor  g2438 (n2329, n1842, n1576, n1776, n1967);
and  g2439 (n2420, n1976, n1721, n968, n1516);
or   g2440 (n2520, n2043, n2003, n1571, n933);
and  g2441 (n2404, n1352, n2052, n1829, n907);
and  g2442 (n2210, n1946, n1260, n1851, n1433);
xor  g2443 (n2443, n2006, n1477, n1798, n1487);
nand g2444 (n2260, n2064, n1531, n1100, n1588);
nand g2445 (n2664, n1412, n2002, n2008, n1768);
nor  g2446 (n2615, n1879, n2030, n1334, n1163);
nand g2447 (n2354, n1893, n1992, n1708, n1985);
xor  g2448 (n2551, n2014, n2062, n1318, n1918);
xor  g2449 (n2694, n1098, n1586, n1920, n1532);
and  g2450 (n2560, n778, n1440, n1254, n1411);
xor  g2451 (n2220, n1703, n1456, n1458, n1874);
or   g2452 (n2278, n1173, n1066, n1274, n1540);
nor  g2453 (n2145, n1412, n942, n1660, n952);
and  g2454 (n2232, n1651, n878, n751, n1454);
xnor g2455 (n2585, n1946, n1623, n1386, n2067);
nor  g2456 (n2268, n832, n782, n1452, n882);
xnor g2457 (n2218, n1981, n1988, n1187, n2026);
nand g2458 (n2380, n1508, n1283, n1418, n1706);
xor  g2459 (n2617, n1873, n1116, n915, n1165);
nor  g2460 (n2582, n858, n1839, n1853, n1913);
and  g2461 (n2174, n1862, n960, n1974, n1987);
xor  g2462 (n2547, n1817, n1604, n2005, n1709);
and  g2463 (n2294, n1909, n1545, n2066, n1959);
nand g2464 (n2344, n1527, n918, n1801, n1626);
xor  g2465 (n2456, n1268, n1964, n1657, n1245);
xnor g2466 (n2104, n1821, n1337, n1849, n2045);
nor  g2467 (n2545, n1221, n948, n1699, n2061);
xnor g2468 (n2481, n715, n1441, n1834, n1343);
xnor g2469 (n2350, n1421, n1318, n2031, n1125);
and  g2470 (n2301, n2066, n860, n2048, n1782);
xor  g2471 (n2407, n859, n1908, n884, n1694);
xor  g2472 (n2605, n1688, n2026, n1593, n845);
nor  g2473 (n2602, n1632, n2042, n1288, n1260);
xor  g2474 (n2422, n2036, n1792, n2018, n787);
nor  g2475 (n2110, n1981, n1549, n1085, n2030);
and  g2476 (n2682, n836, n2033, n1943, n1635);
nand g2477 (n2464, n1797, n1008, n1246, n1190);
and  g2478 (n2211, n1373, n1119, n1536, n1401);
or   g2479 (n2631, n1969, n779, n1931, n1067);
or   g2480 (n2526, n1400, n1546, n1349, n1107);
or   g2481 (n2389, n1444, n1538, n1301, n1917);
xnor g2482 (n2200, n672, n1276, n2021, n1231);
xnor g2483 (n2363, n1948, n1320, n1887, n1736);
and  g2484 (n2557, n2048, n1269, n2070, n1573);
or   g2485 (n2542, n889, n1252, n1690, n1795);
and  g2486 (n2134, n1113, n676, n869, n1966);
nor  g2487 (n2567, n1816, n1203, n850, n1701);
nand g2488 (n2485, n1607, n1359, n2041, n2027);
and  g2489 (n2084, n1574, n1777, n1105, n1787);
xnor g2490 (n2537, n2052, n1049, n1057, n1978);
xnor g2491 (n2318, n1954, n1929, n1796, n1823);
xor  g2492 (n2524, n1996, n1497, n1554, n1566);
xor  g2493 (n2386, n996, n1617, n1531, n1613);
xor  g2494 (n2116, n1460, n1513, n1887, n2014);
nand g2495 (n2710, n1385, n1327, n1215, n1742);
xnor g2496 (n2113, n1813, n861, n1998, n1900);
xnor g2497 (n2495, n1415, n1201, n1264, n981);
nand g2498 (n2668, n1371, n1245, n1150, n2038);
nor  g2499 (n2541, n1270, n763, n1855, n1667);
xnor g2500 (n2198, n1927, n1475, n1791, n825);
nand g2501 (n2633, n1154, n1419, n1263, n1138);
xor  g2502 (n2249, n872, n1279, n1656, n1367);
nor  g2503 (n2418, n1670, n1908, n2069, n1737);
and  g2504 (n2300, n1486, n1904, n1255, n1384);
nand g2505 (n2641, n1277, n2035, n911, n1748);
xnor g2506 (n2291, n2020, n1867, n1342, n1612);
nor  g2507 (n2639, n934, n799, n1256, n1643);
nor  g2508 (n2698, n1691, n1965, n1000, n1266);
xnor g2509 (n2173, n1897, n880, n1828, n1091);
and  g2510 (n2266, n1293, n1980, n1782, n2005);
xnor g2511 (n2308, n1032, n1595, n1757, n1848);
xnor g2512 (n2136, n1078, n1802, n1654, n969);
nor  g2513 (n2415, n1796, n1292, n1614, n1822);
xor  g2514 (n2341, n1312, n1481, n1434, n1671);
nand g2515 (n2597, n723, n2018, n1771, n840);
xor  g2516 (n2180, n1852, n2059, n1976, n834);
xor  g2517 (n2324, n1789, n1082, n1725, n2062);
or   g2518 (n2147, n1672, n1907, n1965, n1875);
nor  g2519 (n2552, n1388, n770, n1256, n1780);
nand g2520 (n2689, n1646, n1465, n1330, n1830);
nand g2521 (n2374, n1807, n1885, n764, n1941);
nor  g2522 (n2240, n804, n1724, n1770, n971);
and  g2523 (n2706, n2069, n1806, n1556, n716);
xnor g2524 (n2334, n1359, n1786, n2012, n1846);
nor  g2525 (n2178, n1441, n2067, n1808, n1734);
nor  g2526 (n2289, n812, n1749, n1773, n919);
or   g2527 (n2378, n1972, n1538, n1365, n800);
or   g2528 (n2298, n1930, n1620, n1992, n2040);
or   g2529 (n2375, n991, n1270, n1611, n1829);
and  g2530 (n2536, n1564, n1398, n1333, n1322);
and  g2531 (n2273, n1555, n1710, n1351, n1170);
nor  g2532 (n2215, n1964, n2058, n1469, n780);
or   g2533 (n2247, n2011, n1330, n1533, n1871);
or   g2534 (n2162, n1819, n1545, n1993, n2013);
xnor g2535 (n2332, n1265, n1732, n1977, n1638);
nand g2536 (n2276, n747, n1772, n784, n1841);
nand g2537 (n2331, n1175, n2036, n1831, n1524);
and  g2538 (n2131, n1308, n1910, n1521, n989);
nand g2539 (n2257, n1798, n1591, n2057, n1636);
xnor g2540 (n2376, n1603, n1047, n1677, n1989);
and  g2541 (n2124, n1372, n1294, n1208, n2056);
nand g2542 (n2087, n1140, n2055, n1751, n1732);
xnor g2543 (n2626, n1959, n1899, n1445, n673);
nor  g2544 (n2530, n1493, n1414, n808, n1741);
and  g2545 (n2160, n1530, n1627, n1526, n1950);
nor  g2546 (n2503, n1648, n842, n1317, n830);
and  g2547 (n2282, n1870, n1453, n1621, n1961);
or   g2548 (n2355, n1669, n1864, n1725, n1663);
nor  g2549 (n2630, n891, n1223, n2034, n1268);
and  g2550 (n2317, n1529, n1879, n987, n1420);
and  g2551 (n2349, n1834, n706, n1544, n1638);
or   g2552 (n2709, n1790, n1087, n1541, n1665);
xor  g2553 (n2440, n1866, n1628, n871, n1472);
and  g2554 (n2544, n1355, n1889, n1696, n1424);
nand g2555 (n2561, n1356, n1753, n1679, n1216);
or   g2556 (n2244, n2029, n1427, n1677, n1826);
nand g2557 (n2566, n1960, n823, n2068, n805);
or   g2558 (n2480, n1876, n1693, n1229, n2069);
and  g2559 (n2666, n1991, n893, n1901, n1701);
and  g2560 (n2392, n1061, n1496, n704, n1552);
nand g2561 (n2446, n1052, n1296, n1438, n1770);
and  g2562 (n2152, n1962, n1728, n1505, n1363);
xnor g2563 (n2473, n691, n1280, n1706, n1712);
and  g2564 (n2287, n1639, n1966, n2067, n937);
xor  g2565 (n2674, n1758, n1716, n1454, n1970);
nand g2566 (n2153, n2051, n1377, n1104, n1991);
nand g2567 (n2121, n1830, n1044, n1592, n785);
or   g2568 (n2119, n1885, n1099, n1939, n1241);
nand g2569 (n2320, n1975, n2064, n1985, n1989);
and  g2570 (n2671, n1843, n883, n1758, n1742);
and  g2571 (n2159, n1506, n1063, n900, n1575);
nor  g2572 (n2099, n1945, n1866, n2006, n1878);
nand g2573 (n2258, n967, n2046, n1663, n1394);
nor  g2574 (n2239, n1522, n1425, n714, n740);
nor  g2575 (n2128, n1498, n1200, n1794, n1361);
nand g2576 (n2307, n2028, n844, n1872, n1619);
nor  g2577 (n2517, n1947, n1507, n1174, n2069);
nand g2578 (n2094, n1446, n838, n679, n1583);
nor  g2579 (n2572, n1198, n1746, n1902, n820);
and  g2580 (n2161, n2017, n2016, n1320, n905);
nor  g2581 (n2612, n1547, n1106, n1433, n921);
nor  g2582 (n2140, n2047, n675, n1992, n2043);
and  g2583 (n2138, n1372, n1227, n999, n1805);
and  g2584 (n2248, n1148, n2041, n1957, n819);
and  g2585 (n2499, n2054, n1282, n1970, n1823);
xnor g2586 (n2381, n2026, n1607, n1299, n973);
nand g2587 (n2224, n938, n727, n1482, n1984);
xnor g2588 (n2192, n1060, n1437, n1328, n1984);
xor  g2589 (n2356, n807, n1021, n1733, n1387);
xnor g2590 (n2419, n1958, n1983, n1944, n1846);
nor  g2591 (n2125, n976, n1956, n1949, n1300);
or   g2592 (n2199, n1347, n1298, n833, n2006);
and  g2593 (n2256, n1023, n729, n1678, n1183);
xnor g2594 (n2579, n1567, n1046, n2038, n1364);
or   g2595 (n2343, n683, n1745, n1281, n1026);
nand g2596 (n2708, n1062, n1572, n2035, n1324);
and  g2597 (n2351, n1789, n2019, n1687, n1787);
nor  g2598 (n2427, n829, n979, n1221, n1845);
nand g2599 (n2417, n1031, n776, n1995, n1976);
xor  g2600 (n2611, n1961, n2011, n1006, n841);
xnor g2601 (n2643, n749, n1931, n1608, n994);
or   g2602 (n2315, n1975, n2015, n1295, n1490);
xor  g2603 (n2462, n2052, n1806, n1092, n1983);
or   g2604 (n2426, n1434, n1906, n1426, n1071);
or   g2605 (n2663, n1028, n908, n1471, n1253);
or   g2606 (n2531, n1780, n1024, n1144, n1966);
and  g2607 (n2569, n2032, n1946, n2063, n1204);
nand g2608 (n2186, n1321, n739, n1896, n695);
xnor g2609 (n2357, n1692, n1856, n1292, n1924);
xnor g2610 (n2484, n1707, n1590, n1494, n1303);
or   g2611 (n2189, n1649, n839, n1208, n1390);
nand g2612 (n2142, n1958, n1768, n1436, n1582);
nor  g2613 (n2562, n1856, n1577, n1662, n1284);
nand g2614 (n2625, n1824, n2016, n1844, n1785);
nand g2615 (n2163, n1609, n1075, n1571, n1687);
or   g2616 (n2083, n1698, n944, n1423, n955);
nor  g2617 (n2512, n700, n1053, n1681, n1814);
xnor g2618 (n2644, n892, n1199, n818, n1627);
nand g2619 (n2337, n1261, n1659, n1448, n1956);
and  g2620 (n2487, n1171, n1459, n1775, n2033);
nand g2621 (n2458, n1522, n1381, n1754, n1240);
and  g2622 (n2101, n1158, n1504, n885, n1717);
nor  g2623 (n2397, n1693, n1259, n1567, n1514);
nor  g2624 (n2640, n1398, n1387, n1813, n1518);
xor  g2625 (n2141, n1468, n870, n2061, n1647);
xnor g2626 (n2118, n1942, n1872, n2032, n1938);
and  g2627 (n2703, n1755, n1185, n1452, n1985);
nand g2628 (n2406, n2061, n822, n1222, n1486);
nand g2629 (n2242, n1346, n1336, n2055, n1689);
nand g2630 (n2203, n1391, n1014, n2014, n1631);
xnor g2631 (n2556, n1753, n1933, n2071, n1801);
and  g2632 (n2699, n709, n1374, n1995, n1469);
xnor g2633 (n2546, n1793, n2034, n1860, n1993);
xor  g2634 (n2604, n1980, n1746, n1838, n1498);
xnor g2635 (n2454, n721, n1652, n1465, n1557);
or   g2636 (n2655, n1108, n1838, n1900, n1539);
and  g2637 (n2431, n1898, n1707, n1719, n1720);
or   g2638 (n2471, n1922, n1803, n1358, n1754);
or   g2639 (n2413, n1700, n1585, n1926, n1396);
nand g2640 (n2528, n1354, n1484, n1547, n1779);
nor  g2641 (n2677, n1715, n1392, n1005, n1820);
or   g2642 (n2452, n1731, n1322, n724, n2048);
nand g2643 (n2225, n2022, n737, n966, n1760);
and  g2644 (n2482, n1450, n789, n1219, n1922);
or   g2645 (n2399, n1122, n993, n1708, n2053);
xnor g2646 (n2100, n1703, n2060, n1578, n1942);
nor  g2647 (n2098, n1491, n1226, n1419, n1102);
nand g2648 (n2472, n1812, n831, n1430, n1244);
nand g2649 (n2660, n1943, n984, n1501, n1263);
xnor g2650 (n2091, n1400, n958, n2065, n1695);
xnor g2651 (n2665, n1204, n1967, n1466, n2013);
and  g2652 (n2326, n1512, n1432, n1997, n1473);
xor  g2653 (n2543, n1406, n1955, n756, n1565);
xor  g2654 (n2196, n1198, n1303, n828, n736);
or   g2655 (n2132, n964, n1258, n1232, n1944);
nor  g2656 (n2190, n1831, n1884, n1748, n1126);
nand g2657 (n2624, n1129, n1500, n1680, n1461);
xnor g2658 (n2447, n1353, n2051, n2021, n1273);
or   g2659 (n2251, n1532, n1612, n1323, n2054);
or   g2660 (n2680, n748, n923, n1565, n1695);
xnor g2661 (n2656, n1432, n1593, n1294, n970);
nor  g2662 (n2713, n1726, n1357, n2045, n1916);
nand g2663 (n2325, n1674, n1905, n1975, n1759);
or   g2664 (n2327, n1542, n1912, n1410, n997);
xnor g2665 (n2676, n1399, n1247, n1094, n1128);
xor  g2666 (n2410, n1149, n1430, n2039, n1153);
nor  g2667 (n2293, n953, n1664, n1553, n1985);
nor  g2668 (n2133, n2008, n2029, n1574, n686);
xor  g2669 (n2283, n1928, n1083, n1641, n1492);
nand g2670 (n2637, n1890, n2040, n1409, n2039);
nand g2671 (n2181, n1895, n1059, n1369, n1713);
and  g2672 (n2353, n1615, n1235, n1007, n1832);
or   g2673 (n2594, n2060, n1987, n1439, n1635);
or   g2674 (n2678, n1941, n681, n1164, n1537);
nand g2675 (n2586, n1321, n1307, n1291, n1243);
xnor g2676 (n2609, n1141, n1971, n1011, n1973);
xor  g2677 (n2269, n1891, n1408, n791);
xor  g2678 (n2253, n1070, n1702, n898, n925);
nor  g2679 (n2610, n767, n1842, n1488, n1310);
nor  g2680 (n2164, n1117, n1445, n1201, n1790);
or   g2681 (n2636, n1744, n974, n1954, n1800);
or   g2682 (n2502, n1362, n1086, n1755, n1423);
and  g2683 (n2492, n1118, n1568, n1854, n1788);
xor  g2684 (n2208, n1156, n1955, n1375, n1882);
nor  g2685 (n2838, n2459, n2119, n2415, n2313);
xor  g2686 (n2777, n2593, n2333, n2660, n2406);
and  g2687 (n2839, n2407, n2591, n2225, n2417);
xnor g2688 (n2797, n2485, n2267, n2128, n2602);
nand g2689 (n2778, n2305, n2255, n2228, n2444);
nand g2690 (n2727, n2588, n2641, n2413, n2293);
or   g2691 (n2825, n2408, n2283, n2546, n2149);
and  g2692 (n2800, n2645, n2087, n2650, n2535);
or   g2693 (n2781, n2322, n2200, n2531, n2093);
and  g2694 (n2834, n2245, n2501, n2506, n2232);
or   g2695 (n2785, n2532, n2102, n2152, n2632);
xor  g2696 (n2842, n2140, n2458, n2321, n2170);
xor  g2697 (n2815, n2375, n2630, n2211, n2499);
xor  g2698 (n2721, n2095, n2190, n2668, n2347);
or   g2699 (n2734, n2442, n2478, n2520, n2303);
or   g2700 (n2789, n2625, n2183, n2278, n2428);
xnor g2701 (n2854, n2577, n2636, n2615, n2503);
nand g2702 (n2749, n2441, n2493, n2560, n2388);
nand g2703 (n2786, n2435, n2171, n2178, n2542);
and  g2704 (n2840, n2513, n2622, n2440, n2304);
xor  g2705 (n2809, n2623, n2184, n2130, n2646);
xnor g2706 (n2771, n2116, n2617, n2374, n2666);
and  g2707 (n2858, n2292, n2248, n2164, n2551);
or   g2708 (n2822, n2567, n2133, n2341, n2165);
nor  g2709 (n2719, n2157, n2421, n2146, n2123);
and  g2710 (n2804, n2371, n2420, n2656, n2181);
and  g2711 (n2843, n2176, n2483, n2271, n2664);
nand g2712 (n2752, n2234, n2576, n2192, n2436);
nor  g2713 (n2799, n2505, n2628, n2174, n2383);
nand g2714 (n2864, n2302, n2151, n2195, n2422);
or   g2715 (n2803, n2318, n2295, n2601, n2574);
xnor g2716 (n2848, n2509, n2162, n2193, n2261);
nand g2717 (n2754, n2541, n2455, n2471, n2522);
or   g2718 (n2783, n2584, n2468, n2312, n2453);
xnor g2719 (n2852, n2543, n2653, n2237, n2160);
nand g2720 (n2790, n2224, n2568, n2284, n2662);
xnor g2721 (n2718, n2308, n2629, n2495, n2398);
nor  g2722 (n2773, n2215, n2605, n2536, n2206);
xor  g2723 (n2757, n2401, n2382, n2640, n2222);
nand g2724 (n2813, n2131, n2434, n2356, n2581);
xnor g2725 (n2782, n2381, n2166, n2239, n2517);
or   g2726 (n2729, n2595, n2296, n2363, n2275);
xor  g2727 (n2796, n2092, n2379, n2502, n2419);
nand g2728 (n2740, n2614, n2547, n2533, n2335);
and  g2729 (n2816, n2571, n2175, n2186, n2583);
or   g2730 (n2821, n2610, n2241, n2085, n2279);
nand g2731 (n2850, n2558, n2418, n2226, n2231);
nand g2732 (n2772, n2639, n2367, n2518, n2187);
xor  g2733 (n2730, n2624, n2243, n2125, n2603);
and  g2734 (n2732, n2438, n2479, n2477, n2212);
nand g2735 (n2831, n2300, n2566, n2462, n2349);
and  g2736 (n2859, n2525, n2516, n2124, n2384);
nor  g2737 (n2792, n2208, n2217, n2665, n2526);
xor  g2738 (n2829, n2557, n2627, n2207, n2270);
xor  g2739 (n2728, n2476, n2613, n2445, n2621);
xnor g2740 (n2806, n2652, n2334, n2142, n2238);
and  g2741 (n2764, n2528, n2262, n2219, n2655);
nor  g2742 (n2794, n2161, n2544, n2562, n2088);
xor  g2743 (n2826, n2463, n2365, n2253, n2553);
and  g2744 (n2725, n2592, n2490, n2556, n2600);
nand g2745 (n2737, n2530, n2108, n2307, n2488);
or   g2746 (n2779, n2514, n2395, n2281, n2089);
xnor g2747 (n2751, n2425, n2537, n2411, n2159);
and  g2748 (n2810, n2129, n2201, n2572, n2106);
xor  g2749 (n2793, n2529, n2155, n2297, n2147);
nor  g2750 (n2780, n2276, n2387, n2214, n2167);
xor  g2751 (n2856, n2378, n2386, n2127, n2635);
nor  g2752 (n2846, n2396, n2429, n2539, n2139);
or   g2753 (n2817, n2109, n2482, n2469, n2179);
or   g2754 (n2862, n2511, n2447, n2575, n2111);
nand g2755 (n2747, n2597, n2115, n2534, n2658);
or   g2756 (n2763, n2230, n2154, n2426, n2240);
nand g2757 (n2759, n2094, n2083, n2194, n2500);
or   g2758 (n2847, n2364, n2180, n2657, n2586);
xor  g2759 (n2860, n2585, n2353, n2389, n2258);
and  g2760 (n2745, n2310, n2663, n2661, n2504);
or   g2761 (n2724, n2216, n2524, n2481, n2096);
xnor g2762 (n2776, n2145, n2590, n2260, n2132);
or   g2763 (n2812, n2323, n2491, n2084, n2596);
nand g2764 (n2832, n2189, n2268, n2366, n2301);
and  g2765 (n2767, n2191, n2474, n2082, n2141);
xnor g2766 (n2723, n2229, n2319, n2105, n2550);
xor  g2767 (n2787, n2579, n2188, n2405, n2545);
and  g2768 (n2731, n2619, n2221, n2608, n2320);
nand g2769 (n2828, n2091, n2654, n2394, n2609);
nor  g2770 (n2805, n2117, n2285, n2570, n2336);
nand g2771 (n2791, n2246, n2594, n2362, n2265);
nand g2772 (n2765, n2327, n2137, n2100, n2134);
xor  g2773 (n2726, n2266, n2598, n2158, n2449);
nor  g2774 (n2849, n2559, n2377, n2252, n2390);
and  g2775 (n2807, n2647, n2642, n2359, n2244);
nor  g2776 (n2855, n2282, n2185, n2345, n2204);
and  g2777 (n2753, n2385, n2317, n2569, n2163);
nand g2778 (n2824, n2487, n2467, n2309, n2450);
or   g2779 (n2798, n2397, n2299, n2565, n2376);
xor  g2780 (n2774, n2330, n2196, n2173, n2393);
nand g2781 (n2857, n2637, n2430, n2644, n2409);
xnor g2782 (n2784, n2242, n2107, n2298, n2431);
nand g2783 (n2738, n2507, n2280, n2315, n2250);
xor  g2784 (n2762, n2669, n2182, n2649, n2348);
and  g2785 (n2770, n2291, n2203, n2472, n2475);
xor  g2786 (n2823, n2263, n2273, n2143, n2168);
xnor g2787 (n2801, n2314, n2099, n2667, n2324);
xor  g2788 (n2739, n2236, n2578, n2209, n2538);
nand g2789 (n2802, n2144, n2373, n2126, n2360);
nand g2790 (n2733, n2492, n2498, n2325, n2573);
nand g2791 (n2833, n2540, n2634, n2519, n2259);
nor  g2792 (n2811, n2361, n2090, n2486, n2549);
xor  g2793 (n2820, n2098, n2156, n2086, n2484);
nor  g2794 (n2844, n2512, n2294, n2424, n2112);
and  g2795 (n2736, n2358, n2523, n2249, n2510);
or   g2796 (n2769, n2494, n2332, n2254, n2172);
xor  g2797 (n2746, n2113, n2337, n2457, n2114);
xor  g2798 (n2835, n2218, n2210, n2552, n2351);
xnor g2799 (n2766, n2264, n2564, n2443, n2399);
xor  g2800 (n2768, n2344, n2412, n2256, n2343);
nand g2801 (n2830, n2150, n2169, n2631, n2451);
or   g2802 (n2722, n2121, n2651, n2439, n2205);
nor  g2803 (n2853, n2326, n2404, n2380, n2198);
xor  g2804 (n2795, n2508, n2247, n2097, n2464);
xor  g2805 (n2836, n2604, n2227, n2616, n2370);
nor  g2806 (n2788, n2311, n2350, n2612, n2354);
nor  g2807 (n2761, n2120, n2611, n2122, n2607);
xnor g2808 (n2744, n2480, n2582, n2177, n2352);
nor  g2809 (n2808, n2286, n2427, n2101, n2456);
xnor g2810 (n2827, n2620, n2233, n2515, n2223);
and  g2811 (n2760, n2497, n2138, n2342, n2153);
or   g2812 (n2742, n2339, n2400, n2432, n2287);
and  g2813 (n2748, n2410, n2606, n2340, n2489);
xnor g2814 (n2841, n2561, n2527, n2328, n2391);
xor  g2815 (n2818, n2460, n2554, n2638, n2355);
or   g2816 (n2720, n2461, n2118, n2466, n2306);
nand g2817 (n2861, n2357, n2496, n2135, n2369);
or   g2818 (n2755, n2288, n2274, n2433, n2437);
and  g2819 (n2743, n2213, n2563, n2220, n2316);
and  g2820 (n2735, n2148, n2103, n2423, n2372);
xnor g2821 (n2814, n2659, n2368, n2648, n2626);
or   g2822 (n2851, n2272, n2257, n2580, n2521);
nor  g2823 (n2845, n2329, n2587, n2465, n2392);
nor  g2824 (n2741, n2548, n2269, n2403, n2633);
or   g2825 (n2775, n2197, n2199, n2599, n2446);
nand g2826 (n2758, n2251, n2454, n2290, n2136);
and  g2827 (n2756, n2346, n2338, n2414, n2555);
and  g2828 (n2863, n2589, n2416, n2277, n2643);
nor  g2829 (n2837, n2331, n2448, n2202, n2402);
and  g2830 (n2819, n2473, n2289, n2104, n2110);
or   g2831 (n2750, n2470, n2618, n2235, n2452);
xor  g2832 (n2868, n2720, n2723, n2725, n2722);
and  g2833 (n2866, n2728, n2732, n2724, n2721);
and  g2834 (n2867, n2731, n2719, n2733, n2726);
nor  g2835 (n2865, n2718, n2730, n2727, n2729);
xor  g2836 (n2873, n2866, n2740, n2735, n2737);
xor  g2837 (n2871, n2671, n2672, n2670, n2674);
or   g2838 (n2870, n2866, n2738, n2865);
or   g2839 (n2869, n2675, n2734, n2739, n2741);
nor  g2840 (n2872, n2867, n2742, n2673, n2736);
nand g2841 (n2882, n2746, n2872, n2871, n2772);
and  g2842 (n2874, n2756, n2745, n2754, n2767);
xnor g2843 (n2883, n2759, n2750, n2762, n2749);
xor  g2844 (n2879, n2771, n2765, n2871, n2753);
xor  g2845 (n2875, n2869, n2764, n2744, n2770);
xnor g2846 (n2880, n2760, n2766, n2769, n2870);
xnor g2847 (n2878, n2747, n2743, n2752, n2872);
xnor g2848 (n2877, n2873, n2748, n2751, n2763);
or   g2849 (n2876, n2755, n2873, n2768, n2761);
nor  g2850 (n2881, n2873, n2873, n2757, n2758);
xor  g2851 (n2887, n2875, n2076, n2079, n2080);
xor  g2852 (n2884, n2078, n2078, n2073, n2072);
xnor g2853 (n2896, n2078, n2077, n2877, n2075);
or   g2854 (n2892, n2074, n2076, n2075, n2071);
xor  g2855 (n2895, n2074, n2073, n2879);
or   g2856 (n2885, n2074, n2080, n2075, n2077);
and  g2857 (n2894, n2080, n2879, n2874, n2072);
nand g2858 (n2891, n2076, n2081, n2878, n2077);
xor  g2859 (n2888, n2078, n2079, n2072, n2881);
xnor g2860 (n2889, n2074, n2878, n2077, n2876);
or   g2861 (n2890, n2080, n2880, n2882, n2079);
xnor g2862 (n2886, n2079, n2076, n2081, n2881);
xor  g2863 (n2893, n2880, n2075, n2072, n2073);
nand g2864 (n2899, n2884, n2888, n2684, n2887);
or   g2865 (n2901, n2681, n2683, n2774, n2688);
xnor g2866 (n2900, n2682, n2689, n2676, n2680);
xor  g2867 (n2902, n2889, n2690, n2886, n2679);
xnor g2868 (n2897, n2687, n2885, n2773, n2686);
nor  g2869 (n2898, n2775, n2678, n2677, n2685);
or   g2870 (n2903, n2902, n2776, n2780, n2777);
or   g2871 (n2904, n2901, n2779, n2781, n2778);
or   g2872 (n2905, n2903, n2693, n2692, n2691);
xor  g2873 (n2906, n2785, n2905, n2784, n2786);
nor  g2874 (n2907, n2783, n2787, n2782, n2905);
buf  g2875 (n2911, n2883);
buf  g2876 (n2909, n2906);
nand g2877 (n2908, n2904, n2907, n2882, n2906);
nor  g2878 (n2910, n2867, n2890, n2907, n2883);
or   g2879 (n2913, n2896, n2911, n2891, n2893);
or   g2880 (n2912, n2894, n2896);
and  g2881 (n2914, n2895, n2892, n2910, n2909);
not  g2882 (n2915, n2913);
buf  g2883 (n2916, n2915);
buf  g2884 (n2917, n2915);
xnor g2885 (n2918, n2914, n2917);
buf  g2886 (n2919, n2918);
buf  g2887 (n2920, n2918);
buf  g2888 (n2923, n2919);
buf  g2889 (n2924, n2920);
not  g2890 (n2922, n2920);
buf  g2891 (n2921, n2919);
not  g2892 (n2930, n2922);
not  g2893 (n2931, n2921);
not  g2894 (n2933, n2922);
buf  g2895 (n2929, n2922);
not  g2896 (n2925, n2923);
buf  g2897 (n2927, n2921);
buf  g2898 (n2926, n2922);
not  g2899 (n2928, n2918);
and  g2900 (n2932, n2918, n2921);
buf  g2901 (n2934, n2925);
buf  g2902 (n2935, n2925);
and  g2903 (n2938, n2924, n2934, n2935, n670);
nor  g2904 (n2939, n670, n669, n2934, n2924);
and  g2905 (n2941, n2924, n668, n669, n2923);
and  g2906 (n2942, n667, n2935, n2934, n669);
or   g2907 (n2937, n2924, n668, n2935);
xor  g2908 (n2940, n2935, n2923, n670);
xnor g2909 (n2936, n668, n2934, n669, n670);
xor  g2910 (n2950, n2938, n2926, n2941, n2700);
nand g2911 (n2946, n2929, n2928, n160, n2940);
or   g2912 (n2955, n2932, n2926, n2927, n2929);
or   g2913 (n2943, n2933, n2931, n2927);
nand g2914 (n2947, n2930, n2697, n2932);
nor  g2915 (n2952, n2929, n2695, n2927, n2931);
nand g2916 (n2944, n2928, n2933, n2936, n2939);
xor  g2917 (n2951, n2940, n2926, n2699, n2930);
xnor g2918 (n2948, n2698, n2933, n2938, n2942);
nor  g2919 (n2954, n2933, n2931, n2941, n160);
or   g2920 (n2945, n2930, n2932, n2927, n2939);
nor  g2921 (n2949, n2928, n2701, n2930, n2942);
nor  g2922 (n2956, n2929, n2694, n2696, n2928);
nand g2923 (n2953, n2937, n2942, n2926);
buf  g2924 (n2957, n2943);
and  g2925 (n2959, n2943, n2945, n2946, n2957);
or   g2926 (n2958, n2957, n2944, n2945);
buf  g2927 (n2962, n2948);
nand g2928 (n2961, n2946, n2958, n2947);
xnor g2929 (n2960, n2958, n2958, n2947, n2948);
nand g2930 (n2964, n2961, n2960, n2962);
xnor g2931 (n2963, n2962, n2961, n2949, n2960);
buf  g2932 (n2965, n2963);
buf  g2933 (n2967, n2965);
not  g2934 (n2966, n2965);
nand g2935 (n2971, n2868, n2950, n2952);
or   g2936 (n2970, n2959, n2949, n2967);
or   g2937 (n2975, n2959, n2868, n2966, n2967);
nor  g2938 (n2973, n2966, n2868, n2953);
xor  g2939 (n2968, n2966, n2953, n2951, n2959);
nor  g2940 (n2974, n2868, n2952, n2966, n2958);
nor  g2941 (n2969, n2951, n2952, n2967, n2959);
xnor g2942 (n2972, n2964, n2951, n2952);
not  g2943 (n2977, n2968);
not  g2944 (n2976, n2968);
buf  g2945 (n2978, n2976);
buf  g2946 (n2979, n2978);
buf  g2947 (n2980, n2978);
nor  g2948 (n2981, n2953, n2954, n2980, n2962);
xor  g2949 (n2983, n2964, n2981);
or   g2950 (n2982, n2968, n2964, n2981);
xor  g2951 (n2984, n2970, n2982, n2969);
xnor g2952 (n2985, n2968, n2970, n2969);
xnor g2953 (n2986, n2970, n2983);
nand g2954 (n2993, n2713, n2977, n2705, n2984);
nor  g2955 (n2996, n2703, n2977, n2984, n2717);
and  g2956 (n2992, n2985, n2986, n2955, n2984);
xor  g2957 (n2991, n2986, n2702, n2977);
xor  g2958 (n2987, n2985, n2715, n2956, n2709);
xor  g2959 (n2988, n2986, n2716, n2955, n2708);
nand g2960 (n2995, n2710, n2984, n2711, n2985);
nand g2961 (n2990, n2706, n2954, n2985, n2712);
and  g2962 (n2997, n2954, n2955, n2976);
and  g2963 (n2989, n2704, n2707, n2956, n2976);
or   g2964 (n2994, n2986, n2714, n2954, n2976);
nand g2965 (n3002, n2975, n2973, n2971, n2972);
nor  g2966 (n3003, n2971, n2974, n2972, n2975);
and  g2967 (n3001, n2972, n2995, n2973, n2974);
nor  g2968 (n3004, n2972, n2992, n2991, n2973);
and  g2969 (n2998, n2788, n2993, n2975);
nand g2970 (n3000, n2973, n2996, n2974);
nand g2971 (n2999, n2994, n2997, n2971);
and  g2972 (n3005, n2956, n3004);
xor  g2973 (n3006, n2789, n2800, n3005);
or   g2974 (n3009, n2790, n2794, n2793, n2795);
xnor g2975 (n3008, n2792, n2799, n3005, n2798);
and  g2976 (n3007, n2791, n2797, n2796, n3005);
nor  g2977 (n3011, n2801, n2810, n3008, n2807);
xor  g2978 (n3020, n2813, n3009, n3007, n2806);
xnor g2979 (n3015, n2818, n2803, n2804, n2827);
and  g2980 (n3014, n2808, n3007, n3009, n2802);
nor  g2981 (n3016, n2817, n2822, n3008, n2824);
nand g2982 (n3010, n2811, n2825, n2823, n2816);
xor  g2983 (n3018, n2831, n2805, n2956, n2821);
or   g2984 (n3013, n2819, n2828, n2830, n2814);
or   g2985 (n3012, n2820, n3008, n2809, n3009);
xnor g2986 (n3017, n3007, n2829, n2826, n2815);
xor  g2987 (n3019, n3009, n3008, n2812, n3007);
xor  g2988 (n3023, n2861, n3020, n3011, n2858);
nor  g2989 (n3026, n2859, n2840, n3013, n2839);
xnor g2990 (n3028, n3020, n2853, n3014, n2836);
and  g2991 (n3022, n2863, n2835, n2864, n3016);
and  g2992 (n3027, n2081, n2837, n2846, n2852);
xnor g2993 (n3029, n2862, n3015, n2841, n2854);
xor  g2994 (n3032, n3012, n2848, n2847, n3017);
nor  g2995 (n3021, n2843, n2845, n2832, n2849);
nor  g2996 (n3025, n2834, n2842, n2856, n2844);
nor  g2997 (n3031, n2833, n2850, n3020);
xor  g2998 (n3030, n3018, n3019, n2860, n2851);
xor  g2999 (n3024, n2081, n2838, n2855, n2857);
endmodule
