// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_183_517 written by SynthGen on 2021/05/24 19:47:14
module Stat_183_517( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26,
 n122, n171, n124, n178, n160, n125, n165, n177,
 n130, n208, n204, n192, n199, n203, n205, n198,
 n200, n197, n201, n195, n196, n209, n194, n207,
 n206, n202, n193);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26;

output n122, n171, n124, n178, n160, n125, n165, n177,
 n130, n208, n204, n192, n199, n203, n205, n198,
 n200, n197, n201, n195, n196, n209, n194, n207,
 n206, n202, n193;

wire n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n123,
 n126, n127, n128, n129, n131, n132, n133, n134,
 n135, n136, n137, n138, n139, n140, n141, n142,
 n143, n144, n145, n146, n147, n148, n149, n150,
 n151, n152, n153, n154, n155, n156, n157, n158,
 n159, n161, n162, n163, n164, n166, n167, n168,
 n169, n170, n172, n173, n174, n175, n176, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n189, n190, n191;

not  g0 (n54, n8);
not  g1 (n61, n23);
not  g2 (n64, n10);
buf  g3 (n72, n1);
buf  g4 (n28, n17);
not  g5 (n73, n9);
not  g6 (n80, n14);
not  g7 (n91, n8);
buf  g8 (n77, n4);
buf  g9 (n79, n19);
buf  g10 (n56, n10);
not  g11 (n57, n11);
buf  g12 (n47, n19);
not  g13 (n50, n7);
not  g14 (n37, n5);
buf  g15 (n90, n20);
not  g16 (n41, n4);
not  g17 (n97, n23);
not  g18 (n55, n7);
not  g19 (n86, n12);
not  g20 (n30, n3);
buf  g21 (n84, n1);
not  g22 (n70, n9);
not  g23 (n78, n20);
buf  g24 (n66, n13);
not  g25 (n69, n14);
not  g26 (n71, n22);
buf  g27 (n32, n24);
not  g28 (n58, n6);
buf  g29 (n53, n20);
not  g30 (n42, n2);
buf  g31 (n76, n11);
buf  g32 (n49, n3);
buf  g33 (n83, n16);
not  g34 (n92, n17);
not  g35 (n40, n22);
not  g36 (n38, n11);
buf  g37 (n59, n6);
buf  g38 (n33, n2);
buf  g39 (n63, n5);
not  g40 (n62, n8);
not  g41 (n36, n14);
buf  g42 (n96, n15);
buf  g43 (n87, n21);
not  g44 (n39, n1);
not  g45 (n29, n6);
not  g46 (n68, n5);
not  g47 (n27, n13);
not  g48 (n44, n13);
buf  g49 (n74, n18);
buf  g50 (n88, n10);
buf  g51 (n34, n7);
buf  g52 (n45, n3);
buf  g53 (n43, n4);
buf  g54 (n60, n9);
not  g55 (n51, n18);
not  g56 (n35, n15);
buf  g57 (n48, n17);
buf  g58 (n52, n16);
not  g59 (n67, n23);
buf  g60 (n75, n16);
buf  g61 (n95, n18);
buf  g62 (n89, n15);
buf  g63 (n82, n12);
not  g64 (n98, n21);
buf  g65 (n81, n12);
buf  g66 (n31, n24);
buf  g67 (n46, n2);
not  g68 (n65, n22);
not  g69 (n94, n21);
not  g70 (n93, n24);
buf  g71 (n85, n19);
not  g72 (n109, n30);
not  g73 (n110, n29);
not  g74 (n111, n33);
buf  g75 (n106, n34);
buf  g76 (n115, n31);
not  g77 (n118, n26);
not  g78 (n108, n28);
buf  g79 (n119, n27);
not  g80 (n114, n25);
not  g81 (n107, n30);
not  g82 (n99, n26);
buf  g83 (n105, n26);
buf  g84 (n102, n29);
buf  g85 (n120, n25);
buf  g86 (n100, n31);
not  g87 (n104, n32);
buf  g88 (n101, n27);
buf  g89 (n117, n31);
buf  g90 (n103, n33);
buf  g91 (n112, n32);
xnor g92 (n116, n30, n27, n32, n28);
nor  g93 (n113, n33, n28, n25, n29);
and  g94 (n128, n49, n116, n95);
or   g95 (n142, n42, n94, n113, n107);
or   g96 (n160, n51, n69, n100, n60);
or   g97 (n138, n83, n60, n79, n42);
xnor g98 (n149, n61, n66, n79, n56);
nor  g99 (n147, n79, n94, n103, n73);
and  g100 (n151, n82, n86, n109, n93);
nor  g101 (n137, n50, n72, n41, n45);
xor  g102 (n124, n51, n55, n57, n117);
nand g103 (n179, n104, n108, n77, n41);
nand g104 (n126, n72, n54, n53, n47);
nor  g105 (n184, n43, n48, n40, n117);
and  g106 (n182, n62, n80, n53, n82);
xnor g107 (n158, n113, n85, n64, n115);
xor  g108 (n125, n36, n72, n78, n89);
or   g109 (n134, n81, n82, n69, n84);
xor  g110 (n172, n46, n114, n115, n108);
or   g111 (n122, n77, n68, n80, n78);
and  g112 (n139, n50, n43, n99, n68);
and  g113 (n157, n93, n110, n100, n92);
nand g114 (n135, n87, n88, n71, n99);
or   g115 (n156, n86, n111, n87, n73);
and  g116 (n178, n96, n76, n36, n52);
nor  g117 (n171, n100, n38, n92, n34);
xor  g118 (n153, n112, n93, n47, n89);
or   g119 (n175, n103, n58, n88, n85);
xnor g120 (n166, n112, n96, n75, n99);
or   g121 (n162, n83, n49, n67, n35);
xnor g122 (n155, n101, n84, n60, n61);
or   g123 (n145, n103, n53, n106, n49);
nand g124 (n130, n59, n54, n62, n104);
nand g125 (n144, n106, n107, n105, n114);
nor  g126 (n133, n78, n120, n70, n59);
xnor g127 (n127, n68, n57, n46, n64);
xnor g128 (n165, n35, n67, n76, n91);
nor  g129 (n164, n111, n39, n63, n44);
xor  g130 (n123, n112, n88, n44, n38);
and  g131 (n152, n81, n71, n111, n65);
nor  g132 (n163, n74, n66, n118, n51);
xor  g133 (n169, n90, n90, n39, n84);
nor  g134 (n143, n59, n104, n118, n63);
nor  g135 (n140, n108, n62, n113, n52);
xnor g136 (n183, n97, n87, n55, n98);
nor  g137 (n180, n58, n63, n119, n55);
nand g138 (n129, n44, n95, n98, n97);
xor  g139 (n141, n102, n75, n71, n45);
nand g140 (n181, n74, n80, n118, n101);
xor  g141 (n168, n102, n95, n61, n40);
or   g142 (n121, n36, n57, n109, n120);
xnor g143 (n185, n90, n86, n47, n117);
nor  g144 (n136, n83, n56, n75, n98);
xnor g145 (n131, n119, n74, n39, n69);
xor  g146 (n177, n64, n35, n38, n34);
xor  g147 (n148, n107, n102, n37, n65);
and  g148 (n176, n54, n94, n45, n89);
xor  g149 (n173, n48, n110, n81);
or   g150 (n170, n76, n97, n92, n109);
or   g151 (n146, n91, n105, n66, n40);
and  g152 (n174, n46, n37, n65, n77);
nand g153 (n159, n67, n50, n115, n91);
and  g154 (n132, n114, n73, n116, n96);
or   g155 (n154, n58, n42, n119, n56);
or   g156 (n161, n101, n37, n70, n106);
nand g157 (n150, n85, n105, n48, n52);
nand g158 (n167, n41, n116, n70, n43);
buf  g159 (n191, n131);
buf  g160 (n186, n132);
buf  g161 (n190, n120);
not  g162 (n189, n134);
buf  g163 (n188, n133);
or   g164 (n187, n135, n130);
nor  g165 (n206, n139, n164, n150, n191);
nand g166 (n208, n190, n143, n159, n191);
xor  g167 (n195, n187, n187, n144, n178);
xor  g168 (n200, n176, n188, n163, n160);
or   g169 (n194, n165, n138, n167, n181);
xnor g170 (n198, n166, n189, n171, n186);
nor  g171 (n207, n172, n157, n151, n174);
or   g172 (n209, n190, n191, n185, n155);
nor  g173 (n205, n187, n145, n190, n149);
or   g174 (n201, n189, n185, n175, n156);
xor  g175 (n202, n148, n184, n146);
or   g176 (n203, n140, n185, n162, n137);
nand g177 (n197, n184, n189, n186, n153);
nor  g178 (n192, n173, n169, n186, n161);
xor  g179 (n196, n188, n136, n147, n177);
xor  g180 (n204, n179, n142, n141, n154);
or   g181 (n199, n158, n182, n170, n152);
nor  g182 (n193, n168, n188, n183, n180);
endmodule
