// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_301 written by SynthGen on 2021/04/05 11:23:27
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_301 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1518, n1517, n1533, n2029, n2025, n2020, n2010, n2031,
 n2008, n2028, n2012, n2027, n2022, n2030, n2006, n2024,
 n2032, n2018, n2009, n2021, n2016, n2013, n2023, n2005,
 n2026, n2014, n2011, n2017, n2004, n2019, n2007, n2015);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1518, n1517, n1533, n2029, n2025, n2020, n2010, n2031,
 n2008, n2028, n2012, n2027, n2022, n2030, n2006, n2024,
 n2032, n2018, n2009, n2021, n2016, n2013, n2023, n2005,
 n2026, n2014, n2011, n2017, n2004, n2019, n2007, n2015;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1534, n1535, n1536, n1537, n1538, n1539,
 n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
 n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
 n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
 n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
 n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
 n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
 n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
 n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
 n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
 n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
 n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
 n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
 n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
 n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
 n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
 n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
 n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
 n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
 n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
 n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
 n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
 n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
 n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
 n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
 n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
 n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
 n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
 n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
 n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
 n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
 n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
 n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
 n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
 n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
 n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
 n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
 n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
 n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
 n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
 n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
 n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
 n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
 n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
 n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
 n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
 n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
 n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
 n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
 n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
 n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
 n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
 n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
 n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
 n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
 n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
 n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
 n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
 n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;

not  g0 (n40, n13);
buf  g1 (n93, n21);
buf  g2 (n83, n29);
not  g3 (n149, n8);
not  g4 (n72, n19);
buf  g5 (n122, n31);
not  g6 (n45, n18);
buf  g7 (n53, n23);
not  g8 (n73, n7);
not  g9 (n139, n25);
not  g10 (n92, n32);
buf  g11 (n87, n32);
not  g12 (n39, n11);
not  g13 (n127, n24);
buf  g14 (n42, n11);
buf  g15 (n134, n11);
not  g16 (n84, n15);
not  g17 (n154, n5);
not  g18 (n75, n16);
buf  g19 (n68, n30);
not  g20 (n88, n25);
buf  g21 (n47, n24);
buf  g22 (n150, n12);
not  g23 (n77, n27);
not  g24 (n36, n14);
not  g25 (n111, n3);
buf  g26 (n58, n26);
buf  g27 (n34, n28);
not  g28 (n144, n10);
buf  g29 (n74, n8);
not  g30 (n104, n9);
not  g31 (n56, n2);
not  g32 (n138, n17);
buf  g33 (n69, n6);
not  g34 (n119, n12);
not  g35 (n136, n11);
not  g36 (n98, n31);
not  g37 (n86, n18);
not  g38 (n35, n7);
buf  g39 (n116, n10);
not  g40 (n153, n25);
not  g41 (n157, n21);
buf  g42 (n85, n31);
buf  g43 (n79, n14);
not  g44 (n33, n22);
not  g45 (n102, n28);
not  g46 (n126, n17);
buf  g47 (n94, n27);
buf  g48 (n140, n23);
not  g49 (n62, n3);
not  g50 (n135, n4);
not  g51 (n55, n29);
not  g52 (n115, n18);
buf  g53 (n108, n30);
buf  g54 (n142, n18);
not  g55 (n123, n10);
buf  g56 (n160, n15);
not  g57 (n89, n5);
not  g58 (n107, n26);
not  g59 (n82, n6);
not  g60 (n132, n22);
not  g61 (n103, n2);
not  g62 (n110, n29);
buf  g63 (n51, n14);
buf  g64 (n120, n5);
not  g65 (n67, n20);
buf  g66 (n97, n2);
buf  g67 (n151, n10);
not  g68 (n60, n1);
buf  g69 (n129, n13);
buf  g70 (n146, n7);
buf  g71 (n99, n4);
not  g72 (n143, n6);
buf  g73 (n91, n16);
not  g74 (n137, n27);
not  g75 (n59, n15);
buf  g76 (n121, n5);
not  g77 (n96, n21);
not  g78 (n61, n17);
buf  g79 (n95, n23);
not  g80 (n57, n16);
buf  g81 (n156, n13);
buf  g82 (n113, n26);
buf  g83 (n125, n16);
not  g84 (n90, n25);
not  g85 (n128, n9);
not  g86 (n152, n22);
not  g87 (n105, n19);
buf  g88 (n41, n13);
not  g89 (n112, n23);
buf  g90 (n117, n4);
buf  g91 (n78, n1);
not  g92 (n106, n6);
not  g93 (n48, n28);
not  g94 (n141, n31);
buf  g95 (n64, n2);
not  g96 (n46, n9);
buf  g97 (n148, n1);
buf  g98 (n101, n3);
buf  g99 (n37, n20);
not  g100 (n65, n19);
not  g101 (n70, n7);
not  g102 (n80, n19);
not  g103 (n50, n24);
buf  g104 (n44, n12);
not  g105 (n118, n30);
not  g106 (n38, n24);
not  g107 (n158, n32);
not  g108 (n71, n12);
not  g109 (n155, n26);
buf  g110 (n130, n20);
buf  g111 (n81, n9);
buf  g112 (n159, n4);
buf  g113 (n43, n14);
buf  g114 (n54, n21);
buf  g115 (n114, n1);
not  g116 (n49, n28);
buf  g117 (n145, n17);
buf  g118 (n124, n20);
not  g119 (n66, n22);
not  g120 (n52, n29);
not  g121 (n147, n8);
not  g122 (n109, n30);
not  g123 (n133, n8);
not  g124 (n76, n3);
not  g125 (n63, n15);
not  g126 (n131, n27);
not  g127 (n100, n32);
buf  g128 (n511, n105);
buf  g129 (n210, n47);
buf  g130 (n394, n41);
buf  g131 (n520, n150);
not  g132 (n221, n65);
not  g133 (n164, n124);
buf  g134 (n633, n89);
not  g135 (n576, n78);
buf  g136 (n339, n114);
buf  g137 (n577, n57);
not  g138 (n224, n138);
not  g139 (n215, n72);
buf  g140 (n338, n66);
not  g141 (n165, n60);
buf  g142 (n312, n116);
not  g143 (n575, n145);
buf  g144 (n260, n100);
not  g145 (n631, n149);
buf  g146 (n421, n97);
not  g147 (n168, n134);
not  g148 (n516, n69);
not  g149 (n550, n124);
buf  g150 (n632, n128);
buf  g151 (n569, n73);
not  g152 (n202, n66);
buf  g153 (n341, n38);
not  g154 (n375, n81);
buf  g155 (n494, n76);
buf  g156 (n248, n130);
buf  g157 (n386, n142);
buf  g158 (n234, n84);
buf  g159 (n324, n136);
not  g160 (n560, n117);
not  g161 (n602, n146);
buf  g162 (n601, n109);
buf  g163 (n505, n99);
not  g164 (n189, n45);
not  g165 (n423, n124);
not  g166 (n586, n144);
buf  g167 (n497, n129);
buf  g168 (n597, n97);
not  g169 (n486, n75);
not  g170 (n384, n107);
buf  g171 (n469, n152);
not  g172 (n618, n52);
buf  g173 (n351, n121);
not  g174 (n363, n142);
not  g175 (n651, n153);
not  g176 (n193, n115);
buf  g177 (n639, n141);
not  g178 (n211, n98);
buf  g179 (n462, n46);
not  g180 (n329, n37);
not  g181 (n173, n42);
buf  g182 (n258, n42);
buf  g183 (n171, n105);
not  g184 (n656, n116);
buf  g185 (n416, n91);
not  g186 (n245, n33);
buf  g187 (n181, n128);
not  g188 (n251, n82);
not  g189 (n587, n63);
buf  g190 (n540, n122);
buf  g191 (n395, n111);
buf  g192 (n390, n149);
not  g193 (n368, n86);
not  g194 (n412, n82);
buf  g195 (n238, n160);
not  g196 (n428, n152);
not  g197 (n549, n48);
buf  g198 (n242, n119);
not  g199 (n222, n99);
not  g200 (n317, n103);
buf  g201 (n273, n43);
buf  g202 (n272, n129);
buf  g203 (n647, n127);
buf  g204 (n567, n37);
not  g205 (n483, n36);
buf  g206 (n356, n88);
buf  g207 (n225, n85);
not  g208 (n182, n78);
buf  g209 (n452, n126);
buf  g210 (n485, n155);
not  g211 (n546, n86);
buf  g212 (n169, n123);
buf  g213 (n366, n34);
not  g214 (n642, n98);
not  g215 (n187, n41);
buf  g216 (n596, n49);
not  g217 (n345, n148);
not  g218 (n545, n74);
not  g219 (n233, n158);
not  g220 (n209, n54);
not  g221 (n568, n159);
not  g222 (n410, n57);
buf  g223 (n574, n144);
buf  g224 (n229, n106);
not  g225 (n327, n47);
buf  g226 (n179, n76);
buf  g227 (n319, n146);
buf  g228 (n203, n72);
buf  g229 (n277, n121);
buf  g230 (n358, n90);
not  g231 (n623, n79);
buf  g232 (n406, n140);
not  g233 (n611, n143);
buf  g234 (n279, n81);
buf  g235 (n268, n126);
not  g236 (n479, n88);
buf  g237 (n243, n106);
buf  g238 (n544, n125);
buf  g239 (n393, n80);
not  g240 (n638, n56);
buf  g241 (n609, n61);
not  g242 (n409, n113);
buf  g243 (n400, n41);
buf  g244 (n493, n87);
not  g245 (n509, n59);
not  g246 (n401, n71);
buf  g247 (n612, n38);
buf  g248 (n561, n45);
buf  g249 (n335, n150);
not  g250 (n413, n64);
buf  g251 (n392, n58);
buf  g252 (n526, n66);
buf  g253 (n298, n121);
buf  g254 (n269, n68);
not  g255 (n630, n88);
not  g256 (n590, n100);
not  g257 (n192, n127);
buf  g258 (n304, n123);
not  g259 (n226, n110);
not  g260 (n257, n50);
buf  g261 (n278, n55);
not  g262 (n201, n113);
not  g263 (n517, n48);
not  g264 (n283, n140);
buf  g265 (n239, n80);
not  g266 (n220, n118);
not  g267 (n660, n128);
not  g268 (n266, n93);
buf  g269 (n364, n87);
buf  g270 (n637, n149);
buf  g271 (n309, n37);
buf  g272 (n478, n39);
not  g273 (n342, n83);
buf  g274 (n161, n79);
not  g275 (n482, n101);
buf  g276 (n628, n93);
not  g277 (n391, n113);
buf  g278 (n565, n153);
not  g279 (n538, n69);
buf  g280 (n223, n112);
buf  g281 (n326, n133);
not  g282 (n383, n75);
buf  g283 (n484, n39);
not  g284 (n252, n139);
buf  g285 (n417, n48);
buf  g286 (n519, n117);
not  g287 (n175, n61);
not  g288 (n167, n53);
not  g289 (n343, n108);
not  g290 (n284, n70);
buf  g291 (n186, n40);
buf  g292 (n573, n135);
not  g293 (n231, n147);
not  g294 (n206, n100);
not  g295 (n228, n102);
buf  g296 (n473, n156);
not  g297 (n426, n152);
buf  g298 (n359, n156);
not  g299 (n434, n82);
buf  g300 (n604, n94);
buf  g301 (n330, n36);
not  g302 (n552, n66);
buf  g303 (n463, n96);
not  g304 (n293, n131);
not  g305 (n634, n125);
not  g306 (n619, n130);
buf  g307 (n643, n136);
buf  g308 (n502, n158);
not  g309 (n177, n92);
not  g310 (n652, n115);
buf  g311 (n296, n44);
buf  g312 (n444, n86);
not  g313 (n608, n60);
buf  g314 (n297, n138);
buf  g315 (n461, n96);
buf  g316 (n584, n94);
not  g317 (n344, n59);
not  g318 (n610, n45);
buf  g319 (n666, n131);
not  g320 (n476, n146);
buf  g321 (n453, n136);
buf  g322 (n492, n152);
not  g323 (n616, n155);
buf  g324 (n571, n39);
not  g325 (n454, n98);
not  g326 (n564, n89);
not  g327 (n337, n116);
buf  g328 (n289, n93);
not  g329 (n340, n125);
buf  g330 (n503, n157);
buf  g331 (n440, n131);
not  g332 (n262, n40);
not  g333 (n558, n62);
not  g334 (n504, n133);
not  g335 (n166, n74);
not  g336 (n606, n39);
not  g337 (n163, n64);
not  g338 (n559, n79);
buf  g339 (n301, n52);
not  g340 (n362, n43);
not  g341 (n305, n124);
not  g342 (n599, n44);
not  g343 (n236, n76);
buf  g344 (n665, n34);
buf  g345 (n667, n59);
buf  g346 (n672, n42);
buf  g347 (n589, n61);
buf  g348 (n240, n65);
buf  g349 (n331, n48);
not  g350 (n350, n64);
not  g351 (n532, n111);
buf  g352 (n582, n38);
buf  g353 (n622, n93);
buf  g354 (n276, n62);
not  g355 (n663, n145);
not  g356 (n365, n73);
buf  g357 (n661, n103);
buf  g358 (n255, n141);
buf  g359 (n649, n55);
buf  g360 (n199, n125);
not  g361 (n624, n104);
not  g362 (n464, n150);
buf  g363 (n196, n145);
buf  g364 (n399, n126);
buf  g365 (n183, n135);
buf  g366 (n653, n123);
not  g367 (n377, n36);
not  g368 (n581, n78);
buf  g369 (n264, n35);
not  g370 (n360, n108);
not  g371 (n515, n95);
not  g372 (n411, n52);
buf  g373 (n455, n108);
not  g374 (n443, n102);
buf  g375 (n398, n84);
not  g376 (n379, n135);
not  g377 (n306, n133);
not  g378 (n372, n64);
buf  g379 (n354, n49);
buf  g380 (n184, n77);
not  g381 (n525, n103);
not  g382 (n274, n88);
not  g383 (n530, n111);
not  g384 (n570, n49);
not  g385 (n408, n122);
buf  g386 (n265, n55);
buf  g387 (n563, n70);
not  g388 (n430, n138);
buf  g389 (n427, n107);
not  g390 (n246, n153);
not  g391 (n562, n65);
not  g392 (n466, n107);
buf  g393 (n543, n117);
not  g394 (n437, n130);
not  g395 (n635, n41);
not  g396 (n446, n109);
buf  g397 (n664, n37);
buf  g398 (n244, n35);
not  g399 (n347, n147);
not  g400 (n669, n67);
not  g401 (n627, n81);
not  g402 (n321, n72);
buf  g403 (n621, n127);
buf  g404 (n172, n103);
buf  g405 (n442, n65);
buf  g406 (n275, n157);
not  g407 (n548, n50);
not  g408 (n227, n54);
buf  g409 (n620, n78);
buf  g410 (n551, n135);
not  g411 (n303, n151);
not  g412 (n217, n140);
not  g413 (n374, n33);
not  g414 (n299, n120);
not  g415 (n605, n63);
buf  g416 (n369, n50);
buf  g417 (n332, n62);
buf  g418 (n650, n156);
buf  g419 (n470, n122);
buf  g420 (n598, n100);
not  g421 (n388, n34);
not  g422 (n370, n81);
not  g423 (n316, n95);
buf  g424 (n495, n159);
buf  g425 (n381, n95);
not  g426 (n445, n97);
buf  g427 (n522, n58);
not  g428 (n518, n115);
not  g429 (n194, n118);
not  g430 (n180, n160);
not  g431 (n636, n80);
buf  g432 (n472, n59);
not  g433 (n198, n54);
not  g434 (n349, n102);
buf  g435 (n389, n57);
buf  g436 (n310, n110);
not  g437 (n378, n102);
buf  g438 (n448, n76);
not  g439 (n555, n94);
not  g440 (n547, n154);
not  g441 (n415, n106);
not  g442 (n190, n49);
not  g443 (n241, n43);
buf  g444 (n314, n33);
buf  g445 (n407, n85);
not  g446 (n467, n77);
not  g447 (n556, n154);
buf  g448 (n441, n61);
buf  g449 (n281, n114);
buf  g450 (n334, n91);
not  g451 (n254, n84);
not  g452 (n641, n143);
not  g453 (n625, n153);
not  g454 (n496, n44);
not  g455 (n539, n150);
buf  g456 (n487, n85);
buf  g457 (n237, n95);
not  g458 (n500, n33);
not  g459 (n583, n87);
not  g460 (n655, n40);
not  g461 (n480, n101);
buf  g462 (n593, n77);
not  g463 (n535, n131);
buf  g464 (n528, n158);
buf  g465 (n458, n36);
buf  g466 (n536, n122);
not  g467 (n396, n132);
buf  g468 (n670, n129);
not  g469 (n318, n84);
buf  g470 (n585, n99);
not  g471 (n253, n155);
not  g472 (n195, n101);
buf  g473 (n214, n90);
buf  g474 (n307, n62);
buf  g475 (n527, n57);
buf  g476 (n501, n53);
buf  g477 (n270, n82);
buf  g478 (n449, n101);
buf  g479 (n475, n58);
not  g480 (n617, n109);
not  g481 (n197, n155);
buf  g482 (n510, n116);
buf  g483 (n592, n151);
buf  g484 (n422, n132);
buf  g485 (n591, n160);
buf  g486 (n282, n83);
buf  g487 (n603, n151);
not  g488 (n292, n112);
buf  g489 (n300, n47);
not  g490 (n185, n104);
not  g491 (n208, n104);
buf  g492 (n424, n99);
not  g493 (n235, n96);
buf  g494 (n512, n110);
buf  g495 (n523, n77);
buf  g496 (n267, n159);
buf  g497 (n419, n106);
buf  g498 (n614, n120);
buf  g499 (n213, n140);
buf  g500 (n320, n51);
not  g501 (n451, n114);
not  g502 (n465, n113);
not  g503 (n323, n115);
buf  g504 (n348, n46);
not  g505 (n205, n128);
buf  g506 (n600, n68);
not  g507 (n325, n44);
not  g508 (n506, n142);
not  g509 (n477, n96);
not  g510 (n657, n120);
buf  g511 (n488, n136);
buf  g512 (n554, n67);
buf  g513 (n380, n85);
not  g514 (n219, n141);
buf  g515 (n645, n92);
buf  g516 (n191, n138);
not  g517 (n468, n147);
not  g518 (n207, n132);
buf  g519 (n459, n79);
not  g520 (n566, n56);
not  g521 (n481, n154);
not  g522 (n382, n43);
not  g523 (n200, n137);
buf  g524 (n615, n119);
not  g525 (n346, n118);
buf  g526 (n230, n83);
buf  g527 (n232, n110);
not  g528 (n658, n120);
buf  g529 (n668, n108);
not  g530 (n218, n139);
buf  g531 (n367, n111);
buf  g532 (n439, n92);
not  g533 (n287, n35);
buf  g534 (n402, n119);
buf  g535 (n263, n52);
buf  g536 (n286, n134);
buf  g537 (n285, n149);
not  g538 (n542, n127);
buf  g539 (n537, n86);
buf  g540 (n435, n73);
buf  g541 (n438, n75);
buf  g542 (n403, n141);
buf  g543 (n302, n71);
buf  g544 (n534, n132);
buf  g545 (n216, n75);
buf  g546 (n397, n156);
buf  g547 (n414, n54);
buf  g548 (n328, n105);
buf  g549 (n271, n139);
buf  g550 (n170, n112);
not  g551 (n259, n90);
buf  g552 (n256, n134);
not  g553 (n294, n46);
not  g554 (n640, n143);
not  g555 (n489, n134);
buf  g556 (n204, n90);
buf  g557 (n429, n71);
buf  g558 (n247, n51);
not  g559 (n572, n89);
not  g560 (n514, n137);
buf  g561 (n280, n60);
buf  g562 (n595, n146);
not  g563 (n376, n118);
buf  g564 (n553, n91);
buf  g565 (n662, n87);
not  g566 (n594, n148);
not  g567 (n471, n105);
buf  g568 (n521, n157);
not  g569 (n433, n89);
buf  g570 (n371, n70);
not  g571 (n578, n55);
buf  g572 (n654, n158);
buf  g573 (n250, n104);
buf  g574 (n420, n139);
not  g575 (n533, n72);
not  g576 (n405, n50);
not  g577 (n557, n35);
not  g578 (n507, n68);
not  g579 (n425, n71);
not  g580 (n490, n63);
buf  g581 (n513, n42);
not  g582 (n322, n129);
not  g583 (n648, n56);
buf  g584 (n646, n114);
buf  g585 (n531, n51);
not  g586 (n404, n69);
buf  g587 (n671, n144);
buf  g588 (n541, n83);
not  g589 (n431, n73);
buf  g590 (n291, n46);
not  g591 (n607, n69);
buf  g592 (n188, n80);
not  g593 (n588, n40);
not  g594 (n353, n154);
not  g595 (n311, n112);
buf  g596 (n212, n68);
buf  g597 (n333, n67);
not  g598 (n176, n97);
not  g599 (n290, n53);
not  g600 (n474, n51);
not  g601 (n357, n91);
not  g602 (n460, n92);
not  g603 (n288, n117);
not  g604 (n456, n142);
not  g605 (n373, n45);
buf  g606 (n313, n126);
not  g607 (n315, n137);
not  g608 (n450, n159);
buf  g609 (n336, n123);
buf  g610 (n457, n133);
not  g611 (n436, n34);
buf  g612 (n174, n143);
buf  g613 (n629, n47);
buf  g614 (n644, n38);
buf  g615 (n579, n58);
not  g616 (n613, n145);
not  g617 (n361, n60);
not  g618 (n261, n160);
buf  g619 (n162, n98);
buf  g620 (n580, n63);
buf  g621 (n498, n74);
not  g622 (n355, n119);
not  g623 (n508, n137);
buf  g624 (n249, n147);
not  g625 (n418, n130);
buf  g626 (n659, n67);
not  g627 (n352, n148);
not  g628 (n499, n74);
buf  g629 (n295, n157);
buf  g630 (n447, n94);
buf  g631 (n524, n151);
not  g632 (n308, n144);
not  g633 (n387, n148);
not  g634 (n626, n109);
buf  g635 (n178, n70);
buf  g636 (n529, n107);
not  g637 (n385, n121);
not  g638 (n491, n56);
buf  g639 (n432, n53);
nand g640 (n695, n397, n518, n426, n668);
and  g641 (n1066, n331, n231, n435, n629);
xnor g642 (n777, n198, n655, n639, n621);
and  g643 (n778, n576, n422, n233, n183);
xor  g644 (n995, n662, n645, n171, n297);
nand g645 (n1121, n465, n351, n325, n355);
and  g646 (n979, n347, n554, n444, n252);
xor  g647 (n742, n620, n428, n484, n575);
xor  g648 (n679, n356, n608, n387, n571);
nand g649 (n826, n498, n478, n602, n212);
nor  g650 (n911, n524, n544, n355, n395);
or   g651 (n868, n275, n381, n436, n604);
nor  g652 (n1007, n444, n316, n261, n204);
xnor g653 (n1045, n480, n300, n605, n630);
nand g654 (n1146, n575, n457, n251, n553);
or   g655 (n727, n278, n665, n190, n549);
and  g656 (n1052, n495, n256, n552, n493);
and  g657 (n1006, n201, n410, n350, n525);
xnor g658 (n1009, n191, n381, n580, n211);
xor  g659 (n1119, n176, n477, n333, n256);
xor  g660 (n717, n417, n358, n479, n596);
xnor g661 (n1161, n265, n416, n590, n496);
nand g662 (n903, n643, n659, n258, n450);
xnor g663 (n1054, n412, n494, n491, n177);
xor  g664 (n1053, n573, n494, n589, n331);
nor  g665 (n1152, n338, n471, n506);
nand g666 (n867, n269, n472, n516, n356);
and  g667 (n1100, n200, n447, n585, n455);
xor  g668 (n1117, n260, n554, n656, n346);
xnor g669 (n988, n432, n416, n407, n300);
and  g670 (n896, n468, n469, n470, n345);
nand g671 (n949, n567, n472, n238, n549);
and  g672 (n714, n450, n436, n578, n236);
xor  g673 (n1167, n378, n611, n250, n565);
xnor g674 (n1068, n545, n164, n450, n182);
xnor g675 (n977, n364, n605, n543, n621);
xnor g676 (n1180, n575, n186, n667, n480);
nand g677 (n786, n397, n172, n349, n304);
and  g678 (n1005, n454, n270, n443, n595);
xnor g679 (n997, n322, n492, n458, n486);
xor  g680 (n1129, n510, n349, n548, n402);
nand g681 (n893, n617, n194, n546, n332);
nand g682 (n722, n361, n213, n339, n262);
nor  g683 (n836, n276, n499, n628, n342);
nor  g684 (n890, n305, n465, n164, n601);
or   g685 (n673, n569, n531, n178, n233);
or   g686 (n992, n642, n462, n165, n339);
nand g687 (n734, n451, n622, n543, n578);
or   g688 (n1091, n470, n593, n216, n498);
or   g689 (n966, n551, n600, n294, n412);
or   g690 (n1151, n555, n294, n420, n379);
xnor g691 (n1039, n359, n484, n537, n659);
or   g692 (n1124, n288, n570, n383, n429);
nor  g693 (n685, n263, n534, n303, n569);
and  g694 (n955, n318, n413, n489, n380);
or   g695 (n989, n191, n648, n595, n219);
or   g696 (n923, n490, n409, n451, n477);
or   g697 (n1042, n432, n389, n204, n227);
nand g698 (n858, n265, n603, n565, n248);
xor  g699 (n969, n418, n622, n660, n296);
xnor g700 (n716, n257, n234, n432, n291);
or   g701 (n880, n258, n162, n271, n603);
nand g702 (n701, n409, n566, n551, n405);
and  g703 (n1174, n416, n325, n601, n339);
xnor g704 (n985, n360, n444, n533, n542);
or   g705 (n784, n321, n240, n179, n613);
or   g706 (n747, n611, n415, n502, n404);
xnor g707 (n1093, n364, n267, n457, n613);
and  g708 (n1128, n618, n194, n469, n432);
nand g709 (n1157, n525, n579, n334, n578);
nand g710 (n774, n524, n522, n558, n466);
nand g711 (n807, n207, n476, n399, n170);
or   g712 (n901, n427, n661, n509, n277);
and  g713 (n1130, n447, n667, n414, n616);
nand g714 (n864, n319, n590, n548, n564);
nor  g715 (n1025, n601, n299, n391, n576);
nor  g716 (n1024, n165, n184, n248, n252);
xor  g717 (n908, n586, n533, n582, n296);
xnor g718 (n682, n611, n622, n405, n557);
and  g719 (n1164, n257, n402, n417, n306);
xor  g720 (n756, n255, n588, n281, n309);
xor  g721 (n741, n480, n367, n473, n422);
nor  g722 (n1016, n510, n415, n624, n301);
xnor g723 (n761, n298, n441, n494, n547);
and  g724 (n1044, n219, n328, n214, n199);
nor  g725 (n866, n414, n172, n250, n427);
nor  g726 (n1060, n396, n373, n323, n421);
nand g727 (n793, n443, n236, n251, n313);
nand g728 (n764, n506, n337, n517, n361);
xnor g729 (n721, n530, n641, n564, n492);
and  g730 (n849, n232, n599, n475, n662);
nand g731 (n1020, n651, n285, n348, n618);
xnor g732 (n1163, n585, n338, n527, n330);
or   g733 (n938, n281, n612, n249, n561);
xor  g734 (n1059, n375, n188, n410, n222);
or   g735 (n863, n195, n567, n248, n302);
and  g736 (n677, n247, n394, n218);
nor  g737 (n1023, n368, n538, n589, n280);
nor  g738 (n841, n457, n557, n363, n621);
or   g739 (n944, n560, n576, n475, n306);
nand g740 (n800, n375, n194, n265, n550);
or   g741 (n848, n529, n544, n186, n522);
xnor g742 (n990, n505, n352, n515, n260);
xnor g743 (n1101, n467, n663, n419, n536);
nor  g744 (n1033, n297, n654, n493, n507);
and  g745 (n986, n590, n539, n201, n350);
xor  g746 (n1051, n259, n164, n360, n518);
xor  g747 (n776, n165, n601, n442, n592);
xnor g748 (n1031, n633, n516, n289, n237);
nand g749 (n810, n354, n455, n587, n536);
nand g750 (n902, n508, n400, n434, n203);
nand g751 (n891, n396, n516, n649, n332);
xor  g752 (n998, n220, n347, n307, n462);
and  g753 (n1126, n206, n311, n545, n524);
xnor g754 (n770, n523, n197, n340, n525);
nor  g755 (n924, n631, n500, n267, n600);
xnor g756 (n823, n364, n312, n493, n512);
and  g757 (n1021, n227, n225, n484, n430);
xor  g758 (n1115, n513, n304, n253, n174);
nand g759 (n811, n284, n650, n563, n225);
and  g760 (n967, n352, n666, n372, n242);
nand g761 (n932, n366, n596, n363, n665);
xnor g762 (n1181, n492, n512, n639, n599);
xnor g763 (n1047, n283, n301, n282, n452);
nor  g764 (n771, n539, n544, n319, n615);
nand g765 (n905, n253, n301, n230, n597);
nor  g766 (n1062, n495, n429, n482, n490);
nor  g767 (n785, n205, n418, n619, n416);
and  g768 (n1084, n414, n342, n434, n395);
or   g769 (n1102, n376, n518, n401, n185);
nor  g770 (n1170, n344, n202, n477, n600);
xnor g771 (n1154, n626, n439, n501, n381);
and  g772 (n851, n614, n254, n603, n461);
and  g773 (n936, n341, n309, n239, n255);
nand g774 (n728, n334, n501, n295, n239);
or   g775 (n820, n647, n378, n622, n431);
nor  g776 (n888, n490, n665, n644, n352);
xnor g777 (n1141, n446, n221, n502, n385);
nor  g778 (n762, n663, n250, n612, n438);
xor  g779 (n853, n668, n658, n610, n452);
xnor g780 (n931, n209, n223, n308, n302);
and  g781 (n1136, n167, n161, n386, n336);
xnor g782 (n1148, n237, n319, n435, n229);
nor  g783 (n675, n226, n321, n391, n401);
nand g784 (n974, n310, n388, n430, n369);
xor  g785 (n999, n557, n273, n554, n167);
xnor g786 (n837, n462, n562, n344, n315);
and  g787 (n1008, n609, n418, n666, n560);
xnor g788 (n754, n184, n166, n564, n636);
or   g789 (n797, n185, n288, n394, n365);
and  g790 (n1109, n583, n487, n217, n351);
xor  g791 (n831, n242, n184, n487, n572);
nor  g792 (n945, n215, n539, n579, n489);
xnor g793 (n686, n406, n441, n438, n629);
xnor g794 (n1160, n358, n666, n424, n485);
and  g795 (n930, n384, n392, n527, n425);
xor  g796 (n731, n367, n445, n392, n597);
nand g797 (n711, n263, n315, n168, n526);
and  g798 (n947, n591, n411, n533, n637);
xor  g799 (n1153, n483, n567, n508, n655);
nor  g800 (n828, n608, n284, n439, n293);
nor  g801 (n812, n235, n396, n278, n173);
or   g802 (n916, n612, n399, n486, n198);
xor  g803 (n912, n317, n541, n292, n403);
nand g804 (n732, n404, n163, n169, n632);
and  g805 (n697, n183, n389, n552, n175);
xnor g806 (n1057, n542, n323, n226, n395);
xnor g807 (n755, n176, n390, n650, n550);
and  g808 (n879, n627, n633, n244, n236);
xor  g809 (n681, n210, n230, n411, n508);
xnor g810 (n1081, n610, n492, n635, n583);
nand g811 (n1094, n429, n239, n631, n257);
nand g812 (n744, n629, n495, n383, n447);
or   g813 (n758, n467, n524, n497, n625);
and  g814 (n1166, n205, n628, n284, n191);
and  g815 (n918, n592, n565, n348, n630);
nor  g816 (n1026, n567, n620, n479, n414);
and  g817 (n688, n606, n227, n272, n266);
nor  g818 (n739, n581, n192, n636, n276);
xor  g819 (n1122, n320, n308, n507, n582);
nor  g820 (n946, n606, n640, n404, n207);
or   g821 (n907, n199, n236, n647, n626);
xor  g822 (n987, n179, n163, n658, n259);
xnor g823 (n809, n575, n317, n201, n410);
and  g824 (n1076, n553, n220, n515, n393);
nand g825 (n782, n633, n451, n660, n552);
nand g826 (n787, n327, n548, n608, n360);
nor  g827 (n935, n193, n402, n374, n425);
nor  g828 (n680, n508, n473, n448, n260);
nand g829 (n1074, n610, n268, n189, n206);
xnor g830 (n933, n219, n585, n565, n235);
xor  g831 (n753, n607, n196, n362, n316);
and  g832 (n982, n592, n330, n530, n474);
xnor g833 (n887, n545, n405, n383, n290);
nor  g834 (n886, n222, n440, n176, n568);
xnor g835 (n1137, n314, n517, n359, n448);
nor  g836 (n862, n185, n450, n472, n510);
or   g837 (n704, n663, n536, n545, n585);
or   g838 (n833, n302, n548, n386, n598);
and  g839 (n759, n289, n497, n653, n199);
nor  g840 (n1120, n382, n511, n657, n576);
and  g841 (n876, n291, n302, n408, n631);
or   g842 (n1065, n437, n371, n348, n239);
nor  g843 (n801, n408, n424, n409, n453);
xor  g844 (n1095, n235, n652, n231, n194);
nor  g845 (n840, n412, n549, n460, n428);
or   g846 (n1070, n327, n556, n495, n469);
nor  g847 (n825, n528, n280, n377);
nor  g848 (n1041, n247, n262, n449, n466);
or   g849 (n708, n623, n400, n214, n547);
xnor g850 (n1088, n531, n568, n294, n275);
nand g851 (n1149, n354, n644, n546, n571);
nand g852 (n1171, n365, n339, n332, n367);
or   g853 (n942, n471, n445, n657, n356);
xnor g854 (n789, n198, n357, n477, n334);
nor  g855 (n1035, n398, n323, n209, n343);
nand g856 (n1037, n543, n361, n329, n358);
xor  g857 (n964, n491, n511, n270, n282);
nand g858 (n1001, n277, n593, n616, n522);
or   g859 (n1144, n193, n254, n192, n168);
or   g860 (n1133, n226, n628, n447, n563);
xor  g861 (n808, n276, n609, n208, n273);
and  g862 (n751, n366, n443, n417, n441);
nor  g863 (n804, n308, n384, n518, n172);
and  g864 (n1032, n384, n439, n520, n423);
and  g865 (n795, n645, n335, n225, n329);
nor  g866 (n1106, n459, n266, n324, n444);
xor  g867 (n906, n270, n361, n470, n396);
nand g868 (n861, n431, n668, n163, n594);
nand g869 (n1107, n400, n461, n258, n512);
or   g870 (n683, n594, n169, n605, n655);
nor  g871 (n1017, n561, n223, n190, n382);
nand g872 (n1118, n180, n643, n557, n490);
nand g873 (n730, n344, n648, n230, n405);
and  g874 (n1058, n433, n163, n429, n581);
and  g875 (n790, n609, n232, n388, n182);
or   g876 (n940, n617, n547, n291, n187);
or   g877 (n709, n295, n470, n166, n233);
and  g878 (n1159, n449, n322, n463, n293);
xor  g879 (n766, n606, n242, n181, n204);
or   g880 (n698, n245, n393, n654, n517);
xor  g881 (n894, n549, n566, n562, n169);
or   g882 (n746, n534, n387, n544, n561);
nor  g883 (n1108, n656, n499, n572, n556);
nand g884 (n951, n540, n268, n483, n203);
or   g885 (n715, n207, n442, n288, n569);
nand g886 (n1175, n357, n202, n271, n219);
xnor g887 (n1105, n503, n421, n533, n188);
xor  g888 (n871, n563, n248, n558, n530);
xor  g889 (n1064, n471, n161, n553, n453);
xor  g890 (n687, n638, n178, n403, n663);
nand g891 (n760, n555, n213, n371, n190);
xor  g892 (n1090, n203, n384, n353, n602);
and  g893 (n691, n591, n398, n468, n623);
xnor g894 (n956, n496, n198, n491, n526);
xor  g895 (n1077, n283, n259, n425, n404);
xnor g896 (n719, n211, n505, n192, n473);
xnor g897 (n1158, n399, n527, n664, n340);
nand g898 (n928, n222, n397, n638, n461);
nand g899 (n978, n209, n428, n652, n561);
and  g900 (n872, n420, n528, n535, n174);
nand g901 (n1173, n476, n427, n306, n347);
xor  g902 (n696, n595, n376, n598);
xnor g903 (n1092, n515, n300, n604, n628);
xor  g904 (n1027, n377, n366, n238, n167);
nand g905 (n1103, n597, n309, n624, n591);
nor  g906 (n814, n644, n521, n642, n220);
nand g907 (n1139, n619, n355, n443, n408);
and  g908 (n1003, n206, n235, n161, n282);
and  g909 (n856, n360, n242, n318, n173);
or   g910 (n950, n238, n210, n428, n423);
xor  g911 (n976, n456, n275, n169, n279);
nand g912 (n748, n359, n181, n253, n667);
or   g913 (n743, n193, n371, n649, n572);
xor  g914 (n1056, n181, n329, n458, n326);
nand g915 (n962, n500, n261, n476, n607);
and  g916 (n1022, n320, n200, n392, n285);
and  g917 (n684, n266, n298, n237, n243);
nor  g918 (n961, n181, n253, n372, n602);
nand g919 (n726, n377, n409, n311, n433);
or   g920 (n937, n417, n535, n532, n335);
or   g921 (n1177, n166, n261, n205, n448);
or   g922 (n818, n180, n357, n192, n595);
xor  g923 (n957, n162, n458, n649, n574);
xor  g924 (n773, n569, n639, n333, n337);
xnor g925 (n984, n614, n607, n489, n657);
nand g926 (n1082, n499, n512, n295, n623);
xnor g927 (n830, n208, n554, n243, n170);
nand g928 (n958, n442, n287, n592, n204);
xnor g929 (n737, n619, n252, n357, n173);
xnor g930 (n819, n621, n397, n210, n223);
nand g931 (n815, n271, n449, n273, n573);
xor  g932 (n860, n195, n582, n380, n645);
xnor g933 (n798, n637, n640, n407, n331);
or   g934 (n972, n351, n221, n454, n627);
xor  g935 (n1172, n231, n333, n262, n464);
xor  g936 (n725, n529, n187, n293, n486);
xnor g937 (n794, n272, n251, n586, n424);
nor  g938 (n980, n303, n646, n260, n459);
nor  g939 (n874, n191, n625, n642, n313);
and  g940 (n775, n426, n190, n324, n172);
or   g941 (n909, n342, n316, n286, n321);
or   g942 (n724, n370, n597, n550, n462);
nor  g943 (n884, n513, n581, n311, n614);
and  g944 (n835, n217, n476, n391, n406);
or   g945 (n788, n460, n424, n177, n620);
and  g946 (n1055, n343, n336, n408, n307);
or   g947 (n713, n370, n555, n288, n579);
or   g948 (n921, n596, n504, n326, n421);
nor  g949 (n1048, n531, n463, n504, n459);
xor  g950 (n1086, n646, n286, n528);
xnor g951 (n842, n632, n299, n382, n279);
or   g952 (n847, n651, n334, n243, n345);
xor  g953 (n1096, n485, n267, n385, n625);
nand g954 (n824, n486, n202, n281, n661);
nor  g955 (n707, n244, n209, n497, n240);
nand g956 (n839, n513, n376, n662, n529);
and  g957 (n1176, n464, n437, n653, n489);
xnor g958 (n1049, n487, n660, n329, n237);
nand g959 (n1015, n306, n251, n374, n266);
and  g960 (n803, n208, n643, n426, n487);
xnor g961 (n735, n522, n425, n615, n244);
xor  g962 (n1000, n307, n273, n304, n285);
xnor g963 (n1142, n234, n527, n540, n639);
xor  g964 (n703, n615, n652, n578, n488);
and  g965 (n736, n650, n478, n584, n534);
nor  g966 (n875, n665, n385, n542, n228);
and  g967 (n1063, n316, n482, n587, n274);
and  g968 (n720, n264, n661, n267, n368);
and  g969 (n1002, n315, n358, n215, n394);
nand g970 (n1078, n174, n580, n211, n411);
nand g971 (n859, n230, n180, n456, n573);
nand g972 (n1127, n325, n349, n662, n542);
xor  g973 (n821, n178, n372, n531, n461);
nand g974 (n692, n418, n278, n293, n201);
or   g975 (n702, n634, n494, n496, n515);
xor  g976 (n843, n175, n634, n465, n324);
or   g977 (n712, n175, n229, n457, n582);
nand g978 (n846, n481, n342, n296, n403);
xnor g979 (n805, n331, n187, n246, n223);
and  g980 (n749, n398, n350, n530, n373);
or   g981 (n993, n453, n284, n249, n337);
nor  g982 (n898, n299, n474, n560, n309);
xor  g983 (n885, n247, n653, n228, n426);
xnor g984 (n834, n627, n587, n667, n543);
xnor g985 (n892, n415, n187, n216, n474);
xor  g986 (n1029, n303, n333, n643, n604);
xnor g987 (n806, n534, n287, n256, n584);
and  g988 (n852, n287, n332, n600, n617);
nand g989 (n791, n195, n488, n648, n373);
nor  g990 (n981, n241, n660, n289, n602);
nand g991 (n926, n619, n328, n510, n589);
nor  g992 (n878, n535, n231, n584, n277);
xnor g993 (n915, n381, n528, n319, n212);
xor  g994 (n817, n336, n215, n170, n594);
nand g995 (n939, n474, n636, n348, n353);
or   g996 (n1013, n218, n340, n499, n507);
xor  g997 (n802, n570, n322, n176, n390);
xor  g998 (n904, n338, n391, n179, n378);
xnor g999 (n1134, n649, n435, n213, n368);
nand g1000 (n816, n519, n394, n354, n382);
nand g1001 (n780, n483, n580, n214, n186);
xnor g1002 (n971, n166, n496, n420, n226);
and  g1003 (n1110, n593, n593, n653, n603);
nor  g1004 (n745, n503, n613, n471, n311);
nand g1005 (n870, n326, n343, n481, n498);
nand g1006 (n963, n604, n442, n466, n558);
nor  g1007 (n1030, n255, n485, n505, n519);
and  g1008 (n917, n162, n634, n389, n553);
xor  g1009 (n973, n546, n314, n577, n410);
xnor g1010 (n838, n301, n246, n541, n379);
or   g1011 (n996, n327, n255, n504, n547);
nor  g1012 (n1099, n368, n614, n386, n599);
or   g1013 (n1004, n599, n314, n188, n484);
xnor g1014 (n952, n413, n199, n568, n274);
and  g1015 (n1050, n423, n238, n363, n523);
and  g1016 (n1073, n184, n264, n330, n589);
nand g1017 (n910, n271, n558, n657, n281);
or   g1018 (n994, n355, n491, n503, n328);
and  g1019 (n822, n283, n196, n587, n616);
and  g1020 (n1143, n341, n436, n440, n581);
nand g1021 (n941, n240, n655, n541, n245);
and  g1022 (n883, n317, n356, n205, n203);
xnor g1023 (n750, n566, n246, n630, n262);
nand g1024 (n1104, n200, n340, n272, n217);
and  g1025 (n1132, n501, n310, n407, n481);
nand g1026 (n900, n338, n537, n430, n388);
xnor g1027 (n718, n535, n326, n189, n164);
xor  g1028 (n1071, n298, n521, n658, n261);
xor  g1029 (n1087, n609, n577, n228, n529);
and  g1030 (n1169, n661, n509, n473, n591);
xor  g1031 (n1069, n598, n454, n272, n606);
and  g1032 (n792, n483, n167, n380, n289);
xnor g1033 (n873, n320, n480, n636, n656);
xnor g1034 (n914, n440, n298, n588, n162);
xnor g1035 (n1028, n654, n475, n347, n320);
nor  g1036 (n1179, n437, n419, n168, n218);
and  g1037 (n850, n285, n514, n625, n224);
nand g1038 (n970, n612, n290, n263, n627);
nand g1039 (n920, n264, n214, n479, n336);
nand g1040 (n913, n637, n171, n227, n177);
or   g1041 (n991, n540, n497, n556, n245);
xnor g1042 (n975, n400, n631, n182, n350);
and  g1043 (n763, n264, n434, n406, n455);
or   g1044 (n1114, n638, n514, n182, n411);
xnor g1045 (n1168, n161, n618, n526, n224);
and  g1046 (n844, n392, n383, n559, n390);
xor  g1047 (n740, n229, n516, n183, n556);
xor  g1048 (n700, n580, n640, n559, n506);
xnor g1049 (n676, n365, n468, n165, n560);
and  g1050 (n1038, n500, n637, n464, n629);
nand g1051 (n1147, n193, n546, n669, n579);
and  g1052 (n1116, n519, n588, n247, n433);
nand g1053 (n689, n268, n168, n318, n666);
xnor g1054 (n882, n536, n280, n183, n312);
xnor g1055 (n779, n313, n467, n197);
nor  g1056 (n1112, n296, n224, n406, n177);
nor  g1057 (n1080, n359, n299, n586, n454);
xnor g1058 (n752, n493, n526, n574, n275);
or   g1059 (n729, n559, n292, n438, n335);
nor  g1060 (n1018, n312, n633, n387, n290);
nor  g1061 (n948, n353, n616, n171, n322);
and  g1062 (n1034, n566, n195, n475, n310);
xnor g1063 (n1123, n439, n647, n669, n456);
xor  g1064 (n965, n385, n305, n469, n403);
xor  g1065 (n783, n504, n171, n590, n520);
xor  g1066 (n678, n521, n341, n291, n270);
nand g1067 (n1083, n446, n646, n583, n365);
nor  g1068 (n765, n507, n328, n244, n422);
nor  g1069 (n877, n213, n353, n314, n647);
nand g1070 (n1145, n305, n521, n537, n460);
nand g1071 (n922, n393, n335, n626, n635);
nand g1072 (n927, n297, n346, n481, n369);
and  g1073 (n1165, n646, n197, n279, n555);
or   g1074 (n1085, n668, n252, n202, n511);
xnor g1075 (n699, n626, n233, n574, n472);
nor  g1076 (n1098, n541, n290, n584, n377);
xnor g1077 (n1014, n441, n283, n485, n257);
nor  g1078 (n1135, n452, n303, n217, n500);
nand g1079 (n934, n294, n234, n189, n641);
and  g1080 (n1075, n211, n520, n517, n449);
or   g1081 (n723, n279, n378, n246, n540);
nand g1082 (n827, n373, n669, n398, n376);
or   g1083 (n857, n664, n618, n249, n479);
xor  g1084 (n1036, n438, n434, n623, n451);
or   g1085 (n929, n605, n523, n174, n312);
or   g1086 (n674, n341, n346, n488, n206);
xor  g1087 (n968, n455, n362, n551, n617);
xor  g1088 (n1155, n330, n656, n509, n562);
xnor g1089 (n694, n511, n370, n287, n185);
and  g1090 (n925, n588, n221, n379, n220);
nor  g1091 (n769, n232, n188, n509, n362);
xnor g1092 (n690, n412, n630, n374, n372);
xnor g1093 (n897, n624, n401, n610, n532);
xor  g1094 (n983, n254, n644, n523, n482);
or   g1095 (n799, n399, n380, n387, n583);
and  g1096 (n1178, n402, n641, n634, n292);
nand g1097 (n733, n364, n648, n440, n321);
or   g1098 (n943, n551, n658, n514, n563);
xor  g1099 (n767, n478, n216, n245, n446);
xor  g1100 (n1113, n241, n415, n664, n620);
and  g1101 (n1131, n577, n395, n652, n207);
nand g1102 (n705, n502, n651, n254, n363);
and  g1103 (n1067, n550, n232, n210, n325);
nor  g1104 (n1150, n352, n460, n249, n645);
and  g1105 (n768, n577, n532, n179, n349);
nand g1106 (n1046, n393, n346, n297, n437);
nand g1107 (n693, n208, n224, n505, n315);
nor  g1108 (n1162, n197, n343, n221, n498);
and  g1109 (n855, n324, n196, n635, n427);
or   g1110 (n960, n379, n362, n292, n642);
nor  g1111 (n889, n389, n659, n265, n222);
xnor g1112 (n1043, n453, n229, n502, n390);
and  g1113 (n1019, n635, n274, n574, n459);
xnor g1114 (n796, n369, n615, n456, n256);
and  g1115 (n953, n241, n370, n212, n519);
or   g1116 (n832, n215, n304, n607, n422);
xor  g1117 (n738, n624, n269, n228, n268);
and  g1118 (n829, n532, n337, n354, n375);
nand g1119 (n865, n445, n659, n559, n419);
or   g1120 (n1138, n436, n638, n513, n216);
nor  g1121 (n1072, n468, n664, n407, n520);
nor  g1122 (n706, n596, n317, n367, n445);
xor  g1123 (n899, n240, n300, n323, n258);
xnor g1124 (n959, n570, n452, n243, n488);
or   g1125 (n869, n478, n263, n277, n537);
xor  g1126 (n895, n278, n501, n463, n175);
nor  g1127 (n1012, n344, n388, n259, n570);
or   g1128 (n1079, n538, n276, n269, n651);
xnor g1129 (n772, n514, n431, n386, n241);
nor  g1130 (n710, n465, n594, n310, n482);
xor  g1131 (n1011, n466, n369, n307, n250);
nor  g1132 (n919, n178, n413, n640, n173);
nor  g1133 (n1111, n433, n374, n413, n571);
xor  g1134 (n1156, n305, n538, n269, n286);
nor  g1135 (n854, n586, n345, n608);
xor  g1136 (n1040, n525, n423, n650, n170);
nand g1137 (n1061, n503, n421, n464, n573);
xor  g1138 (n781, n564, n446, n552, n539);
xor  g1139 (n813, n186, n654, n431, n613);
xnor g1140 (n1010, n282, n572, n419, n371);
nand g1141 (n954, n274, n568, n430, n401);
xor  g1142 (n845, n295, n351, n375, n327);
nand g1143 (n1089, n632, n571, n308, n212);
xor  g1144 (n1097, n420, n189, n611, n435);
nor  g1145 (n757, n225, n632, n313, n458);
nand g1146 (n1140, n366, n641, n538, n196);
nor  g1147 (n1125, n669, n562, n180, n200);
nor  g1148 (n881, n448, n318, n463, n234);
not  g1149 (n1184, n698);
not  g1150 (n1191, n700);
not  g1151 (n1188, n692);
buf  g1152 (n1193, n693);
buf  g1153 (n1185, n677);
buf  g1154 (n1195, n689);
buf  g1155 (n1187, n679);
buf  g1156 (n1199, n690);
not  g1157 (n1186, n678);
not  g1158 (n1194, n675);
not  g1159 (n1198, n684);
buf  g1160 (n1202, n694);
not  g1161 (n1192, n688);
buf  g1162 (n1190, n695);
not  g1163 (n1182, n699);
not  g1164 (n1189, n682);
not  g1165 (n1197, n687);
not  g1166 (n1200, n683);
nand g1167 (n1183, n680, n691);
and  g1168 (n1196, n674, n681, n685, n697);
nand g1169 (n1201, n696, n686, n673, n676);
buf  g1170 (n1203, n1182);
buf  g1171 (n1204, n1182);
not  g1172 (n1212, n1203);
buf  g1173 (n1206, n1204);
buf  g1174 (n1210, n1203);
not  g1175 (n1205, n1204);
buf  g1176 (n1209, n1204);
not  g1177 (n1211, n701);
not  g1178 (n1207, n1203);
or   g1179 (n1208, n1204, n1203, n702);
buf  g1180 (n1244, n1206);
buf  g1181 (n1215, n1208);
buf  g1182 (n1241, n1206);
buf  g1183 (n1227, n1207);
buf  g1184 (n1225, n1208);
not  g1185 (n1218, n1207);
buf  g1186 (n1242, n1211);
not  g1187 (n1216, n1209);
buf  g1188 (n1230, n1208);
buf  g1189 (n1234, n1212);
buf  g1190 (n1213, n1205);
not  g1191 (n1222, n1209);
not  g1192 (n1232, n1212);
not  g1193 (n1214, n1205);
buf  g1194 (n1224, n1210);
buf  g1195 (n1243, n1205);
buf  g1196 (n1235, n1211);
not  g1197 (n1217, n1212);
buf  g1198 (n1220, n1207);
buf  g1199 (n1238, n1210);
not  g1200 (n1240, n1209);
buf  g1201 (n1226, n1207);
not  g1202 (n1233, n1209);
buf  g1203 (n1219, n1210);
buf  g1204 (n1237, n1206);
not  g1205 (n1229, n1211);
not  g1206 (n1228, n1210);
not  g1207 (n1239, n1206);
not  g1208 (n1236, n1211);
not  g1209 (n1231, n1208);
not  g1210 (n1221, n1205);
buf  g1211 (n1223, n1212);
not  g1212 (n1245, n1216);
buf  g1213 (n1253, n1216);
not  g1214 (n1252, n1216);
not  g1215 (n1248, n1214);
buf  g1216 (n1251, n1215);
buf  g1217 (n1254, n1214);
not  g1218 (n1247, n1213);
buf  g1219 (n1246, n1216);
buf  g1220 (n1249, n1213);
not  g1221 (n1250, n1215);
not  g1222 (n1262, n1249);
buf  g1223 (n1264, n1249);
buf  g1224 (n1266, n1247);
not  g1225 (n1268, n1250);
not  g1226 (n1277, n1250);
not  g1227 (n1260, n1246);
not  g1228 (n1261, n1248);
buf  g1229 (n1263, n1246);
not  g1230 (n1273, n1249);
buf  g1231 (n1278, n1247);
not  g1232 (n1275, n1250);
not  g1233 (n1276, n1248);
not  g1234 (n1256, n1248);
buf  g1235 (n1269, n1245);
not  g1236 (n1272, n1246);
not  g1237 (n1257, n1248);
buf  g1238 (n1270, n1245);
not  g1239 (n1255, n1247);
buf  g1240 (n1271, n1245);
buf  g1241 (n1259, n1249);
buf  g1242 (n1258, n1246);
buf  g1243 (n1274, n1245);
not  g1244 (n1267, n1247);
not  g1245 (n1265, n1250);
not  g1246 (n1290, n1255);
not  g1247 (n1293, n1255);
buf  g1248 (n1283, n1255);
buf  g1249 (n1296, n1261);
not  g1250 (n1302, n1261);
not  g1251 (n1295, n1258);
buf  g1252 (n1304, n1258);
not  g1253 (n1306, n1257);
not  g1254 (n1279, n1262);
buf  g1255 (n1280, n1256);
not  g1256 (n1282, n1257);
buf  g1257 (n1297, n1261);
not  g1258 (n1281, n1262);
not  g1259 (n1289, n1255);
buf  g1260 (n1294, n1256);
buf  g1261 (n1284, n1260);
not  g1262 (n1303, n1259);
not  g1263 (n1307, n1256);
buf  g1264 (n1286, n1259);
buf  g1265 (n1305, n1256);
not  g1266 (n1287, n1260);
buf  g1267 (n1298, n1260);
buf  g1268 (n1299, n1258);
not  g1269 (n1301, n1260);
buf  g1270 (n1300, n1259);
buf  g1271 (n1308, n1258);
not  g1272 (n1291, n1257);
not  g1273 (n1292, n1259);
buf  g1274 (n1288, n1257);
not  g1275 (n1285, n1261);
xor  g1276 (n1309, n703, n704, n705, n1279);
buf  g1277 (n1310, n1309);
not  g1278 (n1311, n1309);
or   g1279 (n1313, n1311, n706, n712, n1251);
xnor g1280 (n1312, n708, n1251);
xnor g1281 (n1315, n711, n714, n1253, n1310);
or   g1282 (n1314, n1252, n1252, n1311, n1310);
and  g1283 (n1317, n707, n710, n1252, n1253);
and  g1284 (n1318, n713, n1253, n715, n709);
xnor g1285 (n1316, n1311, n1311, n1252, n1310);
not  g1286 (n1327, n1312);
buf  g1287 (n1328, n1313);
buf  g1288 (n1325, n1313);
not  g1289 (n1324, n1312);
not  g1290 (n1322, n1314);
buf  g1291 (n1320, n1315);
not  g1292 (n1319, n1315);
buf  g1293 (n1323, n1315);
buf  g1294 (n1321, n1315);
buf  g1295 (n1326, n1314);
nor  g1296 (n1360, n734, n766, n1324);
xnor g1297 (n1357, n805, n756, n822, n754);
nor  g1298 (n1365, n1326, n1325, n828, n719);
xnor g1299 (n1364, n1321, n731, n777, n797);
nand g1300 (n1330, n832, n1322, n816, n1326);
and  g1301 (n1359, n736, n831, n818, n774);
and  g1302 (n1340, n727, n765, n1321, n1328);
or   g1303 (n1346, n770, n746, n758, n739);
nor  g1304 (n1354, n1319, n763, n771, n761);
xor  g1305 (n1347, n809, n718, n823, n716);
or   g1306 (n1336, n721, n751, n795, n800);
and  g1307 (n1352, n740, n729, n1328, n819);
nor  g1308 (n1334, n742, n1323, n1324, n1320);
or   g1309 (n1358, n829, n775, n807, n748);
xnor g1310 (n1333, n738, n735, n798, n1320);
xnor g1311 (n1338, n1325, n757, n722, n782);
and  g1312 (n1335, n813, n737, n835, n827);
nand g1313 (n1368, n790, n785, n755, n783);
or   g1314 (n1345, n744, n724, n747, n1327);
xnor g1315 (n1341, n825, n787, n812, n804);
xnor g1316 (n1353, n802, n814, n834, n1325);
and  g1317 (n1356, n799, n817, n792, n801);
and  g1318 (n1351, n796, n810, n1321, n1323);
or   g1319 (n1332, n793, n772, n1327, n788);
and  g1320 (n1329, n1322, n778, n1319, n1323);
xnor g1321 (n1344, n820, n1320, n773, n745);
nor  g1322 (n1355, n764, n759, n743, n1319);
or   g1323 (n1366, n768, n794, n833, n760);
and  g1324 (n1363, n1321, n826, n1320, n1322);
nor  g1325 (n1348, n769, n1327, n723, n803);
xnor g1326 (n1331, n815, n791, n780, n776);
nand g1327 (n1337, n1325, n730, n786, n779);
xnor g1328 (n1350, n789, n1327, n784, n1319);
xor  g1329 (n1343, n1326, n749, n808, n753);
xor  g1330 (n1342, n1324, n1322, n1326, n750);
nor  g1331 (n1362, n1328, n811, n732, n830);
nor  g1332 (n1361, n741, n733, n821, n781);
xor  g1333 (n1349, n767, n806, n762, n717);
and  g1334 (n1367, n752, n1328, n725, n728);
xor  g1335 (n1339, n720, n726, n1323, n824);
not  g1336 (n1370, n1330);
not  g1337 (n1369, n1329);
or   g1338 (n1371, n837, n836);
and  g1339 (n1372, n849, n1369, n842, n845);
xor  g1340 (n1373, n848, n847, n838, n843);
and  g1341 (n1375, n1370, n844, n846, n841);
xnor g1342 (n1374, n839, n1371, n840);
nor  g1343 (n1377, n670, n672, n860, n854);
or   g1344 (n1385, n1375, n1373, n852);
xor  g1345 (n1381, n670, n1372, n850, n1279);
xnor g1346 (n1384, n670, n1316, n857, n1375);
xor  g1347 (n1379, n864, n1374, n670);
xnor g1348 (n1382, n671, n855, n1375, n1373);
and  g1349 (n1386, n862, n1317, n1316, n1318);
or   g1350 (n1376, n853, n671, n863, n1374);
nand g1351 (n1383, n1372, n1317, n858);
and  g1352 (n1380, n1375, n672, n861, n1317);
and  g1353 (n1378, n671, n859, n1374, n1316);
xnor g1354 (n1387, n1316, n851, n671, n856);
not  g1355 (n1388, n1377);
buf  g1356 (n1390, n1378);
not  g1357 (n1392, n1380);
not  g1358 (n1391, n1376);
buf  g1359 (n1393, n1379);
not  g1360 (n1389, n1381);
not  g1361 (n1400, n1392);
not  g1362 (n1413, n872);
buf  g1363 (n1407, n1389);
not  g1364 (n1409, n874);
not  g1365 (n1401, n1390);
not  g1366 (n1404, n1391);
not  g1367 (n1396, n1392);
buf  g1368 (n1405, n875);
buf  g1369 (n1403, n871);
buf  g1370 (n1416, n865);
buf  g1371 (n1411, n1390);
xor  g1372 (n1395, n901, n1391, n900);
nand g1373 (n1417, n866, n897, n1391, n882);
and  g1374 (n1406, n1389, n881, n885, n889);
and  g1375 (n1415, n888, n1388, n891, n1391);
or   g1376 (n1399, n869, n1389, n1392, n1393);
xor  g1377 (n1402, n902, n1390, n892, n880);
xor  g1378 (n1412, n884, n873, n1393, n877);
nor  g1379 (n1397, n870, n1388, n1390, n883);
and  g1380 (n1398, n896, n1393, n887, n898);
or   g1381 (n1410, n890, n878, n879, n867);
xor  g1382 (n1408, n868, n886, n899, n876);
nor  g1383 (n1394, n1393, n893, n1389, n895);
nor  g1384 (n1414, n894, n1392, n1388);
buf  g1385 (n1438, n1402);
not  g1386 (n1506, n1400);
buf  g1387 (n1468, n1404);
buf  g1388 (n1502, n1201);
not  g1389 (n1510, n1190);
not  g1390 (n1507, n1197);
not  g1391 (n1501, n1414);
buf  g1392 (n1462, n1275);
buf  g1393 (n1491, n1269);
buf  g1394 (n1423, n1193);
buf  g1395 (n1434, n1192);
buf  g1396 (n1421, n1417);
buf  g1397 (n1467, n1331);
not  g1398 (n1483, n1273);
not  g1399 (n1444, n1267);
buf  g1400 (n1459, n1332);
not  g1401 (n1500, n1196);
not  g1402 (n1429, n1263);
not  g1403 (n1439, n1195);
buf  g1404 (n1498, n1412);
buf  g1405 (n1503, n1399);
not  g1406 (n1418, n1274);
not  g1407 (n1494, n1333);
not  g1408 (n1422, n1416);
not  g1409 (n1505, n1411);
buf  g1410 (n1458, n1415);
not  g1411 (n1447, n1386);
buf  g1412 (n1442, n1277);
not  g1413 (n1497, n1271);
buf  g1414 (n1449, n1200);
not  g1415 (n1490, n1187);
not  g1416 (n1476, n1200);
buf  g1417 (n1493, n1409);
not  g1418 (n1424, n1275);
buf  g1419 (n1441, n1412);
buf  g1420 (n1477, n1264);
buf  g1421 (n1445, n1383);
not  g1422 (n1482, n1398);
buf  g1423 (n1457, n1218);
not  g1424 (n1486, n1413);
not  g1425 (n1426, n1272);
not  g1426 (n1463, n1200);
not  g1427 (n1443, n1335);
xnor g1428 (n1487, n1272, n1264);
and  g1429 (n1455, n1403, n1191, n1264);
and  g1430 (n1479, n1269, n1384, n1218);
and  g1431 (n1472, n1267, n1275, n1218, n1406);
and  g1432 (n1450, n1413, n1274, n1415, n1411);
xor  g1433 (n1428, n1269, n1268, n1270, n1334);
nand g1434 (n1469, n1187, n1273, n1399, n1411);
xnor g1435 (n1478, n1395, n1401, n1417, n1382);
xor  g1436 (n1466, n1184, n1334, n1412, n1395);
xor  g1437 (n1465, n1394, n1401, n1272, n1269);
and  g1438 (n1508, n1404, n1394, n1278, n1414);
and  g1439 (n1437, n1404, n1263, n1202, n1417);
or   g1440 (n1475, n1333, n1278, n1411, n1194);
xor  g1441 (n1499, n1266, n1268, n1414, n1399);
xor  g1442 (n1456, n1277, n1405, n1414, n1416);
nand g1443 (n1511, n1273, n1408, n1270, n1195);
nor  g1444 (n1430, n1398, n1405, n1409, n1272);
xor  g1445 (n1473, n1189, n1274, n1402, n1266);
nand g1446 (n1509, n1406, n1271, n1397, n1410);
or   g1447 (n1420, n1413, n1413, n1202, n1416);
or   g1448 (n1464, n1405, n1407, n1186, n1382);
or   g1449 (n1454, n1188, n1267, n1217, n1394);
xor  g1450 (n1432, n1186, n1276, n1397, n1396);
or   g1451 (n1496, n1397, n1201, n1415, n1412);
xnor g1452 (n1433, n1194, n1266, n1398, n1415);
xnor g1453 (n1485, n1385, n1198, n1408, n1407);
nand g1454 (n1440, n1271, n1264, n1410, n1394);
xnor g1455 (n1481, n1263, n1265, n1318, n1266);
nor  g1456 (n1446, n1200, n1403, n1278, n1400);
and  g1457 (n1448, n1386, n1185, n1268, n1183);
xnor g1458 (n1480, n1401, n1196, n1277, n1397);
and  g1459 (n1419, n1400, n1184, n1403, n1395);
xor  g1460 (n1461, n1335, n1263, n1330, n1318);
nor  g1461 (n1427, n1402, n1383, n1267, n1202);
nand g1462 (n1425, n1417, n1185, n1406, n1201);
xor  g1463 (n1488, n1265, n1193, n1396, n1407);
nor  g1464 (n1435, n1268, n1199, n1262);
xor  g1465 (n1453, n1183, n1402, n1410, n1273);
nor  g1466 (n1451, n1270, n1331, n1387, n1318);
nor  g1467 (n1460, n1399, n1197, n1409, n1188);
and  g1468 (n1484, n1262, n1407, n1332, n1192);
nand g1469 (n1431, n1409, n1265, n1189, n903);
nand g1470 (n1504, n1387, n1385, n1278, n1217);
nand g1471 (n1492, n1191, n1408, n1190, n1410);
or   g1472 (n1436, n1217, n1416, n1276, n1274);
xor  g1473 (n1489, n1395, n1270, n1217, n1276);
xor  g1474 (n1495, n1398, n1275, n1271, n1406);
xnor g1475 (n1471, n1396, n1384, n1401, n1405);
or   g1476 (n1452, n1218, n1404, n1408, n1265);
nor  g1477 (n1474, n1396, n1403, n1198, n1276);
nor  g1478 (n1470, n1202, n1400, n1277, n1201);
xnor g1479 (n1528, n907, n917, n1433, n921);
xor  g1480 (n1525, n1430, n1421, n1426, n1447);
xnor g1481 (n1513, n923, n1418, n1423, n1443);
nand g1482 (n1526, n920, n925, n1442, n1428);
nand g1483 (n1523, n1432, n928, n1441, n1443);
xnor g1484 (n1518, n1429, n1431, n1446, n1436);
or   g1485 (n1522, n1427, n1437, n1422);
xnor g1486 (n1527, n904, n1421, n1439, n1419);
and  g1487 (n1514, n909, n1442, n911, n1438);
xnor g1488 (n1520, n1438, n1445, n1447, n931);
or   g1489 (n1521, n1428, n1420, n1430, n1444);
xor  g1490 (n1516, n924, n922, n1419, n1440);
nor  g1491 (n1524, n1422, n1434, n905, n935);
or   g1492 (n1515, n916, n1434, n1440, n919);
xor  g1493 (n1533, n1446, n1431, n1436, n1445);
and  g1494 (n1531, n1418, n906, n1420, n1435);
xnor g1495 (n1534, n1435, n913, n915, n1423);
or   g1496 (n1512, n926, n1424, n908);
xor  g1497 (n1517, n932, n912, n1427, n927);
xnor g1498 (n1529, n934, n1426, n1439, n933);
or   g1499 (n1519, n910, n930, n1444, n918);
xnor g1500 (n1532, n1432, n1441, n914, n1425);
nand g1501 (n1530, n929, n1433, n1425, n1429);
nand g1502 (n1549, n972, n965, n959, n1523);
nor  g1503 (n1547, n961, n950, n1534, n968);
nand g1504 (n1552, n1517, n1522, n980, n968);
xnor g1505 (n1536, n1532, n963, n967, n949);
and  g1506 (n1542, n975, n1521, n943, n941);
nor  g1507 (n1548, n1520, n971, n964, n979);
nand g1508 (n1545, n969, n955, n1525, n945);
nor  g1509 (n1540, n948, n956, n962, n1529);
xnor g1510 (n1553, n944, n958, n1533, n1527);
xnor g1511 (n1539, n1526, n969, n1524, n967);
nand g1512 (n1535, n966, n978, n972, n975);
and  g1513 (n1544, n946, n938, n942, n976);
xnor g1514 (n1537, n1530, n977, n954, n1518);
xor  g1515 (n1554, n966, n952, n939, n937);
nand g1516 (n1551, n940, n957, n976, n1531);
xnor g1517 (n1538, n947, n974, n978, n960);
nand g1518 (n1550, n977, n953, n970, n1515);
xor  g1519 (n1546, n979, n1528, n973, n1516);
nand g1520 (n1543, n971, n965, n936, n973);
or   g1521 (n1541, n1519, n974, n970, n951);
xnor g1522 (n1583, n1488, n1504, n1535, n1546);
nor  g1523 (n1602, n1458, n1238, n1490, n1497);
nand g1524 (n1564, n1493, n1464, n1219, n1536);
or   g1525 (n1556, n1280, n1220, n1552, n1239);
xor  g1526 (n1629, n1237, n1231, n1451, n1537);
and  g1527 (n1620, n1470, n1230, n1550, n1448);
or   g1528 (n1569, n1228, n1541, n1238, n981);
or   g1529 (n1597, n1242, n1491, n1234, n1504);
or   g1530 (n1580, n1225, n1465, n1461, n1227);
xor  g1531 (n1560, n1473, n1501, n1228, n1225);
nand g1532 (n1598, n1455, n1243, n1454, n1551);
nand g1533 (n1603, n1487, n1550, n1229, n1462);
or   g1534 (n1558, n1237, n1486, n1541, n1496);
xnor g1535 (n1586, n1552, n980, n1449, n1497);
xnor g1536 (n1605, n1236, n1551, n1550, n1337);
or   g1537 (n1613, n1453, n1341, n1222, n1485);
xnor g1538 (n1610, n1234, n1474, n1336, n1468);
xnor g1539 (n1594, n1553, n1463, n1465, n1538);
xnor g1540 (n1608, n1220, n1547, n1242, n1552);
and  g1541 (n1557, n1539, n1241, n1552, n1225);
or   g1542 (n1596, n1503, n1229, n1494, n1538);
xnor g1543 (n1599, n1478, n1222, n1230, n1542);
and  g1544 (n1614, n1535, n1478, n1543, n1233);
or   g1545 (n1606, n1501, n1486, n1549, n1230);
nor  g1546 (n1567, n1479, n1457, n1240, n1336);
xor  g1547 (n1615, n1241, n1545, n1455, n1338);
nor  g1548 (n1621, n1548, n1544, n1240);
and  g1549 (n1625, n1541, n1448, n1227, n1468);
and  g1550 (n1585, n1343, n1237, n1540, n1227);
xnor g1551 (n1633, n1224, n1461, n1537, n1547);
and  g1552 (n1588, n1537, n1231, n1500, n1471);
nand g1553 (n1563, n1545, n1467, n1498, n1243);
and  g1554 (n1581, n1543, n1475, n1459, n1240);
nand g1555 (n1611, n1484, n1229, n1554, n1502);
nor  g1556 (n1626, n1449, n1537, n1238, n1477);
nor  g1557 (n1573, n1499, n1340, n1226, n1221);
nor  g1558 (n1570, n1502, n1219, n1551, n1340);
xnor g1559 (n1582, n1543, n1554, n1244, n1553);
xor  g1560 (n1619, n1343, n1554, n1234, n1452);
nand g1561 (n1562, n1472, n1540, n1232, n1490);
and  g1562 (n1577, n1550, n1223, n1231);
xnor g1563 (n1624, n1495, n1541, n1244, n1496);
nor  g1564 (n1631, n1542, n1228, n1222, n1500);
or   g1565 (n1604, n1548, n1482, n1227, n1236);
xor  g1566 (n1571, n1339, n1456, n1481, n1548);
nand g1567 (n1575, n1458, n1553, n1491, n1239);
or   g1568 (n1616, n1456, n1547, n1224, n1538);
xnor g1569 (n1600, n1549, n1228, n1476, n1232);
xor  g1570 (n1630, n1244, n1553, n1235, n1453);
xor  g1571 (n1555, n1536, n1235, n1244, n1494);
or   g1572 (n1618, n1538, n1452, n1549, n1220);
and  g1573 (n1609, n1482, n1457, n1239, n1226);
and  g1574 (n1634, n1226, n1466, n1549, n1475);
nand g1575 (n1559, n1454, n1471, n1542);
nand g1576 (n1632, n1466, n1544, n1480, n1505);
nand g1577 (n1576, n1242, n1451, n1503, n1243);
nor  g1578 (n1593, n1235, n1460, n1243, n1484);
xor  g1579 (n1574, n1545, n1535, n1342, n1474);
xnor g1580 (n1622, n1221, n1477, n1223, n1495);
nor  g1581 (n1565, n1535, n1498, n1479, n1222);
nor  g1582 (n1578, n1470, n1551, n1480, n1539);
and  g1583 (n1579, n1499, n1229, n672, n1337);
nand g1584 (n1584, n1536, n1242, n1492, n1221);
xor  g1585 (n1572, n1493, n1546, n1232, n1224);
nand g1586 (n1623, n1489, n1241, n1481, n1544);
and  g1587 (n1607, n1540, n1240, n1543, n1230);
or   g1588 (n1591, n1232, n1459, n1338, n1223);
or   g1589 (n1601, n1467, n1241, n1539, n1341);
and  g1590 (n1592, n1473, n1239, n1476, n1463);
or   g1591 (n1589, n1236, n1548, n1342, n1546);
xnor g1592 (n1568, n1536, n1483, n1238, n1450);
and  g1593 (n1627, n1450, n1233, n1539, n1483);
and  g1594 (n1628, n1487, n1488, n1221, n1231);
and  g1595 (n1595, n1472, n1545, n1464, n1460);
and  g1596 (n1590, n1219, n1492, n1462, n1220);
and  g1597 (n1561, n1469, n1234, n1489, n1485);
nand g1598 (n1587, n1469, n1225, n1219, n1233);
and  g1599 (n1612, n1546, n672, n1554, n1233);
and  g1600 (n1566, n1224, n1236, n1540, n1226);
nand g1601 (n1617, n1547, n1339, n1235, n1237);
not  g1602 (n1656, n1569);
not  g1603 (n1660, n986);
not  g1604 (n1671, n981);
buf  g1605 (n1648, n1557);
not  g1606 (n1642, n1562);
not  g1607 (n1658, n1556);
buf  g1608 (n1677, n1572);
not  g1609 (n1649, n1570);
buf  g1610 (n1657, n1555);
not  g1611 (n1667, n1559);
not  g1612 (n1652, n1573);
buf  g1613 (n1636, n988);
buf  g1614 (n1666, n1561);
buf  g1615 (n1672, n1564);
not  g1616 (n1640, n1571);
not  g1617 (n1646, n989);
not  g1618 (n1674, n1566);
buf  g1619 (n1668, n1565);
not  g1620 (n1654, n1558);
buf  g1621 (n1673, n984);
not  g1622 (n1639, n990);
buf  g1623 (n1661, n987);
not  g1624 (n1635, n986);
not  g1625 (n1675, n1555);
not  g1626 (n1647, n988);
buf  g1627 (n1664, n1569);
not  g1628 (n1645, n1558);
not  g1629 (n1651, n1562);
not  g1630 (n1659, n982);
not  g1631 (n1637, n1574);
buf  g1632 (n1663, n989);
buf  g1633 (n1655, n983);
buf  g1634 (n1641, n987);
not  g1635 (n1669, n1576);
not  g1636 (n1665, n1568);
nand g1637 (n1670, n1575, n1574, n1567);
and  g1638 (n1676, n1567, n1572, n1571);
xor  g1639 (n1650, n1573, n985, n1557);
xor  g1640 (n1678, n984, n1575, n1576);
nor  g1641 (n1638, n1563, n1565, n1564);
nor  g1642 (n1644, n1568, n1570, n983);
nand g1643 (n1643, n982, n1563, n1560);
nor  g1644 (n1653, n1556, n985, n1566);
xor  g1645 (n1662, n1560, n1559, n1561);
nand g1646 (n1692, n1644, n1026, n1009, n993);
nor  g1647 (n1694, n1036, n992, n1649, n994);
and  g1648 (n1691, n1040, n1648, n994, n1022);
xnor g1649 (n1690, n1013, n1038, n1650, n1002);
nor  g1650 (n1704, n1017, n1020, n1015, n1016);
xnor g1651 (n1703, n1639, n999, n1039, n997);
xor  g1652 (n1710, n1003, n1642, n1008, n1640);
xnor g1653 (n1687, n1640, n1642, n1008, n1003);
nand g1654 (n1701, n1024, n1649, n1036, n1646);
xor  g1655 (n1712, n993, n1002, n1010, n1037);
xnor g1656 (n1683, n1031, n999, n1636, n1011);
nand g1657 (n1679, n1012, n1647, n1022, n1637);
xor  g1658 (n1707, n1035, n1032, n998);
nand g1659 (n1711, n1024, n1007, n1019, n1006);
nand g1660 (n1695, n1027, n990, n1011, n1641);
nor  g1661 (n1686, n1001, n1643, n1021, n1030);
nor  g1662 (n1682, n1016, n996, n1649, n1033);
or   g1663 (n1684, n1031, n1018, n1004, n1015);
xor  g1664 (n1689, n1006, n1635, n1010, n1644);
nand g1665 (n1681, n1638, n1001, n997, n1000);
xnor g1666 (n1702, n991, n1005, n1034, n1028);
xnor g1667 (n1700, n1636, n1637, n991, n1012);
nand g1668 (n1709, n1035, n1014, n1643, n995);
nand g1669 (n1708, n1041, n992, n1019, n1039);
xnor g1670 (n1685, n1026, n1000, n1025);
and  g1671 (n1693, n1645, n1649, n1639, n1032);
or   g1672 (n1688, n1021, n1638, n1005, n1028);
xor  g1673 (n1680, n1650, n1017, n1029, n1645);
or   g1674 (n1698, n1648, n1029, n1641, n995);
xor  g1675 (n1706, n1004, n1635, n1009, n1646);
xor  g1676 (n1705, n1027, n1007, n1023, n1034);
nand g1677 (n1699, n1038, n1023, n1040, n1033);
nand g1678 (n1696, n996, n1037, n1647, n1020);
xor  g1679 (n1697, n1030, n1018, n1013, n1014);
and  g1680 (n1719, n1685, n1358, n1290, n1712);
and  g1681 (n1730, n1683, n1691, n1706, n1353);
and  g1682 (n1723, n1352, n1298, n1346, n1702);
nor  g1683 (n1714, n1297, n1303, n1357, n1286);
xor  g1684 (n1721, n1682, n1346, n1301, n1306);
xor  g1685 (n1727, n1351, n1284, n1359, n1293);
or   g1686 (n1732, n1292, n1681, n1290, n1709);
nand g1687 (n1725, n1304, n1288, n1306, n1308);
nor  g1688 (n1720, n1361, n1299, n1689, n1697);
or   g1689 (n1737, n1042, n1345, n1308, n1693);
nand g1690 (n1746, n1304, n1284, n1291, n1345);
xnor g1691 (n1716, n1679, n1347, n1043, n1344);
nand g1692 (n1736, n1360, n1298, n1359, n1355);
or   g1693 (n1739, n1291, n1686, n1353, n1280);
xor  g1694 (n1741, n1043, n1283, n1699, n1297);
nor  g1695 (n1743, n1688, n1700, n1349, n1306);
nand g1696 (n1731, n1687, n1293, n1710, n1360);
xnor g1697 (n1728, n1287, n1354, n1307);
xor  g1698 (n1729, n1283, n1684, n1305, n1348);
nor  g1699 (n1718, n1707, n1692, n1344, n1350);
xor  g1700 (n1742, n1303, n1300, n1296, n1695);
xnor g1701 (n1747, n1705, n1650, n1711, n1042);
nor  g1702 (n1745, n1351, n1289, n1282, n1307);
nand g1703 (n1744, n1281, n1302, n1294, n1295);
nand g1704 (n1740, n1289, n1305, n1698, n1299);
or   g1705 (n1738, n1708, n1690, n1307, n1308);
nand g1706 (n1726, n1350, n1357, n1358, n1282);
and  g1707 (n1713, n1712, n1704, n1696, n1286);
nand g1708 (n1715, n1292, n1356, n1285, n1348);
xor  g1709 (n1717, n1349, n1044, n1356, n1703);
and  g1710 (n1724, n1307, n1694, n1288, n1302);
xor  g1711 (n1722, n1295, n1300, n1355, n1308);
xnor g1712 (n1734, n1352, n1281, n1294, n1347);
nand g1713 (n1733, n1287, n1701, n1044, n1285);
and  g1714 (n1735, n1301, n1041, n1680, n1296);
not  g1715 (n1872, n1659);
buf  g1716 (n1815, n1731);
buf  g1717 (n1881, n1672);
buf  g1718 (n1852, n1621);
buf  g1719 (n1846, n1584);
not  g1720 (n1874, n1599);
not  g1721 (n1779, n1725);
not  g1722 (n1788, n1585);
not  g1723 (n1842, n1362);
not  g1724 (n1825, n1596);
buf  g1725 (n1835, n1740);
not  g1726 (n1878, n1737);
not  g1727 (n1887, n1677);
not  g1728 (n1804, n1660);
buf  g1729 (n1829, n1594);
not  g1730 (n1850, n1746);
buf  g1731 (n1860, n1734);
buf  g1732 (n1773, n1724);
not  g1733 (n1751, n1593);
buf  g1734 (n1856, n1579);
buf  g1735 (n1799, n1580);
not  g1736 (n1843, n1665);
buf  g1737 (n1752, n1737);
buf  g1738 (n1851, n1598);
buf  g1739 (n1783, n1677);
buf  g1740 (n1778, n1731);
not  g1741 (n1816, n1659);
not  g1742 (n1823, n1583);
not  g1743 (n1848, n1667);
buf  g1744 (n1865, n1590);
and  g1745 (n1784, n1747, n1722, n1728, n1614);
nand g1746 (n1828, n1670, n1656, n1621, n1619);
or   g1747 (n1885, n1598, n1585, n1673, n1593);
nand g1748 (n1786, n1584, n1651, n1599, n1594);
or   g1749 (n1834, n1726, n1599, n1678, n1658);
nand g1750 (n1847, n1617, n1579, n1656, n1253);
nand g1751 (n1830, n1722, n1746, n1591, n1656);
and  g1752 (n1812, n1622, n1612, n1587, n1590);
xor  g1753 (n1871, n1740, n1673, n1666, n1587);
xor  g1754 (n1781, n1723, n1605, n1604, n1603);
xnor g1755 (n1798, n1715, n1602, n1723, n1719);
and  g1756 (n1800, n1739, n1601, n1604, n1738);
nor  g1757 (n1775, n1595, n1652, n1593, n1713);
xnor g1758 (n1782, n1511, n1651, n1668, n1587);
nor  g1759 (n1749, n1659, n1595, n1657, n1728);
nor  g1760 (n1765, n1611, n1669, n1605, n1725);
xnor g1761 (n1794, n1653, n1615, n1743, n1597);
or   g1762 (n1755, n1661, n1738, n1510, n1735);
xor  g1763 (n1787, n1661, n1670, n1595, n1591);
or   g1764 (n1813, n1721, n1651, n1731, n1677);
and  g1765 (n1753, n1587, n1678, n1722, n1578);
or   g1766 (n1831, n1719, n1589, n1361, n1577);
and  g1767 (n1771, n1729, n1721, n1741, n1601);
nor  g1768 (n1760, n1717, n1730, n1665, n1668);
nand g1769 (n1803, n1662, n1720, n1617, n1603);
xnor g1770 (n1886, n1579, n1667, n1670, n1606);
xor  g1771 (n1821, n1592, n1658, n1650, n1713);
xnor g1772 (n1818, n1618, n1662, n1596, n1742);
xor  g1773 (n1868, n1254, n1506, n1593, n1608);
and  g1774 (n1777, n1724, n1677, n1582, n1590);
xor  g1775 (n1884, n1715, n1599, n1655, n1718);
xor  g1776 (n1845, n1617, n1747, n1676, n1507);
nand g1777 (n1750, n1662, n1715, n1586, n1727);
xor  g1778 (n1841, n1747, n1601, n1734, n1727);
xor  g1779 (n1795, n1616, n1663, n1747, n1364);
and  g1780 (n1807, n1368, n1730, n1576, n1745);
nand g1781 (n1748, n1675, n1620, n1612, n1591);
and  g1782 (n1801, n1718, n1743, n1717, n1746);
xor  g1783 (n1849, n1676, n1611, n1608, n1509);
or   g1784 (n1822, n1669, n1673, n1652, n1720);
or   g1785 (n1776, n1713, n1744, n1607, n1254);
and  g1786 (n1767, n1675, n1620, n1728, n1589);
or   g1787 (n1817, n1614, n1589, n1676, n1714);
xor  g1788 (n1757, n1672, n1727, n1740, n1678);
xnor g1789 (n1802, n1675, n1724, n1585, n1657);
nor  g1790 (n1855, n1674, n1595, n1733, n1613);
xnor g1791 (n1797, n1662, n1658, n1580, n1741);
and  g1792 (n1863, n1672, n1735, n1665, n1600);
xor  g1793 (n1873, n1612, n1654, n1576, n1603);
xor  g1794 (n1811, n1605, n1718, n1732, n1582);
xor  g1795 (n1769, n1732, n1602, n1586, n1610);
xor  g1796 (n1870, n1742, n1584, n1716, n1664);
nor  g1797 (n1770, n1606, n1583, n1659);
nor  g1798 (n1754, n1509, n1734, n1668, n1735);
and  g1799 (n1790, n1602, n1658, n1678, n1508);
xor  g1800 (n1862, n1724, n1614, n1620, n1507);
or   g1801 (n1761, n1582, n1738, n1667, n1741);
xor  g1802 (n1858, n1739, n1668, n1725, n1652);
and  g1803 (n1806, n1588, n1745, n1616, n1729);
nor  g1804 (n1796, n1666, n1592, n1598, n1743);
or   g1805 (n1789, n1620, n1714, n1590, n1676);
xor  g1806 (n1772, n1666, n1674, n1723, n1510);
nor  g1807 (n1762, n1739, n1610, n1716);
nor  g1808 (n1808, n1600, n1669, n1609, n1592);
or   g1809 (n1832, n1664, n1743, n1615, n1657);
and  g1810 (n1759, n1365, n1718, n1651, n1655);
and  g1811 (n1861, n1733, n1732, n1614, n1586);
nand g1812 (n1864, n1671, n1654, n1665, n1669);
xnor g1813 (n1866, n1720, n1744, n1730, n1663);
xor  g1814 (n1814, n1254, n1580, n1654, n1602);
nand g1815 (n1844, n1588, n1729, n1578, n1736);
xnor g1816 (n1826, n1745, n1615, n1732);
xnor g1817 (n1791, n1608, n1616, n1715, n1594);
or   g1818 (n1840, n1672, n1613, n1674, n1621);
and  g1819 (n1877, n1742, n1663, n1577, n1604);
nand g1820 (n1879, n1363, n1365, n1596, n1674);
and  g1821 (n1763, n1607, n1612, n1606, n1740);
nor  g1822 (n1827, n1581, n1607, n1654, n1652);
nand g1823 (n1854, n1733, n1661, n1577, n1585);
nand g1824 (n1766, n1577, n1367, n1363, n1741);
and  g1825 (n1824, n1622, n1609, n1616, n1619);
nor  g1826 (n1756, n1734, n1597, n1656, n1746);
and  g1827 (n1838, n1738, n1719, n1739, n1609);
and  g1828 (n1867, n1671, n1725, n1619, n1714);
or   g1829 (n1792, n1506, n1610, n1663, n1660);
nor  g1830 (n1880, n1596, n1254, n1736, n1597);
xnor g1831 (n1768, n1366, n1720, n1717, n1726);
nor  g1832 (n1857, n1613, n1611, n1664, n1737);
and  g1833 (n1819, n1600, n1723, n1735, n1714);
xnor g1834 (n1810, n1660, n1716, n1584, n1582);
nand g1835 (n1883, n1727, n1675, n1671, n1655);
and  g1836 (n1809, n1673, n1578, n1744, n1742);
xnor g1837 (n1837, n1717, n1736, n1728, n1716);
nor  g1838 (n1836, n1364, n1609, n1591, n1597);
xnor g1839 (n1820, n1580, n1617, n1729, n1598);
xor  g1840 (n1882, n1594, n1621, n1653, n1613);
or   g1841 (n1793, n1606, n1670, n1588, n1737);
nand g1842 (n1876, n1511, n1618, n1603, n1721);
xor  g1843 (n1785, n1588, n1730, n1721, n1736);
and  g1844 (n1869, n1666, n1618, n1719, n1722);
xor  g1845 (n1780, n1367, n1592, n1726, n1366);
nand g1846 (n1853, n1661, n1508, n1586, n1505);
or   g1847 (n1833, n1733, n1660, n1657, n1604);
and  g1848 (n1764, n1745, n1671, n1619, n1368);
and  g1849 (n1875, n1608, n1653, n1601, n1605);
nor  g1850 (n1758, n1726, n1744, n1581, n1362);
nor  g1851 (n1774, n1618, n1600, n1667, n1611);
nor  g1852 (n1859, n1713, n1589, n1731, n1653);
xor  g1853 (n1839, n1664, n1578, n1581);
nor  g1854 (n1805, n1607, n1655, n1583, n1579);
xor  g1855 (n1952, n1080, n1153, n1143, n1772);
nand g1856 (n1998, n1627, n1816, n1855, n1045);
xor  g1857 (n1979, n1828, n1082, n1124, n1080);
xor  g1858 (n1934, n1622, n1172, n1860, n1760);
nand g1859 (n1955, n1156, n1624, n1754, n1084);
nor  g1860 (n1961, n1761, n1096, n1178, n1633);
nand g1861 (n1903, n1046, n1858, n1105, n1058);
nand g1862 (n1974, n1112, n1623, n1804, n1628);
and  g1863 (n1990, n1166, n1775, n1631, n1849);
or   g1864 (n1969, n1148, n1123, n1070, n1054);
nand g1865 (n1892, n1848, n1865, n1845, n1843);
and  g1866 (n2001, n1134, n1164, n1630, n1048);
and  g1867 (n1931, n1078, n1148, n1140, n1066);
or   g1868 (n1929, n1814, n1624, n1864, n1626);
and  g1869 (n2002, n1752, n1048, n1130, n1116);
and  g1870 (n1935, n1085, n1881, n1629, n1105);
or   g1871 (n1973, n1057, n1052, n1759, n1132);
nor  g1872 (n1893, n1630, n1162, n1099, n1807);
xnor g1873 (n1991, n1825, n1079, n1126, n1869);
xor  g1874 (n1959, n1076, n1175, n1832, n1120);
nor  g1875 (n1986, n1853, n1096, n1846, n1109);
or   g1876 (n1971, n1111, n1115, n1072, n1103);
xor  g1877 (n1904, n1632, n1753, n1107, n1145);
xnor g1878 (n1932, n1762, n1049, n1167, n1854);
xor  g1879 (n1949, n1113, n1622, n1070, n1075);
nor  g1880 (n1890, n1887, n1780, n1133, n1122);
xnor g1881 (n1977, n1632, n1836, n1179, n1131);
and  g1882 (n1916, n1063, n1093, n1626, n1176);
or   g1883 (n1924, n1794, n1824, n1068, n1155);
and  g1884 (n1936, n1058, n1169, n1086, n1758);
xor  g1885 (n1976, n1790, n1177, n1136, n1059);
nor  g1886 (n1941, n1776, n1162, n1090, n1151);
xor  g1887 (n1913, n1088, n1050, n1630, n1808);
xnor g1888 (n1911, n1119, n1629, n1118, n1114);
xor  g1889 (n1888, n1095, n1047, n1128, n1066);
and  g1890 (n1915, n1628, n1781, n1081, n1885);
nand g1891 (n1899, n1166, n1108, n1065, n1149);
nand g1892 (n1950, n1053, n1139, n1101, n1176);
nor  g1893 (n1997, n1763, n1160, n1073, n1154);
and  g1894 (n1953, n1822, n1144, n1173, n1632);
xnor g1895 (n1962, n1631, n1099, n1883, n1076);
nand g1896 (n1920, n1631, n1150, n1815, n1056);
nand g1897 (n1907, n1121, n1056, n1112, n1633);
and  g1898 (n1943, n1051, n1094, n1135, n1626);
xnor g1899 (n1895, n1168, n1059, n1634, n1764);
or   g1900 (n1933, n1625, n1805, n1046, n1870);
and  g1901 (n1967, n1767, n1175, n1130, n1095);
or   g1902 (n1926, n1097, n1793, n1084, n1788);
nand g1903 (n1984, n1092, n1068, n1127, n1077);
and  g1904 (n1921, n1871, n1147, n1629, n1069);
xor  g1905 (n1958, n1072, n1167, n1135, n1139);
nand g1906 (n1889, n1839, n1784, n1811, n1057);
xnor g1907 (n1891, n1078, n1168, n1796, n1134);
xor  g1908 (n1988, n1124, n1777, n1109, n1180);
xor  g1909 (n1945, n1089, n1623, n1110, n1091);
xnor g1910 (n1951, n1097, n1876, n1129, n1170);
xor  g1911 (n1939, n1165, n1868, n1633, n1768);
nand g1912 (n1938, n1053, n1098, n1144, n1074);
xor  g1913 (n1906, n1634, n1071, n1102, n1833);
nor  g1914 (n1937, n1067, n1156, n1789, n1061);
and  g1915 (n1994, n1077, n1857, n1838, n1089);
nor  g1916 (n2000, n1114, n1091, n1157, n1104);
xnor g1917 (n1970, n1803, n1823, n1634, n1103);
or   g1918 (n2003, n1136, n1062, n1785, n1120);
or   g1919 (n1894, n1625, n1161, n1791, n1840);
nor  g1920 (n1946, n1797, n1131, n1141, n1847);
or   g1921 (n1930, n1631, n1145, n1875, n1111);
and  g1922 (n1978, n1169, n1122, n1164, n1809);
or   g1923 (n1897, n1094, n1118, n1163, n1137);
xor  g1924 (n1987, n1799, n1877, n1143, n1866);
and  g1925 (n1908, n1829, n1123, n1770, n1159);
and  g1926 (n1964, n1060, n1101, n1882, n1831);
xnor g1927 (n1914, n1082, n1125, n1117, n1088);
xor  g1928 (n1972, n1750, n1792, n1063, n1627);
and  g1929 (n1923, n1756, n1093, n1632, n1774);
and  g1930 (n1960, n1142, n1087, n1100, n1121);
and  g1931 (n1965, n1065, n1817, n1126, n1782);
xnor g1932 (n1925, n1152, n1067, n1051, n1138);
and  g1933 (n1901, n1117, n1771, n1623, n1787);
nor  g1934 (n1948, n1623, n1630, n1830, n1073);
xor  g1935 (n1956, n1769, n1173, n1062, n1075);
or   g1936 (n1980, n1624, n1872, n1826, n1625);
nand g1937 (n1902, n1874, n1154, n1060, n1172);
nand g1938 (n1968, n1102, n1125, n1628, n1174);
and  g1939 (n1975, n1813, n1786, n1779, n1844);
xnor g1940 (n1989, n1879, n1778, n1810, n1146);
and  g1941 (n1905, n1171, n1626, n1884, n1054);
and  g1942 (n1940, n1069, n1064, n1147, n1106);
nand g1943 (n1900, n1087, n1064, n1181, n1174);
and  g1944 (n1957, n1127, n1079, n1106, n1055);
or   g1945 (n1954, n1100, n1842, n1783, n1165);
nor  g1946 (n1942, n1812, n1146, n1878, n1170);
nor  g1947 (n1985, n1798, n1801, n1757, n1116);
or   g1948 (n1996, n1795, n1171, n1629, n1104);
xor  g1949 (n1917, n1049, n1083, n1625, n1863);
or   g1950 (n1898, n1153, n1110, n1755, n1841);
xor  g1951 (n1928, n1634, n1806, n1050, n1862);
or   g1952 (n1966, n1155, n1074, n1835, n1128);
nand g1953 (n1999, n1098, n1047, n1867, n1802);
nor  g1954 (n1918, n1129, n1142, n1873, n1071);
or   g1955 (n1912, n1751, n1137, n1819, n1851);
xor  g1956 (n1963, n1800, n1765, n1119, n1180);
nand g1957 (n1927, n1179, n1856, n1820, n1052);
and  g1958 (n1983, n1766, n1108, n1859, n1045);
xnor g1959 (n1919, n1083, n1627, n1161, n1749);
xnor g1960 (n1922, n1834, n1821, n1149, n1627);
or   g1961 (n1982, n1886, n1133, n1132, n1138);
xor  g1962 (n1944, n1055, n1141, n1061, n1178);
nor  g1963 (n1947, n1090, n1181, n1151, n1818);
xor  g1964 (n1981, n1850, n1107, n1159, n1773);
nand g1965 (n1909, n1086, n1633, n1092, n1628);
and  g1966 (n1910, n1163, n1113, n1081, n1880);
and  g1967 (n1993, n1150, n1152, n1748, n1158);
nand g1968 (n1992, n1160, n1827, n1115, n1861);
and  g1969 (n1896, n1158, n1852, n1177, n1085);
xnor g1970 (n1995, n1837, n1624, n1140, n1157);
xor  g1971 (n2030, n1991, n1897, n1893, n1894);
or   g1972 (n2008, n1984, n1961, n1949, n1934);
xnor g1973 (n2032, n1924, n1977, n1923, n2002);
xnor g1974 (n2027, n1992, n1953, n1936, n1922);
and  g1975 (n2025, n1948, n1963, n1909, n1969);
nor  g1976 (n2020, n1906, n1929, n1890, n1899);
or   g1977 (n2004, n1937, n1965, n1892, n1968);
nor  g1978 (n2024, n1966, n1938, n1927, n1939);
xnor g1979 (n2022, n1935, n1970, n1898, n1981);
xnor g1980 (n2013, n1987, n1913, n1996, n1914);
and  g1981 (n2023, n1978, n1976, n1955, n1960);
nor  g1982 (n2016, n1990, n1988, n1904, n1905);
nor  g1983 (n2012, n1980, n1989, n1896, n1926);
nand g1984 (n2006, n1907, n1947, n1908, n1903);
and  g1985 (n2005, n1888, n1986, n1917, n1925);
xor  g1986 (n2021, n1999, n1982, n1958, n1933);
and  g1987 (n2010, n1891, n1983, n1997, n1956);
nor  g1988 (n2026, n1943, n1951, n1971, n1920);
xor  g1989 (n2017, n1889, n1918, n1952, n1957);
and  g1990 (n2031, n1919, n1942, n1912, n1915);
nand g1991 (n2029, n1972, n1901, n2000, n1973);
and  g1992 (n2009, n1946, n1979, n1944, n1985);
xor  g1993 (n2015, n1967, n1998, n1930, n1964);
xnor g1994 (n2019, n1959, n1975, n1902, n1921);
or   g1995 (n2018, n2003, n1932, n1974, n1940);
nand g1996 (n2014, n1931, n1995, n2001, n1916);
nor  g1997 (n2007, n1910, n1950, n1962, n1994);
nand g1998 (n2011, n1928, n1945, n1954, n1941);
xnor g1999 (n2028, n1993, n1911, n1895, n1900);
endmodule
