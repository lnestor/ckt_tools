

module Stat_3000_305
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1538,
  n2983,
  n2981,
  n2989,
  n2980,
  n2986,
  n2985,
  n2988,
  n2982,
  n2984,
  n3019,
  n3026,
  n3013,
  n3032,
  n3020,
  n3018,
  n3022,
  n3015,
  n3027,
  n3017,
  n3012,
  n3024,
  n3021,
  n3016,
  n3029,
  n3011,
  n3025,
  n3014,
  n3028,
  n3023,
  n3031,
  n3030,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1538;output n2983;output n2981;output n2989;output n2980;output n2986;output n2985;output n2988;output n2982;output n2984;output n3019;output n3026;output n3013;output n3032;output n3020;output n3018;output n3022;output n3015;output n3027;output n3017;output n3012;output n3024;output n3021;output n3016;output n3029;output n3011;output n3025;output n3014;output n3028;output n3023;output n3031;output n3030;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2987;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n74,
    n13
  );


  not
  g1
  (
    n56,
    n8
  );


  not
  g2
  (
    n52,
    n1
  );


  not
  g3
  (
    n55,
    n2
  );


  not
  g4
  (
    n79,
    n1
  );


  buf
  g5
  (
    n92,
    n7
  );


  buf
  g6
  (
    n82,
    n17
  );


  buf
  g7
  (
    n36,
    n3
  );


  buf
  g8
  (
    n85,
    n2
  );


  buf
  g9
  (
    n95,
    n13
  );


  not
  g10
  (
    n46,
    n10
  );


  not
  g11
  (
    n66,
    n3
  );


  buf
  g12
  (
    n65,
    n16
  );


  not
  g13
  (
    n96,
    n15
  );


  not
  g14
  (
    n60,
    n16
  );


  not
  g15
  (
    n70,
    n10
  );


  not
  g16
  (
    n86,
    n7
  );


  buf
  g17
  (
    n48,
    n17
  );


  buf
  g18
  (
    n83,
    n12
  );


  buf
  g19
  (
    n64,
    n13
  );


  not
  g20
  (
    n37,
    n1
  );


  buf
  g21
  (
    n59,
    n10
  );


  not
  g22
  (
    n87,
    n2
  );


  not
  g23
  (
    n51,
    n3
  );


  buf
  g24
  (
    n54,
    n4
  );


  buf
  g25
  (
    n98,
    n13
  );


  not
  g26
  (
    n97,
    n6
  );


  buf
  g27
  (
    n80,
    n14
  );


  buf
  g28
  (
    n40,
    n2
  );


  not
  g29
  (
    n71,
    n11
  );


  buf
  g30
  (
    n76,
    n5
  );


  buf
  g31
  (
    n49,
    n3
  );


  buf
  g32
  (
    n63,
    n7
  );


  buf
  g33
  (
    n43,
    n6
  );


  buf
  g34
  (
    n90,
    n12
  );


  not
  g35
  (
    n39,
    n5
  );


  buf
  g36
  (
    n45,
    n14
  );


  buf
  g37
  (
    n69,
    n8
  );


  not
  g38
  (
    n75,
    n6
  );


  not
  g39
  (
    n73,
    n9
  );


  not
  g40
  (
    n34,
    n4
  );


  not
  g41
  (
    n38,
    n12
  );


  not
  g42
  (
    n77,
    n16
  );


  buf
  g43
  (
    n47,
    n16
  );


  buf
  g44
  (
    n57,
    n9
  );


  buf
  g45
  (
    n41,
    n9
  );


  not
  g46
  (
    n33,
    n4
  );


  not
  g47
  (
    n78,
    n14
  );


  buf
  g48
  (
    n67,
    n4
  );


  buf
  g49
  (
    n62,
    n14
  );


  not
  g50
  (
    n91,
    n5
  );


  buf
  g51
  (
    n58,
    n8
  );


  not
  g52
  (
    n35,
    n12
  );


  buf
  g53
  (
    n61,
    n10
  );


  buf
  g54
  (
    n42,
    n11
  );


  buf
  g55
  (
    n84,
    n15
  );


  not
  g56
  (
    n72,
    n7
  );


  buf
  g57
  (
    n94,
    n5
  );


  buf
  g58
  (
    n81,
    n15
  );


  buf
  g59
  (
    n89,
    n8
  );


  not
  g60
  (
    n68,
    n11
  );


  not
  g61
  (
    n50,
    n6
  );


  buf
  g62
  (
    n44,
    n15
  );


  not
  g63
  (
    n53,
    n1
  );


  not
  g64
  (
    n88,
    n9
  );


  not
  g65
  (
    n93,
    n11
  );


  not
  g66
  (
    n172,
    n44
  );


  not
  g67
  (
    n275,
    n48
  );


  buf
  g68
  (
    n244,
    n60
  );


  buf
  g69
  (
    n139,
    n33
  );


  not
  g70
  (
    n138,
    n75
  );


  not
  g71
  (
    n196,
    n64
  );


  buf
  g72
  (
    n214,
    n67
  );


  buf
  g73
  (
    n204,
    n49
  );


  not
  g74
  (
    n140,
    n34
  );


  not
  g75
  (
    n248,
    n77
  );


  not
  g76
  (
    n199,
    n47
  );


  not
  g77
  (
    n239,
    n45
  );


  not
  g78
  (
    n185,
    n74
  );


  buf
  g79
  (
    n187,
    n71
  );


  buf
  g80
  (
    n141,
    n55
  );


  not
  g81
  (
    n205,
    n74
  );


  not
  g82
  (
    n175,
    n53
  );


  buf
  g83
  (
    n206,
    n72
  );


  buf
  g84
  (
    n266,
    n76
  );


  buf
  g85
  (
    n112,
    n46
  );


  buf
  g86
  (
    n170,
    n61
  );


  buf
  g87
  (
    n146,
    n47
  );


  buf
  g88
  (
    n237,
    n55
  );


  buf
  g89
  (
    n260,
    n63
  );


  not
  g90
  (
    n166,
    n36
  );


  buf
  g91
  (
    n182,
    n37
  );


  not
  g92
  (
    n270,
    n50
  );


  not
  g93
  (
    n156,
    n36
  );


  buf
  g94
  (
    n122,
    n39
  );


  buf
  g95
  (
    n202,
    n41
  );


  not
  g96
  (
    n251,
    n63
  );


  buf
  g97
  (
    n176,
    n69
  );


  buf
  g98
  (
    n255,
    n38
  );


  buf
  g99
  (
    n119,
    n65
  );


  buf
  g100
  (
    n236,
    n52
  );


  not
  g101
  (
    n179,
    n63
  );


  not
  g102
  (
    n133,
    n78
  );


  buf
  g103
  (
    n144,
    n60
  );


  not
  g104
  (
    n128,
    n45
  );


  buf
  g105
  (
    n274,
    n47
  );


  buf
  g106
  (
    n190,
    n73
  );


  buf
  g107
  (
    n269,
    n34
  );


  buf
  g108
  (
    n117,
    n77
  );


  not
  g109
  (
    n136,
    n73
  );


  not
  g110
  (
    n225,
    n70
  );


  not
  g111
  (
    n167,
    n43
  );


  not
  g112
  (
    n178,
    n61
  );


  not
  g113
  (
    n118,
    n38
  );


  buf
  g114
  (
    n265,
    n71
  );


  buf
  g115
  (
    n183,
    n68
  );


  buf
  g116
  (
    n177,
    n42
  );


  not
  g117
  (
    n189,
    n76
  );


  buf
  g118
  (
    n252,
    n65
  );


  buf
  g119
  (
    n249,
    n33
  );


  not
  g120
  (
    n180,
    n66
  );


  buf
  g121
  (
    n173,
    n51
  );


  not
  g122
  (
    n123,
    n75
  );


  not
  g123
  (
    n147,
    n37
  );


  buf
  g124
  (
    n273,
    n54
  );


  not
  g125
  (
    n134,
    n43
  );


  buf
  g126
  (
    n235,
    n58
  );


  buf
  g127
  (
    n191,
    n36
  );


  not
  g128
  (
    n253,
    n69
  );


  not
  g129
  (
    n192,
    n45
  );


  buf
  g130
  (
    n105,
    n77
  );


  not
  g131
  (
    n127,
    n65
  );


  not
  g132
  (
    n151,
    n39
  );


  not
  g133
  (
    n233,
    n50
  );


  not
  g134
  (
    n109,
    n42
  );


  buf
  g135
  (
    n110,
    n48
  );


  buf
  g136
  (
    n230,
    n51
  );


  buf
  g137
  (
    n115,
    n78
  );


  buf
  g138
  (
    n247,
    n70
  );


  buf
  g139
  (
    n242,
    n46
  );


  not
  g140
  (
    n164,
    n52
  );


  buf
  g141
  (
    n238,
    n33
  );


  not
  g142
  (
    n174,
    n36
  );


  not
  g143
  (
    n203,
    n38
  );


  not
  g144
  (
    n113,
    n52
  );


  buf
  g145
  (
    n246,
    n58
  );


  not
  g146
  (
    n223,
    n38
  );


  not
  g147
  (
    n227,
    n63
  );


  not
  g148
  (
    n121,
    n70
  );


  not
  g149
  (
    n142,
    n74
  );


  not
  g150
  (
    n220,
    n62
  );


  buf
  g151
  (
    n217,
    n56
  );


  not
  g152
  (
    n152,
    n76
  );


  not
  g153
  (
    n163,
    n37
  );


  buf
  g154
  (
    n207,
    n68
  );


  not
  g155
  (
    n259,
    n46
  );


  buf
  g156
  (
    n268,
    n71
  );


  not
  g157
  (
    n278,
    n35
  );


  not
  g158
  (
    n150,
    n53
  );


  not
  g159
  (
    n194,
    n45
  );


  buf
  g160
  (
    n120,
    n76
  );


  not
  g161
  (
    n267,
    n66
  );


  buf
  g162
  (
    n261,
    n75
  );


  not
  g163
  (
    n102,
    n41
  );


  not
  g164
  (
    n100,
    n35
  );


  not
  g165
  (
    n201,
    n46
  );


  buf
  g166
  (
    n271,
    n72
  );


  not
  g167
  (
    n245,
    n71
  );


  not
  g168
  (
    n221,
    n48
  );


  buf
  g169
  (
    n155,
    n54
  );


  buf
  g170
  (
    n148,
    n68
  );


  not
  g171
  (
    n211,
    n62
  );


  buf
  g172
  (
    n103,
    n39
  );


  buf
  g173
  (
    n243,
    n42
  );


  buf
  g174
  (
    n209,
    n67
  );


  buf
  g175
  (
    n130,
    n73
  );


  not
  g176
  (
    n162,
    n54
  );


  buf
  g177
  (
    n272,
    n35
  );


  not
  g178
  (
    n250,
    n47
  );


  not
  g179
  (
    n226,
    n66
  );


  not
  g180
  (
    n215,
    n58
  );


  not
  g181
  (
    n108,
    n41
  );


  buf
  g182
  (
    n143,
    n59
  );


  not
  g183
  (
    n281,
    n64
  );


  buf
  g184
  (
    n213,
    n69
  );


  buf
  g185
  (
    n137,
    n34
  );


  buf
  g186
  (
    n101,
    n57
  );


  buf
  g187
  (
    n193,
    n64
  );


  not
  g188
  (
    n234,
    n34
  );


  not
  g189
  (
    n208,
    n59
  );


  buf
  g190
  (
    n228,
    n57
  );


  buf
  g191
  (
    n241,
    n78
  );


  not
  g192
  (
    n184,
    n42
  );


  not
  g193
  (
    n212,
    n43
  );


  not
  g194
  (
    n124,
    n74
  );


  not
  g195
  (
    n181,
    n62
  );


  buf
  g196
  (
    n104,
    n64
  );


  not
  g197
  (
    n231,
    n48
  );


  not
  g198
  (
    n129,
    n59
  );


  buf
  g199
  (
    n279,
    n37
  );


  not
  g200
  (
    n111,
    n54
  );


  not
  g201
  (
    n264,
    n51
  );


  not
  g202
  (
    n145,
    n50
  );


  not
  g203
  (
    n126,
    n73
  );


  buf
  g204
  (
    n276,
    n70
  );


  buf
  g205
  (
    n216,
    n57
  );


  not
  g206
  (
    n280,
    n69
  );


  buf
  g207
  (
    n149,
    n41
  );


  buf
  g208
  (
    n263,
    n52
  );


  not
  g209
  (
    n218,
    n44
  );


  not
  g210
  (
    n200,
    n58
  );


  buf
  g211
  (
    n107,
    n60
  );


  buf
  g212
  (
    n169,
    n56
  );


  buf
  g213
  (
    n198,
    n43
  );


  buf
  g214
  (
    n116,
    n77
  );


  not
  g215
  (
    n186,
    n33
  );


  not
  g216
  (
    n258,
    n57
  );


  not
  g217
  (
    n114,
    n44
  );


  buf
  g218
  (
    n229,
    n68
  );


  not
  g219
  (
    n240,
    n40
  );


  not
  g220
  (
    n224,
    n39
  );


  not
  g221
  (
    n135,
    n50
  );


  buf
  g222
  (
    n153,
    n40
  );


  not
  g223
  (
    n106,
    n72
  );


  not
  g224
  (
    n262,
    n40
  );


  not
  g225
  (
    n171,
    n56
  );


  buf
  g226
  (
    n232,
    n53
  );


  buf
  g227
  (
    n159,
    n59
  );


  buf
  g228
  (
    n277,
    n35
  );


  buf
  g229
  (
    n188,
    n72
  );


  buf
  g230
  (
    n254,
    n44
  );


  buf
  g231
  (
    n158,
    n75
  );


  not
  g232
  (
    n131,
    n66
  );


  not
  g233
  (
    n195,
    n65
  );


  buf
  g234
  (
    n168,
    n60
  );


  buf
  g235
  (
    n125,
    n40
  );


  not
  g236
  (
    n99,
    n51
  );


  buf
  g237
  (
    n210,
    n55
  );


  not
  g238
  (
    n165,
    n49
  );


  buf
  g239
  (
    n197,
    n62
  );


  not
  g240
  (
    n222,
    n55
  );


  not
  g241
  (
    n256,
    n49
  );


  buf
  g242
  (
    n161,
    n53
  );


  not
  g243
  (
    n160,
    n56
  );


  not
  g244
  (
    n157,
    n61
  );


  buf
  g245
  (
    n154,
    n67
  );


  not
  g246
  (
    n219,
    n61
  );


  not
  g247
  (
    n132,
    n67
  );


  not
  g248
  (
    n257,
    n49
  );


  not
  g249
  (
    n851,
    n164
  );


  not
  g250
  (
    n798,
    n107
  );


  not
  g251
  (
    n536,
    n204
  );


  not
  g252
  (
    n677,
    n142
  );


  buf
  g253
  (
    n881,
    n137
  );


  buf
  g254
  (
    n746,
    n101
  );


  buf
  g255
  (
    n491,
    n184
  );


  not
  g256
  (
    n443,
    n200
  );


  buf
  g257
  (
    n825,
    n223
  );


  not
  g258
  (
    n291,
    n126
  );


  buf
  g259
  (
    n815,
    n207
  );


  not
  g260
  (
    n880,
    n208
  );


  not
  g261
  (
    n644,
    n178
  );


  buf
  g262
  (
    n841,
    n173
  );


  buf
  g263
  (
    n460,
    n237
  );


  not
  g264
  (
    n831,
    n119
  );


  not
  g265
  (
    n296,
    n162
  );


  buf
  g266
  (
    n767,
    n238
  );


  not
  g267
  (
    n415,
    n207
  );


  buf
  g268
  (
    n540,
    n170
  );


  buf
  g269
  (
    n305,
    n203
  );


  not
  g270
  (
    n956,
    n255
  );


  not
  g271
  (
    n959,
    n120
  );


  buf
  g272
  (
    n449,
    n148
  );


  buf
  g273
  (
    n522,
    n138
  );


  buf
  g274
  (
    n393,
    n174
  );


  not
  g275
  (
    n555,
    n179
  );


  buf
  g276
  (
    n696,
    n145
  );


  not
  g277
  (
    n930,
    n214
  );


  not
  g278
  (
    n572,
    n105
  );


  not
  g279
  (
    n423,
    n130
  );


  buf
  g280
  (
    n576,
    n248
  );


  not
  g281
  (
    n725,
    n187
  );


  not
  g282
  (
    n863,
    n175
  );


  buf
  g283
  (
    n949,
    n240
  );


  not
  g284
  (
    n721,
    n239
  );


  buf
  g285
  (
    n727,
    n216
  );


  buf
  g286
  (
    n285,
    n138
  );


  not
  g287
  (
    n699,
    n100
  );


  not
  g288
  (
    n665,
    n176
  );


  not
  g289
  (
    n331,
    n218
  );


  buf
  g290
  (
    n704,
    n131
  );


  not
  g291
  (
    n861,
    n227
  );


  not
  g292
  (
    n361,
    n181
  );


  not
  g293
  (
    n712,
    n255
  );


  buf
  g294
  (
    n913,
    n231
  );


  buf
  g295
  (
    n312,
    n177
  );


  buf
  g296
  (
    n821,
    n249
  );


  buf
  g297
  (
    n806,
    n106
  );


  not
  g298
  (
    n934,
    n197
  );


  buf
  g299
  (
    n364,
    n232
  );


  buf
  g300
  (
    n655,
    n263
  );


  not
  g301
  (
    n669,
    n110
  );


  buf
  g302
  (
    n664,
    n102
  );


  buf
  g303
  (
    n474,
    n250
  );


  buf
  g304
  (
    n805,
    n123
  );


  not
  g305
  (
    n390,
    n135
  );


  buf
  g306
  (
    n611,
    n165
  );


  not
  g307
  (
    n420,
    n260
  );


  not
  g308
  (
    n589,
    n163
  );


  not
  g309
  (
    n952,
    n135
  );


  buf
  g310
  (
    n330,
    n163
  );


  buf
  g311
  (
    n634,
    n253
  );


  buf
  g312
  (
    n919,
    n158
  );


  buf
  g313
  (
    n747,
    n216
  );


  not
  g314
  (
    n594,
    n243
  );


  not
  g315
  (
    n631,
    n154
  );


  buf
  g316
  (
    n528,
    n106
  );


  not
  g317
  (
    n609,
    n137
  );


  not
  g318
  (
    n450,
    n186
  );


  not
  g319
  (
    n297,
    n219
  );


  not
  g320
  (
    n355,
    n250
  );


  buf
  g321
  (
    n288,
    n225
  );


  buf
  g322
  (
    n958,
    n165
  );


  buf
  g323
  (
    n516,
    n175
  );


  buf
  g324
  (
    n541,
    n102
  );


  buf
  g325
  (
    n463,
    n185
  );


  buf
  g326
  (
    n652,
    n118
  );


  not
  g327
  (
    n781,
    n264
  );


  buf
  g328
  (
    n858,
    n178
  );


  buf
  g329
  (
    n695,
    n166
  );


  buf
  g330
  (
    n636,
    n160
  );


  not
  g331
  (
    n846,
    n256
  );


  buf
  g332
  (
    n398,
    n242
  );


  buf
  g333
  (
    n283,
    n238
  );


  buf
  g334
  (
    n549,
    n235
  );


  buf
  g335
  (
    n809,
    n252
  );


  not
  g336
  (
    n627,
    n151
  );


  buf
  g337
  (
    n584,
    n263
  );


  buf
  g338
  (
    n345,
    n152
  );


  not
  g339
  (
    n910,
    n203
  );


  buf
  g340
  (
    n748,
    n133
  );


  not
  g341
  (
    n726,
    n196
  );


  not
  g342
  (
    n843,
    n124
  );


  not
  g343
  (
    n466,
    n167
  );


  not
  g344
  (
    n356,
    n150
  );


  not
  g345
  (
    n803,
    n148
  );


  not
  g346
  (
    n388,
    n121
  );


  buf
  g347
  (
    n744,
    n260
  );


  not
  g348
  (
    n922,
    n142
  );


  not
  g349
  (
    n828,
    n233
  );


  buf
  g350
  (
    n383,
    n221
  );


  buf
  g351
  (
    n945,
    n150
  );


  buf
  g352
  (
    n392,
    n173
  );


  buf
  g353
  (
    n898,
    n144
  );


  not
  g354
  (
    n893,
    n142
  );


  not
  g355
  (
    n412,
    n144
  );


  not
  g356
  (
    n947,
    n250
  );


  not
  g357
  (
    n710,
    n210
  );


  not
  g358
  (
    n943,
    n253
  );


  not
  g359
  (
    n944,
    n207
  );


  not
  g360
  (
    n292,
    n209
  );


  not
  g361
  (
    n562,
    n99
  );


  not
  g362
  (
    n658,
    n146
  );


  not
  g363
  (
    n765,
    n262
  );


  buf
  g364
  (
    n926,
    n145
  );


  not
  g365
  (
    n857,
    n132
  );


  buf
  g366
  (
    n351,
    n199
  );


  not
  g367
  (
    n845,
    n254
  );


  not
  g368
  (
    n328,
    n241
  );


  not
  g369
  (
    n534,
    n147
  );


  not
  g370
  (
    n564,
    n146
  );


  buf
  g371
  (
    n946,
    n194
  );


  buf
  g372
  (
    n810,
    n101
  );


  not
  g373
  (
    n539,
    n130
  );


  not
  g374
  (
    n569,
    n120
  );


  buf
  g375
  (
    n357,
    n179
  );


  not
  g376
  (
    n754,
    n175
  );


  buf
  g377
  (
    n801,
    n253
  );


  not
  g378
  (
    n384,
    n251
  );


  buf
  g379
  (
    n618,
    n140
  );


  not
  g380
  (
    n724,
    n208
  );


  not
  g381
  (
    n509,
    n164
  );


  buf
  g382
  (
    n406,
    n243
  );


  buf
  g383
  (
    n366,
    n247
  );


  buf
  g384
  (
    n577,
    n161
  );


  not
  g385
  (
    n855,
    n259
  );


  buf
  g386
  (
    n619,
    n166
  );


  buf
  g387
  (
    n788,
    n190
  );


  not
  g388
  (
    n447,
    n139
  );


  not
  g389
  (
    n394,
    n187
  );


  not
  g390
  (
    n313,
    n157
  );


  buf
  g391
  (
    n344,
    n128
  );


  buf
  g392
  (
    n306,
    n115
  );


  not
  g393
  (
    n827,
    n99
  );


  not
  g394
  (
    n349,
    n170
  );


  not
  g395
  (
    n775,
    n100
  );


  buf
  g396
  (
    n853,
    n202
  );


  buf
  g397
  (
    n340,
    n135
  );


  buf
  g398
  (
    n322,
    n125
  );


  not
  g399
  (
    n593,
    n152
  );


  not
  g400
  (
    n896,
    n213
  );


  not
  g401
  (
    n751,
    n161
  );


  not
  g402
  (
    n914,
    n231
  );


  buf
  g403
  (
    n650,
    n174
  );


  buf
  g404
  (
    n335,
    n182
  );


  buf
  g405
  (
    n923,
    n113
  );


  not
  g406
  (
    n703,
    n265
  );


  buf
  g407
  (
    n583,
    n226
  );


  buf
  g408
  (
    n647,
    n232
  );


  not
  g409
  (
    n396,
    n177
  );


  not
  g410
  (
    n755,
    n226
  );


  not
  g411
  (
    n282,
    n217
  );


  not
  g412
  (
    n284,
    n116
  );


  not
  g413
  (
    n342,
    n259
  );


  buf
  g414
  (
    n370,
    n190
  );


  not
  g415
  (
    n502,
    n176
  );


  not
  g416
  (
    n659,
    n201
  );


  buf
  g417
  (
    n505,
    n248
  );


  buf
  g418
  (
    n918,
    n214
  );


  not
  g419
  (
    n615,
    n200
  );


  buf
  g420
  (
    n854,
    n252
  );


  buf
  g421
  (
    n741,
    n262
  );


  buf
  g422
  (
    n503,
    n199
  );


  not
  g423
  (
    n738,
    n121
  );


  not
  g424
  (
    n362,
    n105
  );


  buf
  g425
  (
    n425,
    n256
  );


  not
  g426
  (
    n911,
    n212
  );


  buf
  g427
  (
    n929,
    n227
  );


  not
  g428
  (
    n433,
    n223
  );


  not
  g429
  (
    n544,
    n228
  );


  buf
  g430
  (
    n360,
    n217
  );


  not
  g431
  (
    n909,
    n163
  );


  not
  g432
  (
    n777,
    n102
  );


  buf
  g433
  (
    n641,
    n149
  );


  not
  g434
  (
    n599,
    n157
  );


  not
  g435
  (
    n849,
    n137
  );


  not
  g436
  (
    n739,
    n248
  );


  buf
  g437
  (
    n906,
    n242
  );


  not
  g438
  (
    n728,
    n188
  );


  buf
  g439
  (
    n617,
    n103
  );


  not
  g440
  (
    n596,
    n205
  );


  buf
  g441
  (
    n445,
    n107
  );


  buf
  g442
  (
    n733,
    n194
  );


  buf
  g443
  (
    n882,
    n118
  );


  not
  g444
  (
    n640,
    n249
  );


  not
  g445
  (
    n796,
    n246
  );


  buf
  g446
  (
    n490,
    n249
  );


  buf
  g447
  (
    n471,
    n123
  );


  not
  g448
  (
    n878,
    n216
  );


  not
  g449
  (
    n797,
    n157
  );


  not
  g450
  (
    n686,
    n108
  );


  not
  g451
  (
    n737,
    n149
  );


  buf
  g452
  (
    n614,
    n197
  );


  not
  g453
  (
    n424,
    n214
  );


  not
  g454
  (
    n916,
    n225
  );


  not
  g455
  (
    n713,
    n126
  );


  not
  g456
  (
    n921,
    n206
  );


  not
  g457
  (
    n558,
    n104
  );


  buf
  g458
  (
    n729,
    n265
  );


  not
  g459
  (
    n604,
    n127
  );


  buf
  g460
  (
    n864,
    n244
  );


  not
  g461
  (
    n711,
    n168
  );


  buf
  g462
  (
    n592,
    n206
  );


  buf
  g463
  (
    n512,
    n178
  );


  buf
  g464
  (
    n761,
    n105
  );


  not
  g465
  (
    n568,
    n111
  );


  not
  g466
  (
    n338,
    n169
  );


  buf
  g467
  (
    n648,
    n200
  );


  not
  g468
  (
    n465,
    n147
  );


  buf
  g469
  (
    n308,
    n126
  );


  not
  g470
  (
    n417,
    n264
  );


  buf
  g471
  (
    n680,
    n136
  );


  not
  g472
  (
    n481,
    n248
  );


  not
  g473
  (
    n295,
    n144
  );


  buf
  g474
  (
    n377,
    n172
  );


  not
  g475
  (
    n674,
    n140
  );


  buf
  g476
  (
    n920,
    n268
  );


  not
  g477
  (
    n372,
    n211
  );


  buf
  g478
  (
    n877,
    n158
  );


  not
  g479
  (
    n553,
    n178
  );


  buf
  g480
  (
    n839,
    n244
  );


  not
  g481
  (
    n936,
    n132
  );


  not
  g482
  (
    n753,
    n205
  );


  not
  g483
  (
    n286,
    n117
  );


  not
  g484
  (
    n673,
    n158
  );


  buf
  g485
  (
    n879,
    n167
  );


  not
  g486
  (
    n298,
    n268
  );


  buf
  g487
  (
    n687,
    n241
  );


  not
  g488
  (
    n832,
    n115
  );


  buf
  g489
  (
    n942,
    n128
  );


  not
  g490
  (
    n698,
    n159
  );


  buf
  g491
  (
    n875,
    n144
  );


  not
  g492
  (
    n459,
    n226
  );


  buf
  g493
  (
    n679,
    n108
  );


  buf
  g494
  (
    n381,
    n268
  );


  not
  g495
  (
    n787,
    n245
  );


  buf
  g496
  (
    n758,
    n217
  );


  buf
  g497
  (
    n626,
    n215
  );


  not
  g498
  (
    n535,
    n259
  );


  not
  g499
  (
    n409,
    n242
  );


  buf
  g500
  (
    n657,
    n258
  );


  buf
  g501
  (
    n666,
    n233
  );


  buf
  g502
  (
    n578,
    n191
  );


  buf
  g503
  (
    n817,
    n133
  );


  buf
  g504
  (
    n427,
    n142
  );


  buf
  g505
  (
    n354,
    n154
  );


  buf
  g506
  (
    n760,
    n103
  );


  buf
  g507
  (
    n551,
    n235
  );


  buf
  g508
  (
    n435,
    n247
  );


  not
  g509
  (
    n925,
    n136
  );


  buf
  g510
  (
    n519,
    n174
  );


  not
  g511
  (
    n421,
    n146
  );


  buf
  g512
  (
    n337,
    n180
  );


  not
  g513
  (
    n570,
    n172
  );


  not
  g514
  (
    n763,
    n205
  );


  buf
  g515
  (
    n780,
    n173
  );


  not
  g516
  (
    n649,
    n130
  );


  not
  g517
  (
    n363,
    n215
  );


  not
  g518
  (
    n499,
    n154
  );


  buf
  g519
  (
    n823,
    n184
  );


  not
  g520
  (
    n902,
    n217
  );


  not
  g521
  (
    n319,
    n112
  );


  not
  g522
  (
    n542,
    n202
  );


  not
  g523
  (
    n772,
    n160
  );


  buf
  g524
  (
    n957,
    n129
  );


  buf
  g525
  (
    n579,
    n229
  );


  buf
  g526
  (
    n822,
    n168
  );


  buf
  g527
  (
    n932,
    n247
  );


  not
  g528
  (
    n660,
    n193
  );


  buf
  g529
  (
    n489,
    n106
  );


  not
  g530
  (
    n903,
    n102
  );


  buf
  g531
  (
    n715,
    n236
  );


  buf
  g532
  (
    n327,
    n254
  );


  not
  g533
  (
    n667,
    n181
  );


  buf
  g534
  (
    n613,
    n183
  );


  buf
  g535
  (
    n847,
    n103
  );


  not
  g536
  (
    n299,
    n147
  );


  buf
  g537
  (
    n938,
    n261
  );


  buf
  g538
  (
    n560,
    n235
  );


  not
  g539
  (
    n386,
    n183
  );


  buf
  g540
  (
    n812,
    n169
  );


  buf
  g541
  (
    n718,
    n186
  );


  not
  g542
  (
    n336,
    n182
  );


  buf
  g543
  (
    n480,
    n114
  );


  buf
  g544
  (
    n301,
    n175
  );


  not
  g545
  (
    n819,
    n212
  );


  buf
  g546
  (
    n820,
    n195
  );


  buf
  g547
  (
    n454,
    n198
  );


  buf
  g548
  (
    n643,
    n241
  );


  buf
  g549
  (
    n402,
    n107
  );


  buf
  g550
  (
    n961,
    n215
  );


  buf
  g551
  (
    n411,
    n156
  );


  not
  g552
  (
    n483,
    n187
  );


  buf
  g553
  (
    n353,
    n141
  );


  not
  g554
  (
    n482,
    n143
  );


  buf
  g555
  (
    n374,
    n189
  );


  buf
  g556
  (
    n321,
    n187
  );


  not
  g557
  (
    n689,
    n148
  );


  not
  g558
  (
    n743,
    n171
  );


  buf
  g559
  (
    n380,
    n199
  );


  not
  g560
  (
    n639,
    n199
  );


  buf
  g561
  (
    n397,
    n149
  );


  not
  g562
  (
    n468,
    n239
  );


  buf
  g563
  (
    n529,
    n192
  );


  not
  g564
  (
    n448,
    n197
  );


  buf
  g565
  (
    n808,
    n208
  );


  not
  g566
  (
    n456,
    n229
  );


  buf
  g567
  (
    n838,
    n134
  );


  not
  g568
  (
    n317,
    n254
  );


  not
  g569
  (
    n559,
    n143
  );


  buf
  g570
  (
    n789,
    n218
  );


  not
  g571
  (
    n430,
    n161
  );


  not
  g572
  (
    n418,
    n246
  );


  not
  g573
  (
    n874,
    n214
  );


  not
  g574
  (
    n759,
    n132
  );


  buf
  g575
  (
    n314,
    n140
  );


  buf
  g576
  (
    n813,
    n128
  );


  buf
  g577
  (
    n811,
    n127
  );


  not
  g578
  (
    n757,
    n237
  );


  buf
  g579
  (
    n690,
    n234
  );


  buf
  g580
  (
    n414,
    n211
  );


  buf
  g581
  (
    n464,
    n166
  );


  not
  g582
  (
    n734,
    n250
  );


  buf
  g583
  (
    n642,
    n151
  );


  buf
  g584
  (
    n469,
    n227
  );


  not
  g585
  (
    n325,
    n222
  );


  buf
  g586
  (
    n706,
    n236
  );


  buf
  g587
  (
    n586,
    n252
  );


  buf
  g588
  (
    n300,
    n111
  );


  not
  g589
  (
    n403,
    n182
  );


  buf
  g590
  (
    n735,
    n246
  );


  not
  g591
  (
    n511,
    n186
  );


  not
  g592
  (
    n622,
    n244
  );


  not
  g593
  (
    n740,
    n202
  );


  not
  g594
  (
    n520,
    n136
  );


  buf
  g595
  (
    n745,
    n258
  );


  buf
  g596
  (
    n441,
    n129
  );


  not
  g597
  (
    n561,
    n239
  );


  not
  g598
  (
    n782,
    n123
  );


  not
  g599
  (
    n645,
    n117
  );


  not
  g600
  (
    n473,
    n172
  );


  buf
  g601
  (
    n897,
    n267
  );


  buf
  g602
  (
    n694,
    n205
  );


  buf
  g603
  (
    n341,
    n222
  );


  buf
  g604
  (
    n701,
    n218
  );


  buf
  g605
  (
    n506,
    n161
  );


  not
  g606
  (
    n510,
    n213
  );


  buf
  g607
  (
    n707,
    n193
  );


  not
  g608
  (
    n543,
    n186
  );


  buf
  g609
  (
    n307,
    n195
  );


  buf
  g610
  (
    n426,
    n172
  );


  not
  g611
  (
    n367,
    n154
  );


  not
  g612
  (
    n554,
    n204
  );


  not
  g613
  (
    n462,
    n231
  );


  buf
  g614
  (
    n868,
    n156
  );


  not
  g615
  (
    n401,
    n109
  );


  not
  g616
  (
    n799,
    n174
  );


  buf
  g617
  (
    n479,
    n198
  );


  buf
  g618
  (
    n610,
    n245
  );


  buf
  g619
  (
    n895,
    n254
  );


  buf
  g620
  (
    n369,
    n155
  );


  not
  g621
  (
    n742,
    n147
  );


  not
  g622
  (
    n530,
    n165
  );


  not
  g623
  (
    n478,
    n156
  );


  buf
  g624
  (
    n873,
    n107
  );


  buf
  g625
  (
    n883,
    n150
  );


  buf
  g626
  (
    n311,
    n251
  );


  buf
  g627
  (
    n507,
    n188
  );


  buf
  g628
  (
    n616,
    n169
  );


  not
  g629
  (
    n612,
    n234
  );


  not
  g630
  (
    n867,
    n141
  );


  buf
  g631
  (
    n457,
    n213
  );


  not
  g632
  (
    n783,
    n134
  );


  buf
  g633
  (
    n395,
    n256
  );


  not
  g634
  (
    n623,
    n166
  );


  not
  g635
  (
    n842,
    n219
  );


  buf
  g636
  (
    n684,
    n188
  );


  buf
  g637
  (
    n598,
    n244
  );


  buf
  g638
  (
    n807,
    n110
  );


  buf
  g639
  (
    n571,
    n264
  );


  not
  g640
  (
    n485,
    n140
  );


  buf
  g641
  (
    n630,
    n245
  );


  not
  g642
  (
    n440,
    n201
  );


  not
  g643
  (
    n635,
    n221
  );


  buf
  g644
  (
    n702,
    n104
  );


  not
  g645
  (
    n859,
    n208
  );


  not
  g646
  (
    n316,
    n153
  );


  not
  g647
  (
    n872,
    n218
  );


  buf
  g648
  (
    n527,
    n141
  );


  not
  g649
  (
    n494,
    n101
  );


  not
  g650
  (
    n590,
    n139
  );


  buf
  g651
  (
    n442,
    n111
  );


  buf
  g652
  (
    n359,
    n192
  );


  not
  g653
  (
    n347,
    n230
  );


  not
  g654
  (
    n829,
    n157
  );


  not
  g655
  (
    n912,
    n249
  );


  not
  g656
  (
    n683,
    n266
  );


  buf
  g657
  (
    n682,
    n176
  );


  buf
  g658
  (
    n416,
    n143
  );


  not
  g659
  (
    n840,
    n151
  );


  not
  g660
  (
    n455,
    n130
  );


  not
  g661
  (
    n472,
    n225
  );


  not
  g662
  (
    n470,
    n189
  );


  not
  g663
  (
    n632,
    n203
  );


  not
  g664
  (
    n352,
    n257
  );


  buf
  g665
  (
    n885,
    n204
  );


  not
  g666
  (
    n939,
    n238
  );


  buf
  g667
  (
    n672,
    n266
  );


  not
  g668
  (
    n904,
    n189
  );


  not
  g669
  (
    n884,
    n104
  );


  not
  g670
  (
    n488,
    n209
  );


  buf
  g671
  (
    n582,
    n128
  );


  buf
  g672
  (
    n324,
    n201
  );


  buf
  g673
  (
    n575,
    n264
  );


  not
  g674
  (
    n818,
    n183
  );


  buf
  g675
  (
    n770,
    n112
  );


  buf
  g676
  (
    n326,
    n159
  );


  not
  g677
  (
    n792,
    n265
  );


  not
  g678
  (
    n567,
    n262
  );


  not
  g679
  (
    n786,
    n223
  );


  buf
  g680
  (
    n638,
    n184
  );


  not
  g681
  (
    n907,
    n100
  );


  buf
  g682
  (
    n670,
    n190
  );


  not
  g683
  (
    n302,
    n192
  );


  not
  g684
  (
    n439,
    n230
  );


  buf
  g685
  (
    n931,
    n118
  );


  buf
  g686
  (
    n685,
    n253
  );


  not
  g687
  (
    n368,
    n153
  );


  not
  g688
  (
    n581,
    n194
  );


  buf
  g689
  (
    n793,
    n197
  );


  buf
  g690
  (
    n869,
    n262
  );


  not
  g691
  (
    n515,
    n220
  );


  buf
  g692
  (
    n557,
    n221
  );


  not
  g693
  (
    n804,
    n160
  );


  buf
  g694
  (
    n941,
    n139
  );


  buf
  g695
  (
    n764,
    n260
  );


  not
  g696
  (
    n940,
    n222
  );


  buf
  g697
  (
    n310,
    n133
  );


  not
  g698
  (
    n496,
    n256
  );


  buf
  g699
  (
    n816,
    n258
  );


  not
  g700
  (
    n476,
    n233
  );


  buf
  g701
  (
    n732,
    n185
  );


  buf
  g702
  (
    n436,
    n206
  );


  buf
  g703
  (
    n661,
    n149
  );


  not
  g704
  (
    n376,
    n124
  );


  buf
  g705
  (
    n607,
    n236
  );


  buf
  g706
  (
    n837,
    n101
  );


  not
  g707
  (
    n891,
    n226
  );


  buf
  g708
  (
    n834,
    n242
  );


  buf
  g709
  (
    n960,
    n203
  );


  buf
  g710
  (
    n814,
    n234
  );


  not
  g711
  (
    n538,
    n160
  );


  buf
  g712
  (
    n752,
    n171
  );


  not
  g713
  (
    n563,
    n237
  );


  buf
  g714
  (
    n924,
    n243
  );


  not
  g715
  (
    n784,
    n230
  );


  not
  g716
  (
    n526,
    n131
  );


  not
  g717
  (
    n651,
    n195
  );


  buf
  g718
  (
    n730,
    n169
  );


  buf
  g719
  (
    n768,
    n117
  );


  not
  g720
  (
    n603,
    n252
  );


  not
  g721
  (
    n444,
    n105
  );


  buf
  g722
  (
    n332,
    n191
  );


  buf
  g723
  (
    n315,
    n127
  );


  buf
  g724
  (
    n866,
    n119
  );


  not
  g725
  (
    n320,
    n236
  );


  buf
  g726
  (
    n550,
    n180
  );


  buf
  g727
  (
    n573,
    n261
  );


  buf
  g728
  (
    n547,
    n162
  );


  buf
  g729
  (
    n856,
    n228
  );


  not
  g730
  (
    n766,
    n193
  );


  not
  g731
  (
    n446,
    n230
  );


  not
  g732
  (
    n387,
    n200
  );


  not
  g733
  (
    n654,
    n131
  );


  not
  g734
  (
    n408,
    n145
  );


  buf
  g735
  (
    n844,
    n198
  );


  not
  g736
  (
    n717,
    n167
  );


  buf
  g737
  (
    n373,
    n126
  );


  buf
  g738
  (
    n574,
    n221
  );


  buf
  g739
  (
    n750,
    n224
  );


  not
  g740
  (
    n776,
    n152
  );


  not
  g741
  (
    n705,
    n122
  );


  not
  g742
  (
    n605,
    n210
  );


  buf
  g743
  (
    n375,
    n116
  );


  buf
  g744
  (
    n871,
    n246
  );


  not
  g745
  (
    n899,
    n158
  );


  buf
  g746
  (
    n693,
    n257
  );


  buf
  g747
  (
    n517,
    n251
  );


  buf
  g748
  (
    n365,
    n191
  );


  buf
  g749
  (
    n431,
    n258
  );


  buf
  g750
  (
    n467,
    n193
  );


  not
  g751
  (
    n865,
    n133
  );


  buf
  g752
  (
    n722,
    n117
  );


  not
  g753
  (
    n429,
    n150
  );


  buf
  g754
  (
    n399,
    n159
  );


  buf
  g755
  (
    n692,
    n148
  );


  not
  g756
  (
    n495,
    n211
  );


  not
  g757
  (
    n438,
    n247
  );


  buf
  g758
  (
    n954,
    n109
  );


  buf
  g759
  (
    n587,
    n112
  );


  buf
  g760
  (
    n769,
    n119
  );


  buf
  g761
  (
    n346,
    n240
  );


  buf
  g762
  (
    n836,
    n177
  );


  buf
  g763
  (
    n452,
    n224
  );


  buf
  g764
  (
    n537,
    n121
  );


  buf
  g765
  (
    n802,
    n104
  );


  buf
  g766
  (
    n791,
    n103
  );


  buf
  g767
  (
    n477,
    n257
  );


  not
  g768
  (
    n566,
    n155
  );


  buf
  g769
  (
    n458,
    n196
  );


  buf
  g770
  (
    n546,
    n198
  );


  not
  g771
  (
    n716,
    n227
  );


  buf
  g772
  (
    n329,
    n204
  );


  buf
  g773
  (
    n422,
    n216
  );


  not
  g774
  (
    n620,
    n220
  );


  buf
  g775
  (
    n790,
    n261
  );


  not
  g776
  (
    n628,
    n116
  );


  not
  g777
  (
    n862,
    n196
  );


  buf
  g778
  (
    n714,
    n191
  );


  buf
  g779
  (
    n876,
    n113
  );


  not
  g780
  (
    n900,
    n263
  );


  not
  g781
  (
    n432,
    n241
  );


  buf
  g782
  (
    n545,
    n164
  );


  not
  g783
  (
    n889,
    n145
  );


  not
  g784
  (
    n595,
    n125
  );


  buf
  g785
  (
    n531,
    n225
  );


  not
  g786
  (
    n892,
    n163
  );


  buf
  g787
  (
    n826,
    n109
  );


  not
  g788
  (
    n294,
    n219
  );


  buf
  g789
  (
    n585,
    n210
  );


  buf
  g790
  (
    n629,
    n106
  );


  not
  g791
  (
    n933,
    n189
  );


  not
  g792
  (
    n548,
    n115
  );


  not
  g793
  (
    n498,
    n156
  );


  not
  g794
  (
    n400,
    n112
  );


  buf
  g795
  (
    n835,
    n220
  );


  not
  g796
  (
    n608,
    n170
  );


  not
  g797
  (
    n289,
    n215
  );


  buf
  g798
  (
    n407,
    n267
  );


  not
  g799
  (
    n688,
    n232
  );


  not
  g800
  (
    n475,
    n229
  );


  not
  g801
  (
    n624,
    n125
  );


  not
  g802
  (
    n580,
    n129
  );


  not
  g803
  (
    n334,
    n164
  );


  not
  g804
  (
    n637,
    n232
  );


  buf
  g805
  (
    n795,
    n108
  );


  buf
  g806
  (
    n908,
    n211
  );


  buf
  g807
  (
    n556,
    n136
  );


  buf
  g808
  (
    n833,
    n195
  );


  buf
  g809
  (
    n600,
    n132
  );


  not
  g810
  (
    n830,
    n155
  );


  buf
  g811
  (
    n656,
    n113
  );


  not
  g812
  (
    n762,
    n179
  );


  buf
  g813
  (
    n385,
    n182
  );


  not
  g814
  (
    n453,
    n100
  );


  buf
  g815
  (
    n410,
    n229
  );


  not
  g816
  (
    n736,
    n176
  );


  not
  g817
  (
    n333,
    n114
  );


  not
  g818
  (
    n662,
    n228
  );


  not
  g819
  (
    n779,
    n259
  );


  not
  g820
  (
    n513,
    n124
  );


  buf
  g821
  (
    n287,
    n235
  );


  buf
  g822
  (
    n532,
    n180
  );


  not
  g823
  (
    n708,
    n238
  );


  not
  g824
  (
    n824,
    n194
  );


  not
  g825
  (
    n887,
    n138
  );


  not
  g826
  (
    n497,
    n231
  );


  not
  g827
  (
    n437,
    n240
  );


  not
  g828
  (
    n675,
    n113
  );


  buf
  g829
  (
    n773,
    n121
  );


  not
  g830
  (
    n565,
    n224
  );


  not
  g831
  (
    n723,
    n129
  );


  buf
  g832
  (
    n493,
    n152
  );


  not
  g833
  (
    n697,
    n228
  );


  not
  g834
  (
    n886,
    n170
  );


  not
  g835
  (
    n653,
    n131
  );


  not
  g836
  (
    n428,
    n181
  );


  buf
  g837
  (
    n621,
    n179
  );


  not
  g838
  (
    n800,
    n138
  );


  not
  g839
  (
    n434,
    n224
  );


  not
  g840
  (
    n348,
    n108
  );


  buf
  g841
  (
    n293,
    n266
  );


  not
  g842
  (
    n749,
    n141
  );


  buf
  g843
  (
    n518,
    n135
  );


  not
  g844
  (
    n358,
    n168
  );


  buf
  g845
  (
    n785,
    n257
  );


  not
  g846
  (
    n860,
    n122
  );


  buf
  g847
  (
    n552,
    n114
  );


  not
  g848
  (
    n484,
    n122
  );


  buf
  g849
  (
    n591,
    n151
  );


  buf
  g850
  (
    n486,
    n209
  );


  not
  g851
  (
    n413,
    n155
  );


  not
  g852
  (
    n720,
    n109
  );


  not
  g853
  (
    n508,
    n124
  );


  buf
  g854
  (
    n523,
    n118
  );


  not
  g855
  (
    n848,
    n99
  );


  buf
  g856
  (
    n774,
    n219
  );


  buf
  g857
  (
    n597,
    n223
  );


  buf
  g858
  (
    n378,
    n139
  );


  buf
  g859
  (
    n382,
    n237
  );


  buf
  g860
  (
    n905,
    n99
  );


  buf
  g861
  (
    n935,
    n266
  );


  not
  g862
  (
    n888,
    n213
  );


  not
  g863
  (
    n678,
    n180
  );


  not
  g864
  (
    n951,
    n212
  );


  buf
  g865
  (
    n700,
    n267
  );


  buf
  g866
  (
    n343,
    n120
  );


  buf
  g867
  (
    n461,
    n122
  );


  buf
  g868
  (
    n756,
    n255
  );


  not
  g869
  (
    n487,
    n159
  );


  buf
  g870
  (
    n709,
    n162
  );


  not
  g871
  (
    n524,
    n134
  );


  buf
  g872
  (
    n691,
    n206
  );


  not
  g873
  (
    n318,
    n123
  );


  not
  g874
  (
    n719,
    n167
  );


  buf
  g875
  (
    n339,
    n201
  );


  buf
  g876
  (
    n602,
    n125
  );


  not
  g877
  (
    n500,
    n261
  );


  buf
  g878
  (
    n501,
    n267
  );


  buf
  g879
  (
    n633,
    n268
  );


  buf
  g880
  (
    n955,
    n165
  );


  not
  g881
  (
    n304,
    n234
  );


  buf
  g882
  (
    n405,
    n134
  );


  buf
  g883
  (
    n950,
    n220
  );


  buf
  g884
  (
    n915,
    n177
  );


  buf
  g885
  (
    n371,
    n190
  );


  buf
  g886
  (
    n379,
    n185
  );


  not
  g887
  (
    n668,
    n260
  );


  not
  g888
  (
    n525,
    n114
  );


  buf
  g889
  (
    n601,
    n240
  );


  buf
  g890
  (
    n533,
    n153
  );


  not
  g891
  (
    n350,
    n110
  );


  buf
  g892
  (
    n937,
    n239
  );


  buf
  g893
  (
    n917,
    n162
  );


  buf
  g894
  (
    n389,
    n181
  );


  not
  g895
  (
    n521,
    n127
  );


  not
  g896
  (
    n492,
    n184
  );


  not
  g897
  (
    n778,
    n222
  );


  not
  g898
  (
    n681,
    n110
  );


  not
  g899
  (
    n504,
    n183
  );


  buf
  g900
  (
    n391,
    n196
  );


  not
  g901
  (
    n309,
    n146
  );


  not
  g902
  (
    n928,
    n116
  );


  buf
  g903
  (
    n303,
    n171
  );


  not
  g904
  (
    n870,
    n137
  );


  not
  g905
  (
    n514,
    n120
  );


  buf
  g906
  (
    n290,
    n251
  );


  not
  g907
  (
    n588,
    n115
  );


  not
  g908
  (
    n890,
    n255
  );


  buf
  g909
  (
    n850,
    n168
  );


  not
  g910
  (
    n323,
    n111
  );


  not
  g911
  (
    n771,
    n265
  );


  buf
  g912
  (
    n663,
    n207
  );


  buf
  g913
  (
    n927,
    n119
  );


  buf
  g914
  (
    n451,
    n210
  );


  not
  g915
  (
    n953,
    n192
  );


  not
  g916
  (
    n901,
    n263
  );


  not
  g917
  (
    n404,
    n245
  );


  buf
  g918
  (
    n794,
    n212
  );


  not
  g919
  (
    n852,
    n153
  );


  buf
  g920
  (
    n894,
    n143
  );


  buf
  g921
  (
    n625,
    n185
  );


  buf
  g922
  (
    n948,
    n171
  );


  buf
  g923
  (
    n671,
    n243
  );


  not
  g924
  (
    n606,
    n233
  );


  not
  g925
  (
    n676,
    n188
  );


  not
  g926
  (
    n646,
    n202
  );


  not
  g927
  (
    n419,
    n209
  );


  not
  g928
  (
    n731,
    n173
  );


  xnor
  g929
  (
    n1052,
    n791,
    n793,
    n792,
    n432
  );


  xnor
  g930
  (
    n1241,
    n331,
    n828,
    n461,
    n579
  );


  xor
  g931
  (
    n975,
    n901,
    n397,
    n825,
    n730
  );


  nand
  g932
  (
    n1267,
    n746,
    n327,
    n924,
    n323
  );


  or
  g933
  (
    n993,
    n758,
    n894,
    n936,
    n875
  );


  nor
  g934
  (
    n1323,
    n695,
    n342,
    n626,
    n913
  );


  and
  g935
  (
    n990,
    n472,
    n895,
    n707,
    n911
  );


  and
  g936
  (
    n1132,
    n479,
    n317,
    n846,
    n935
  );


  xnor
  g937
  (
    n1125,
    n672,
    n724,
    n919,
    n584
  );


  nor
  g938
  (
    n1047,
    n916,
    n463,
    n471,
    n943
  );


  and
  g939
  (
    n1246,
    n802,
    n741,
    n695,
    n591
  );


  nor
  g940
  (
    n1135,
    n897,
    n763,
    n853,
    n911
  );


  or
  g941
  (
    n1143,
    n877,
    n818,
    n382,
    n808
  );


  xnor
  g942
  (
    n983,
    n865,
    n577,
    n784,
    n765
  );


  nor
  g943
  (
    n1328,
    n357,
    n734,
    n779,
    n856
  );


  and
  g944
  (
    n1302,
    n941,
    n343,
    n711,
    n908
  );


  or
  g945
  (
    n1096,
    n467,
    n878,
    n812,
    n893
  );


  or
  g946
  (
    n1128,
    n745,
    n598,
    n942,
    n685
  );


  nand
  g947
  (
    n1129,
    n326,
    n418,
    n557,
    n908
  );


  or
  g948
  (
    n1330,
    n858,
    n283,
    n771,
    n820
  );


  xnor
  g949
  (
    n1153,
    n482,
    n572,
    n541,
    n699
  );


  and
  g950
  (
    n1083,
    n516,
    n606,
    n402,
    n387
  );


  and
  g951
  (
    n1119,
    n440,
    n766,
    n459,
    n840
  );


  nand
  g952
  (
    n1259,
    n467,
    n813,
    n389,
    n344
  );


  and
  g953
  (
    n1090,
    n688,
    n892,
    n633,
    n391
  );


  xnor
  g954
  (
    n1173,
    n582,
    n405,
    n855,
    n625
  );


  xor
  g955
  (
    n1053,
    n934,
    n929,
    n719,
    n485
  );


  xnor
  g956
  (
    n985,
    n513,
    n901,
    n407,
    n898
  );


  and
  g957
  (
    n1284,
    n514,
    n806,
    n887,
    n392
  );


  xnor
  g958
  (
    n1195,
    n656,
    n603,
    n943,
    n925
  );


  xnor
  g959
  (
    n1237,
    n892,
    n933,
    n514,
    n828
  );


  nor
  g960
  (
    n1326,
    n503,
    n589,
    n418,
    n308
  );


  nor
  g961
  (
    n1170,
    n372,
    n833,
    n653,
    n603
  );


  nand
  g962
  (
    n1198,
    n740,
    n400,
    n838,
    n886
  );


  xnor
  g963
  (
    n1130,
    n317,
    n721,
    n383,
    n345
  );


  xnor
  g964
  (
    n1319,
    n596,
    n369,
    n673,
    n493
  );


  xnor
  g965
  (
    n1234,
    n350,
    n687,
    n359,
    n473
  );


  xnor
  g966
  (
    n963,
    n913,
    n748,
    n507,
    n298
  );


  or
  g967
  (
    n966,
    n848,
    n301,
    n484,
    n727
  );


  or
  g968
  (
    n968,
    n878,
    n947,
    n509,
    n302
  );


  xnor
  g969
  (
    n1276,
    n940,
    n666,
    n368,
    n702
  );


  xor
  g970
  (
    n1278,
    n346,
    n656,
    n515,
    n904
  );


  xor
  g971
  (
    n1308,
    n503,
    n399,
    n365,
    n919
  );


  and
  g972
  (
    n1050,
    n755,
    n639,
    n526,
    n558
  );


  and
  g973
  (
    n1268,
    n940,
    n768,
    n915,
    n735
  );


  and
  g974
  (
    n1254,
    n930,
    n677,
    n652,
    n636
  );


  xnor
  g975
  (
    n1188,
    n783,
    n611,
    n825,
    n502
  );


  xnor
  g976
  (
    n1157,
    n699,
    n832,
    n751,
    n932
  );


  and
  g977
  (
    n1131,
    n856,
    n419,
    n642,
    n664
  );


  nand
  g978
  (
    n1318,
    n294,
    n906,
    n829,
    n632
  );


  and
  g979
  (
    n1035,
    n445,
    n443,
    n413,
    n714
  );


  xor
  g980
  (
    n1257,
    n573,
    n920,
    n415,
    n702
  );


  xor
  g981
  (
    n1235,
    n316,
    n333,
    n399,
    n332
  );


  xor
  g982
  (
    n1048,
    n737,
    n456,
    n653,
    n460
  );


  nand
  g983
  (
    n1098,
    n874,
    n466,
    n551,
    n906
  );


  or
  g984
  (
    n1008,
    n640,
    n852,
    n923,
    n760
  );


  xor
  g985
  (
    n1043,
    n615,
    n704,
    n804,
    n926
  );


  xor
  g986
  (
    n1317,
    n380,
    n629,
    n532,
    n396
  );


  nor
  g987
  (
    n1097,
    n906,
    n686,
    n403,
    n290
  );


  and
  g988
  (
    n1179,
    n482,
    n608,
    n321,
    n668
  );


  xnor
  g989
  (
    n987,
    n663,
    n618,
    n512,
    n710
  );


  and
  g990
  (
    n1189,
    n383,
    n464,
    n705,
    n886
  );


  xor
  g991
  (
    n1113,
    n761,
    n554,
    n469,
    n487
  );


  xor
  g992
  (
    n1309,
    n388,
    n291,
    n858,
    n701
  );


  nor
  g993
  (
    n1068,
    n847,
    n738,
    n506,
    n854
  );


  nand
  g994
  (
    n1277,
    n942,
    n841,
    n934,
    n463
  );


  nor
  g995
  (
    n1306,
    n620,
    n434,
    n876,
    n379
  );


  and
  g996
  (
    n1218,
    n569,
    n867,
    n406,
    n470
  );


  and
  g997
  (
    n1071,
    n422,
    n904,
    n564,
    n842
  );


  nand
  g998
  (
    n1212,
    n893,
    n849,
    n426,
    n674
  );


  and
  g999
  (
    n1169,
    n824,
    n877,
    n841,
    n917
  );


  nor
  g1000
  (
    n1226,
    n813,
    n769,
    n511,
    n632
  );


  or
  g1001
  (
    n1031,
    n911,
    n922,
    n935,
    n421
  );


  and
  g1002
  (
    n1185,
    n946,
    n629,
    n574,
    n690
  );


  and
  g1003
  (
    n1066,
    n822,
    n914,
    n519,
    n559
  );


  nor
  g1004
  (
    n1209,
    n348,
    n700,
    n854,
    n926
  );


  xnor
  g1005
  (
    n1229,
    n901,
    n910,
    n410,
    n387
  );


  and
  g1006
  (
    n1332,
    n707,
    n788,
    n661,
    n453
  );


  nand
  g1007
  (
    n1089,
    n769,
    n293,
    n394,
    n592
  );


  nor
  g1008
  (
    n1099,
    n742,
    n344,
    n759,
    n377
  );


  xnor
  g1009
  (
    n1194,
    n433,
    n912,
    n924,
    n933
  );


  and
  g1010
  (
    n965,
    n698,
    n891,
    n823,
    n648
  );


  xnor
  g1011
  (
    n1263,
    n771,
    n351,
    n663,
    n808
  );


  or
  g1012
  (
    n1206,
    n430,
    n926,
    n568,
    n680
  );


  nor
  g1013
  (
    n1281,
    n893,
    n805,
    n307,
    n874
  );


  or
  g1014
  (
    n1296,
    n749,
    n594,
    n869,
    n907
  );


  or
  g1015
  (
    n1011,
    n447,
    n930,
    n845,
    n875
  );


  xor
  g1016
  (
    n1165,
    n554,
    n921,
    n339,
    n403
  );


  or
  g1017
  (
    n1149,
    n581,
    n341,
    n907,
    n883
  );


  xor
  g1018
  (
    n1145,
    n733,
    n936,
    n730,
    n433
  );


  or
  g1019
  (
    n972,
    n728,
    n376,
    n325,
    n303
  );


  xor
  g1020
  (
    n1019,
    n920,
    n648,
    n543,
    n923
  );


  xor
  g1021
  (
    n973,
    n853,
    n367,
    n406,
    n366
  );


  xor
  g1022
  (
    n1168,
    n349,
    n907,
    n558,
    n539
  );


  xor
  g1023
  (
    n1134,
    n944,
    n782,
    n835,
    n912
  );


  nand
  g1024
  (
    n1193,
    n660,
    n807,
    n889,
    n703
  );


  and
  g1025
  (
    n1091,
    n819,
    n505,
    n453,
    n634
  );


  nand
  g1026
  (
    n1018,
    n347,
    n932,
    n490,
    n676
  );


  or
  g1027
  (
    n1010,
    n884,
    n805,
    n659,
    n547
  );


  xnor
  g1028
  (
    n967,
    n583,
    n551,
    n913,
    n521
  );


  xor
  g1029
  (
    n1270,
    n887,
    n465,
    n798,
    n462
  );


  and
  g1030
  (
    n1126,
    n502,
    n476,
    n946,
    n927
  );


  xor
  g1031
  (
    n1067,
    n376,
    n786,
    n824,
    n292
  );


  xnor
  g1032
  (
    n1311,
    n939,
    n290,
    n927,
    n649
  );


  xor
  g1033
  (
    n1219,
    n549,
    n938,
    n322,
    n839
  );


  and
  g1034
  (
    n1022,
    n915,
    n510,
    n809,
    n429
  );


  xnor
  g1035
  (
    n1070,
    n869,
    n362,
    n896,
    n488
  );


  nor
  g1036
  (
    n1014,
    n799,
    n356,
    n526,
    n887
  );


  nor
  g1037
  (
    n1073,
    n651,
    n299,
    n597,
    n712
  );


  xor
  g1038
  (
    n1217,
    n720,
    n422,
    n739,
    n889
  );


  and
  g1039
  (
    n1211,
    n303,
    n844,
    n607,
    n309
  );


  and
  g1040
  (
    n1002,
    n899,
    n829,
    n888,
    n325
  );


  and
  g1041
  (
    n1294,
    n716,
    n935,
    n790,
    n696
  );


  and
  g1042
  (
    n1264,
    n581,
    n507,
    n834,
    n555
  );


  xnor
  g1043
  (
    n964,
    n661,
    n739,
    n896,
    n615
  );


  or
  g1044
  (
    n1285,
    n937,
    n938,
    n452,
    n857
  );


  xnor
  g1045
  (
    n1140,
    n548,
    n747,
    n600,
    n449
  );


  and
  g1046
  (
    n1141,
    n416,
    n870,
    n884,
    n887
  );


  and
  g1047
  (
    n1147,
    n381,
    n620,
    n334,
    n420
  );


  nand
  g1048
  (
    n1148,
    n647,
    n322,
    n448,
    n614
  );


  xor
  g1049
  (
    n1144,
    n340,
    n677,
    n878,
    n882
  );


  and
  g1050
  (
    n986,
    n518,
    n566,
    n890,
    n571
  );


  or
  g1051
  (
    n1292,
    n836,
    n381,
    n886,
    n590
  );


  nor
  g1052
  (
    n978,
    n300,
    n535,
    n922,
    n773
  );


  or
  g1053
  (
    n1085,
    n587,
    n691,
    n608,
    n349
  );


  and
  g1054
  (
    n1321,
    n872,
    n338,
    n457,
    n818
  );


  xnor
  g1055
  (
    n1046,
    n757,
    n832,
    n791,
    n684
  );


  or
  g1056
  (
    n1075,
    n304,
    n394,
    n880,
    n756
  );


  nor
  g1057
  (
    n1327,
    n427,
    n560,
    n764,
    n901
  );


  nand
  g1058
  (
    n1081,
    n888,
    n793,
    n670,
    n881
  );


  and
  g1059
  (
    n1286,
    n446,
    n770,
    n500,
    n426
  );


  or
  g1060
  (
    n1084,
    n857,
    n546,
    n943,
    n754
  );


  nand
  g1061
  (
    n1183,
    n937,
    n566,
    n800,
    n814
  );


  nor
  g1062
  (
    n1177,
    n944,
    n908,
    n869,
    n922
  );


  or
  g1063
  (
    n1271,
    n401,
    n836,
    n811,
    n543
  );


  nand
  g1064
  (
    n1005,
    n594,
    n391,
    n649,
    n537
  );


  and
  g1065
  (
    n1182,
    n936,
    n643,
    n909,
    n517
  );


  xor
  g1066
  (
    n1248,
    n882,
    n302,
    n741,
    n917
  );


  nor
  g1067
  (
    n1155,
    n652,
    n900,
    n843,
    n395
  );


  xnor
  g1068
  (
    n1110,
    n714,
    n816,
    n918,
    n930
  );


  or
  g1069
  (
    n1095,
    n569,
    n419,
    n497,
    n540
  );


  and
  g1070
  (
    n1315,
    n870,
    n922,
    n413,
    n794
  );


  and
  g1071
  (
    n1262,
    n619,
    n464,
    n868,
    n664
  );


  or
  g1072
  (
    n1100,
    n390,
    n844,
    n693,
    n885
  );


  nand
  g1073
  (
    n1162,
    n942,
    n535,
    n438,
    n301
  );


  nor
  g1074
  (
    n1175,
    n339,
    n328,
    n885,
    n903
  );


  xnor
  g1075
  (
    n1205,
    n866,
    n720,
    n564,
    n616
  );


  xor
  g1076
  (
    n1251,
    n428,
    n533,
    n732,
    n436
  );


  nand
  g1077
  (
    n1334,
    n506,
    n444,
    n921,
    n319
  );


  nor
  g1078
  (
    n1051,
    n855,
    n318,
    n667,
    n492
  );


  xor
  g1079
  (
    n1108,
    n536,
    n811,
    n884,
    n890
  );


  or
  g1080
  (
    n1054,
    n420,
    n903,
    n585,
    n284
  );


  xor
  g1081
  (
    n1304,
    n495,
    n446,
    n777,
    n670
  );


  nor
  g1082
  (
    n1045,
    n423,
    n635,
    n774,
    n488
  );


  and
  g1083
  (
    n1214,
    n560,
    n571,
    n417,
    n723
  );


  nor
  g1084
  (
    n1142,
    n897,
    n368,
    n561,
    n874
  );


  or
  g1085
  (
    n1191,
    n886,
    n683,
    n402,
    n788
  );


  and
  g1086
  (
    n1106,
    n941,
    n912,
    n938,
    n404
  );


  or
  g1087
  (
    n998,
    n545,
    n852,
    n925,
    n645
  );


  nor
  g1088
  (
    n1015,
    n414,
    n424,
    n873,
    n489
  );


  nand
  g1089
  (
    n1065,
    n498,
    n477,
    n550,
    n519
  );


  or
  g1090
  (
    n1289,
    n431,
    n712,
    n528,
    n792
  );


  xor
  g1091
  (
    n1228,
    n545,
    n644,
    n817,
    n487
  );


  xnor
  g1092
  (
    n1138,
    n665,
    n523,
    n425,
    n331
  );


  nor
  g1093
  (
    n1210,
    n647,
    n917,
    n916,
    n679
  );


  or
  g1094
  (
    n979,
    n579,
    n530,
    n354,
    n480
  );


  nand
  g1095
  (
    n1017,
    n946,
    n787,
    n342,
    n561
  );


  xnor
  g1096
  (
    n962,
    n917,
    n745,
    n537,
    n782
  );


  nand
  g1097
  (
    n1024,
    n444,
    n588,
    n622,
    n496
  );


  xnor
  g1098
  (
    n1056,
    n891,
    n622,
    n845,
    n689
  );


  nor
  g1099
  (
    n1030,
    n304,
    n449,
    n364,
    n341
  );


  and
  g1100
  (
    n1290,
    n731,
    n565,
    n905,
    n732
  );


  or
  g1101
  (
    n1034,
    n481,
    n333,
    n868,
    n915
  );


  and
  g1102
  (
    n1023,
    n610,
    n327,
    n797,
    n762
  );


  nor
  g1103
  (
    n988,
    n599,
    n531,
    n296,
    n686
  );


  nor
  g1104
  (
    n1280,
    n758,
    n640,
    n870,
    n826
  );


  nand
  g1105
  (
    n1049,
    n688,
    n931,
    n678,
    n725
  );


  and
  g1106
  (
    n1080,
    n491,
    n578,
    n708,
    n434
  );


  xor
  g1107
  (
    n991,
    n362,
    n534,
    n754,
    n542
  );


  nor
  g1108
  (
    n1061,
    n763,
    n822,
    n837,
    n892
  );


  xnor
  g1109
  (
    n971,
    n582,
    n697,
    n624,
    n494
  );


  xnor
  g1110
  (
    n1305,
    n334,
    n515,
    n628,
    n494
  );


  and
  g1111
  (
    n1094,
    n382,
    n455,
    n466,
    n616
  );


  and
  g1112
  (
    n996,
    n925,
    n862,
    n430,
    n803
  );


  and
  g1113
  (
    n1310,
    n945,
    n477,
    n892,
    n736
  );


  nand
  g1114
  (
    n1301,
    n873,
    n484,
    n459,
    n722
  );


  nand
  g1115
  (
    n1320,
    n617,
    n796,
    n881,
    n934
  );


  nand
  g1116
  (
    n994,
    n796,
    n363,
    n777,
    n923
  );


  or
  g1117
  (
    n1322,
    n842,
    n861,
    n612,
    n838
  );


  xnor
  g1118
  (
    n1295,
    n693,
    n929,
    n447,
    n520
  );


  xnor
  g1119
  (
    n1006,
    n914,
    n921,
    n289,
    n475
  );


  nor
  g1120
  (
    n1167,
    n440,
    n312,
    n690,
    n789
  );


  nand
  g1121
  (
    n1037,
    n809,
    n562,
    n940,
    n883
  );


  xor
  g1122
  (
    n1112,
    n784,
    n912,
    n438,
    n872
  );


  and
  g1123
  (
    n995,
    n933,
    n723,
    n814,
    n356
  );


  or
  g1124
  (
    n1032,
    n641,
    n867,
    n348,
    n744
  );


  nor
  g1125
  (
    n1044,
    n860,
    n637,
    n575,
    n884
  );


  xnor
  g1126
  (
    n1057,
    n384,
    n709,
    n743,
    n539
  );


  xor
  g1127
  (
    n1062,
    n337,
    n945,
    n498,
    n553
  );


  nor
  g1128
  (
    n1275,
    n928,
    n896,
    n345,
    n889
  );


  nor
  g1129
  (
    n1216,
    n340,
    n445,
    n871,
    n898
  );


  nand
  g1130
  (
    n1256,
    n850,
    n454,
    n657,
    n928
  );


  nand
  g1131
  (
    n1039,
    n613,
    n933,
    n353,
    n305
  );


  or
  g1132
  (
    n1076,
    n363,
    n920,
    n885,
    n937
  );


  and
  g1133
  (
    n977,
    n454,
    n735,
    n683,
    n655
  );


  xnor
  g1134
  (
    n1184,
    n897,
    n409,
    n696,
    n417
  );


  nand
  g1135
  (
    n1133,
    n563,
    n567,
    n767,
    n821
  );


  and
  g1136
  (
    n1250,
    n353,
    n311,
    n801,
    n902
  );


  and
  g1137
  (
    n1324,
    n481,
    n778,
    n352,
    n429
  );


  nor
  g1138
  (
    n1004,
    n877,
    n604,
    n587,
    n531
  );


  xor
  g1139
  (
    n1215,
    n727,
    n329,
    n654,
    n918
  );


  and
  g1140
  (
    n1137,
    n914,
    n728,
    n586,
    n337
  );


  or
  g1141
  (
    n1114,
    n726,
    n442,
    n874,
    n937
  );


  nor
  g1142
  (
    n1000,
    n715,
    n504,
    n918,
    n324
  );


  xor
  g1143
  (
    n1291,
    n635,
    n837,
    n516,
    n634
  );


  and
  g1144
  (
    n1158,
    n680,
    n380,
    n588,
    n352
  );


  xor
  g1145
  (
    n974,
    n785,
    n803,
    n609,
    n525
  );


  nor
  g1146
  (
    n1058,
    n493,
    n909,
    n592,
    n295
  );


  and
  g1147
  (
    n1253,
    n815,
    n896,
    n485,
    n807
  );


  nor
  g1148
  (
    n1120,
    n606,
    n398,
    n734,
    n604
  );


  xnor
  g1149
  (
    n1020,
    n324,
    n500,
    n935,
    n736
  );


  nand
  g1150
  (
    n1252,
    n889,
    n880,
    n673,
    n795
  );


  and
  g1151
  (
    n1087,
    n760,
    n330,
    n717,
    n575
  );


  xnor
  g1152
  (
    n992,
    n655,
    n768,
    n873,
    n666
  );


  xor
  g1153
  (
    n1163,
    n522,
    n725,
    n369,
    n450
  );


  nor
  g1154
  (
    n1104,
    n492,
    n715,
    n878,
    n286
  );


  xnor
  g1155
  (
    n1124,
    n806,
    n286,
    n416,
    n318
  );


  nand
  g1156
  (
    n1118,
    n607,
    n724,
    n678,
    n552
  );


  or
  g1157
  (
    n1203,
    n659,
    n567,
    n495,
    n326
  );


  nor
  g1158
  (
    n1026,
    n871,
    n310,
    n396,
    n752
  );


  nand
  g1159
  (
    n1016,
    n512,
    n532,
    n877,
    n800
  );


  xor
  g1160
  (
    n976,
    n827,
    n895,
    n389,
    n457
  );


  nand
  g1161
  (
    n1260,
    n627,
    n718,
    n578,
    n573
  );


  or
  g1162
  (
    n1176,
    n753,
    n287,
    n315,
    n713
  );


  nand
  g1163
  (
    n1266,
    n522,
    n795,
    n883,
    n411
  );


  and
  g1164
  (
    n1060,
    n848,
    n704,
    n370,
    n291
  );


  xnor
  g1165
  (
    n1078,
    n431,
    n859,
    n562,
    n586
  );


  and
  g1166
  (
    n1288,
    n755,
    n443,
    n613,
    n521
  );


  and
  g1167
  (
    n1220,
    n472,
    n833,
    n802,
    n684
  );


  nand
  g1168
  (
    n1086,
    n870,
    n625,
    n305,
    n407
  );


  and
  g1169
  (
    n999,
    n650,
    n930,
    n751,
    n733
  );


  nand
  g1170
  (
    n1072,
    n785,
    n395,
    n513,
    n703
  );


  nand
  g1171
  (
    n1159,
    n478,
    n415,
    n750,
    n942
  );


  and
  g1172
  (
    n1204,
    n692,
    n293,
    n595,
    n458
  );


  nand
  g1173
  (
    n1160,
    n524,
    n929,
    n523,
    n408
  );


  xnor
  g1174
  (
    n1283,
    n633,
    n491,
    n421,
    n423
  );


  xnor
  g1175
  (
    n1223,
    n336,
    n682,
    n830,
    n306
  );


  or
  g1176
  (
    n1021,
    n899,
    n576,
    n905,
    n546
  );


  or
  g1177
  (
    n1154,
    n602,
    n474,
    n820,
    n898
  );


  nor
  g1178
  (
    n1139,
    n501,
    n789,
    n931,
    n910
  );


  xnor
  g1179
  (
    n1093,
    n919,
    n536,
    n772,
    n471
  );


  xnor
  g1180
  (
    n1064,
    n913,
    n907,
    n939,
    n614
  );


  xnor
  g1181
  (
    n1303,
    n372,
    n469,
    n580,
    n583
  );


  or
  g1182
  (
    n1101,
    n883,
    n740,
    n359,
    n367
  );


  nor
  g1183
  (
    n1146,
    n297,
    n497,
    n478,
    n888
  );


  or
  g1184
  (
    n1238,
    n748,
    n486,
    n691,
    n294
  );


  xnor
  g1185
  (
    n1115,
    n462,
    n780,
    n749,
    n315
  );


  nor
  g1186
  (
    n1233,
    n511,
    n903,
    n412,
    n335
  );


  and
  g1187
  (
    n1243,
    n787,
    n375,
    n669,
    n746
  );


  xnor
  g1188
  (
    n1186,
    n282,
    n400,
    n328,
    n672
  );


  and
  g1189
  (
    n1261,
    n876,
    n631,
    n894,
    n350
  );


  xnor
  g1190
  (
    n1029,
    n398,
    n557,
    n320,
    n931
  );


  xnor
  g1191
  (
    n1293,
    n427,
    n726,
    n899,
    n593
  );


  xnor
  g1192
  (
    n1152,
    n773,
    n761,
    n776,
    n743
  );


  nor
  g1193
  (
    n1279,
    n530,
    n504,
    n489,
    n774
  );


  xnor
  g1194
  (
    n1282,
    n881,
    n775,
    n864,
    n890
  );


  nand
  g1195
  (
    n1009,
    n770,
    n297,
    n520,
    n534
  );


  and
  g1196
  (
    n1249,
    n364,
    n849,
    n347,
    n882
  );


  xnor
  g1197
  (
    n1213,
    n641,
    n627,
    n517,
    n801
  );


  nand
  g1198
  (
    n1069,
    n668,
    n601,
    n645,
    n939
  );


  xnor
  g1199
  (
    n1123,
    n451,
    n458,
    n924,
    n414
  );


  or
  g1200
  (
    n1240,
    n941,
    n388,
    n541,
    n810
  );


  nand
  g1201
  (
    n1150,
    n871,
    n742,
    n288,
    n374
  );


  xor
  g1202
  (
    n1105,
    n750,
    n900,
    n729,
    n411
  );


  xnor
  g1203
  (
    n1221,
    n863,
    n909,
    n626,
    n437
  );


  or
  g1204
  (
    n1325,
    n378,
    n623,
    n639,
    n624
  );


  xnor
  g1205
  (
    n1127,
    n658,
    n692,
    n804,
    n556
  );


  nand
  g1206
  (
    n1224,
    n306,
    n775,
    n361,
    n570
  );


  xor
  g1207
  (
    n1231,
    n358,
    n835,
    n599,
    n916
  );


  xnor
  g1208
  (
    n1027,
    n662,
    n617,
    n335,
    n605
  );


  nand
  g1209
  (
    n1273,
    n872,
    n373,
    n483,
    n563
  );


  or
  g1210
  (
    n1181,
    n662,
    n450,
    n799,
    n932
  );


  nand
  g1211
  (
    n1225,
    n529,
    n729,
    n611,
    n598
  );


  and
  g1212
  (
    n1007,
    n898,
    n860,
    n851,
    n397
  );


  xnor
  g1213
  (
    n969,
    n766,
    n840,
    n357,
    n947
  );


  or
  g1214
  (
    n1025,
    n374,
    n393,
    n320,
    n580
  );


  or
  g1215
  (
    n1088,
    n638,
    n867,
    n709,
    n671
  );


  nand
  g1216
  (
    n1180,
    n285,
    n867,
    n694,
    n918
  );


  or
  g1217
  (
    n1190,
    n527,
    n631,
    n900,
    n931
  );


  nor
  g1218
  (
    n1274,
    n378,
    n473,
    n881,
    n612
  );


  nand
  g1219
  (
    n1297,
    n605,
    n559,
    n810,
    n321
  );


  nand
  g1220
  (
    n982,
    n392,
    n865,
    n819,
    n895
  );


  or
  g1221
  (
    n1079,
    n584,
    n409,
    n821,
    n719
  );


  xor
  g1222
  (
    n1255,
    n371,
    n448,
    n437,
    n283
  );


  or
  g1223
  (
    n1116,
    n425,
    n570,
    n548,
    n910
  );


  nor
  g1224
  (
    n1202,
    n675,
    n474,
    n650,
    n556
  );


  or
  g1225
  (
    n1196,
    n676,
    n547,
    n934,
    n718
  );


  or
  g1226
  (
    n1156,
    n946,
    n816,
    n851,
    n897
  );


  xor
  g1227
  (
    n1111,
    n879,
    n314,
    n875,
    n385
  );


  xor
  g1228
  (
    n1329,
    n783,
    n284,
    n373,
    n839
  );


  nor
  g1229
  (
    n1207,
    n486,
    n895,
    n823,
    n916
  );


  xor
  g1230
  (
    n984,
    n772,
    n619,
    n894,
    n921
  );


  xor
  g1231
  (
    n1287,
    n314,
    n442,
    n928,
    n738
  );


  nand
  g1232
  (
    n1316,
    n651,
    n282,
    n831,
    n424
  );


  and
  g1233
  (
    n1121,
    n843,
    n377,
    n550,
    n596
  );


  or
  g1234
  (
    n1299,
    n929,
    n576,
    n759,
    n681
  );


  and
  g1235
  (
    n1313,
    n891,
    n875,
    n379,
    n872
  );


  nor
  g1236
  (
    n1122,
    n358,
    n927,
    n386,
    n371
  );


  xor
  g1237
  (
    n1222,
    n906,
    n628,
    n757,
    n831
  );


  xnor
  g1238
  (
    n1172,
    n295,
    n595,
    n289,
    n879
  );


  nor
  g1239
  (
    n1300,
    n885,
    n710,
    n568,
    n764
  );


  xor
  g1240
  (
    n997,
    n939,
    n574,
    n441,
    n744
  );


  nor
  g1241
  (
    n1033,
    n540,
    n846,
    n553,
    n296
  );


  xnor
  g1242
  (
    n1117,
    n452,
    n470,
    n786,
    n682
  );


  nand
  g1243
  (
    n1164,
    n351,
    n610,
    n700,
    n869
  );


  xnor
  g1244
  (
    n1187,
    n412,
    n890,
    n637,
    n309
  );


  nor
  g1245
  (
    n1208,
    n355,
    n505,
    n509,
    n313
  );


  nor
  g1246
  (
    n1001,
    n826,
    n847,
    n319,
    n904
  );


  nand
  g1247
  (
    n1244,
    n941,
    n667,
    n508,
    n589
  );


  xor
  g1248
  (
    n1236,
    n671,
    n902,
    n882,
    n393
  );


  xnor
  g1249
  (
    n1171,
    n924,
    n893,
    n657,
    n873
  );


  xnor
  g1250
  (
    n1227,
    n490,
    n479,
    n797,
    n602
  );


  or
  g1251
  (
    n989,
    n375,
    n465,
    n527,
    n518
  );


  and
  g1252
  (
    n1109,
    n863,
    n868,
    n287,
    n879
  );


  nor
  g1253
  (
    n1103,
    n945,
    n944,
    n790,
    n850
  );


  xor
  g1254
  (
    n1200,
    n765,
    n756,
    n601,
    n830
  );


  nor
  g1255
  (
    n1232,
    n525,
    n630,
    n310,
    n336
  );


  nand
  g1256
  (
    n981,
    n798,
    n646,
    n880,
    n544
  );


  xnor
  g1257
  (
    n1063,
    n642,
    n476,
    n905,
    n552
  );


  nand
  g1258
  (
    n1242,
    n538,
    n544,
    n524,
    n355
  );


  xor
  g1259
  (
    n1272,
    n292,
    n674,
    n323,
    n542
  );


  nand
  g1260
  (
    n1245,
    n915,
    n685,
    n410,
    n779
  );


  or
  g1261
  (
    n1042,
    n468,
    n722,
    n711,
    n689
  );


  xnor
  g1262
  (
    n1013,
    n827,
    n914,
    n386,
    n834
  );


  nand
  g1263
  (
    n1036,
    n299,
    n909,
    n899,
    n721
  );


  nand
  g1264
  (
    n1201,
    n572,
    n555,
    n902,
    n565
  );


  and
  g1265
  (
    n1178,
    n920,
    n288,
    n585,
    n330
  );


  xnor
  g1266
  (
    n1077,
    n577,
    n591,
    n510,
    n903
  );


  nand
  g1267
  (
    n1230,
    n908,
    n940,
    n864,
    n496
  );


  and
  g1268
  (
    n1247,
    n475,
    n499,
    n675,
    n483
  );


  xnor
  g1269
  (
    n1074,
    n436,
    n747,
    n285,
    n638
  );


  nor
  g1270
  (
    n1239,
    n752,
    n919,
    n621,
    n900
  );


  xor
  g1271
  (
    n1174,
    n461,
    n776,
    n538,
    n354
  );


  nand
  g1272
  (
    n1055,
    n932,
    n817,
    n346,
    n928
  );


  xnor
  g1273
  (
    n1258,
    n902,
    n360,
    n658,
    n366
  );


  xor
  g1274
  (
    n1028,
    n300,
    n508,
    n911,
    n861
  );


  or
  g1275
  (
    n1333,
    n435,
    n528,
    n643,
    n868
  );


  xnor
  g1276
  (
    n1298,
    n938,
    n307,
    n439,
    n600
  );


  xnor
  g1277
  (
    n1161,
    n338,
    n706,
    n549,
    n456
  );


  and
  g1278
  (
    n1041,
    n439,
    n298,
    n862,
    n501
  );


  nor
  g1279
  (
    n980,
    n390,
    n737,
    n408,
    n316
  );


  or
  g1280
  (
    n1082,
    n687,
    n361,
    n708,
    n329
  );


  and
  g1281
  (
    n970,
    n694,
    n894,
    n891,
    n468
  );


  nand
  g1282
  (
    n1059,
    n480,
    n405,
    n313,
    n879
  );


  xor
  g1283
  (
    n1038,
    n597,
    n451,
    n701,
    n384
  );


  xor
  g1284
  (
    n1312,
    n880,
    n762,
    n753,
    n593
  );


  nand
  g1285
  (
    n1102,
    n665,
    n630,
    n590,
    n697
  );


  xnor
  g1286
  (
    n1107,
    n660,
    n654,
    n778,
    n428
  );


  xor
  g1287
  (
    n1003,
    n716,
    n781,
    n888,
    n529
  );


  or
  g1288
  (
    n1265,
    n717,
    n432,
    n876,
    n360
  );


  or
  g1289
  (
    n1166,
    n623,
    n401,
    n370,
    n926
  );


  xnor
  g1290
  (
    n1012,
    n646,
    n332,
    n441,
    n943
  );


  and
  g1291
  (
    n1040,
    n343,
    n644,
    n910,
    n871
  );


  or
  g1292
  (
    n1269,
    n308,
    n927,
    n669,
    n713
  );


  nand
  g1293
  (
    n1197,
    n618,
    n767,
    n904,
    n812
  );


  xnor
  g1294
  (
    n1199,
    n533,
    n945,
    n780,
    n876
  );


  or
  g1295
  (
    n1307,
    n731,
    n636,
    n621,
    n460
  );


  nor
  g1296
  (
    n1092,
    n925,
    n706,
    n385,
    n866
  );


  nor
  g1297
  (
    n1331,
    n923,
    n311,
    n365,
    n499
  );


  xor
  g1298
  (
    n1151,
    n435,
    n781,
    n794,
    n815
  );


  nor
  g1299
  (
    n1314,
    n698,
    n905,
    n609,
    n681
  );


  and
  g1300
  (
    n1136,
    n936,
    n404,
    n705,
    n455
  );


  and
  g1301
  (
    n1192,
    n859,
    n944,
    n679,
    n312
  );


  nand
  g1302
  (
    n1340,
    n982,
    n1023,
    n974,
    n1005
  );


  xor
  g1303
  (
    n1336,
    n969,
    n986,
    n1031,
    n981
  );


  or
  g1304
  (
    n1345,
    n1010,
    n991,
    n1014,
    n966
  );


  or
  g1305
  (
    n1335,
    n979,
    n1026,
    n985,
    n1000
  );


  xnor
  g1306
  (
    n1350,
    n1018,
    n1020,
    n983,
    n1006
  );


  xor
  g1307
  (
    n1348,
    n964,
    n1007,
    n977,
    n1016
  );


  xnor
  g1308
  (
    n1343,
    n992,
    n1012,
    n1025,
    n976
  );


  and
  g1309
  (
    n1344,
    n989,
    n1009,
    n980,
    n995
  );


  or
  g1310
  (
    n1352,
    n1029,
    n1001,
    n963,
    n1022
  );


  xnor
  g1311
  (
    n1339,
    n997,
    n1003,
    n971,
    n962
  );


  or
  g1312
  (
    n1337,
    n987,
    n993,
    n1024,
    n968
  );


  nor
  g1313
  (
    n1342,
    n1019,
    n1015,
    n984,
    n996
  );


  xor
  g1314
  (
    n1341,
    n978,
    n1011,
    n988,
    n994
  );


  xor
  g1315
  (
    n1338,
    n967,
    n1032,
    n972,
    n1027
  );


  or
  g1316
  (
    n1347,
    n973,
    n998,
    n1030,
    n975
  );


  nor
  g1317
  (
    n1346,
    n990,
    n999,
    n1017,
    n1002
  );


  nor
  g1318
  (
    n1351,
    n1033,
    n1004,
    n970,
    n1028
  );


  nor
  g1319
  (
    n1349,
    n1021,
    n1008,
    n1013,
    n965
  );


  buf
  g1320
  (
    n1358,
    n1342
  );


  buf
  g1321
  (
    n1356,
    n1341
  );


  not
  g1322
  (
    n1354,
    n1339
  );


  not
  g1323
  (
    n1353,
    n1348
  );


  buf
  g1324
  (
    n1363,
    n1343
  );


  not
  g1325
  (
    n1355,
    n1336
  );


  not
  g1326
  (
    n1366,
    n269
  );


  not
  g1327
  (
    n1362,
    n1346
  );


  buf
  g1328
  (
    n1359,
    n1338
  );


  not
  g1329
  (
    n1357,
    n269
  );


  buf
  g1330
  (
    n1365,
    n1344
  );


  buf
  g1331
  (
    n1364,
    n1347
  );


  or
  g1332
  (
    n1361,
    n1340,
    n1335
  );


  nand
  g1333
  (
    n1360,
    n1345,
    n1337,
    n269
  );


  buf
  g1334
  (
    n1377,
    n1354
  );


  not
  g1335
  (
    n1371,
    n1358
  );


  buf
  g1336
  (
    n1379,
    n1359
  );


  buf
  g1337
  (
    n1372,
    n1353
  );


  buf
  g1338
  (
    n1380,
    n1357
  );


  buf
  g1339
  (
    n1368,
    n1356
  );


  buf
  g1340
  (
    n1382,
    n1355
  );


  not
  g1341
  (
    n1383,
    n1355
  );


  not
  g1342
  (
    n1381,
    n1359
  );


  not
  g1343
  (
    n1386,
    n1357
  );


  buf
  g1344
  (
    n1374,
    n1358
  );


  buf
  g1345
  (
    n1373,
    n1358
  );


  buf
  g1346
  (
    n1367,
    n1357
  );


  buf
  g1347
  (
    n1369,
    n1359
  );


  buf
  g1348
  (
    n1370,
    n1359
  );


  not
  g1349
  (
    n1375,
    n1357
  );


  not
  g1350
  (
    n1384,
    n1354
  );


  buf
  g1351
  (
    n1385,
    n1353
  );


  buf
  g1352
  (
    n1376,
    n1358
  );


  buf
  g1353
  (
    n1378,
    n1356
  );


  or
  g1354
  (
    n1456,
    n1173,
    n1369,
    n1241,
    n1270
  );


  xnor
  g1355
  (
    n1462,
    n1368,
    n1236,
    n1232,
    n1071
  );


  and
  g1356
  (
    n1443,
    n1145,
    n1378,
    n1374,
    n1182
  );


  nor
  g1357
  (
    n1450,
    n1062,
    n1257,
    n1226,
    n1197
  );


  nor
  g1358
  (
    n1455,
    n1181,
    n1227,
    n1177,
    n1120
  );


  nand
  g1359
  (
    n1444,
    n1101,
    n1104,
    n1114,
    n1382
  );


  xnor
  g1360
  (
    n1440,
    n1386,
    n1235,
    n1196,
    n1269
  );


  xnor
  g1361
  (
    n1417,
    n1133,
    n1155,
    n1371,
    n1213
  );


  nand
  g1362
  (
    n1405,
    n1260,
    n1147,
    n1249,
    n1386
  );


  or
  g1363
  (
    n1449,
    n1372,
    n1384,
    n1050,
    n1191
  );


  xor
  g1364
  (
    n1411,
    n1125,
    n1262,
    n1385,
    n1228
  );


  xnor
  g1365
  (
    n1453,
    n1080,
    n1201,
    n1045,
    n1156
  );


  nor
  g1366
  (
    n1421,
    n1242,
    n1383,
    n1251,
    n1246
  );


  xnor
  g1367
  (
    n1427,
    n1074,
    n1183,
    n1381,
    n1141
  );


  xor
  g1368
  (
    n1437,
    n1167,
    n1069,
    n1384,
    n1377
  );


  and
  g1369
  (
    n1429,
    n1038,
    n1068,
    n1093,
    n1157
  );


  xnor
  g1370
  (
    n1424,
    n1385,
    n1189,
    n1130,
    n1134
  );


  nor
  g1371
  (
    n1412,
    n1372,
    n1371,
    n1165,
    n1253
  );


  nor
  g1372
  (
    n1413,
    n1161,
    n1057,
    n1188,
    n1386
  );


  and
  g1373
  (
    n1396,
    n1267,
    n1090,
    n1209,
    n1218
  );


  nand
  g1374
  (
    n1409,
    n1273,
    n1124,
    n1210,
    n1233
  );


  nor
  g1375
  (
    n1401,
    n1138,
    n1372,
    n1265,
    n1162
  );


  xnor
  g1376
  (
    n1419,
    n1149,
    n1375,
    n1166,
    n1059
  );


  xnor
  g1377
  (
    n1416,
    n1041,
    n1373,
    n1383,
    n1217
  );


  or
  g1378
  (
    n1394,
    n1216,
    n1136,
    n1379,
    n1077
  );


  nor
  g1379
  (
    n1432,
    n1386,
    n1179,
    n1103,
    n1379
  );


  xor
  g1380
  (
    n1447,
    n1252,
    n1144,
    n1040,
    n1194
  );


  or
  g1381
  (
    n1466,
    n1370,
    n1374,
    n1375,
    n1271
  );


  nor
  g1382
  (
    n1457,
    n1369,
    n1231,
    n1368,
    n1079
  );


  xnor
  g1383
  (
    n1403,
    n1121,
    n1107,
    n1379,
    n1072
  );


  nor
  g1384
  (
    n1465,
    n1087,
    n1139,
    n1172,
    n1272
  );


  xor
  g1385
  (
    n1398,
    n1369,
    n1203,
    n1099,
    n1094
  );


  nand
  g1386
  (
    n1441,
    n1381,
    n1110,
    n1206,
    n1065
  );


  and
  g1387
  (
    n1423,
    n1067,
    n1381,
    n1176,
    n1380
  );


  or
  g1388
  (
    n1387,
    n1132,
    n1192,
    n1234,
    n1160
  );


  xor
  g1389
  (
    n1436,
    n1108,
    n1106,
    n1143,
    n1053
  );


  nand
  g1390
  (
    n1404,
    n1111,
    n1381,
    n1046,
    n1034
  );


  nand
  g1391
  (
    n1393,
    n1150,
    n1043,
    n1223,
    n1054
  );


  xor
  g1392
  (
    n1418,
    n1086,
    n1377,
    n1075,
    n1088
  );


  nand
  g1393
  (
    n1428,
    n1118,
    n1367,
    n1247,
    n1230
  );


  xor
  g1394
  (
    n1452,
    n1174,
    n1140,
    n1225,
    n1255
  );


  nand
  g1395
  (
    n1431,
    n1379,
    n1168,
    n1212,
    n1367
  );


  xnor
  g1396
  (
    n1407,
    n1055,
    n1219,
    n1187,
    n1229
  );


  or
  g1397
  (
    n1420,
    n1371,
    n1078,
    n1119,
    n1044
  );


  or
  g1398
  (
    n1392,
    n1100,
    n1142,
    n1238,
    n1244
  );


  nand
  g1399
  (
    n1425,
    n1169,
    n1377,
    n1215,
    n1385
  );


  xnor
  g1400
  (
    n1395,
    n1383,
    n1035,
    n1378
  );


  xor
  g1401
  (
    n1446,
    n1070,
    n1186,
    n1175,
    n1375
  );


  or
  g1402
  (
    n1430,
    n1367,
    n1049,
    n1259,
    n1116
  );


  and
  g1403
  (
    n1410,
    n1250,
    n1066,
    n1131,
    n1063
  );


  xnor
  g1404
  (
    n1458,
    n1370,
    n1254,
    n1221,
    n1185
  );


  xor
  g1405
  (
    n1426,
    n1380,
    n1170,
    n1383,
    n1064
  );


  nand
  g1406
  (
    n1454,
    n1382,
    n1266,
    n1037,
    n1243
  );


  xnor
  g1407
  (
    n1445,
    n1105,
    n1039,
    n1091,
    n1369
  );


  nor
  g1408
  (
    n1415,
    n1089,
    n1085,
    n1384
  );


  xor
  g1409
  (
    n1463,
    n1372,
    n1382,
    n1220,
    n1098
  );


  nand
  g1410
  (
    n1389,
    n1152,
    n1268,
    n1258,
    n1052
  );


  and
  g1411
  (
    n1399,
    n1109,
    n1199,
    n1204,
    n1153
  );


  xnor
  g1412
  (
    n1397,
    n1135,
    n1376,
    n1081,
    n1158
  );


  or
  g1413
  (
    n1461,
    n1373,
    n1073,
    n1375,
    n1083
  );


  xor
  g1414
  (
    n1435,
    n1163,
    n1123,
    n1376,
    n1082
  );


  xnor
  g1415
  (
    n1434,
    n1382,
    n1126,
    n1048,
    n1127
  );


  xor
  g1416
  (
    n1422,
    n1190,
    n1376,
    n1198,
    n1151
  );


  xor
  g1417
  (
    n1459,
    n1148,
    n1261,
    n1237,
    n1373
  );


  or
  g1418
  (
    n1460,
    n1096,
    n1211,
    n1154,
    n1263
  );


  nor
  g1419
  (
    n1406,
    n1092,
    n1380,
    n1368,
    n1222
  );


  nor
  g1420
  (
    n1433,
    n1245,
    n1129,
    n1380,
    n1180
  );


  or
  g1421
  (
    n1390,
    n1264,
    n1117,
    n1239,
    n1195
  );


  xnor
  g1422
  (
    n1402,
    n1047,
    n1256,
    n1368,
    n1128
  );


  nor
  g1423
  (
    n1451,
    n1208,
    n1376,
    n1373,
    n1171
  );


  xnor
  g1424
  (
    n1391,
    n1371,
    n1112,
    n1370,
    n1248
  );


  or
  g1425
  (
    n1408,
    n1200,
    n1060,
    n1178,
    n1122
  );


  xnor
  g1426
  (
    n1448,
    n1370,
    n1137,
    n1056,
    n1385
  );


  and
  g1427
  (
    n1439,
    n1042,
    n1207,
    n1193,
    n1084
  );


  and
  g1428
  (
    n1388,
    n1240,
    n1377,
    n1214,
    n1097
  );


  xor
  g1429
  (
    n1414,
    n1374,
    n1367,
    n1115,
    n1146
  );


  nor
  g1430
  (
    n1438,
    n1374,
    n1378,
    n1061,
    n1224
  );


  or
  g1431
  (
    n1400,
    n1051,
    n1159,
    n1184,
    n1058
  );


  nor
  g1432
  (
    n1464,
    n1113,
    n1202,
    n1076,
    n1095
  );


  xor
  g1433
  (
    n1442,
    n1036,
    n1164,
    n1205,
    n1102
  );


  not
  g1434
  (
    n1467,
    n1387
  );


  not
  g1435
  (
    n1468,
    n1387
  );


  not
  g1436
  (
    n1470,
    n1387
  );


  buf
  g1437
  (
    n1469,
    n1387
  );


  buf
  g1438
  (
    n1477,
    n1362
  );


  not
  g1439
  (
    n1472,
    n1467
  );


  nor
  g1440
  (
    n1478,
    n1467,
    n1280,
    n1363,
    n1468
  );


  xnor
  g1441
  (
    n1476,
    n1363,
    n1276,
    n1360
  );


  and
  g1442
  (
    n1473,
    n1361,
    n1360,
    n1275,
    n1362
  );


  or
  g1443
  (
    n1475,
    n1362,
    n1467,
    n1468
  );


  or
  g1444
  (
    n1471,
    n1468,
    n1277,
    n1469,
    n1360
  );


  xnor
  g1445
  (
    n1474,
    n1362,
    n1274,
    n1361,
    n1279
  );


  xnor
  g1446
  (
    n1479,
    n1278,
    n1361,
    n1468
  );


  buf
  g1447
  (
    n1484,
    n1473
  );


  buf
  g1448
  (
    n1493,
    n1471
  );


  not
  g1449
  (
    n1487,
    n1474
  );


  buf
  g1450
  (
    n1489,
    n1472
  );


  not
  g1451
  (
    n1480,
    n1471
  );


  not
  g1452
  (
    n1485,
    n1473
  );


  buf
  g1453
  (
    n1495,
    n1471
  );


  buf
  g1454
  (
    n1481,
    n1472
  );


  not
  g1455
  (
    n1494,
    n1474
  );


  buf
  g1456
  (
    n1491,
    n1473
  );


  not
  g1457
  (
    n1482,
    n1474
  );


  not
  g1458
  (
    n1492,
    n1474
  );


  not
  g1459
  (
    n1483,
    n1472
  );


  buf
  g1460
  (
    n1488,
    n1472
  );


  buf
  g1461
  (
    n1486,
    n1471
  );


  not
  g1462
  (
    n1490,
    n1473
  );


  xor
  g1463
  (
    n1543,
    n1390,
    n1401
  );


  nor
  g1464
  (
    n1522,
    n1394,
    n1483
  );


  xnor
  g1465
  (
    n1540,
    n1487,
    n1397,
    n1396,
    n1489
  );


  nor
  g1466
  (
    n1536,
    n1487,
    n1389,
    n1416,
    n1415
  );


  xor
  g1467
  (
    n1496,
    n1480,
    n1416,
    n1402,
    n1418
  );


  or
  g1468
  (
    n1535,
    n1481,
    n1424,
    n1389,
    n1409
  );


  nor
  g1469
  (
    n1519,
    n1486,
    n1402,
    n1415,
    n1406
  );


  xnor
  g1470
  (
    n1542,
    n1420,
    n1409,
    n1413,
    n1423
  );


  nand
  g1471
  (
    n1499,
    n1424,
    n1488,
    n1413,
    n1421
  );


  or
  g1472
  (
    n1548,
    n1400,
    n1426,
    n1412,
    n1401
  );


  xor
  g1473
  (
    n1529,
    n1484,
    n1401,
    n1392,
    n1490
  );


  nand
  g1474
  (
    n1504,
    n1407,
    n1490,
    n1417,
    n1418
  );


  nand
  g1475
  (
    n1538,
    n1400,
    n1397,
    n1414,
    n1491
  );


  xnor
  g1476
  (
    n1526,
    n1420,
    n1408,
    n1391
  );


  nand
  g1477
  (
    n1505,
    n1486,
    n1487,
    n1392,
    n1388
  );


  nand
  g1478
  (
    n1516,
    n1413,
    n1420,
    n1492,
    n1402
  );


  or
  g1479
  (
    n1518,
    n1411,
    n1481,
    n1491,
    n1393
  );


  nor
  g1480
  (
    n1501,
    n1482,
    n1485
  );


  xor
  g1481
  (
    n1531,
    n1416,
    n1488,
    n1412,
    n1398
  );


  xnor
  g1482
  (
    n1506,
    n1489,
    n1423,
    n1491,
    n1481
  );


  xnor
  g1483
  (
    n1527,
    n1417,
    n1421,
    n1422,
    n1426
  );


  or
  g1484
  (
    n1503,
    n1395,
    n1417,
    n1413,
    n1406
  );


  nand
  g1485
  (
    n1515,
    n1425,
    n1419,
    n1426,
    n1395
  );


  xor
  g1486
  (
    n1517,
    n1410,
    n1402,
    n1419,
    n1398
  );


  or
  g1487
  (
    n1544,
    n1483,
    n1421,
    n1492,
    n1404
  );


  xnor
  g1488
  (
    n1547,
    n1405,
    n1412,
    n1411,
    n1418
  );


  and
  g1489
  (
    n1546,
    n1483,
    n1425,
    n1396,
    n1410
  );


  xnor
  g1490
  (
    n1500,
    n1403,
    n1399,
    n1480,
    n1391
  );


  xnor
  g1491
  (
    n1502,
    n1486,
    n1392,
    n1412,
    n1485
  );


  or
  g1492
  (
    n1534,
    n1398,
    n1422,
    n1405,
    n1484
  );


  xor
  g1493
  (
    n1514,
    n1425,
    n1489,
    n1391,
    n1388
  );


  nor
  g1494
  (
    n1507,
    n1408,
    n1482,
    n1394,
    n1400
  );


  xor
  g1495
  (
    n1508,
    n1492,
    n1480,
    n1484,
    n1406
  );


  xnor
  g1496
  (
    n1523,
    n1396,
    n1425,
    n1400,
    n1390
  );


  xnor
  g1497
  (
    n1509,
    n1422,
    n1489,
    n1420,
    n1394
  );


  xnor
  g1498
  (
    n1545,
    n1417,
    n1492,
    n1423,
    n1406
  );


  nor
  g1499
  (
    n1537,
    n1486,
    n1396,
    n1415,
    n1407
  );


  or
  g1500
  (
    n1497,
    n1424,
    n1403,
    n1405,
    n1388
  );


  nand
  g1501
  (
    n1530,
    n1482,
    n1399,
    n1401,
    n1421
  );


  nand
  g1502
  (
    n1511,
    n1408,
    n1393,
    n1488,
    n1480
  );


  or
  g1503
  (
    n1521,
    n1410,
    n1393,
    n1414,
    n1394
  );


  nand
  g1504
  (
    n1512,
    n1397,
    n1483,
    n1399,
    n1391
  );


  nor
  g1505
  (
    n1524,
    n1393,
    n1414,
    n1399,
    n1423
  );


  xnor
  g1506
  (
    n1541,
    n1424,
    n1411,
    n1487,
    n1490
  );


  xor
  g1507
  (
    n1539,
    n1397,
    n1407,
    n1404,
    n1410
  );


  xnor
  g1508
  (
    n1533,
    n1403,
    n1398,
    n1411,
    n1390
  );


  xor
  g1509
  (
    n1510,
    n1419,
    n1409,
    n1392,
    n1488
  );


  nor
  g1510
  (
    n1520,
    n1390,
    n1404,
    n1389,
    n1409
  );


  nor
  g1511
  (
    n1513,
    n1490,
    n1407,
    n1395,
    n1493
  );


  and
  g1512
  (
    n1498,
    n1419,
    n1416,
    n1405,
    n1491
  );


  and
  g1513
  (
    n1525,
    n1422,
    n1484,
    n1485,
    n1418
  );


  and
  g1514
  (
    n1532,
    n1389,
    n1404,
    n1403,
    n1414
  );


  nor
  g1515
  (
    n1528,
    n1481,
    n1415,
    n1388,
    n1395
  );


  and
  g1516
  (
    n1582,
    n1432,
    n950,
    n1469,
    n1296
  );


  nor
  g1517
  (
    n1560,
    n1438,
    n948,
    n1493,
    n1508
  );


  nor
  g1518
  (
    n1585,
    n274,
    n1517,
    n1526,
    n949
  );


  xnor
  g1519
  (
    n1565,
    n1527,
    n271,
    n1497,
    n1520
  );


  nand
  g1520
  (
    n1562,
    n1441,
    n1435,
    n1439,
    n270
  );


  or
  g1521
  (
    n1594,
    n1288,
    n1547,
    n272,
    n1427
  );


  and
  g1522
  (
    n1584,
    n1430,
    n1364,
    n1516,
    n1284
  );


  nor
  g1523
  (
    n1579,
    n271,
    n1429,
    n273,
    n270
  );


  xor
  g1524
  (
    n1592,
    n1428,
    n1365,
    n1293,
    n1431
  );


  nand
  g1525
  (
    n1598,
    n950,
    n270,
    n1433,
    n1427
  );


  nand
  g1526
  (
    n1570,
    n1470,
    n1535,
    n1503,
    n1439
  );


  or
  g1527
  (
    n1596,
    n274,
    n1430,
    n1439,
    n1499
  );


  nor
  g1528
  (
    n1549,
    n1429,
    n1437,
    n271,
    n1442
  );


  xor
  g1529
  (
    n1587,
    n270,
    n1532,
    n949,
    n1443
  );


  or
  g1530
  (
    n1571,
    n1438,
    n1364,
    n79,
    n1510
  );


  or
  g1531
  (
    n1595,
    n1435,
    n952,
    n950,
    n1436
  );


  nand
  g1532
  (
    n1589,
    n1506,
    n1282,
    n1544,
    n1364
  );


  xnor
  g1533
  (
    n1553,
    n1285,
    n1430,
    n1438,
    n950
  );


  nor
  g1534
  (
    n1593,
    n1530,
    n1437,
    n1513,
    n1469
  );


  or
  g1535
  (
    n1550,
    n951,
    n1435,
    n949,
    n1363
  );


  or
  g1536
  (
    n1563,
    n1540,
    n1433,
    n1294,
    n1502
  );


  nand
  g1537
  (
    n1578,
    n1507,
    n1439,
    n275
  );


  nand
  g1538
  (
    n1559,
    n1546,
    n1519,
    n272,
    n1529
  );


  and
  g1539
  (
    n1590,
    n79,
    n1289,
    n1543,
    n951
  );


  nor
  g1540
  (
    n1574,
    n1469,
    n1434,
    n1426,
    n274
  );


  nand
  g1541
  (
    n1557,
    n1537,
    n1363,
    n1524,
    n1431
  );


  xnor
  g1542
  (
    n1575,
    n1435,
    n1433,
    n947,
    n1440
  );


  xnor
  g1543
  (
    n1558,
    n1545,
    n1470,
    n79
  );


  nor
  g1544
  (
    n1581,
    n1440,
    n1505,
    n273,
    n1427
  );


  xnor
  g1545
  (
    n1586,
    n1523,
    n1290,
    n1428,
    n1538
  );


  xnor
  g1546
  (
    n1597,
    n1522,
    n1500,
    n1365,
    n1350
  );


  and
  g1547
  (
    n1568,
    n1432,
    n1364,
    n1531,
    n1440
  );


  nand
  g1548
  (
    n1577,
    n1352,
    n272,
    n1436,
    n1509
  );


  or
  g1549
  (
    n1573,
    n1501,
    n1431,
    n949,
    n273
  );


  nor
  g1550
  (
    n1564,
    n1287,
    n1470,
    n1431,
    n1514
  );


  xor
  g1551
  (
    n1566,
    n1281,
    n1541,
    n1512,
    n1365
  );


  and
  g1552
  (
    n1555,
    n1441,
    n1428,
    n951
  );


  xor
  g1553
  (
    n1599,
    n1351,
    n1434,
    n1436,
    n1536
  );


  xor
  g1554
  (
    n1583,
    n276,
    n273,
    n1432,
    n1442
  );


  xnor
  g1555
  (
    n1556,
    n1441,
    n1493,
    n1427,
    n1498
  );


  xnor
  g1556
  (
    n1561,
    n1292,
    n1525,
    n1434,
    n1438
  );


  xnor
  g1557
  (
    n1569,
    n1286,
    n1440,
    n271,
    n1542
  );


  xor
  g1558
  (
    n1591,
    n948,
    n1295,
    n1548,
    n1518
  );


  or
  g1559
  (
    n1572,
    n1429,
    n1437,
    n948,
    n1494
  );


  nand
  g1560
  (
    n1551,
    n947,
    n1442,
    n274,
    n1430
  );


  xor
  g1561
  (
    n1552,
    n1349,
    n1442,
    n1429,
    n1493
  );


  nand
  g1562
  (
    n1580,
    n1534,
    n1515,
    n275,
    n78
  );


  or
  g1563
  (
    n1600,
    n272,
    n1432,
    n1437,
    n1521
  );


  and
  g1564
  (
    n1576,
    n1433,
    n948,
    n951,
    n1434
  );


  xnor
  g1565
  (
    n1554,
    n275,
    n1365,
    n1511,
    n1436
  );


  nor
  g1566
  (
    n1567,
    n1283,
    n79,
    n1504,
    n1528
  );


  or
  g1567
  (
    n1588,
    n1533,
    n1291,
    n1441,
    n1539
  );


  buf
  g1568
  (
    n1626,
    n1570
  );


  not
  g1569
  (
    n1672,
    n1575
  );


  buf
  g1570
  (
    n1794,
    n1593
  );


  buf
  g1571
  (
    n1690,
    n1551
  );


  buf
  g1572
  (
    n1748,
    n1586
  );


  buf
  g1573
  (
    n1782,
    n1559
  );


  buf
  g1574
  (
    n1606,
    n1553
  );


  not
  g1575
  (
    n1753,
    n1597
  );


  buf
  g1576
  (
    n1714,
    n1587
  );


  buf
  g1577
  (
    n1670,
    n1557
  );


  not
  g1578
  (
    n1668,
    n1571
  );


  not
  g1579
  (
    n1736,
    n1565
  );


  not
  g1580
  (
    n1603,
    n1579
  );


  buf
  g1581
  (
    n1750,
    n1560
  );


  not
  g1582
  (
    n1702,
    n1596
  );


  buf
  g1583
  (
    n1747,
    n1572
  );


  buf
  g1584
  (
    n1665,
    n1568
  );


  buf
  g1585
  (
    n1757,
    n1569
  );


  not
  g1586
  (
    n1646,
    n1575
  );


  buf
  g1587
  (
    n1725,
    n1597
  );


  not
  g1588
  (
    n1790,
    n1588
  );


  not
  g1589
  (
    n1696,
    n1579
  );


  not
  g1590
  (
    n1742,
    n1575
  );


  buf
  g1591
  (
    n1614,
    n1584
  );


  not
  g1592
  (
    n1629,
    n1554
  );


  not
  g1593
  (
    n1662,
    n1585
  );


  not
  g1594
  (
    n1632,
    n1558
  );


  not
  g1595
  (
    n1608,
    n1551
  );


  not
  g1596
  (
    n1723,
    n1479
  );


  not
  g1597
  (
    n1621,
    n1554
  );


  buf
  g1598
  (
    n1617,
    n1600
  );


  not
  g1599
  (
    n1688,
    n1567
  );


  buf
  g1600
  (
    n1805,
    n1476
  );


  buf
  g1601
  (
    n1631,
    n1479
  );


  buf
  g1602
  (
    n1795,
    n1566
  );


  buf
  g1603
  (
    n1746,
    n1592
  );


  buf
  g1604
  (
    n1800,
    n1562
  );


  not
  g1605
  (
    n1735,
    n1476
  );


  not
  g1606
  (
    n1673,
    n1600
  );


  buf
  g1607
  (
    n1604,
    n1560
  );


  buf
  g1608
  (
    n1793,
    n1561
  );


  buf
  g1609
  (
    n1726,
    n1577
  );


  buf
  g1610
  (
    n1781,
    n1598
  );


  not
  g1611
  (
    n1756,
    n1599
  );


  buf
  g1612
  (
    n1709,
    n1576
  );


  not
  g1613
  (
    n1738,
    n1580
  );


  buf
  g1614
  (
    n1787,
    n1571
  );


  buf
  g1615
  (
    n1745,
    n1583
  );


  buf
  g1616
  (
    n1763,
    n1590
  );


  buf
  g1617
  (
    n1715,
    n1584
  );


  buf
  g1618
  (
    n1737,
    n1552
  );


  not
  g1619
  (
    n1788,
    n1574
  );


  buf
  g1620
  (
    n1661,
    n1580
  );


  not
  g1621
  (
    n1642,
    n1478
  );


  buf
  g1622
  (
    n1773,
    n1557
  );


  not
  g1623
  (
    n1767,
    n1598
  );


  not
  g1624
  (
    n1752,
    n1569
  );


  not
  g1625
  (
    n1691,
    n1567
  );


  buf
  g1626
  (
    n1612,
    n1562
  );


  not
  g1627
  (
    n1644,
    n1552
  );


  not
  g1628
  (
    n1601,
    n1591
  );


  buf
  g1629
  (
    n1666,
    n1592
  );


  not
  g1630
  (
    n1679,
    n1550
  );


  buf
  g1631
  (
    n1743,
    n1589
  );


  not
  g1632
  (
    n1692,
    n1563
  );


  not
  g1633
  (
    n1807,
    n1549
  );


  not
  g1634
  (
    n1769,
    n1598
  );


  buf
  g1635
  (
    n1766,
    n1590
  );


  buf
  g1636
  (
    n1719,
    n1566
  );


  buf
  g1637
  (
    n1609,
    n1561
  );


  not
  g1638
  (
    n1799,
    n1561
  );


  not
  g1639
  (
    n1657,
    n1585
  );


  not
  g1640
  (
    n1768,
    n1597
  );


  not
  g1641
  (
    n1624,
    n1588
  );


  not
  g1642
  (
    n1703,
    n1574
  );


  not
  g1643
  (
    n1710,
    n1567
  );


  not
  g1644
  (
    n1754,
    n1572
  );


  buf
  g1645
  (
    n1681,
    n1564
  );


  buf
  g1646
  (
    n1802,
    n1596
  );


  buf
  g1647
  (
    n1722,
    n1589
  );


  buf
  g1648
  (
    n1732,
    n1569
  );


  not
  g1649
  (
    n1650,
    n1581
  );


  not
  g1650
  (
    n1651,
    n1558
  );


  buf
  g1651
  (
    n1783,
    n1564
  );


  buf
  g1652
  (
    n1697,
    n1551
  );


  buf
  g1653
  (
    n1700,
    n1576
  );


  buf
  g1654
  (
    n1640,
    n1557
  );


  not
  g1655
  (
    n1694,
    n1475
  );


  not
  g1656
  (
    n1716,
    n1573
  );


  buf
  g1657
  (
    n1731,
    n1568
  );


  buf
  g1658
  (
    n1762,
    n1577
  );


  buf
  g1659
  (
    n1619,
    n1567
  );


  not
  g1660
  (
    n1605,
    n1577
  );


  not
  g1661
  (
    n1647,
    n1556
  );


  not
  g1662
  (
    n1622,
    n1565
  );


  buf
  g1663
  (
    n1695,
    n1560
  );


  not
  g1664
  (
    n1680,
    n1478
  );


  not
  g1665
  (
    n1740,
    n1478
  );


  buf
  g1666
  (
    n1765,
    n1556
  );


  buf
  g1667
  (
    n1789,
    n1593
  );


  not
  g1668
  (
    n1777,
    n1582
  );


  buf
  g1669
  (
    n1685,
    n1560
  );


  not
  g1670
  (
    n1636,
    n1568
  );


  not
  g1671
  (
    n1620,
    n1599
  );


  not
  g1672
  (
    n1751,
    n1477
  );


  buf
  g1673
  (
    n1669,
    n1594
  );


  buf
  g1674
  (
    n1711,
    n1591
  );


  buf
  g1675
  (
    n1728,
    n1581
  );


  not
  g1676
  (
    n1659,
    n1600
  );


  not
  g1677
  (
    n1638,
    n1563
  );


  buf
  g1678
  (
    n1775,
    n1591
  );


  buf
  g1679
  (
    n1618,
    n1565
  );


  buf
  g1680
  (
    n1734,
    n1578
  );


  not
  g1681
  (
    n1804,
    n1593
  );


  not
  g1682
  (
    n1806,
    n1570
  );


  not
  g1683
  (
    n1607,
    n1558
  );


  buf
  g1684
  (
    n1671,
    n1551
  );


  buf
  g1685
  (
    n1796,
    n1595
  );


  not
  g1686
  (
    n1760,
    n1578
  );


  buf
  g1687
  (
    n1724,
    n1577
  );


  not
  g1688
  (
    n1705,
    n1591
  );


  not
  g1689
  (
    n1641,
    n1549
  );


  not
  g1690
  (
    n1625,
    n1479
  );


  buf
  g1691
  (
    n1759,
    n1574
  );


  not
  g1692
  (
    n1771,
    n1555
  );


  not
  g1693
  (
    n1602,
    n1571
  );


  not
  g1694
  (
    n1718,
    n1552
  );


  not
  g1695
  (
    n1613,
    n1477
  );


  not
  g1696
  (
    n1678,
    n1596
  );


  not
  g1697
  (
    n1634,
    n1593
  );


  not
  g1698
  (
    n1628,
    n1565
  );


  not
  g1699
  (
    n1676,
    n1581
  );


  not
  g1700
  (
    n1664,
    n1595
  );


  buf
  g1701
  (
    n1761,
    n1554
  );


  buf
  g1702
  (
    n1713,
    n1588
  );


  buf
  g1703
  (
    n1675,
    n1581
  );


  not
  g1704
  (
    n1656,
    n1582
  );


  buf
  g1705
  (
    n1798,
    n1562
  );


  buf
  g1706
  (
    n1610,
    n1475
  );


  buf
  g1707
  (
    n1635,
    n1573
  );


  buf
  g1708
  (
    n1730,
    n1552
  );


  buf
  g1709
  (
    n1706,
    n1590
  );


  not
  g1710
  (
    n1776,
    n1583
  );


  buf
  g1711
  (
    n1755,
    n1550
  );


  not
  g1712
  (
    n1654,
    n1600
  );


  not
  g1713
  (
    n1689,
    n1555
  );


  not
  g1714
  (
    n1683,
    n1597
  );


  not
  g1715
  (
    n1637,
    n1590
  );


  buf
  g1716
  (
    n1686,
    n1578
  );


  buf
  g1717
  (
    n1648,
    n1476
  );


  not
  g1718
  (
    n1627,
    n1575
  );


  buf
  g1719
  (
    n1733,
    n1587
  );


  buf
  g1720
  (
    n1785,
    n1477
  );


  buf
  g1721
  (
    n1797,
    n1599
  );


  buf
  g1722
  (
    n1630,
    n1550
  );


  buf
  g1723
  (
    n1687,
    n1475
  );


  buf
  g1724
  (
    n1720,
    n1569
  );


  buf
  g1725
  (
    n1643,
    n1563
  );


  not
  g1726
  (
    n1653,
    n1598
  );


  not
  g1727
  (
    n1698,
    n1579
  );


  not
  g1728
  (
    n1774,
    n1555
  );


  buf
  g1729
  (
    n1803,
    n1572
  );


  buf
  g1730
  (
    n1633,
    n1587
  );


  buf
  g1731
  (
    n1699,
    n1596
  );


  buf
  g1732
  (
    n1704,
    n1595
  );


  buf
  g1733
  (
    n1749,
    n1559
  );


  not
  g1734
  (
    n1727,
    n1586
  );


  buf
  g1735
  (
    n1663,
    n1566
  );


  buf
  g1736
  (
    n1615,
    n1561
  );


  buf
  g1737
  (
    n1729,
    n1583
  );


  not
  g1738
  (
    n1721,
    n1573
  );


  buf
  g1739
  (
    n1791,
    n1564
  );


  not
  g1740
  (
    n1712,
    n1579
  );


  not
  g1741
  (
    n1707,
    n1571
  );


  not
  g1742
  (
    n1677,
    n1586
  );


  not
  g1743
  (
    n1652,
    n1554
  );


  buf
  g1744
  (
    n1764,
    n1568
  );


  not
  g1745
  (
    n1779,
    n1559
  );


  not
  g1746
  (
    n1684,
    n1594
  );


  not
  g1747
  (
    n1801,
    n1595
  );


  not
  g1748
  (
    n1772,
    n1576
  );


  buf
  g1749
  (
    n1744,
    n1564
  );


  buf
  g1750
  (
    n1616,
    n1553
  );


  not
  g1751
  (
    n1649,
    n1563
  );


  buf
  g1752
  (
    n1784,
    n1588
  );


  buf
  g1753
  (
    n1778,
    n1592
  );


  not
  g1754
  (
    n1758,
    n1553
  );


  buf
  g1755
  (
    n1739,
    n1592
  );


  buf
  g1756
  (
    n1658,
    n1599
  );


  buf
  g1757
  (
    n1682,
    n1562
  );


  buf
  g1758
  (
    n1741,
    n1570
  );


  not
  g1759
  (
    n1693,
    n1594
  );


  not
  g1760
  (
    n1717,
    n1550
  );


  not
  g1761
  (
    n1780,
    n1585
  );


  buf
  g1762
  (
    n1611,
    n1589
  );


  not
  g1763
  (
    n1667,
    n1478
  );


  not
  g1764
  (
    n1808,
    n1584
  );


  buf
  g1765
  (
    n1792,
    n1589
  );


  not
  g1766
  (
    n1701,
    n1576
  );


  not
  g1767
  (
    n1623,
    n1574
  );


  not
  g1768
  (
    n1786,
    n1479
  );


  or
  g1769
  (
    n1645,
    n1582,
    n1573,
    n1557
  );


  xor
  g1770
  (
    n1674,
    n1558,
    n1475,
    n1559,
    n1549
  );


  and
  g1771
  (
    n1639,
    n1549,
    n1584,
    n1594,
    n1578
  );


  nor
  g1772
  (
    n1708,
    n1476,
    n1587,
    n1585,
    n1580
  );


  and
  g1773
  (
    n1660,
    n1582,
    n1583,
    n1566,
    n1570
  );


  xor
  g1774
  (
    n1655,
    n1553,
    n1555,
    n1580,
    n1572
  );


  nand
  g1775
  (
    n1770,
    n1477,
    n1556,
    n1586
  );


  buf
  g1776
  (
    n1853,
    n1650
  );


  not
  g1777
  (
    n2134,
    n1646
  );


  buf
  g1778
  (
    n2092,
    n1715
  );


  not
  g1779
  (
    n2375,
    n1695
  );


  not
  g1780
  (
    n2244,
    n1668
  );


  not
  g1781
  (
    n2069,
    n1693
  );


  not
  g1782
  (
    n2296,
    n1726
  );


  buf
  g1783
  (
    n1887,
    n1792
  );


  buf
  g1784
  (
    n2107,
    n1763
  );


  buf
  g1785
  (
    n1996,
    n1730
  );


  buf
  g1786
  (
    n2185,
    n1778
  );


  not
  g1787
  (
    n2288,
    n1729
  );


  not
  g1788
  (
    n1925,
    n1495
  );


  buf
  g1789
  (
    n2114,
    n1728
  );


  not
  g1790
  (
    n1992,
    n1723
  );


  not
  g1791
  (
    n2062,
    n1684
  );


  not
  g1792
  (
    n2262,
    n1714
  );


  not
  g1793
  (
    n1895,
    n1673
  );


  buf
  g1794
  (
    n1972,
    n1763
  );


  not
  g1795
  (
    n2111,
    n1632
  );


  not
  g1796
  (
    n1981,
    n1671
  );


  not
  g1797
  (
    n2106,
    n1603
  );


  buf
  g1798
  (
    n1826,
    n1776
  );


  buf
  g1799
  (
    n2089,
    n1696
  );


  buf
  g1800
  (
    n1913,
    n1678
  );


  not
  g1801
  (
    n1933,
    n1737
  );


  not
  g1802
  (
    n2316,
    n1794
  );


  buf
  g1803
  (
    n2327,
    n1637
  );


  not
  g1804
  (
    n2266,
    n1658
  );


  not
  g1805
  (
    n2036,
    n1715
  );


  not
  g1806
  (
    n2238,
    n1629
  );


  not
  g1807
  (
    n2030,
    n1724
  );


  buf
  g1808
  (
    n2359,
    n1807
  );


  buf
  g1809
  (
    n2142,
    n1724
  );


  not
  g1810
  (
    n2085,
    n1749
  );


  not
  g1811
  (
    n2053,
    n1750
  );


  not
  g1812
  (
    n2306,
    n1638
  );


  not
  g1813
  (
    n2381,
    n1665
  );


  buf
  g1814
  (
    n1898,
    n1682
  );


  buf
  g1815
  (
    n2127,
    n1746
  );


  buf
  g1816
  (
    n2215,
    n1735
  );


  not
  g1817
  (
    n1849,
    n1644
  );


  buf
  g1818
  (
    n1980,
    n1705
  );


  not
  g1819
  (
    n2105,
    n1746
  );


  buf
  g1820
  (
    n2044,
    n1792
  );


  not
  g1821
  (
    n2257,
    n1655
  );


  not
  g1822
  (
    n2251,
    n1608
  );


  buf
  g1823
  (
    n1984,
    n1724
  );


  buf
  g1824
  (
    n2309,
    n1748
  );


  buf
  g1825
  (
    n2050,
    n1623
  );


  buf
  g1826
  (
    n2035,
    n1748
  );


  buf
  g1827
  (
    n2122,
    n1767
  );


  buf
  g1828
  (
    n2297,
    n1694
  );


  not
  g1829
  (
    n1985,
    n1603
  );


  buf
  g1830
  (
    n2131,
    n1608
  );


  not
  g1831
  (
    n2322,
    n1667
  );


  not
  g1832
  (
    n1882,
    n1661
  );


  not
  g1833
  (
    n1840,
    n1798
  );


  buf
  g1834
  (
    n2038,
    n1806
  );


  buf
  g1835
  (
    n2292,
    n1629
  );


  buf
  g1836
  (
    n2370,
    n1785
  );


  buf
  g1837
  (
    n2263,
    n1716
  );


  not
  g1838
  (
    n2135,
    n1627
  );


  not
  g1839
  (
    n2249,
    n1745
  );


  not
  g1840
  (
    n2016,
    n1634
  );


  not
  g1841
  (
    n2311,
    n1640
  );


  not
  g1842
  (
    n2214,
    n1764
  );


  buf
  g1843
  (
    n2285,
    n1690
  );


  not
  g1844
  (
    n2002,
    n1791
  );


  not
  g1845
  (
    n1909,
    n1746
  );


  not
  g1846
  (
    n1944,
    n1770
  );


  buf
  g1847
  (
    n1920,
    n1736
  );


  buf
  g1848
  (
    n2197,
    n1783
  );


  not
  g1849
  (
    n2243,
    n1646
  );


  buf
  g1850
  (
    n2178,
    n1754
  );


  buf
  g1851
  (
    n2155,
    n1770
  );


  buf
  g1852
  (
    n2293,
    n1753
  );


  buf
  g1853
  (
    n1934,
    n1677
  );


  buf
  g1854
  (
    n1941,
    n1778
  );


  not
  g1855
  (
    n2174,
    n1715
  );


  buf
  g1856
  (
    n1998,
    n1620
  );


  not
  g1857
  (
    n2103,
    n1719
  );


  not
  g1858
  (
    n1891,
    n1647
  );


  buf
  g1859
  (
    n1879,
    n1666
  );


  not
  g1860
  (
    n2290,
    n1756
  );


  buf
  g1861
  (
    n2113,
    n1625
  );


  buf
  g1862
  (
    n2312,
    n1621
  );


  buf
  g1863
  (
    n2136,
    n1695
  );


  not
  g1864
  (
    n2310,
    n1685
  );


  buf
  g1865
  (
    n1931,
    n1777
  );


  not
  g1866
  (
    n1819,
    n1611
  );


  buf
  g1867
  (
    n1923,
    n1621
  );


  buf
  g1868
  (
    n1885,
    n1793
  );


  buf
  g1869
  (
    n2137,
    n1772
  );


  buf
  g1870
  (
    n1912,
    n1755
  );


  not
  g1871
  (
    n1864,
    n1673
  );


  not
  g1872
  (
    n2330,
    n1709
  );


  not
  g1873
  (
    n2274,
    n1640
  );


  buf
  g1874
  (
    n2203,
    n1643
  );


  not
  g1875
  (
    n2331,
    n1757
  );


  buf
  g1876
  (
    n1815,
    n1804
  );


  not
  g1877
  (
    n2216,
    n1638
  );


  buf
  g1878
  (
    n1971,
    n1725
  );


  buf
  g1879
  (
    n2004,
    n1663
  );


  not
  g1880
  (
    n2321,
    n1787
  );


  not
  g1881
  (
    n2011,
    n1751
  );


  not
  g1882
  (
    n2065,
    n1681
  );


  buf
  g1883
  (
    n1940,
    n1607
  );


  buf
  g1884
  (
    n2273,
    n1667
  );


  not
  g1885
  (
    n2230,
    n1765
  );


  not
  g1886
  (
    n2098,
    n1495
  );


  buf
  g1887
  (
    n2080,
    n1776
  );


  not
  g1888
  (
    n1862,
    n1606
  );


  buf
  g1889
  (
    n1818,
    n1649
  );


  buf
  g1890
  (
    n1926,
    n1631
  );


  not
  g1891
  (
    n2032,
    n1774
  );


  buf
  g1892
  (
    n1850,
    n1765
  );


  not
  g1893
  (
    n2110,
    n1622
  );


  not
  g1894
  (
    n1869,
    n1784
  );


  not
  g1895
  (
    n1811,
    n1603
  );


  buf
  g1896
  (
    n1835,
    n1684
  );


  buf
  g1897
  (
    n1861,
    n1768
  );


  buf
  g1898
  (
    n2099,
    n1779
  );


  not
  g1899
  (
    n2350,
    n1712
  );


  not
  g1900
  (
    n2094,
    n1618
  );


  not
  g1901
  (
    n2188,
    n1619
  );


  not
  g1902
  (
    n1969,
    n1750
  );


  buf
  g1903
  (
    n1859,
    n1792
  );


  not
  g1904
  (
    n2121,
    n1679
  );


  buf
  g1905
  (
    n2328,
    n1665
  );


  not
  g1906
  (
    n2169,
    n1699
  );


  buf
  g1907
  (
    n2353,
    n1793
  );


  buf
  g1908
  (
    n1899,
    n1658
  );


  buf
  g1909
  (
    n1883,
    n1762
  );


  not
  g1910
  (
    n1950,
    n1639
  );


  buf
  g1911
  (
    n1884,
    n1617
  );


  buf
  g1912
  (
    n2366,
    n1760
  );


  buf
  g1913
  (
    n2100,
    n1660
  );


  buf
  g1914
  (
    n2138,
    n1619
  );


  buf
  g1915
  (
    n2021,
    n1639
  );


  not
  g1916
  (
    n2252,
    n1709
  );


  not
  g1917
  (
    n2338,
    n1655
  );


  not
  g1918
  (
    n2160,
    n1625
  );


  buf
  g1919
  (
    n2031,
    n1603
  );


  not
  g1920
  (
    n1994,
    n1732
  );


  not
  g1921
  (
    n2242,
    n1723
  );


  not
  g1922
  (
    n2182,
    n1737
  );


  buf
  g1923
  (
    n2084,
    n1721
  );


  not
  g1924
  (
    n2347,
    n1610
  );


  not
  g1925
  (
    n1823,
    n1762
  );


  buf
  g1926
  (
    n2161,
    n1674
  );


  not
  g1927
  (
    n1977,
    n1722
  );


  buf
  g1928
  (
    n2170,
    n1790
  );


  not
  g1929
  (
    n2333,
    n1636
  );


  not
  g1930
  (
    n1962,
    n1628
  );


  buf
  g1931
  (
    n1852,
    n1787
  );


  buf
  g1932
  (
    n1890,
    n1768
  );


  not
  g1933
  (
    n2248,
    n1686
  );


  not
  g1934
  (
    n2298,
    n1673
  );


  not
  g1935
  (
    n2097,
    n1648
  );


  buf
  g1936
  (
    n1902,
    n1651
  );


  buf
  g1937
  (
    n2163,
    n1795
  );


  buf
  g1938
  (
    n2219,
    n1777
  );


  not
  g1939
  (
    n2074,
    n1741
  );


  not
  g1940
  (
    n1824,
    n1792
  );


  not
  g1941
  (
    n2237,
    n1615
  );


  not
  g1942
  (
    n2229,
    n1781
  );


  buf
  g1943
  (
    n2010,
    n1715
  );


  not
  g1944
  (
    n2042,
    n1782
  );


  not
  g1945
  (
    n2017,
    n1732
  );


  buf
  g1946
  (
    n2264,
    n1707
  );


  not
  g1947
  (
    n2102,
    n1683
  );


  not
  g1948
  (
    n2341,
    n1741
  );


  not
  g1949
  (
    n1841,
    n1666
  );


  not
  g1950
  (
    n1905,
    n1689
  );


  buf
  g1951
  (
    n2019,
    n1602
  );


  buf
  g1952
  (
    n1914,
    n1743
  );


  buf
  g1953
  (
    n2172,
    n1730
  );


  not
  g1954
  (
    n2192,
    n1711
  );


  not
  g1955
  (
    n1903,
    n1727
  );


  not
  g1956
  (
    n2008,
    n1720
  );


  not
  g1957
  (
    n2077,
    n1663
  );


  not
  g1958
  (
    n1873,
    n1602
  );


  not
  g1959
  (
    n2014,
    n1636
  );


  buf
  g1960
  (
    n2147,
    n1801
  );


  buf
  g1961
  (
    n1911,
    n1776
  );


  buf
  g1962
  (
    n1904,
    n1684
  );


  buf
  g1963
  (
    n2057,
    n1655
  );


  not
  g1964
  (
    n1893,
    n1739
  );


  not
  g1965
  (
    n2278,
    n1734
  );


  not
  g1966
  (
    n2360,
    n1614
  );


  buf
  g1967
  (
    n2261,
    n1801
  );


  not
  g1968
  (
    n2159,
    n1601
  );


  buf
  g1969
  (
    n2104,
    n1806
  );


  not
  g1970
  (
    n1888,
    n1699
  );


  buf
  g1971
  (
    n2209,
    n1652
  );


  buf
  g1972
  (
    n2168,
    n1670
  );


  buf
  g1973
  (
    n2270,
    n1678
  );


  not
  g1974
  (
    n2046,
    n1648
  );


  not
  g1975
  (
    n2294,
    n1765
  );


  buf
  g1976
  (
    n2060,
    n1702
  );


  buf
  g1977
  (
    n1810,
    n1691
  );


  not
  g1978
  (
    n1922,
    n1620
  );


  buf
  g1979
  (
    n2139,
    n1622
  );


  not
  g1980
  (
    n2018,
    n1788
  );


  not
  g1981
  (
    n1851,
    n1766
  );


  not
  g1982
  (
    n1907,
    n1664
  );


  buf
  g1983
  (
    n2207,
    n1780
  );


  not
  g1984
  (
    n1865,
    n1738
  );


  buf
  g1985
  (
    n2167,
    n1760
  );


  buf
  g1986
  (
    n1866,
    n1775
  );


  buf
  g1987
  (
    n2211,
    n1805
  );


  not
  g1988
  (
    n2049,
    n1644
  );


  not
  g1989
  (
    n2090,
    n1687
  );


  not
  g1990
  (
    n1896,
    n1721
  );


  not
  g1991
  (
    n2007,
    n1642
  );


  buf
  g1992
  (
    n2256,
    n1781
  );


  not
  g1993
  (
    n1827,
    n1706
  );


  buf
  g1994
  (
    n2279,
    n1743
  );


  buf
  g1995
  (
    n2189,
    n1797
  );


  not
  g1996
  (
    n2344,
    n1771
  );


  buf
  g1997
  (
    n1820,
    n1655
  );


  buf
  g1998
  (
    n2096,
    n1677
  );


  not
  g1999
  (
    n2054,
    n1646
  );


  not
  g2000
  (
    n2156,
    n1656
  );


  buf
  g2001
  (
    n2283,
    n1675
  );


  buf
  g2002
  (
    n2368,
    n1613
  );


  buf
  g2003
  (
    n2003,
    n1728
  );


  not
  g2004
  (
    n1863,
    n1768
  );


  buf
  g2005
  (
    n2371,
    n1617
  );


  buf
  g2006
  (
    n2220,
    n1747
  );


  not
  g2007
  (
    n2227,
    n1748
  );


  not
  g2008
  (
    n2233,
    n1656
  );


  not
  g2009
  (
    n2115,
    n1728
  );


  not
  g2010
  (
    n1976,
    n1630
  );


  not
  g2011
  (
    n2040,
    n1748
  );


  buf
  g2012
  (
    n2091,
    n1662
  );


  buf
  g2013
  (
    n2141,
    n1691
  );


  buf
  g2014
  (
    n1844,
    n1745
  );


  not
  g2015
  (
    n2145,
    n1807
  );


  not
  g2016
  (
    n2171,
    n1740
  );


  buf
  g2017
  (
    n2028,
    n1758
  );


  buf
  g2018
  (
    n2340,
    n1785
  );


  not
  g2019
  (
    n1966,
    n1767
  );


  not
  g2020
  (
    n2128,
    n1799
  );


  buf
  g2021
  (
    n2276,
    n1649
  );


  not
  g2022
  (
    n1817,
    n1494
  );


  not
  g2023
  (
    n2346,
    n1646
  );


  not
  g2024
  (
    n1886,
    n1724
  );


  not
  g2025
  (
    n2314,
    n1644
  );


  not
  g2026
  (
    n1952,
    n1704
  );


  buf
  g2027
  (
    n2177,
    n1806
  );


  not
  g2028
  (
    n2058,
    n1612
  );


  buf
  g2029
  (
    n1943,
    n1604
  );


  not
  g2030
  (
    n2152,
    n1774
  );


  buf
  g2031
  (
    n1982,
    n1638
  );


  buf
  g2032
  (
    n2223,
    n1788
  );


  buf
  g2033
  (
    n1834,
    n1691
  );


  buf
  g2034
  (
    n2006,
    n1756
  );


  buf
  g2035
  (
    n1878,
    n1690
  );


  buf
  g2036
  (
    n2318,
    n1668
  );


  buf
  g2037
  (
    n1937,
    n1690
  );


  buf
  g2038
  (
    n2076,
    n1669
  );


  not
  g2039
  (
    n2175,
    n1674
  );


  buf
  g2040
  (
    n2225,
    n1672
  );


  not
  g2041
  (
    n1857,
    n1776
  );


  not
  g2042
  (
    n1874,
    n1681
  );


  buf
  g2043
  (
    n2180,
    n1630
  );


  not
  g2044
  (
    n1845,
    n1751
  );


  buf
  g2045
  (
    n2260,
    n1701
  );


  buf
  g2046
  (
    n1870,
    n1624
  );


  not
  g2047
  (
    n1846,
    n1628
  );


  buf
  g2048
  (
    n1921,
    n1742
  );


  buf
  g2049
  (
    n2315,
    n1789
  );


  buf
  g2050
  (
    n2123,
    n1636
  );


  not
  g2051
  (
    n2253,
    n1761
  );


  not
  g2052
  (
    n2001,
    n1752
  );


  buf
  g2053
  (
    n2281,
    n1773
  );


  not
  g2054
  (
    n2027,
    n1781
  );


  buf
  g2055
  (
    n1954,
    n1630
  );


  not
  g2056
  (
    n2358,
    n1758
  );


  buf
  g2057
  (
    n1945,
    n1794
  );


  not
  g2058
  (
    n2117,
    n1711
  );


  buf
  g2059
  (
    n1928,
    n1772
  );


  buf
  g2060
  (
    n1961,
    n1676
  );


  buf
  g2061
  (
    n2034,
    n1804
  );


  buf
  g2062
  (
    n2070,
    n1714
  );


  not
  g2063
  (
    n2047,
    n1685
  );


  buf
  g2064
  (
    n2342,
    n1659
  );


  buf
  g2065
  (
    n2277,
    n1606
  );


  buf
  g2066
  (
    n2250,
    n1641
  );


  buf
  g2067
  (
    n1831,
    n1606
  );


  not
  g2068
  (
    n1892,
    n1788
  );


  not
  g2069
  (
    n2148,
    n1805
  );


  not
  g2070
  (
    n2164,
    n1726
  );


  not
  g2071
  (
    n1848,
    n1667
  );


  not
  g2072
  (
    n2267,
    n1619
  );


  not
  g2073
  (
    n2140,
    n1766
  );


  buf
  g2074
  (
    n2205,
    n1673
  );


  not
  g2075
  (
    n2324,
    n1752
  );


  buf
  g2076
  (
    n2093,
    n1624
  );


  buf
  g2077
  (
    n1986,
    n1743
  );


  not
  g2078
  (
    n2120,
    n1694
  );


  buf
  g2079
  (
    n1953,
    n1689
  );


  buf
  g2080
  (
    n1894,
    n1747
  );


  buf
  g2081
  (
    n1935,
    n1632
  );


  buf
  g2082
  (
    n2023,
    n1664
  );


  buf
  g2083
  (
    n2087,
    n1769
  );


  not
  g2084
  (
    n1919,
    n1754
  );


  buf
  g2085
  (
    n2239,
    n1649
  );


  not
  g2086
  (
    n2146,
    n1635
  );


  not
  g2087
  (
    n2291,
    n1702
  );


  not
  g2088
  (
    n2334,
    n1637
  );


  buf
  g2089
  (
    n2116,
    n1651
  );


  buf
  g2090
  (
    n2025,
    n1612
  );


  not
  g2091
  (
    n2201,
    n1733
  );


  not
  g2092
  (
    n2247,
    n1651
  );


  buf
  g2093
  (
    n2235,
    n1744
  );


  buf
  g2094
  (
    n1938,
    n1756
  );


  not
  g2095
  (
    n2063,
    n1706
  );


  not
  g2096
  (
    n2218,
    n1722
  );


  buf
  g2097
  (
    n2165,
    n1610
  );


  not
  g2098
  (
    n1814,
    n1763
  );


  buf
  g2099
  (
    n1897,
    n1688
  );


  buf
  g2100
  (
    n2191,
    n1761
  );


  not
  g2101
  (
    n1880,
    n1602
  );


  buf
  g2102
  (
    n1837,
    n1800
  );


  not
  g2103
  (
    n1833,
    n1767
  );


  buf
  g2104
  (
    n2039,
    n1620
  );


  not
  g2105
  (
    n2304,
    n1601
  );


  buf
  g2106
  (
    n2383,
    n1739
  );


  not
  g2107
  (
    n2108,
    n1648
  );


  buf
  g2108
  (
    n1990,
    n1800
  );


  buf
  g2109
  (
    n2020,
    n1708
  );


  not
  g2110
  (
    n1989,
    n1678
  );


  not
  g2111
  (
    n2269,
    n1757
  );


  buf
  g2112
  (
    n2012,
    n1803
  );


  not
  g2113
  (
    n1936,
    n1666
  );


  not
  g2114
  (
    n2367,
    n1802
  );


  buf
  g2115
  (
    n1918,
    n1641
  );


  not
  g2116
  (
    n2061,
    n1749
  );


  not
  g2117
  (
    n2086,
    n1745
  );


  buf
  g2118
  (
    n2119,
    n1678
  );


  buf
  g2119
  (
    n1963,
    n1626
  );


  not
  g2120
  (
    n1917,
    n1618
  );


  not
  g2121
  (
    n2326,
    n1624
  );


  buf
  g2122
  (
    n1856,
    n1744
  );


  not
  g2123
  (
    n1939,
    n1789
  );


  not
  g2124
  (
    n2271,
    n1706
  );


  buf
  g2125
  (
    n1958,
    n1746
  );


  buf
  g2126
  (
    n1974,
    n1793
  );


  buf
  g2127
  (
    n2037,
    n1659
  );


  buf
  g2128
  (
    n2213,
    n1738
  );


  not
  g2129
  (
    n2287,
    n1623
  );


  not
  g2130
  (
    n2190,
    n1736
  );


  not
  g2131
  (
    n2289,
    n1616
  );


  not
  g2132
  (
    n2362,
    n1719
  );


  buf
  g2133
  (
    n2354,
    n1791
  );


  buf
  g2134
  (
    n1900,
    n1606
  );


  buf
  g2135
  (
    n1983,
    n1692
  );


  buf
  g2136
  (
    n1999,
    n1679
  );


  not
  g2137
  (
    n1838,
    n1687
  );


  buf
  g2138
  (
    n2335,
    n1726
  );


  not
  g2139
  (
    n1942,
    n1692
  );


  not
  g2140
  (
    n2282,
    n1689
  );


  not
  g2141
  (
    n2343,
    n1702
  );


  buf
  g2142
  (
    n1965,
    n1727
  );


  not
  g2143
  (
    n2373,
    n1779
  );


  not
  g2144
  (
    n1924,
    n1714
  );


  not
  g2145
  (
    n1951,
    n1645
  );


  buf
  g2146
  (
    n2319,
    n1791
  );


  buf
  g2147
  (
    n2272,
    n1798
  );


  buf
  g2148
  (
    n2206,
    n1798
  );


  not
  g2149
  (
    n2355,
    n1607
  );


  buf
  g2150
  (
    n2245,
    n1763
  );


  not
  g2151
  (
    n2382,
    n1676
  );


  not
  g2152
  (
    n1988,
    n1668
  );


  buf
  g2153
  (
    n1855,
    n1716
  );


  buf
  g2154
  (
    n2313,
    n1661
  );


  buf
  g2155
  (
    n2064,
    n1731
  );


  not
  g2156
  (
    n2345,
    n1650
  );


  not
  g2157
  (
    n2051,
    n1657
  );


  not
  g2158
  (
    n1967,
    n1654
  );


  not
  g2159
  (
    n1872,
    n1682
  );


  buf
  g2160
  (
    n2194,
    n1680
  );


  buf
  g2161
  (
    n2236,
    n1663
  );


  not
  g2162
  (
    n2079,
    n1657
  );


  not
  g2163
  (
    n1847,
    n1701
  );


  not
  g2164
  (
    n2153,
    n1708
  );


  not
  g2165
  (
    n2255,
    n1712
  );


  not
  g2166
  (
    n2348,
    n1642
  );


  buf
  g2167
  (
    n2339,
    n1796
  );


  not
  g2168
  (
    n2082,
    n1604
  );


  not
  g2169
  (
    n1816,
    n1679
  );


  not
  g2170
  (
    n2379,
    n1605
  );


  buf
  g2171
  (
    n2055,
    n1653
  );


  buf
  g2172
  (
    n1927,
    n1667
  );


  buf
  g2173
  (
    n2176,
    n1635
  );


  not
  g2174
  (
    n2222,
    n1695
  );


  not
  g2175
  (
    n2349,
    n1697
  );


  not
  g2176
  (
    n2217,
    n1618
  );


  not
  g2177
  (
    n2068,
    n1685
  );


  not
  g2178
  (
    n2181,
    n1764
  );


  not
  g2179
  (
    n2284,
    n1773
  );


  not
  g2180
  (
    n1829,
    n1607
  );


  buf
  g2181
  (
    n2200,
    n1634
  );


  buf
  g2182
  (
    n1975,
    n1656
  );


  buf
  g2183
  (
    n2369,
    n1752
  );


  buf
  g2184
  (
    n2000,
    n1710
  );


  not
  g2185
  (
    n2024,
    n1664
  );


  not
  g2186
  (
    n2081,
    n1654
  );


  buf
  g2187
  (
    n2118,
    n1783
  );


  not
  g2188
  (
    n1906,
    n1633
  );


  buf
  g2189
  (
    n1868,
    n1643
  );


  buf
  g2190
  (
    n1915,
    n1669
  );


  not
  g2191
  (
    n1860,
    n1725
  );


  buf
  g2192
  (
    n1991,
    n1604
  );


  not
  g2193
  (
    n2124,
    n1653
  );


  not
  g2194
  (
    n1959,
    n1660
  );


  buf
  g2195
  (
    n1960,
    n1784
  );


  not
  g2196
  (
    n2212,
    n1801
  );


  buf
  g2197
  (
    n2356,
    n1802
  );


  buf
  g2198
  (
    n1987,
    n1750
  );


  not
  g2199
  (
    n1875,
    n1707
  );


  buf
  g2200
  (
    n1854,
    n1622
  );


  buf
  g2201
  (
    n1955,
    n1613
  );


  not
  g2202
  (
    n2022,
    n1637
  );


  buf
  g2203
  (
    n2363,
    n1742
  );


  not
  g2204
  (
    n2158,
    n1607
  );


  not
  g2205
  (
    n1948,
    n1722
  );


  not
  g2206
  (
    n1947,
    n1615
  );


  buf
  g2207
  (
    n1932,
    n1743
  );


  buf
  g2208
  (
    n1809,
    n1711
  );


  not
  g2209
  (
    n1901,
    n1622
  );


  not
  g2210
  (
    n2029,
    n1784
  );


  not
  g2211
  (
    n1949,
    n1777
  );


  not
  g2212
  (
    n2378,
    n1774
  );


  buf
  g2213
  (
    n2320,
    n1718
  );


  not
  g2214
  (
    n2280,
    n1796
  );


  buf
  g2215
  (
    n2196,
    n1632
  );


  not
  g2216
  (
    n1889,
    n1771
  );


  buf
  g2217
  (
    n2073,
    n1740
  );


  not
  g2218
  (
    n2183,
    n1609
  );


  buf
  g2219
  (
    n1970,
    n1787
  );


  buf
  g2220
  (
    n1842,
    n1757
  );


  not
  g2221
  (
    n1836,
    n1681
  );


  buf
  g2222
  (
    n2202,
    n1762
  );


  not
  g2223
  (
    n1916,
    n1658
  );


  buf
  g2224
  (
    n2009,
    n1627
  );


  buf
  g2225
  (
    n1964,
    n1705
  );


  not
  g2226
  (
    n2208,
    n1601
  );


  buf
  g2227
  (
    n2224,
    n1616
  );


  not
  g2228
  (
    n1973,
    n1778
  );


  not
  g2229
  (
    n2275,
    n1697
  );


  not
  g2230
  (
    n1979,
    n1680
  );


  not
  g2231
  (
    n2286,
    n1728
  );


  not
  g2232
  (
    n2240,
    n1674
  );


  not
  g2233
  (
    n2336,
    n1675
  );


  not
  g2234
  (
    n1812,
    n1719
  );


  not
  g2235
  (
    n2154,
    n1713
  );


  buf
  g2236
  (
    n1968,
    n1739
  );


  not
  g2237
  (
    n2365,
    n1796
  );


  buf
  g2238
  (
    n2337,
    n1789
  );


  not
  g2239
  (
    n2048,
    n1717
  );


  buf
  g2240
  (
    n2162,
    n1608
  );


  buf
  g2241
  (
    n2083,
    n1770
  );


  not
  g2242
  (
    n1858,
    n1804
  );


  buf
  g2243
  (
    n2072,
    n1692
  );


  buf
  g2244
  (
    n2013,
    n1744
  );


  not
  g2245
  (
    n1821,
    n1720
  );


  buf
  g2246
  (
    n2317,
    n1805
  );


  not
  g2247
  (
    n2043,
    n1790
  );


  not
  g2248
  (
    n2268,
    n1775
  );


  not
  g2249
  (
    n2130,
    n1786
  );


  buf
  g2250
  (
    n1813,
    n1704
  );


  not
  g2251
  (
    n2352,
    n1621
  );


  not
  g2252
  (
    n2198,
    n1664
  );


  not
  g2253
  (
    n1871,
    n1653
  );


  not
  g2254
  (
    n2125,
    n1722
  );


  buf
  g2255
  (
    n2143,
    n1653
  );


  not
  g2256
  (
    n2033,
    n1617
  );


  not
  g2257
  (
    n2151,
    n1702
  );


  buf
  g2258
  (
    n2150,
    n1761
  );


  not
  g2259
  (
    n2231,
    n1623
  );


  not
  g2260
  (
    n2026,
    n1712
  );


  buf
  g2261
  (
    n2308,
    n1703
  );


  buf
  g2262
  (
    n2210,
    n1785
  );


  xnor
  g2263
  (
    n2259,
    n1609,
    n1613,
    n1684,
    n1805
  );


  nand
  g2264
  (
    n2015,
    n1700,
    n1707,
    n1494,
    n1657
  );


  and
  g2265
  (
    n2364,
    n1780,
    n1495,
    n1726,
    n1803
  );


  or
  g2266
  (
    n2246,
    n1661,
    n1688,
    n1654
  );


  and
  g2267
  (
    n2075,
    n1753,
    n1786,
    n1740,
    n1700
  );


  xor
  g2268
  (
    n2195,
    n1734,
    n1671,
    n1619,
    n1700
  );


  nand
  g2269
  (
    n2301,
    n1708,
    n1808,
    n1755,
    n1769
  );


  nor
  g2270
  (
    n2193,
    n1808,
    n1662,
    n1645,
    n1677
  );


  and
  g2271
  (
    n2041,
    n1716,
    n1672,
    n1723,
    n1804
  );


  or
  g2272
  (
    n2173,
    n1638,
    n1808,
    n1701,
    n1794
  );


  xnor
  g2273
  (
    n2095,
    n1698,
    n1627,
    n1799,
    n1682
  );


  nand
  g2274
  (
    n2234,
    n1797,
    n1758,
    n1775,
    n1676
  );


  xor
  g2275
  (
    n2226,
    n1759,
    n1745,
    n1741,
    n1610
  );


  nand
  g2276
  (
    n2052,
    n1661,
    n1760,
    n1685,
    n1624
  );


  xor
  g2277
  (
    n2241,
    n1742,
    n1634,
    n1635,
    n1800
  );


  xnor
  g2278
  (
    n2179,
    n1688,
    n1733,
    n1693,
    n1658
  );


  and
  g2279
  (
    n2299,
    n1633,
    n1790,
    n1800,
    n1629
  );


  xor
  g2280
  (
    n2129,
    n1696,
    n1697,
    n1744,
    n1615
  );


  and
  g2281
  (
    n1978,
    n1761,
    n1747,
    n1771,
    n1694
  );


  xor
  g2282
  (
    n1828,
    n1793,
    n1611,
    n1635,
    n1705
  );


  xnor
  g2283
  (
    n2204,
    n1647,
    n1704,
    n1730,
    n1618
  );


  nor
  g2284
  (
    n2071,
    n1682,
    n1713,
    n1650,
    n1773
  );


  and
  g2285
  (
    n2067,
    n1628,
    n1758,
    n1614,
    n1799
  );


  xnor
  g2286
  (
    n1956,
    n1768,
    n1778,
    n1640,
    n1698
  );


  and
  g2287
  (
    n2066,
    n1672,
    n1747,
    n1753,
    n1795
  );


  nor
  g2288
  (
    n1881,
    n1791,
    n1721,
    n1626,
    n1713
  );


  nand
  g2289
  (
    n2109,
    n1704,
    n1641,
    n1495,
    n1628
  );


  or
  g2290
  (
    n2059,
    n1601,
    n1656,
    n1643,
    n1755
  );


  or
  g2291
  (
    n2133,
    n1639,
    n1672,
    n1634,
    n1679
  );


  xnor
  g2292
  (
    n2254,
    n1762,
    n1786,
    n1612,
    n1771
  );


  or
  g2293
  (
    n2005,
    n1799,
    n1604,
    n1764,
    n1788
  );


  nand
  g2294
  (
    n2332,
    n1759,
    n1693,
    n1610,
    n1803
  );


  xor
  g2295
  (
    n2258,
    n1654,
    n1641,
    n1719,
    n1696
  );


  xnor
  g2296
  (
    n2157,
    n1782,
    n1705,
    n1769,
    n1707
  );


  nand
  g2297
  (
    n2228,
    n1738,
    n1730,
    n1689,
    n1754
  );


  xnor
  g2298
  (
    n1930,
    n1650,
    n1720,
    n1725,
    n1659
  );


  or
  g2299
  (
    n1822,
    n1670,
    n1727,
    n1644,
    n1657
  );


  xnor
  g2300
  (
    n2325,
    n1637,
    n1605,
    n1642,
    n1611
  );


  nand
  g2301
  (
    n2144,
    n1766,
    n1611,
    n1765,
    n1782
  );


  nor
  g2302
  (
    n2361,
    n1671,
    n1602,
    n1736,
    n1700
  );


  nand
  g2303
  (
    n2303,
    n1716,
    n1732,
    n1779,
    n1665
  );


  and
  g2304
  (
    n2166,
    n1701,
    n1647,
    n1731,
    n1677
  );


  nor
  g2305
  (
    n1946,
    n1723,
    n1621,
    n1683,
    n1735
  );


  or
  g2306
  (
    n2088,
    n1750,
    n1609,
    n1642,
    n1652
  );


  xor
  g2307
  (
    n2186,
    n1749,
    n1784,
    n1627,
    n1797
  );


  nand
  g2308
  (
    n2149,
    n1692,
    n1729,
    n1698,
    n1735
  );


  xnor
  g2309
  (
    n1867,
    n1652,
    n1615,
    n1608,
    n1710
  );


  xor
  g2310
  (
    n2045,
    n1660,
    n1721,
    n1733,
    n1645
  );


  and
  g2311
  (
    n2132,
    n1731,
    n1751,
    n1753,
    n1680
  );


  or
  g2312
  (
    n1877,
    n1687,
    n1703,
    n1787,
    n1669
  );


  xnor
  g2313
  (
    n1830,
    n1737,
    n1742,
    n1752,
    n1494
  );


  and
  g2314
  (
    n2372,
    n1648,
    n1749,
    n1633,
    n1803
  );


  xor
  g2315
  (
    n1997,
    n1782,
    n1785,
    n1786,
    n1760
  );


  or
  g2316
  (
    n1832,
    n1740,
    n1614,
    n1790,
    n1717
  );


  xor
  g2317
  (
    n2329,
    n1739,
    n1732,
    n1625,
    n1623
  );


  or
  g2318
  (
    n2302,
    n1796,
    n1645,
    n1683,
    n1718
  );


  xor
  g2319
  (
    n1995,
    n1706,
    n1717,
    n1783,
    n1686
  );


  xnor
  g2320
  (
    n1839,
    n1759,
    n1777,
    n1639,
    n1681
  );


  nand
  g2321
  (
    n1825,
    n1731,
    n1769,
    n1620,
    n1725
  );


  xnor
  g2322
  (
    n2126,
    n1659,
    n1662,
    n1729,
    n1691
  );


  or
  g2323
  (
    n1876,
    n1718,
    n1798,
    n1647,
    n1770
  );


  xnor
  g2324
  (
    n2199,
    n1712,
    n1708,
    n1767,
    n1697
  );


  xor
  g2325
  (
    n2112,
    n1773,
    n1616,
    n1808,
    n1714
  );


  and
  g2326
  (
    n1843,
    n1737,
    n1698,
    n1780,
    n1806
  );


  xnor
  g2327
  (
    n2265,
    n1690,
    n1687,
    n1713,
    n1631
  );


  nand
  g2328
  (
    n2232,
    n1674,
    n1801,
    n1751,
    n1670
  );


  nor
  g2329
  (
    n1908,
    n1640,
    n1669,
    n1802,
    n1703
  );


  and
  g2330
  (
    n2295,
    n1631,
    n1613,
    n1626
  );


  xnor
  g2331
  (
    n2307,
    n1676,
    n1660,
    n1652,
    n1757
  );


  nand
  g2332
  (
    n2056,
    n1675,
    n1605,
    n1754,
    n1699
  );


  xnor
  g2333
  (
    n2357,
    n1703,
    n1631,
    n1633,
    n1614
  );


  and
  g2334
  (
    n2300,
    n1780,
    n1774,
    n1709,
    n1741
  );


  xor
  g2335
  (
    n1957,
    n1797,
    n1665,
    n1779,
    n1617
  );


  and
  g2336
  (
    n2351,
    n1663,
    n1710,
    n1795,
    n1772
  );


  or
  g2337
  (
    n2184,
    n1695,
    n1729,
    n1783,
    n1781
  );


  xor
  g2338
  (
    n2380,
    n1605,
    n1759,
    n1693,
    n1775
  );


  nor
  g2339
  (
    n1929,
    n1794,
    n1756,
    n1720,
    n1643
  );


  or
  g2340
  (
    n2187,
    n1651,
    n1807,
    n1764,
    n1680
  );


  nor
  g2341
  (
    n2323,
    n1670,
    n1694,
    n1649,
    n1807
  );


  xnor
  g2342
  (
    n2221,
    n1636,
    n1662,
    n1735,
    n1625
  );


  xnor
  g2343
  (
    n2377,
    n1696,
    n1734,
    n1717,
    n1699
  );


  and
  g2344
  (
    n2101,
    n1686,
    n1711,
    n1789,
    n1612
  );


  and
  g2345
  (
    n1910,
    n1772,
    n1727,
    n1630,
    n1738
  );


  xnor
  g2346
  (
    n2376,
    n1755,
    n1616,
    n1718,
    n1686
  );


  xnor
  g2347
  (
    n2374,
    n1736,
    n1802,
    n1733,
    n1666
  );


  xor
  g2348
  (
    n1993,
    n1675,
    n1632,
    n1683,
    n1734
  );


  nor
  g2349
  (
    n2305,
    n1766,
    n1629,
    n1710,
    n1609
  );


  nand
  g2350
  (
    n2078,
    n1671,
    n1709,
    n1795,
    n1668
  );


  and
  g2351
  (
    n2495,
    n2210,
    n1838,
    n1945,
    n2181
  );


  nand
  g2352
  (
    n2443,
    n1987,
    n2342,
    n2308,
    n2171
  );


  nand
  g2353
  (
    n2388,
    n2080,
    n2045,
    n1990,
    n2085
  );


  xor
  g2354
  (
    n2561,
    n2170,
    n1995,
    n2275,
    n2050
  );


  or
  g2355
  (
    n2488,
    n2321,
    n2262,
    n2309,
    n1973
  );


  and
  g2356
  (
    n2420,
    n2278,
    n2355,
    n2037,
    n2146
  );


  or
  g2357
  (
    n2585,
    n1823,
    n1912,
    n2254,
    n2202
  );


  and
  g2358
  (
    n2427,
    n2359,
    n2169,
    n2086,
    n2082
  );


  xor
  g2359
  (
    n2541,
    n2326,
    n2336,
    n2292,
    n1937
  );


  xnor
  g2360
  (
    n2515,
    n2047,
    n2214,
    n2111,
    n1989
  );


  xnor
  g2361
  (
    n2554,
    n2182,
    n2168,
    n2293,
    n2268
  );


  and
  g2362
  (
    n2481,
    n1870,
    n2230,
    n2134,
    n2255
  );


  xor
  g2363
  (
    n2456,
    n2006,
    n2160,
    n2204,
    n2180
  );


  nand
  g2364
  (
    n2405,
    n2215,
    n2314,
    n2216,
    n2284
  );


  xor
  g2365
  (
    n2549,
    n2228,
    n2157,
    n2295,
    n2294
  );


  and
  g2366
  (
    n2398,
    n1896,
    n2126,
    n2360,
    n2075
  );


  xor
  g2367
  (
    n2417,
    n2288,
    n2218,
    n2090,
    n2344
  );


  xnor
  g2368
  (
    n2499,
    n1891,
    n2235,
    n2145,
    n2194
  );


  or
  g2369
  (
    n2565,
    n2361,
    n2356,
    n1983,
    n1934
  );


  or
  g2370
  (
    n2451,
    n2128,
    n1956,
    n2274,
    n2163
  );


  nor
  g2371
  (
    n2454,
    n2276,
    n2107,
    n2296,
    n2188
  );


  nor
  g2372
  (
    n2513,
    n2277,
    n2265,
    n2186,
    n1910
  );


  nand
  g2373
  (
    n2446,
    n2341,
    n2265,
    n2191,
    n2288
  );


  nor
  g2374
  (
    n2489,
    n2089,
    n2201,
    n2254,
    n2085
  );


  xnor
  g2375
  (
    n2544,
    n2312,
    n2325,
    n1994,
    n2327
  );


  xnor
  g2376
  (
    n2396,
    n2334,
    n1841,
    n2026,
    n1924
  );


  and
  g2377
  (
    n2466,
    n2173,
    n1890,
    n2305,
    n2055
  );


  nand
  g2378
  (
    n2505,
    n1913,
    n2348,
    n2116,
    n2337
  );


  xor
  g2379
  (
    n2556,
    n2034,
    n2137,
    n2226,
    n2328
  );


  and
  g2380
  (
    n2385,
    n2078,
    n2205,
    n2190,
    n2120
  );


  or
  g2381
  (
    n2453,
    n1970,
    n2202,
    n2149,
    n1862
  );


  xor
  g2382
  (
    n2403,
    n2287,
    n2358,
    n2255,
    n1820
  );


  nand
  g2383
  (
    n2461,
    n1878,
    n1980,
    n2244,
    n2191
  );


  nor
  g2384
  (
    n2529,
    n2290,
    n2118,
    n2147,
    n2151
  );


  and
  g2385
  (
    n2416,
    n2101,
    n2269,
    n1968,
    n2276
  );


  xor
  g2386
  (
    n2412,
    n2156,
    n1887,
    n2100,
    n2221
  );


  nand
  g2387
  (
    n2389,
    n2271,
    n2308,
    n2115,
    n2131
  );


  xor
  g2388
  (
    n2437,
    n2187,
    n2148,
    n1986,
    n1926
  );


  xor
  g2389
  (
    n2525,
    n2110,
    n2220,
    n1984,
    n1822
  );


  xor
  g2390
  (
    n2479,
    n2302,
    n1837,
    n2014,
    n2063
  );


  nor
  g2391
  (
    n2474,
    n2186,
    n2043,
    n1908,
    n1828
  );


  and
  g2392
  (
    n2575,
    n1825,
    n2246,
    n2136,
    n1849
  );


  nor
  g2393
  (
    n2587,
    n2183,
    n2062,
    n2230,
    n2135
  );


  nand
  g2394
  (
    n2462,
    n1900,
    n1819,
    n2140,
    n1836
  );


  xor
  g2395
  (
    n2573,
    n2168,
    n2198,
    n2227,
    n2209
  );


  xnor
  g2396
  (
    n2586,
    n2263,
    n2017,
    n1954,
    n2097
  );


  nor
  g2397
  (
    n2480,
    n1875,
    n2133,
    n2121,
    n1907
  );


  nor
  g2398
  (
    n2563,
    n2253,
    n2099,
    n1960,
    n1903
  );


  and
  g2399
  (
    n2524,
    n2112,
    n2155,
    n2015,
    n2243
  );


  nand
  g2400
  (
    n2478,
    n2259,
    n2301,
    n2176,
    n2125
  );


  xor
  g2401
  (
    n2472,
    n2077,
    n2005,
    n2028,
    n2161
  );


  nor
  g2402
  (
    n2557,
    n1949,
    n2183,
    n2358,
    n2256
  );


  nor
  g2403
  (
    n2533,
    n1917,
    n1873,
    n1948,
    n2101
  );


  xor
  g2404
  (
    n2387,
    n2356,
    n2152,
    n1932,
    n2172
  );


  xor
  g2405
  (
    n2476,
    n1978,
    n1943,
    n2088,
    n2149
  );


  and
  g2406
  (
    n2506,
    n2161,
    n2221,
    n2318,
    n2353
  );


  nor
  g2407
  (
    n2568,
    n2169,
    n1952,
    n2263,
    n2129
  );


  nor
  g2408
  (
    n2564,
    n2162,
    n1893,
    n2330,
    n2136
  );


  xor
  g2409
  (
    n2426,
    n2080,
    n2106,
    n2320,
    n2258
  );


  and
  g2410
  (
    n2455,
    n2289,
    n1992,
    n2270,
    n2122
  );


  or
  g2411
  (
    n2503,
    n2199,
    n2350,
    n2339,
    n2257
  );


  xnor
  g2412
  (
    n2395,
    n2319,
    n2331,
    n2192,
    n1827
  );


  and
  g2413
  (
    n2532,
    n2067,
    n2206,
    n2158,
    n1815
  );


  nand
  g2414
  (
    n2452,
    n2079,
    n2133,
    n2245,
    n2208
  );


  and
  g2415
  (
    n2519,
    n2317,
    n2346,
    n2152,
    n2351
  );


  or
  g2416
  (
    n2578,
    n2142,
    n2238,
    n1976
  );


  and
  g2417
  (
    n2439,
    n1914,
    n2292,
    n1920,
    n2189
  );


  and
  g2418
  (
    n2577,
    n1839,
    n2329,
    n2018,
    n2299
  );


  and
  g2419
  (
    n2408,
    n2347,
    n2182,
    n2158,
    n2035
  );


  nor
  g2420
  (
    n2468,
    n2140,
    n2210,
    n2128,
    n2179
  );


  nand
  g2421
  (
    n2516,
    n2181,
    n1899,
    n2326,
    n2156
  );


  nor
  g2422
  (
    n2401,
    n2009,
    n1911,
    n1957,
    n1824
  );


  nor
  g2423
  (
    n2580,
    n2025,
    n2317,
    n2138,
    n2076
  );


  nand
  g2424
  (
    n2440,
    n2040,
    n2195,
    n2150,
    n2021
  );


  nor
  g2425
  (
    n2393,
    n2041,
    n1946,
    n2159,
    n2125
  );


  xor
  g2426
  (
    n2402,
    n2096,
    n1919,
    n2144,
    n2245
  );


  nand
  g2427
  (
    n2407,
    n1951,
    n2341,
    n2170,
    n2222
  );


  nor
  g2428
  (
    n2491,
    n2258,
    n1940,
    n2273,
    n2131
  );


  and
  g2429
  (
    n2507,
    n2344,
    n2323,
    n2081,
    n2331
  );


  nand
  g2430
  (
    n2566,
    n2348,
    n2298,
    n1826,
    n2165
  );


  xor
  g2431
  (
    n2435,
    n2357,
    n1857,
    n1889,
    n2108
  );


  xor
  g2432
  (
    n2404,
    n2240,
    n2004,
    n2218,
    n1982
  );


  or
  g2433
  (
    n2444,
    n2196,
    n1964,
    n2316,
    n1821
  );


  xor
  g2434
  (
    n2477,
    n2173,
    n2211,
    n2212,
    n2209
  );


  nor
  g2435
  (
    n2409,
    n2077,
    n1996,
    n2082,
    n2338
  );


  xnor
  g2436
  (
    n2588,
    n2109,
    n2114,
    n2307,
    n2283
  );


  or
  g2437
  (
    n2501,
    n2232,
    n1999,
    n2318,
    n2117
  );


  nor
  g2438
  (
    n2482,
    n1866,
    n1988,
    n1835,
    n1953
  );


  xnor
  g2439
  (
    n2540,
    n2180,
    n2030,
    n2242,
    n2144
  );


  nand
  g2440
  (
    n2530,
    n1901,
    n2330,
    n1955,
    n2219
  );


  xor
  g2441
  (
    n2460,
    n2162,
    n2234,
    n2197,
    n1981
  );


  nor
  g2442
  (
    n2464,
    n2075,
    n2112,
    n1869,
    n1929
  );


  nor
  g2443
  (
    n2422,
    n2332,
    n2095,
    n1925,
    n1985
  );


  xnor
  g2444
  (
    n2433,
    n2281,
    n2360,
    n2102,
    n2118
  );


  nand
  g2445
  (
    n2441,
    n2247,
    n2086,
    n2165,
    n2175
  );


  and
  g2446
  (
    n2560,
    n2220,
    n2107,
    n2244,
    n2307
  );


  xnor
  g2447
  (
    n2527,
    n1892,
    n2066,
    n1856,
    n2184
  );


  nand
  g2448
  (
    n2411,
    n2290,
    n2332,
    n2334,
    n2146
  );


  xor
  g2449
  (
    n2486,
    n2349,
    n2324,
    n2248,
    n2363
  );


  xnor
  g2450
  (
    n2421,
    n2325,
    n2365,
    n2232,
    n1833
  );


  xnor
  g2451
  (
    n2591,
    n2148,
    n1977,
    n2108,
    n2257
  );


  xor
  g2452
  (
    n2518,
    n2088,
    n2123,
    n2310,
    n2083
  );


  xnor
  g2453
  (
    n2509,
    n2203,
    n1923,
    n2306,
    n2011
  );


  nor
  g2454
  (
    n2429,
    n2100,
    n2294,
    n2225,
    n2293
  );


  nand
  g2455
  (
    n2579,
    n2003,
    n2224,
    n2147,
    n2177
  );


  and
  g2456
  (
    n2448,
    n1814,
    n2083,
    n2189,
    n1832
  );


  xnor
  g2457
  (
    n2418,
    n2187,
    n1867,
    n1885,
    n2116
  );


  xor
  g2458
  (
    n2490,
    n1905,
    n2250,
    n2121,
    n2321
  );


  xor
  g2459
  (
    n2553,
    n2188,
    n2247,
    n2104,
    n1935
  );


  or
  g2460
  (
    n2559,
    n1927,
    n2207,
    n2231,
    n2167
  );


  or
  g2461
  (
    n2582,
    n1939,
    n2279,
    n2340,
    n2145
  );


  or
  g2462
  (
    n2457,
    n2091,
    n2057,
    n2051,
    n2105
  );


  or
  g2463
  (
    n2494,
    n1897,
    n2184,
    n1931,
    n2058
  );


  xor
  g2464
  (
    n2425,
    n2038,
    n1997,
    n1854,
    n1902
  );


  and
  g2465
  (
    n2517,
    n2000,
    n2216,
    n2022,
    n2241
  );


  xor
  g2466
  (
    n2526,
    n2251,
    n2282,
    n2027,
    n2239
  );


  or
  g2467
  (
    n2595,
    n2127,
    n2124,
    n2020,
    n2343
  );


  xor
  g2468
  (
    n2465,
    n2223,
    n2235,
    n2090,
    n2260
  );


  and
  g2469
  (
    n2500,
    n2081,
    n2286,
    n2141,
    n2093
  );


  xnor
  g2470
  (
    n2423,
    n2355,
    n1872,
    n2319,
    n2354
  );


  xnor
  g2471
  (
    n2546,
    n2142,
    n2291,
    n2249,
    n2141
  );


  xor
  g2472
  (
    n2391,
    n1941,
    n2217,
    n2163,
    n1816
  );


  xor
  g2473
  (
    n2576,
    n2032,
    n1846,
    n1962,
    n2102
  );


  xnor
  g2474
  (
    n2569,
    n2060,
    n2124,
    n2347,
    n2266
  );


  and
  g2475
  (
    n2543,
    n2059,
    n2091,
    n2335,
    n2049
  );


  or
  g2476
  (
    n2535,
    n2048,
    n2069,
    n1936,
    n2272
  );


  xnor
  g2477
  (
    n2434,
    n1898,
    n2214,
    n1906,
    n1852
  );


  nand
  g2478
  (
    n2548,
    n2110,
    n1847,
    n2073,
    n1969
  );


  nor
  g2479
  (
    n2400,
    n2013,
    n1991,
    n2164,
    n2333
  );


  and
  g2480
  (
    n2583,
    n1933,
    n2267,
    n1861,
    n2007
  );


  or
  g2481
  (
    n2536,
    n2178,
    n2229,
    n2304,
    n2119
  );


  nor
  g2482
  (
    n2463,
    n2064,
    n1883,
    n2300,
    n2094
  );


  nor
  g2483
  (
    n2534,
    n2179,
    n2284,
    n2260,
    n2196
  );


  nor
  g2484
  (
    n2550,
    n2302,
    n2106,
    n1855,
    n2076
  );


  xnor
  g2485
  (
    n2386,
    n2211,
    n2084,
    n2153,
    n2104
  );


  nand
  g2486
  (
    n2390,
    n2251,
    n2117,
    n2203,
    n2252
  );


  and
  g2487
  (
    n2510,
    n1965,
    n2291,
    n2315,
    n2174
  );


  xnor
  g2488
  (
    n2520,
    n2237,
    n2016,
    n1881,
    n1882
  );


  nor
  g2489
  (
    n2410,
    n2193,
    n2310,
    n2249,
    n1812
  );


  xor
  g2490
  (
    n2485,
    n2079,
    n1813,
    n2243,
    n2357
  );


  and
  g2491
  (
    n2581,
    n2087,
    n1918,
    n2120,
    n1963
  );


  nor
  g2492
  (
    n2470,
    n2143,
    n2199,
    n2008,
    n2264
  );


  xor
  g2493
  (
    n2528,
    n2233,
    n2270,
    n2177,
    n2364
  );


  xnor
  g2494
  (
    n2496,
    n2296,
    n2217,
    n2264,
    n1817
  );


  xor
  g2495
  (
    n2431,
    n1853,
    n1904,
    n2099,
    n2031
  );


  xnor
  g2496
  (
    n2537,
    n2335,
    n2103,
    n2208,
    n2150
  );


  nand
  g2497
  (
    n2572,
    n1865,
    n2215,
    n2213,
    n2287
  );


  nand
  g2498
  (
    n2521,
    n2250,
    n1930,
    n2095,
    n2010
  );


  xor
  g2499
  (
    n2450,
    n2351,
    n2002,
    n2153,
    n2349
  );


  xnor
  g2500
  (
    n2504,
    n2139,
    n2143,
    n2042,
    n2023
  );


  xnor
  g2501
  (
    n2483,
    n1950,
    n2001,
    n2113,
    n1974
  );


  xnor
  g2502
  (
    n2512,
    n2278,
    n2313,
    n2098,
    n1871
  );


  nor
  g2503
  (
    n2487,
    n2070,
    n2309,
    n2138,
    n2224
  );


  and
  g2504
  (
    n2399,
    n2074,
    n2267,
    n2024,
    n2033
  );


  xor
  g2505
  (
    n2592,
    n2094,
    n2333,
    n2345,
    n2092
  );


  xor
  g2506
  (
    n2414,
    n1851,
    n2313,
    n2115,
    n2052
  );


  and
  g2507
  (
    n2567,
    n2363,
    n2134,
    n1975,
    n2213
  );


  xnor
  g2508
  (
    n2471,
    n2301,
    n1928,
    n2300,
    n2200
  );


  or
  g2509
  (
    n2449,
    n2322,
    n2127,
    n2248,
    n2185
  );


  and
  g2510
  (
    n2397,
    n2289,
    n2212,
    n2241,
    n2151
  );


  nand
  g2511
  (
    n2458,
    n1966,
    n2114,
    n2336,
    n2343
  );


  and
  g2512
  (
    n2590,
    n2337,
    n2315,
    n2084,
    n1947
  );


  xnor
  g2513
  (
    n2406,
    n2364,
    n2266,
    n1829,
    n2236
  );


  and
  g2514
  (
    n2475,
    n1834,
    n2053,
    n2071,
    n1868
  );


  nor
  g2515
  (
    n2545,
    n2338,
    n1967,
    n2353,
    n2029
  );


  and
  g2516
  (
    n2469,
    n2275,
    n2231,
    n1809,
    n2253
  );


  and
  g2517
  (
    n2547,
    n2039,
    n2154,
    n2362,
    n2192
  );


  or
  g2518
  (
    n2508,
    n2159,
    n2297,
    n2119,
    n1886
  );


  and
  g2519
  (
    n2523,
    n2303,
    n2365,
    n2185,
    n1848
  );


  nor
  g2520
  (
    n2428,
    n2087,
    n2272,
    n2252,
    n2166
  );


  or
  g2521
  (
    n2392,
    n2036,
    n1916,
    n2044,
    n2103
  );


  and
  g2522
  (
    n2413,
    n2155,
    n2277,
    n2197,
    n1840
  );


  and
  g2523
  (
    n2522,
    n2359,
    n1915,
    n1874,
    n2200
  );


  nor
  g2524
  (
    n2570,
    n2222,
    n2130,
    n2061,
    n2324
  );


  xor
  g2525
  (
    n2497,
    n1850,
    n2176,
    n2065,
    n2135
  );


  nand
  g2526
  (
    n2555,
    n2274,
    n2328,
    n2164,
    n2167
  );


  xnor
  g2527
  (
    n2438,
    n2236,
    n1938,
    n2228,
    n2195
  );


  or
  g2528
  (
    n2430,
    n2172,
    n1979,
    n2194,
    n2280
  );


  and
  g2529
  (
    n2419,
    n1880,
    n2154,
    n2056,
    n1864
  );


  xnor
  g2530
  (
    n2467,
    n2126,
    n2111,
    n2352,
    n2304
  );


  nand
  g2531
  (
    n2436,
    n1863,
    n2242,
    n2096,
    n2137
  );


  nand
  g2532
  (
    n2459,
    n1860,
    n2322,
    n2282,
    n2285
  );


  nand
  g2533
  (
    n2384,
    n1894,
    n2012,
    n1858,
    n1942
  );


  or
  g2534
  (
    n2539,
    n2323,
    n2285,
    n2132,
    n2280
  );


  xnor
  g2535
  (
    n2571,
    n1818,
    n1971,
    n2093,
    n1959
  );


  and
  g2536
  (
    n2538,
    n2178,
    n1884,
    n2240,
    n2219
  );


  xnor
  g2537
  (
    n2442,
    n2295,
    n1961,
    n1859,
    n2068
  );


  xnor
  g2538
  (
    n2424,
    n2097,
    n1888,
    n2098,
    n2246
  );


  or
  g2539
  (
    n2473,
    n2190,
    n2054,
    n2362,
    n2129
  );


  or
  g2540
  (
    n2492,
    n2311,
    n2340,
    n2329,
    n2072
  );


  xnor
  g2541
  (
    n2589,
    n2259,
    n2078,
    n1993,
    n2361
  );


  xnor
  g2542
  (
    n2484,
    n1879,
    n2109,
    n2174,
    n2201
  );


  and
  g2543
  (
    n2552,
    n2350,
    n2262,
    n2019,
    n2342
  );


  and
  g2544
  (
    n2584,
    n1998,
    n2354,
    n2160,
    n1944
  );


  and
  g2545
  (
    n2542,
    n2298,
    n2320,
    n1842,
    n1921
  );


  nor
  g2546
  (
    n2493,
    n1895,
    n2261,
    n2283,
    n2157
  );


  nor
  g2547
  (
    n2511,
    n2256,
    n2206,
    n2286,
    n1831
  );


  or
  g2548
  (
    n2432,
    n2227,
    n2303,
    n2198,
    n2204
  );


  nand
  g2549
  (
    n2558,
    n2089,
    n2312,
    n1845,
    n2352
  );


  nand
  g2550
  (
    n2502,
    n2233,
    n1909,
    n2092,
    n2225
  );


  xor
  g2551
  (
    n2498,
    n1958,
    n1810,
    n2139,
    n2237
  );


  nor
  g2552
  (
    n2593,
    n2226,
    n2234,
    n1876,
    n2105
  );


  and
  g2553
  (
    n2531,
    n1877,
    n1844,
    n2113,
    n2130
  );


  nor
  g2554
  (
    n2562,
    n2166,
    n2327,
    n2269,
    n2279
  );


  xor
  g2555
  (
    n2594,
    n1922,
    n2345,
    n2205,
    n1972
  );


  nand
  g2556
  (
    n2394,
    n2268,
    n2299,
    n2046,
    n2339
  );


  nor
  g2557
  (
    n2447,
    n2207,
    n2171,
    n2132,
    n2314
  );


  xnor
  g2558
  (
    n2415,
    n2271,
    n2316,
    n2346,
    n2239
  );


  nand
  g2559
  (
    n2551,
    n1830,
    n2123,
    n2297,
    n2223
  );


  or
  g2560
  (
    n2514,
    n2122,
    n2273,
    n2281,
    n1811
  );


  xnor
  g2561
  (
    n2574,
    n1843,
    n2311,
    n2305,
    n2229
  );


  or
  g2562
  (
    n2445,
    n2175,
    n2193,
    n2306,
    n2261
  );


  nor
  g2563
  (
    n2608,
    n2486,
    n2453,
    n2415,
    n2424
  );


  nor
  g2564
  (
    n2598,
    n2500,
    n2493,
    n2430,
    n2487
  );


  and
  g2565
  (
    n2612,
    n2465,
    n2400,
    n2483,
    n2404
  );


  or
  g2566
  (
    n2596,
    n2459,
    n2452,
    n2393,
    n2478
  );


  nand
  g2567
  (
    n2625,
    n2392,
    n2429,
    n2475,
    n2451
  );


  xor
  g2568
  (
    n2597,
    n2432,
    n2388,
    n2456,
    n2410
  );


  and
  g2569
  (
    n2601,
    n2420,
    n2494,
    n2448,
    n2398
  );


  nor
  g2570
  (
    n2602,
    n2417,
    n2394,
    n2445,
    n2495
  );


  and
  g2571
  (
    n2618,
    n2454,
    n2396,
    n2476,
    n2403
  );


  nand
  g2572
  (
    n2609,
    n2499,
    n2458,
    n2413,
    n2435
  );


  or
  g2573
  (
    n2616,
    n2480,
    n2431,
    n2385,
    n2389
  );


  or
  g2574
  (
    n2611,
    n2390,
    n2472,
    n2440,
    n2473
  );


  or
  g2575
  (
    n2617,
    n2443,
    n2491,
    n2479,
    n2399
  );


  xor
  g2576
  (
    n2606,
    n2488,
    n2426,
    n2391,
    n2497
  );


  xor
  g2577
  (
    n2599,
    n2409,
    n2384,
    n2464,
    n2418
  );


  nand
  g2578
  (
    n2600,
    n2484,
    n2423,
    n2407,
    n2433
  );


  or
  g2579
  (
    n2622,
    n2462,
    n2466,
    n2455,
    n2439
  );


  or
  g2580
  (
    n2623,
    n2419,
    n2470,
    n2427,
    n2397
  );


  xnor
  g2581
  (
    n2607,
    n2490,
    n2450,
    n2469,
    n2411
  );


  or
  g2582
  (
    n2604,
    n2447,
    n2401,
    n2405,
    n2498
  );


  and
  g2583
  (
    n2610,
    n2428,
    n2449,
    n2460,
    n2422
  );


  xnor
  g2584
  (
    n2615,
    n2485,
    n2461,
    n2442,
    n2395
  );


  xor
  g2585
  (
    n2624,
    n2416,
    n2503,
    n2437,
    n2482
  );


  xnor
  g2586
  (
    n2605,
    n2434,
    n2502,
    n2408,
    n2444
  );


  nor
  g2587
  (
    n2614,
    n2387,
    n2406,
    n2441,
    n2474
  );


  nand
  g2588
  (
    n2613,
    n2438,
    n2457,
    n2412,
    n2468
  );


  or
  g2589
  (
    n2621,
    n2467,
    n2436,
    n2481,
    n2492
  );


  xnor
  g2590
  (
    n2619,
    n2425,
    n2402,
    n2489,
    n2446
  );


  xor
  g2591
  (
    n2620,
    n2496,
    n2386,
    n2463,
    n2477
  );


  xnor
  g2592
  (
    n2603,
    n2471,
    n2414,
    n2421,
    n2501
  );


  buf
  g2593
  (
    n2630,
    n1299
  );


  buf
  g2594
  (
    n2635,
    n1303
  );


  buf
  g2595
  (
    n2632,
    n2606
  );


  not
  g2596
  (
    n2627,
    n2599
  );


  not
  g2597
  (
    n2631,
    n1298
  );


  buf
  g2598
  (
    n2639,
    n2599
  );


  buf
  g2599
  (
    n2626,
    n2606
  );


  not
  g2600
  (
    n2633,
    n2600
  );


  buf
  g2601
  (
    n2628,
    n1304
  );


  not
  g2602
  (
    n2629,
    n2597
  );


  nand
  g2603
  (
    n2634,
    n1310,
    n1305
  );


  xor
  g2604
  (
    n2637,
    n2596,
    n2601,
    n1307,
    n1300
  );


  xor
  g2605
  (
    n2636,
    n2597,
    n2601,
    n2596,
    n2600
  );


  and
  g2606
  (
    n2642,
    n2602,
    n2604,
    n1301,
    n1308
  );


  xnor
  g2607
  (
    n2638,
    n2603,
    n1302,
    n2605
  );


  and
  g2608
  (
    n2641,
    n2602,
    n2603,
    n2604,
    n2598
  );


  nor
  g2609
  (
    n2640,
    n1306,
    n1297,
    n2598,
    n1309
  );


  not
  g2610
  (
    n2661,
    n2370
  );


  buf
  g2611
  (
    n2650,
    n2628
  );


  not
  g2612
  (
    n2651,
    n2374
  );


  not
  g2613
  (
    n2662,
    n2630
  );


  buf
  g2614
  (
    n2649,
    n2633
  );


  buf
  g2615
  (
    n2669,
    n2639
  );


  buf
  g2616
  (
    n2664,
    n2627
  );


  buf
  g2617
  (
    n2659,
    n2369
  );


  buf
  g2618
  (
    n2652,
    n2631
  );


  buf
  g2619
  (
    n2665,
    n2373
  );


  buf
  g2620
  (
    n2660,
    n2636
  );


  not
  g2621
  (
    n2667,
    n2368
  );


  buf
  g2622
  (
    n2668,
    n2375
  );


  buf
  g2623
  (
    n2671,
    n2638
  );


  buf
  g2624
  (
    n2653,
    n2631
  );


  not
  g2625
  (
    n2656,
    n2376
  );


  not
  g2626
  (
    n2644,
    n2639
  );


  nand
  g2627
  (
    n2647,
    n2381,
    n2628,
    n2635
  );


  xor
  g2628
  (
    n2658,
    n2627,
    n2374,
    n2634,
    n2369
  );


  and
  g2629
  (
    n2643,
    n2626,
    n2383,
    n2382,
    n2367
  );


  and
  g2630
  (
    n2648,
    n2378,
    n2640,
    n2379,
    n2634
  );


  or
  g2631
  (
    n2663,
    n2373,
    n2371,
    n2368
  );


  nand
  g2632
  (
    n2666,
    n2630,
    n2378,
    n2629,
    n2638
  );


  nor
  g2633
  (
    n2655,
    n2626,
    n2629,
    n2366,
    n2632
  );


  xor
  g2634
  (
    n2670,
    n2370,
    n2372,
    n2366,
    n2367
  );


  or
  g2635
  (
    n2657,
    n2377,
    n2380,
    n2372,
    n2636
  );


  xnor
  g2636
  (
    n2645,
    n2376,
    n2379,
    n2375,
    n2377
  );


  xnor
  g2637
  (
    n2654,
    n2633,
    n2637,
    n2632
  );


  nand
  g2638
  (
    n2646,
    n2382,
    n2381,
    n2635,
    n2380
  );


  and
  g2639
  (
    n2688,
    n2566,
    n2576,
    n2573,
    n2578
  );


  and
  g2640
  (
    n2679,
    n2648,
    n2518,
    n2587,
    n2519
  );


  nor
  g2641
  (
    n2692,
    n2570,
    n2582,
    n2544,
    n2569
  );


  nand
  g2642
  (
    n2691,
    n2555,
    n2530,
    n2577,
    n2644
  );


  nor
  g2643
  (
    n2676,
    n2539,
    n2564,
    n2644,
    n2532
  );


  or
  g2644
  (
    n2699,
    n2552,
    n2512,
    n2549,
    n2560
  );


  xor
  g2645
  (
    n2693,
    n2507,
    n2643,
    n2648,
    n2529
  );


  and
  g2646
  (
    n2685,
    n2551,
    n2545,
    n2646
  );


  xor
  g2647
  (
    n2694,
    n2649,
    n2647,
    n2583,
    n2585
  );


  and
  g2648
  (
    n2681,
    n2568,
    n2649,
    n2556,
    n2504
  );


  and
  g2649
  (
    n2690,
    n2575,
    n2645,
    n2580,
    n2584
  );


  nor
  g2650
  (
    n2683,
    n2644,
    n2557,
    n2579,
    n2536
  );


  nand
  g2651
  (
    n2677,
    n2644,
    n2517,
    n2533,
    n2506
  );


  xnor
  g2652
  (
    n2689,
    n2572,
    n2565,
    n2510,
    n2650
  );


  xnor
  g2653
  (
    n2680,
    n2515,
    n2646,
    n2521,
    n2650
  );


  nand
  g2654
  (
    n2696,
    n2647,
    n2561,
    n2531,
    n2540
  );


  xor
  g2655
  (
    n2672,
    n2505,
    n2514,
    n2527,
    n2534
  );


  or
  g2656
  (
    n2686,
    n2550,
    n2535,
    n2538,
    n2649
  );


  and
  g2657
  (
    n2698,
    n2523,
    n2649,
    n2558,
    n2516
  );


  nand
  g2658
  (
    n2678,
    n2646,
    n2647,
    n2548,
    n2645
  );


  xor
  g2659
  (
    n2675,
    n2547,
    n2528,
    n2559,
    n2525
  );


  and
  g2660
  (
    n2684,
    n2645,
    n2520,
    n2542,
    n2511
  );


  xor
  g2661
  (
    n2695,
    n2522,
    n2571,
    n2581,
    n2537
  );


  xor
  g2662
  (
    n2682,
    n2643,
    n2567,
    n2563,
    n2562
  );


  and
  g2663
  (
    n2673,
    n2543,
    n2554,
    n2524,
    n2648
  );


  or
  g2664
  (
    n2687,
    n2648,
    n2553,
    n2574,
    n2645
  );


  and
  g2665
  (
    n2697,
    n2513,
    n2509,
    n2546,
    n2508
  );


  or
  g2666
  (
    n2674,
    n2541,
    n2526,
    n2586,
    n2647
  );


  not
  g2667
  (
    n2701,
    n2609
  );


  buf
  g2668
  (
    n2718,
    n2675
  );


  not
  g2669
  (
    n2710,
    n2675
  );


  buf
  g2670
  (
    n2720,
    n2676
  );


  not
  g2671
  (
    n2714,
    n2679
  );


  not
  g2672
  (
    n2702,
    n953
  );


  buf
  g2673
  (
    n2729,
    n2617
  );


  buf
  g2674
  (
    n2723,
    n953
  );


  buf
  g2675
  (
    n2728,
    n2678
  );


  not
  g2676
  (
    n2713,
    n954
  );


  not
  g2677
  (
    n2700,
    n2673
  );


  buf
  g2678
  (
    n2706,
    n2675
  );


  buf
  g2679
  (
    n2705,
    n2613
  );


  xor
  g2680
  (
    n2704,
    n2676,
    n2621,
    n2607
  );


  or
  g2681
  (
    n2707,
    n954,
    n2612,
    n2676,
    n2614
  );


  xor
  g2682
  (
    n2722,
    n952,
    n2608,
    n2624,
    n2622
  );


  or
  g2683
  (
    n2709,
    n2611,
    n2619,
    n2622,
    n2610
  );


  and
  g2684
  (
    n2703,
    n2608,
    n2676,
    n2674,
    n2625
  );


  and
  g2685
  (
    n2727,
    n2617,
    n2673,
    n2677,
    n2678
  );


  xnor
  g2686
  (
    n2715,
    n2672,
    n2674,
    n952
  );


  xnor
  g2687
  (
    n2726,
    n2672,
    n2621,
    n2619,
    n2674
  );


  xor
  g2688
  (
    n2712,
    n2678,
    n2677,
    n2672,
    n2615
  );


  or
  g2689
  (
    n2721,
    n2610,
    n2624,
    n2609,
    n953
  );


  xor
  g2690
  (
    n2724,
    n2620,
    n2677,
    n2613,
    n953
  );


  nand
  g2691
  (
    n2711,
    n2677,
    n2675,
    n954,
    n2673
  );


  xor
  g2692
  (
    n2708,
    n2672,
    n2611,
    n2678,
    n2383
  );


  xnor
  g2693
  (
    n2725,
    n2673,
    n2620,
    n2679,
    n2616
  );


  xnor
  g2694
  (
    n2716,
    n2625,
    n2623,
    n2616,
    n2615
  );


  xnor
  g2695
  (
    n2719,
    n2623,
    n2607,
    n954,
    n2674
  );


  xnor
  g2696
  (
    n2717,
    n2618,
    n2618,
    n2612,
    n2614
  );


  nor
  g2697
  (
    n2738,
    n2722,
    n2714,
    n2721,
    n2704
  );


  nor
  g2698
  (
    n2742,
    n2709,
    n2713,
    n2710,
    n2719
  );


  nor
  g2699
  (
    n2732,
    n2722,
    n2700,
    n2716,
    n2706
  );


  xnor
  g2700
  (
    n2741,
    n2713,
    n2718,
    n2705
  );


  xnor
  g2701
  (
    n2737,
    n2716,
    n2707,
    n2717,
    n2703
  );


  nand
  g2702
  (
    n2731,
    n2720,
    n2724,
    n2721,
    n2711
  );


  nand
  g2703
  (
    n2740,
    n2701,
    n2706,
    n2708,
    n2717
  );


  or
  g2704
  (
    n2730,
    n2724,
    n2719,
    n2714,
    n2704
  );


  nor
  g2705
  (
    n2736,
    n2725,
    n2725,
    n2709,
    n2720
  );


  xnor
  g2706
  (
    n2735,
    n2705,
    n2703,
    n2701,
    n2708
  );


  nand
  g2707
  (
    n2733,
    n2707,
    n2700,
    n2712
  );


  nand
  g2708
  (
    n2734,
    n2711,
    n2715,
    n2723,
    n2702
  );


  and
  g2709
  (
    n2739,
    n2715,
    n2702,
    n2710,
    n2723
  );


  xnor
  g2710
  (
    n2772,
    n2732,
    n2651,
    n2655
  );


  xnor
  g2711
  (
    n2783,
    n2731,
    n2737,
    n2654
  );


  nor
  g2712
  (
    n2762,
    n2658,
    n2669,
    n2662
  );


  and
  g2713
  (
    n2775,
    n2670,
    n2738,
    n2737
  );


  xnor
  g2714
  (
    n2755,
    n2671,
    n1443,
    n2733
  );


  and
  g2715
  (
    n2784,
    n2665,
    n2663,
    n2652
  );


  nor
  g2716
  (
    n2751,
    n2728,
    n2653,
    n2736
  );


  xor
  g2717
  (
    n2753,
    n2668,
    n2656,
    n2732
  );


  or
  g2718
  (
    n2757,
    n2656,
    n2736,
    n2671
  );


  nor
  g2719
  (
    n2773,
    n2734,
    n2728,
    n1444
  );


  nor
  g2720
  (
    n2778,
    n2660,
    n2739,
    n2667
  );


  and
  g2721
  (
    n2764,
    n2662,
    n2734,
    n2655
  );


  xnor
  g2722
  (
    n2766,
    n2661,
    n2740,
    n2659
  );


  nand
  g2723
  (
    n2779,
    n2736,
    n2660
  );


  and
  g2724
  (
    n2759,
    n2661,
    n2739,
    n2662
  );


  or
  g2725
  (
    n2769,
    n2664,
    n2659,
    n2651,
    n2655
  );


  xnor
  g2726
  (
    n2768,
    n2666,
    n2742,
    n1445,
    n2741
  );


  nand
  g2727
  (
    n2748,
    n2657,
    n2653,
    n2665,
    n1314
  );


  xor
  g2728
  (
    n2765,
    n2735,
    n1311,
    n2741,
    n2738
  );


  xnor
  g2729
  (
    n2756,
    n2652,
    n2659,
    n1316,
    n2651
  );


  nor
  g2730
  (
    n2754,
    n2738,
    n2727,
    n2739
  );


  and
  g2731
  (
    n2776,
    n1313,
    n2726,
    n1315,
    n2730
  );


  xnor
  g2732
  (
    n2781,
    n2742,
    n2731,
    n2737,
    n2730
  );


  xnor
  g2733
  (
    n2770,
    n2670,
    n2655,
    n1312,
    n1444
  );


  nor
  g2734
  (
    n2771,
    n2740,
    n2654,
    n2664,
    n2662
  );


  and
  g2735
  (
    n2782,
    n2663,
    n1318,
    n2669,
    n2657
  );


  xor
  g2736
  (
    n2777,
    n2670,
    n2668,
    n2665,
    n2666
  );


  xor
  g2737
  (
    n2746,
    n2671,
    n2651,
    n2741
  );


  nor
  g2738
  (
    n2767,
    n1444,
    n2671,
    n2658,
    n2668
  );


  nand
  g2739
  (
    n2745,
    n2658,
    n2667,
    n2738,
    n2666
  );


  and
  g2740
  (
    n2744,
    n2659,
    n2661,
    n2736,
    n2663
  );


  and
  g2741
  (
    n2750,
    n2664,
    n2654,
    n2650,
    n1319
  );


  xnor
  g2742
  (
    n2780,
    n2737,
    n2661,
    n2667,
    n2658
  );


  or
  g2743
  (
    n2763,
    n2657,
    n2652,
    n1443,
    n2656
  );


  xnor
  g2744
  (
    n2761,
    n2657,
    n2652,
    n2742,
    n2665
  );


  xnor
  g2745
  (
    n2743,
    n2669,
    n2668,
    n2650,
    n2654
  );


  xor
  g2746
  (
    n2758,
    n2726,
    n2742,
    n2653,
    n1317
  );


  xor
  g2747
  (
    n2760,
    n2670,
    n2728,
    n2740,
    n1444
  );


  nor
  g2748
  (
    n2749,
    n1443,
    n2656,
    n2660,
    n2728
  );


  nor
  g2749
  (
    n2752,
    n2740,
    n2669,
    n2735,
    n2664
  );


  nand
  g2750
  (
    n2774,
    n2666,
    n2653,
    n2735
  );


  xor
  g2751
  (
    n2747,
    n2667,
    n2739,
    n2733,
    n2663
  );


  not
  g2752
  (
    n2835,
    n1461
  );


  buf
  g2753
  (
    n2846,
    n1449
  );


  buf
  g2754
  (
    n2898,
    n2776
  );


  buf
  g2755
  (
    n2848,
    n2764
  );


  not
  g2756
  (
    n2852,
    n1466
  );


  buf
  g2757
  (
    n2873,
    n2754
  );


  not
  g2758
  (
    n2795,
    n2683
  );


  not
  g2759
  (
    n2786,
    n279
  );


  buf
  g2760
  (
    n2804,
    n1457
  );


  not
  g2761
  (
    n2794,
    n1323
  );


  not
  g2762
  (
    n2792,
    n280
  );


  not
  g2763
  (
    n2829,
    n2692
  );


  not
  g2764
  (
    n2808,
    n1465
  );


  not
  g2765
  (
    n2904,
    n2691
  );


  buf
  g2766
  (
    n2907,
    n1459
  );


  buf
  g2767
  (
    n2840,
    n955
  );


  not
  g2768
  (
    n2915,
    n2762
  );


  not
  g2769
  (
    n2796,
    n2745
  );


  buf
  g2770
  (
    n2789,
    n1330
  );


  buf
  g2771
  (
    n2924,
    n1455
  );


  not
  g2772
  (
    n2875,
    n2595
  );


  not
  g2773
  (
    n2809,
    n1334
  );


  not
  g2774
  (
    n2903,
    n1449
  );


  not
  g2775
  (
    n2879,
    n2780
  );


  not
  g2776
  (
    n2860,
    n2695
  );


  buf
  g2777
  (
    n2928,
    n2697
  );


  not
  g2778
  (
    n2891,
    n2699
  );


  not
  g2779
  (
    n2830,
    n2697
  );


  buf
  g2780
  (
    n2921,
    n2684
  );


  buf
  g2781
  (
    n2871,
    n2687
  );


  buf
  g2782
  (
    n2837,
    n1460
  );


  buf
  g2783
  (
    n2853,
    n1333
  );


  buf
  g2784
  (
    n2895,
    n2774
  );


  buf
  g2785
  (
    n2888,
    n2592
  );


  not
  g2786
  (
    n2925,
    n2696
  );


  buf
  g2787
  (
    n2920,
    n2748
  );


  buf
  g2788
  (
    n2845,
    n80
  );


  buf
  g2789
  (
    n2843,
    n1465
  );


  buf
  g2790
  (
    n2831,
    n1445
  );


  buf
  g2791
  (
    n2896,
    n956
  );


  not
  g2792
  (
    n2785,
    n1464
  );


  not
  g2793
  (
    n2934,
    n2753
  );


  buf
  g2794
  (
    n2803,
    n2773
  );


  buf
  g2795
  (
    n2890,
    n2771
  );


  not
  g2796
  (
    n2844,
    n2746
  );


  buf
  g2797
  (
    n2828,
    n2690
  );


  not
  g2798
  (
    n2824,
    n2783
  );


  buf
  g2799
  (
    n2936,
    n2749
  );


  buf
  g2800
  (
    n2814,
    n2745
  );


  buf
  g2801
  (
    n2857,
    n2772
  );


  buf
  g2802
  (
    n2894,
    n1458
  );


  not
  g2803
  (
    n2790,
    n2761
  );


  buf
  g2804
  (
    n2869,
    n2695
  );


  buf
  g2805
  (
    n2849,
    n278
  );


  not
  g2806
  (
    n2821,
    n2589
  );


  not
  g2807
  (
    n2932,
    n2759
  );


  buf
  g2808
  (
    n2851,
    n2688
  );


  buf
  g2809
  (
    n2923,
    n2697
  );


  buf
  g2810
  (
    n2867,
    n1458
  );


  not
  g2811
  (
    n2862,
    n1456
  );


  buf
  g2812
  (
    n2842,
    n2684
  );


  buf
  g2813
  (
    n2818,
    n2777
  );


  not
  g2814
  (
    n2900,
    n1446
  );


  buf
  g2815
  (
    n2834,
    n277
  );


  xnor
  g2816
  (
    n2820,
    n2750,
    n1454,
    n1464,
    n277
  );


  xor
  g2817
  (
    n2816,
    n2754,
    n2779,
    n2784,
    n80
  );


  xnor
  g2818
  (
    n2905,
    n1451,
    n1451,
    n2744,
    n1448
  );


  or
  g2819
  (
    n2791,
    n2688,
    n2778,
    n956,
    n1455
  );


  xnor
  g2820
  (
    n2897,
    n1324,
    n2691,
    n2760,
    n80
  );


  and
  g2821
  (
    n2931,
    n2757,
    n2692,
    n2694,
    n1466
  );


  nor
  g2822
  (
    n2918,
    n2779,
    n1331,
    n2640,
    n2686
  );


  and
  g2823
  (
    n2870,
    n2756,
    n2782,
    n957,
    n2774
  );


  xnor
  g2824
  (
    n2807,
    n2767,
    n2752,
    n1454,
    n1456
  );


  nand
  g2825
  (
    n2832,
    n1451,
    n2686,
    n956,
    n2757
  );


  nand
  g2826
  (
    n2910,
    n276,
    n2755,
    n2691
  );


  or
  g2827
  (
    n2864,
    n1446,
    n2688,
    n2764,
    n2689
  );


  or
  g2828
  (
    n2926,
    n2743,
    n2761,
    n1366,
    n1328
  );


  nor
  g2829
  (
    n2806,
    n2641,
    n2764,
    n2753,
    n278
  );


  or
  g2830
  (
    n2868,
    n2766,
    n2762,
    n2768,
    n1320
  );


  or
  g2831
  (
    n2911,
    n2759,
    n2683,
    n1464,
    n1450
  );


  nor
  g2832
  (
    n2863,
    n2777,
    n2780,
    n2753,
    n2771
  );


  xor
  g2833
  (
    n2854,
    n2755,
    n2593,
    n1366,
    n2685
  );


  nand
  g2834
  (
    n2788,
    n2683,
    n2695,
    n2776,
    n278
  );


  nand
  g2835
  (
    n2839,
    n2768,
    n2699,
    n957,
    n1464
  );


  or
  g2836
  (
    n2901,
    n2698,
    n2748,
    n277,
    n2757
  );


  or
  g2837
  (
    n2819,
    n81,
    n280,
    n2751,
    n2763
  );


  xor
  g2838
  (
    n2793,
    n2749,
    n2767,
    n955,
    n2692
  );


  nand
  g2839
  (
    n2880,
    n281,
    n2681,
    n2784,
    n2754
  );


  xnor
  g2840
  (
    n2865,
    n1326,
    n1452,
    n2679,
    n2747
  );


  xnor
  g2841
  (
    n2906,
    n1459,
    n2763,
    n2699,
    n2783
  );


  xor
  g2842
  (
    n2817,
    n1332,
    n2686,
    n2689,
    n2773
  );


  and
  g2843
  (
    n2855,
    n2755,
    n2681,
    n2770,
    n2747
  );


  and
  g2844
  (
    n2833,
    n1321,
    n1462,
    n1446,
    n2642
  );


  xnor
  g2845
  (
    n2876,
    n2760,
    n2746,
    n2590,
    n2745
  );


  xnor
  g2846
  (
    n2877,
    n2689,
    n2775,
    n2758,
    n1449
  );


  or
  g2847
  (
    n2935,
    n2763,
    n1460,
    n1322,
    n2744
  );


  xnor
  g2848
  (
    n2927,
    n2765,
    n2680,
    n2761,
    n958
  );


  xnor
  g2849
  (
    n2885,
    n1463,
    n82,
    n2699,
    n2745
  );


  xnor
  g2850
  (
    n2799,
    n2782,
    n1463,
    n1446,
    n2784
  );


  or
  g2851
  (
    n2850,
    n1447,
    n2766,
    n1450,
    n1458
  );


  xnor
  g2852
  (
    n2827,
    n2682,
    n1447,
    n1366,
    n2743
  );


  xnor
  g2853
  (
    n2859,
    n2778,
    n958,
    n2756,
    n280
  );


  or
  g2854
  (
    n2823,
    n1463,
    n2693,
    n2774,
    n2766
  );


  xor
  g2855
  (
    n2914,
    n1451,
    n1459,
    n2750,
    n2772
  );


  and
  g2856
  (
    n2913,
    n2777,
    n1457,
    n2697,
    n279
  );


  or
  g2857
  (
    n2797,
    n1465,
    n2780,
    n2778,
    n2694
  );


  and
  g2858
  (
    n2893,
    n2747,
    n2779,
    n1366,
    n1462
  );


  or
  g2859
  (
    n2919,
    n2751,
    n2775,
    n2750,
    n2769
  );


  xor
  g2860
  (
    n2902,
    n1452,
    n1453,
    n2783,
    n2758
  );


  nand
  g2861
  (
    n2882,
    n279,
    n2779,
    n2769,
    n276
  );


  xnor
  g2862
  (
    n2922,
    n958,
    n2698,
    n2781,
    n2690
  );


  xor
  g2863
  (
    n2874,
    n2772,
    n1450,
    n2641,
    n2680
  );


  xor
  g2864
  (
    n2802,
    n2771,
    n2756,
    n955,
    n2744
  );


  and
  g2865
  (
    n2841,
    n1457,
    n2769,
    n1455,
    n2770
  );


  nand
  g2866
  (
    n2847,
    n276,
    n2750,
    n2759,
    n1448
  );


  or
  g2867
  (
    n2825,
    n1463,
    n2696,
    n1462
  );


  nand
  g2868
  (
    n2822,
    n2762,
    n2692,
    n2755,
    n2684
  );


  and
  g2869
  (
    n2826,
    n80,
    n2758,
    n2698,
    n1448
  );


  and
  g2870
  (
    n2892,
    n2681,
    n1452,
    n2693,
    n2680
  );


  xor
  g2871
  (
    n2798,
    n2749,
    n957,
    n2751,
    n1453
  );


  nand
  g2872
  (
    n2856,
    n1465,
    n956,
    n2694,
    n2772
  );


  or
  g2873
  (
    n2858,
    n2774,
    n2743,
    n1447
  );


  and
  g2874
  (
    n2912,
    n2749,
    n2758,
    n1459,
    n2729
  );


  nand
  g2875
  (
    n2812,
    n2679,
    n2782,
    n1456,
    n2698
  );


  nor
  g2876
  (
    n2861,
    n1460,
    n1457,
    n2748,
    n1461
  );


  or
  g2877
  (
    n2787,
    n2767,
    n2773,
    n2687,
    n2680
  );


  xor
  g2878
  (
    n2889,
    n2729,
    n2770,
    n1461,
    n2682
  );


  xor
  g2879
  (
    n2930,
    n280,
    n2761,
    n1455,
    n2773
  );


  nand
  g2880
  (
    n2933,
    n2684,
    n2765,
    n2759,
    n1454
  );


  xnor
  g2881
  (
    n2800,
    n1325,
    n1449,
    n2762,
    n2696
  );


  nand
  g2882
  (
    n2884,
    n958,
    n2752,
    n2757,
    n81
  );


  nor
  g2883
  (
    n2916,
    n81,
    n277,
    n1466,
    n1462
  );


  xor
  g2884
  (
    n2838,
    n2746,
    n2766,
    n2771,
    n2690
  );


  or
  g2885
  (
    n2811,
    n1453,
    n2687,
    n2683,
    n2686
  );


  nor
  g2886
  (
    n2908,
    n2765,
    n1453,
    n81,
    n2770
  );


  and
  g2887
  (
    n2866,
    n2642,
    n2765,
    n2694,
    n2682
  );


  xor
  g2888
  (
    n2801,
    n1456,
    n2780,
    n2695,
    n957
  );


  xnor
  g2889
  (
    n2929,
    n2744,
    n1445,
    n1447,
    n2776
  );


  or
  g2890
  (
    n2917,
    n1452,
    n2775,
    n2748
  );


  or
  g2891
  (
    n2881,
    n2776,
    n1461,
    n2752,
    n2693
  );


  or
  g2892
  (
    n2899,
    n2781,
    n2769,
    n2682,
    n2688
  );


  and
  g2893
  (
    n2815,
    n2767,
    n2782,
    n2756,
    n1448
  );


  nor
  g2894
  (
    n2887,
    n2746,
    n2752,
    n2591,
    n2693
  );


  nor
  g2895
  (
    n2878,
    n2760,
    n2687,
    n1445,
    n1460
  );


  or
  g2896
  (
    n2909,
    n2754,
    n2764,
    n1454,
    n1450
  );


  xnor
  g2897
  (
    n2810,
    n2751,
    n2690,
    n2768,
    n2594
  );


  or
  g2898
  (
    n2805,
    n2781,
    n2760,
    n2685,
    n2763
  );


  xor
  g2899
  (
    n2883,
    n1327,
    n2689,
    n2685,
    n278
  );


  nand
  g2900
  (
    n2836,
    n2681,
    n2588,
    n1466,
    n2784
  );


  xnor
  g2901
  (
    n2886,
    n279,
    n2753,
    n2777,
    n2781
  );


  xnor
  g2902
  (
    n2813,
    n2778,
    n955,
    n2685,
    n2747
  );


  xnor
  g2903
  (
    n2872,
    n1458,
    n2783,
    n1329,
    n2768
  );


  xor
  g2904
  (
    n2954,
    n2799,
    n2813,
    n2847,
    n2901
  );


  nor
  g2905
  (
    n2943,
    n2806,
    n2829,
    n2885,
    n2935
  );


  nand
  g2906
  (
    n2969,
    n2851,
    n2830,
    n2878,
    n2870
  );


  xnor
  g2907
  (
    n2952,
    n2845,
    n2865,
    n2869,
    n2820
  );


  nor
  g2908
  (
    n2951,
    n20,
    n2906,
    n2924,
    n2911
  );


  xor
  g2909
  (
    n2947,
    n17,
    n2828,
    n2801,
    n2922
  );


  xnor
  g2910
  (
    n2975,
    n2805,
    n2825,
    n2797,
    n2826
  );


  xor
  g2911
  (
    n2966,
    n2900,
    n2792,
    n2863,
    n2816
  );


  or
  g2912
  (
    n2979,
    n2796,
    n2929,
    n2867,
    n2852
  );


  nor
  g2913
  (
    n2978,
    n2822,
    n2807,
    n2888,
    n2862
  );


  xnor
  g2914
  (
    n2972,
    n2894,
    n2899,
    n2871,
    n2932
  );


  xor
  g2915
  (
    n2956,
    n2819,
    n2927,
    n2883,
    n2858
  );


  nor
  g2916
  (
    n2942,
    n2926,
    n2872,
    n2884,
    n2785
  );


  and
  g2917
  (
    n2941,
    n2879,
    n2896,
    n2890,
    n2902
  );


  nand
  g2918
  (
    n2948,
    n2930,
    n2912,
    n2925,
    n18
  );


  nor
  g2919
  (
    n2959,
    n2920,
    n2812,
    n2895,
    n21
  );


  xor
  g2920
  (
    n2945,
    n2877,
    n2892,
    n2891,
    n21
  );


  nand
  g2921
  (
    n2938,
    n2856,
    n2860,
    n2849,
    n2931
  );


  xnor
  g2922
  (
    n2939,
    n2841,
    n2903,
    n2889,
    n2843
  );


  nand
  g2923
  (
    n2971,
    n2848,
    n82,
    n2803,
    n2850
  );


  or
  g2924
  (
    n2944,
    n2875,
    n2793,
    n2836,
    n2842
  );


  nand
  g2925
  (
    n2953,
    n2923,
    n2802,
    n2918,
    n2853
  );


  xnor
  g2926
  (
    n2940,
    n17,
    n2817,
    n2789,
    n2874
  );


  and
  g2927
  (
    n2965,
    n2839,
    n2790,
    n20,
    n2934
  );


  nand
  g2928
  (
    n2973,
    n2818,
    n2897,
    n2837,
    n2916
  );


  xor
  g2929
  (
    n2960,
    n2846,
    n2855,
    n2913,
    n2905
  );


  nor
  g2930
  (
    n2955,
    n2919,
    n2873,
    n2810,
    n2834
  );


  xnor
  g2931
  (
    n2963,
    n20,
    n2787,
    n2910,
    n2886
  );


  xnor
  g2932
  (
    n2961,
    n19,
    n2887,
    n21,
    n18
  );


  or
  g2933
  (
    n2976,
    n2838,
    n2824,
    n2811,
    n2786
  );


  xnor
  g2934
  (
    n2967,
    n19,
    n2880,
    n2882,
    n2832
  );


  and
  g2935
  (
    n2950,
    n2933,
    n2840,
    n2904,
    n2808
  );


  nand
  g2936
  (
    n2968,
    n2893,
    n2936,
    n2833,
    n2794
  );


  xnor
  g2937
  (
    n2974,
    n2791,
    n2917,
    n2831,
    n2914
  );


  or
  g2938
  (
    n2949,
    n18,
    n2815,
    n2729,
    n2876
  );


  nand
  g2939
  (
    n2937,
    n2798,
    n18,
    n2907,
    n2835
  );


  or
  g2940
  (
    n2958,
    n2868,
    n2821,
    n2844,
    n2800
  );


  and
  g2941
  (
    n2946,
    n2827,
    n2729,
    n19,
    n2921
  );


  or
  g2942
  (
    n2977,
    n2823,
    n2864,
    n2908,
    n19
  );


  nor
  g2943
  (
    n2962,
    n20,
    n2909,
    n2928,
    n2809
  );


  xor
  g2944
  (
    n2964,
    n2795,
    n2788,
    n2814,
    n2854
  );


  xnor
  g2945
  (
    n2957,
    n2881,
    n2804,
    n2857,
    n2861
  );


  xor
  g2946
  (
    n2970,
    n2915,
    n2898,
    n2859,
    n2866
  );


  xnor
  g2947
  (
    n2981,
    n2975,
    n2958,
    n2968,
    n2944
  );


  xor
  g2948
  (
    n2985,
    n2963,
    n2964,
    n2969,
    n2962
  );


  xnor
  g2949
  (
    n2984,
    n2938,
    n2959,
    n2945,
    n2965
  );


  nor
  g2950
  (
    n2983,
    n2941,
    n2951,
    n2947,
    n2956
  );


  nor
  g2951
  (
    n2980,
    n2967,
    n2943,
    n2955,
    n2960
  );


  or
  g2952
  (
    n2986,
    n2949,
    n2937,
    n2950,
    n2952
  );


  or
  g2953
  (
    AntiSAT_key_wire,
    n2954,
    n2948,
    n2976,
    n2972
  );


  or
  g2954
  (
    n2982,
    n2961,
    n2940,
    n2939,
    n2953
  );


  xor
  g2955
  (
    n2987,
    n2971,
    n2970,
    n2957,
    n2973
  );


  nor
  g2956
  (
    n2989,
    n2966,
    n2946,
    n2942,
    n2974
  );


  or
  g2957
  (
    n2990,
    n2989,
    n281
  );


  xor
  g2958
  (
    n2992,
    n961,
    n960
  );


  nor
  g2959
  (
    n2991,
    n959,
    n2990,
    n961
  );


  xnor
  g2960
  (
    n2994,
    n2990,
    n959
  );


  and
  g2961
  (
    n2993,
    n961,
    n961,
    n2990,
    n960
  );


  nand
  g2962
  (
    n2997,
    n2992,
    n27,
    n2991,
    n26
  );


  or
  g2963
  (
    n2996,
    n25,
    n25,
    n30,
    n2994
  );


  nor
  g2964
  (
    n3000,
    n29,
    n28,
    n27,
    n2993
  );


  nor
  g2965
  (
    n3005,
    n32,
    n32,
    n2994,
    n2978
  );


  nand
  g2966
  (
    n3002,
    n2993,
    n2994,
    n2992,
    n28
  );


  nand
  g2967
  (
    n3009,
    n29,
    n26,
    n2992
  );


  or
  g2968
  (
    n2999,
    n32,
    n2993,
    n26,
    n31
  );


  or
  g2969
  (
    n3004,
    n2991,
    n27,
    n24
  );


  nand
  g2970
  (
    n2998,
    n2991,
    n22,
    n2994,
    n26
  );


  and
  g2971
  (
    n3007,
    n32,
    n28,
    n30,
    n23
  );


  xor
  g2972
  (
    n2995,
    n22,
    n24,
    n2993,
    n31
  );


  xor
  g2973
  (
    n3010,
    n21,
    n23,
    n24,
    n22
  );


  or
  g2974
  (
    n3003,
    n2991,
    n30,
    n24
  );


  nand
  g2975
  (
    n3006,
    n2977,
    n29,
    n23,
    n2979
  );


  xor
  g2976
  (
    n3001,
    n31,
    n22,
    n23,
    n29
  );


  and
  g2977
  (
    n3008,
    n31,
    n25,
    n28
  );


  or
  g2978
  (
    n3019,
    n96,
    n3008,
    n2995,
    n86
  );


  xor
  g2979
  (
    n3017,
    n83,
    n86,
    n82,
    n3004
  );


  or
  g2980
  (
    n3027,
    n2996,
    n93,
    n83,
    n92
  );


  xnor
  g2981
  (
    n3026,
    n97,
    n87,
    n3006,
    n92
  );


  nor
  g2982
  (
    n3025,
    n3002,
    n3003,
    n97,
    n82
  );


  xor
  g2983
  (
    n3012,
    n2998,
    n93,
    n96,
    n95
  );


  nor
  g2984
  (
    n3023,
    n89,
    n90,
    n98,
    n85
  );


  nor
  g2985
  (
    n3015,
    n96,
    n94,
    n3007,
    n90
  );


  nor
  g2986
  (
    n3024,
    n85,
    n91,
    n89,
    n86
  );


  nand
  g2987
  (
    n3018,
    n98,
    n90,
    n84,
    n3006
  );


  and
  g2988
  (
    n3011,
    n83,
    n3010,
    n3001,
    n3007
  );


  and
  g2989
  (
    n3028,
    n93,
    n84,
    n3005,
    n83
  );


  xor
  g2990
  (
    n3020,
    n85,
    n84,
    n3008,
    n3009
  );


  xor
  g2991
  (
    n3032,
    n2999,
    n92,
    n90,
    n84
  );


  nor
  g2992
  (
    n3022,
    n87,
    n86,
    n88,
    n94
  );


  nand
  g2993
  (
    n3016,
    n91,
    n3005,
    n98,
    n94
  );


  or
  g2994
  (
    n3013,
    n91,
    n95
  );


  or
  g2995
  (
    n3029,
    n3010,
    n3009,
    n94,
    n89
  );


  nand
  g2996
  (
    n3030,
    n96,
    n93,
    n88,
    n89
  );


  nand
  g2997
  (
    n3014,
    n98,
    n87,
    n97
  );


  or
  g2998
  (
    n3021,
    n91,
    n92,
    n2997,
    n85
  );


  xnor
  g2999
  (
    n3031,
    n3000,
    n88,
    n87
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n2988,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

