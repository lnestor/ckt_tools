

module Stat_2000_312
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n774,
  n765,
  n826,
  n825,
  n828,
  n819,
  n830,
  n818,
  n824,
  n2015,
  n2011,
  n2029,
  n2014,
  n2030,
  n2022,
  n2017,
  n2021,
  n2023,
  n2013,
  n2019,
  n2018,
  n2020,
  n2032,
  n2028,
  n2026,
  n2010,
  n2025,
  n2027,
  n2024,
  n2016,
  n2012,
  n2031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n774;output n765;output n826;output n825;output n828;output n819;output n830;output n818;output n824;output n2015;output n2011;output n2029;output n2014;output n2030;output n2022;output n2017;output n2021;output n2023;output n2013;output n2019;output n2018;output n2020;output n2032;output n2028;output n2026;output n2010;output n2025;output n2027;output n2024;output n2016;output n2012;output n2031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n820;wire n821;wire n822;wire n823;wire n827;wire n829;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n35,
    n1
  );


  buf
  g1
  (
    n45,
    n5
  );


  not
  g2
  (
    n39,
    n5
  );


  buf
  g3
  (
    n34,
    n2
  );


  buf
  g4
  (
    n42,
    n3
  );


  not
  g5
  (
    KeyWire_0_22,
    n1
  );


  buf
  g6
  (
    KeyWire_0_12,
    n3
  );


  buf
  g7
  (
    n38,
    n4
  );


  buf
  g8
  (
    n46,
    n4
  );


  not
  g9
  (
    n40,
    n2
  );


  not
  g10
  (
    n44,
    n4
  );


  buf
  g11
  (
    n33,
    n5
  );


  buf
  g12
  (
    n47,
    n4
  );


  not
  g13
  (
    n37,
    n2
  );


  buf
  g14
  (
    n43,
    n3
  );


  buf
  g15
  (
    n75,
    n43
  );


  not
  g16
  (
    n77,
    n40
  );


  not
  g17
  (
    n82,
    n41
  );


  buf
  g18
  (
    n86,
    n44
  );


  not
  g19
  (
    n92,
    n39
  );


  not
  g20
  (
    n67,
    n43
  );


  not
  g21
  (
    n80,
    n42
  );


  buf
  g22
  (
    n49,
    n35
  );


  buf
  g23
  (
    n79,
    n44
  );


  not
  g24
  (
    n48,
    n42
  );


  not
  g25
  (
    n76,
    n34
  );


  buf
  g26
  (
    n64,
    n36
  );


  buf
  g27
  (
    n90,
    n42
  );


  not
  g28
  (
    n61,
    n33
  );


  not
  g29
  (
    n63,
    n36
  );


  not
  g30
  (
    n52,
    n39
  );


  buf
  g31
  (
    n78,
    n37
  );


  buf
  g32
  (
    n91,
    n40
  );


  buf
  g33
  (
    n50,
    n37
  );


  not
  g34
  (
    n83,
    n41
  );


  not
  g35
  (
    n62,
    n35
  );


  not
  g36
  (
    n53,
    n36
  );


  not
  g37
  (
    n51,
    n38
  );


  buf
  g38
  (
    n56,
    n40
  );


  not
  g39
  (
    n84,
    n34
  );


  buf
  g40
  (
    n72,
    n44
  );


  not
  g41
  (
    n73,
    n38
  );


  buf
  g42
  (
    n89,
    n33
  );


  buf
  g43
  (
    n88,
    n44
  );


  not
  g44
  (
    n87,
    n39
  );


  buf
  g45
  (
    n66,
    n39
  );


  buf
  g46
  (
    n69,
    n33
  );


  buf
  g47
  (
    n85,
    n37
  );


  buf
  g48
  (
    n58,
    n40
  );


  not
  g49
  (
    n68,
    n34
  );


  not
  g50
  (
    n74,
    n35
  );


  buf
  g51
  (
    n81,
    n43
  );


  buf
  g52
  (
    n54,
    n38
  );


  not
  g53
  (
    n57,
    n41
  );


  not
  g54
  (
    n60,
    n37
  );


  buf
  g55
  (
    n59,
    n43
  );


  not
  g56
  (
    n65,
    n41
  );


  not
  g57
  (
    n70,
    n38
  );


  buf
  g58
  (
    n71,
    n42
  );


  buf
  g59
  (
    n55,
    n36
  );


  not
  g60
  (
    n143,
    n74
  );


  not
  g61
  (
    n233,
    n55
  );


  buf
  g62
  (
    n262,
    n51
  );


  not
  g63
  (
    n147,
    n91
  );


  not
  g64
  (
    n234,
    n66
  );


  buf
  g65
  (
    n129,
    n63
  );


  buf
  g66
  (
    n106,
    n59
  );


  not
  g67
  (
    n207,
    n92
  );


  not
  g68
  (
    n134,
    n50
  );


  not
  g69
  (
    n167,
    n72
  );


  buf
  g70
  (
    n109,
    n78
  );


  buf
  g71
  (
    n182,
    n66
  );


  not
  g72
  (
    n214,
    n49
  );


  not
  g73
  (
    n241,
    n84
  );


  not
  g74
  (
    n127,
    n68
  );


  not
  g75
  (
    n261,
    n79
  );


  buf
  g76
  (
    n191,
    n60
  );


  not
  g77
  (
    n126,
    n92
  );


  not
  g78
  (
    n166,
    n89
  );


  not
  g79
  (
    n260,
    n57
  );


  not
  g80
  (
    n146,
    n64
  );


  not
  g81
  (
    n218,
    n76
  );


  not
  g82
  (
    n144,
    n70
  );


  not
  g83
  (
    n231,
    n78
  );


  buf
  g84
  (
    n247,
    n86
  );


  buf
  g85
  (
    n217,
    n87
  );


  not
  g86
  (
    n205,
    n51
  );


  not
  g87
  (
    n152,
    n81
  );


  buf
  g88
  (
    n265,
    n89
  );


  buf
  g89
  (
    n193,
    n60
  );


  buf
  g90
  (
    n200,
    n80
  );


  buf
  g91
  (
    n99,
    n71
  );


  not
  g92
  (
    n169,
    n86
  );


  buf
  g93
  (
    n232,
    n80
  );


  not
  g94
  (
    n229,
    n64
  );


  buf
  g95
  (
    n270,
    n53
  );


  buf
  g96
  (
    n239,
    n48
  );


  buf
  g97
  (
    n245,
    n71
  );


  buf
  g98
  (
    n184,
    n82
  );


  buf
  g99
  (
    n131,
    n88
  );


  buf
  g100
  (
    n158,
    n82
  );


  buf
  g101
  (
    n170,
    n91
  );


  not
  g102
  (
    n257,
    n60
  );


  buf
  g103
  (
    n165,
    n56
  );


  not
  g104
  (
    n151,
    n80
  );


  not
  g105
  (
    n115,
    n88
  );


  buf
  g106
  (
    n135,
    n76
  );


  buf
  g107
  (
    n221,
    n61
  );


  not
  g108
  (
    n112,
    n72
  );


  not
  g109
  (
    n153,
    n92
  );


  not
  g110
  (
    n216,
    n58
  );


  buf
  g111
  (
    n102,
    n56
  );


  not
  g112
  (
    n240,
    n73
  );


  not
  g113
  (
    n180,
    n50
  );


  buf
  g114
  (
    n155,
    n54
  );


  buf
  g115
  (
    n256,
    n69
  );


  buf
  g116
  (
    n246,
    n87
  );


  not
  g117
  (
    n192,
    n68
  );


  buf
  g118
  (
    n157,
    n55
  );


  buf
  g119
  (
    n150,
    n55
  );


  not
  g120
  (
    n111,
    n58
  );


  not
  g121
  (
    n228,
    n75
  );


  not
  g122
  (
    n168,
    n89
  );


  not
  g123
  (
    n138,
    n79
  );


  not
  g124
  (
    n238,
    n61
  );


  not
  g125
  (
    n121,
    n82
  );


  not
  g126
  (
    n142,
    n81
  );


  not
  g127
  (
    n101,
    n52
  );


  buf
  g128
  (
    n195,
    n74
  );


  not
  g129
  (
    n271,
    n48
  );


  buf
  g130
  (
    n227,
    n48
  );


  buf
  g131
  (
    n161,
    n90
  );


  buf
  g132
  (
    n237,
    n89
  );


  not
  g133
  (
    n178,
    n52
  );


  buf
  g134
  (
    n242,
    n70
  );


  not
  g135
  (
    n117,
    n67
  );


  buf
  g136
  (
    n204,
    n54
  );


  not
  g137
  (
    n212,
    n50
  );


  not
  g138
  (
    n176,
    n68
  );


  buf
  g139
  (
    KeyWire_0_28,
    n88
  );


  not
  g140
  (
    n114,
    n49
  );


  buf
  g141
  (
    n213,
    n58
  );


  buf
  g142
  (
    n203,
    n57
  );


  buf
  g143
  (
    n201,
    n63
  );


  buf
  g144
  (
    n268,
    n72
  );


  buf
  g145
  (
    n266,
    n49
  );


  buf
  g146
  (
    n98,
    n71
  );


  not
  g147
  (
    n133,
    n84
  );


  buf
  g148
  (
    n226,
    n61
  );


  not
  g149
  (
    n199,
    n88
  );


  buf
  g150
  (
    n253,
    n50
  );


  buf
  g151
  (
    n97,
    n57
  );


  buf
  g152
  (
    n105,
    n69
  );


  not
  g153
  (
    n194,
    n75
  );


  buf
  g154
  (
    n224,
    n86
  );


  not
  g155
  (
    n250,
    n48
  );


  buf
  g156
  (
    n136,
    n73
  );


  not
  g157
  (
    n190,
    n58
  );


  buf
  g158
  (
    n210,
    n84
  );


  buf
  g159
  (
    n255,
    n81
  );


  not
  g160
  (
    n252,
    n90
  );


  not
  g161
  (
    n244,
    n56
  );


  not
  g162
  (
    n185,
    n91
  );


  buf
  g163
  (
    n179,
    n62
  );


  buf
  g164
  (
    n94,
    n79
  );


  not
  g165
  (
    n107,
    n69
  );


  not
  g166
  (
    n122,
    n78
  );


  not
  g167
  (
    n202,
    n73
  );


  buf
  g168
  (
    n230,
    n62
  );


  not
  g169
  (
    n162,
    n81
  );


  buf
  g170
  (
    n160,
    n80
  );


  buf
  g171
  (
    n243,
    n87
  );


  buf
  g172
  (
    n215,
    n82
  );


  buf
  g173
  (
    n181,
    n74
  );


  not
  g174
  (
    n159,
    n90
  );


  buf
  g175
  (
    n124,
    n66
  );


  buf
  g176
  (
    n140,
    n74
  );


  buf
  g177
  (
    KeyWire_0_23,
    n54
  );


  buf
  g178
  (
    n104,
    n85
  );


  buf
  g179
  (
    n128,
    n62
  );


  not
  g180
  (
    n103,
    n67
  );


  not
  g181
  (
    n220,
    n51
  );


  buf
  g182
  (
    n100,
    n63
  );


  buf
  g183
  (
    n141,
    n69
  );


  not
  g184
  (
    n164,
    n52
  );


  not
  g185
  (
    n236,
    n53
  );


  buf
  g186
  (
    n183,
    n77
  );


  not
  g187
  (
    n148,
    n83
  );


  not
  g188
  (
    n174,
    n70
  );


  not
  g189
  (
    n110,
    n67
  );


  buf
  g190
  (
    n196,
    n83
  );


  not
  g191
  (
    n163,
    n52
  );


  not
  g192
  (
    n258,
    n75
  );


  buf
  g193
  (
    n132,
    n90
  );


  not
  g194
  (
    n264,
    n64
  );


  not
  g195
  (
    n267,
    n59
  );


  buf
  g196
  (
    n108,
    n87
  );


  not
  g197
  (
    n130,
    n51
  );


  not
  g198
  (
    n208,
    n83
  );


  not
  g199
  (
    n154,
    n55
  );


  not
  g200
  (
    n95,
    n73
  );


  buf
  g201
  (
    n177,
    n65
  );


  buf
  g202
  (
    n156,
    n86
  );


  not
  g203
  (
    n123,
    n65
  );


  not
  g204
  (
    n211,
    n77
  );


  not
  g205
  (
    n259,
    n72
  );


  not
  g206
  (
    n197,
    n53
  );


  buf
  g207
  (
    n186,
    n54
  );


  buf
  g208
  (
    n263,
    n84
  );


  buf
  g209
  (
    n113,
    n75
  );


  buf
  g210
  (
    n145,
    n78
  );


  not
  g211
  (
    n173,
    n83
  );


  not
  g212
  (
    n225,
    n71
  );


  buf
  g213
  (
    n116,
    n85
  );


  buf
  g214
  (
    n209,
    n77
  );


  buf
  g215
  (
    n269,
    n68
  );


  not
  g216
  (
    n254,
    n49
  );


  not
  g217
  (
    n219,
    n63
  );


  buf
  g218
  (
    n188,
    n62
  );


  buf
  g219
  (
    n120,
    n59
  );


  buf
  g220
  (
    n172,
    n60
  );


  not
  g221
  (
    n175,
    n79
  );


  not
  g222
  (
    n139,
    n76
  );


  buf
  g223
  (
    n248,
    n56
  );


  not
  g224
  (
    KeyWire_0_2,
    n85
  );


  not
  g225
  (
    n137,
    n59
  );


  not
  g226
  (
    n189,
    n91
  );


  not
  g227
  (
    n96,
    n77
  );


  buf
  g228
  (
    n125,
    n66
  );


  not
  g229
  (
    n249,
    n76
  );


  buf
  g230
  (
    n223,
    n67
  );


  not
  g231
  (
    n119,
    n61
  );


  not
  g232
  (
    n198,
    n57
  );


  not
  g233
  (
    n171,
    n85
  );


  not
  g234
  (
    n206,
    n64
  );


  not
  g235
  (
    n149,
    n53
  );


  not
  g236
  (
    n251,
    n65
  );


  not
  g237
  (
    n187,
    n70
  );


  not
  g238
  (
    n93,
    n65
  );


  not
  g239
  (
    n507,
    n19
  );


  buf
  g240
  (
    n405,
    n143
  );


  not
  g241
  (
    n291,
    n185
  );


  buf
  g242
  (
    n506,
    n11
  );


  buf
  g243
  (
    n314,
    n161
  );


  buf
  g244
  (
    n432,
    n26
  );


  not
  g245
  (
    n329,
    n254
  );


  not
  g246
  (
    n377,
    n217
  );


  buf
  g247
  (
    n439,
    n110
  );


  buf
  g248
  (
    n287,
    n202
  );


  not
  g249
  (
    n488,
    n211
  );


  buf
  g250
  (
    n353,
    n16
  );


  not
  g251
  (
    n486,
    n240
  );


  buf
  g252
  (
    n290,
    n136
  );


  buf
  g253
  (
    n400,
    n110
  );


  buf
  g254
  (
    n311,
    n96
  );


  buf
  g255
  (
    n416,
    n139
  );


  not
  g256
  (
    n478,
    n124
  );


  buf
  g257
  (
    n278,
    n124
  );


  buf
  g258
  (
    n414,
    n112
  );


  buf
  g259
  (
    n497,
    n253
  );


  buf
  g260
  (
    n344,
    n261
  );


  buf
  g261
  (
    n461,
    n256
  );


  not
  g262
  (
    n309,
    n126
  );


  buf
  g263
  (
    n471,
    n25
  );


  not
  g264
  (
    n399,
    n122
  );


  buf
  g265
  (
    n464,
    n214
  );


  not
  g266
  (
    n318,
    n257
  );


  buf
  g267
  (
    n275,
    n107
  );


  not
  g268
  (
    n321,
    n176
  );


  not
  g269
  (
    n304,
    n252
  );


  buf
  g270
  (
    n474,
    n230
  );


  not
  g271
  (
    n482,
    n111
  );


  not
  g272
  (
    n450,
    n241
  );


  buf
  g273
  (
    n494,
    n196
  );


  not
  g274
  (
    n305,
    n22
  );


  buf
  g275
  (
    n342,
    n207
  );


  buf
  g276
  (
    n332,
    n213
  );


  buf
  g277
  (
    n327,
    n118
  );


  buf
  g278
  (
    n480,
    n213
  );


  not
  g279
  (
    n381,
    n179
  );


  not
  g280
  (
    n297,
    n205
  );


  not
  g281
  (
    n288,
    n164
  );


  not
  g282
  (
    n443,
    n110
  );


  not
  g283
  (
    n339,
    n124
  );


  buf
  g284
  (
    n300,
    n153
  );


  not
  g285
  (
    n364,
    n105
  );


  buf
  g286
  (
    n445,
    n204
  );


  buf
  g287
  (
    n387,
    n106
  );


  not
  g288
  (
    n501,
    n266
  );


  buf
  g289
  (
    n324,
    n195
  );


  buf
  g290
  (
    n453,
    n215
  );


  not
  g291
  (
    n352,
    n108
  );


  not
  g292
  (
    n379,
    n171
  );


  and
  g293
  (
    n415,
    n184,
    n199,
    n135
  );


  xnor
  g294
  (
    n365,
    n116,
    n188,
    n235,
    n237
  );


  or
  g295
  (
    n468,
    n248,
    n214,
    n16,
    n153
  );


  nand
  g296
  (
    n282,
    n146,
    n147,
    n127,
    n184
  );


  nand
  g297
  (
    n411,
    n156,
    n94,
    n174,
    n17
  );


  nand
  g298
  (
    n333,
    n255,
    n172,
    n162,
    n167
  );


  or
  g299
  (
    n383,
    n214,
    n118,
    n257,
    n99
  );


  nand
  g300
  (
    n449,
    n152,
    n242,
    n13,
    n155
  );


  nor
  g301
  (
    n407,
    n11,
    n178,
    n118,
    n263
  );


  or
  g302
  (
    n295,
    n267,
    n98,
    n264,
    n171
  );


  or
  g303
  (
    n397,
    n205,
    n109,
    n99,
    n10
  );


  xnor
  g304
  (
    n505,
    n269,
    n105,
    n182,
    n229
  );


  nor
  g305
  (
    n346,
    n106,
    n234,
    n210,
    n215
  );


  xor
  g306
  (
    n292,
    n130,
    n100,
    n135,
    n208
  );


  nor
  g307
  (
    n277,
    n216,
    n268,
    n225,
    n176
  );


  or
  g308
  (
    n463,
    n174,
    n9,
    n252,
    n231
  );


  or
  g309
  (
    n313,
    n259,
    n95,
    n12,
    n246
  );


  or
  g310
  (
    n391,
    n244,
    n10,
    n203,
    n156
  );


  xor
  g311
  (
    n354,
    n125,
    n179,
    n123,
    n104
  );


  xor
  g312
  (
    n472,
    n168,
    n150,
    n149,
    n129
  );


  xor
  g313
  (
    n499,
    n225,
    n235,
    n204,
    n158
  );


  and
  g314
  (
    n476,
    n119,
    n174,
    n189,
    n155
  );


  nor
  g315
  (
    n328,
    n265,
    n191,
    n226,
    n242
  );


  xnor
  g316
  (
    n452,
    n6,
    n189,
    n195,
    n151
  );


  nor
  g317
  (
    n429,
    n251,
    n9,
    n173,
    n15
  );


  nand
  g318
  (
    n487,
    n243,
    n97,
    n21,
    n251
  );


  xor
  g319
  (
    n437,
    n250,
    n15,
    n23,
    n256
  );


  nand
  g320
  (
    n440,
    n210,
    n219,
    n102,
    n22
  );


  nand
  g321
  (
    n441,
    n156,
    n238,
    n26,
    n111
  );


  nand
  g322
  (
    n459,
    n165,
    n158,
    n120,
    n222
  );


  or
  g323
  (
    n279,
    n205,
    n14,
    n213,
    n99
  );


  or
  g324
  (
    n294,
    n148,
    n123,
    n166,
    n200
  );


  xor
  g325
  (
    n317,
    n227,
    n115,
    n16,
    n20
  );


  or
  g326
  (
    n484,
    n214,
    n94,
    n202,
    n119
  );


  nand
  g327
  (
    n496,
    n220,
    n263,
    n144,
    n232
  );


  nand
  g328
  (
    n408,
    n190,
    n211,
    n144,
    n23
  );


  xor
  g329
  (
    n359,
    n207,
    n236,
    n241,
    n224
  );


  xor
  g330
  (
    n308,
    n136,
    n178,
    n248,
    n127
  );


  or
  g331
  (
    n373,
    n5,
    n132,
    n268,
    n203
  );


  xor
  g332
  (
    n375,
    n178,
    n253,
    n180,
    n164
  );


  xor
  g333
  (
    n285,
    n177,
    n149,
    n223,
    n217
  );


  nand
  g334
  (
    n331,
    n170,
    n22,
    n260,
    n177
  );


  nand
  g335
  (
    n418,
    n127,
    n211,
    n223,
    n266
  );


  xor
  g336
  (
    n276,
    n249,
    n127,
    n181,
    n183
  );


  xor
  g337
  (
    n369,
    n210,
    n109,
    n245,
    n113
  );


  nor
  g338
  (
    n508,
    n181,
    n247,
    n137,
    n201
  );


  or
  g339
  (
    n386,
    n258,
    n192,
    n149,
    n161
  );


  and
  g340
  (
    n503,
    n130,
    n9,
    n240,
    n255
  );


  nand
  g341
  (
    n362,
    n247,
    n262,
    n209,
    n134
  );


  nor
  g342
  (
    n372,
    n249,
    n169,
    n232,
    n11
  );


  xnor
  g343
  (
    n492,
    n162,
    n14,
    n154,
    n196
  );


  and
  g344
  (
    n356,
    n181,
    n264,
    n252,
    n166
  );


  and
  g345
  (
    n358,
    n133,
    n100,
    n245,
    n220
  );


  xor
  g346
  (
    n340,
    n143,
    n262,
    n102,
    n173
  );


  nor
  g347
  (
    n433,
    n141,
    n155,
    n234,
    n115
  );


  nand
  g348
  (
    n448,
    n254,
    n209,
    n126,
    n114
  );


  and
  g349
  (
    n500,
    n111,
    n193,
    n95,
    n211
  );


  or
  g350
  (
    n410,
    n142,
    n176,
    n259,
    n27
  );


  or
  g351
  (
    n402,
    n265,
    n175,
    n158,
    n181
  );


  and
  g352
  (
    n401,
    n114,
    n18,
    n109,
    n230
  );


  and
  g353
  (
    n396,
    n253,
    n125,
    n147,
    n170
  );


  nand
  g354
  (
    n296,
    n146,
    n18,
    n198,
    n103
  );


  nand
  g355
  (
    n462,
    n258,
    n142,
    n241,
    n111
  );


  nand
  g356
  (
    n302,
    n7,
    n131,
    n208,
    n267
  );


  xor
  g357
  (
    n335,
    n12,
    n141,
    n194,
    n262
  );


  xnor
  g358
  (
    n419,
    n160,
    n251,
    n169,
    n218
  );


  xnor
  g359
  (
    n322,
    n217,
    n107,
    n105,
    n195
  );


  xnor
  g360
  (
    KeyWire_0_14,
    n163,
    n231,
    n230,
    n139
  );


  xnor
  g361
  (
    n465,
    n97,
    n226,
    n21,
    n242
  );


  and
  g362
  (
    n427,
    n167,
    n19,
    n172,
    n141
  );


  xnor
  g363
  (
    n320,
    n150,
    n185,
    n157,
    n264
  );


  and
  g364
  (
    n510,
    n266,
    n165,
    n135,
    n120
  );


  and
  g365
  (
    n430,
    n172,
    n268,
    n236,
    n148
  );


  xor
  g366
  (
    n436,
    n103,
    n198,
    n163,
    n221
  );


  nand
  g367
  (
    n435,
    n242,
    n101,
    n16,
    n239
  );


  nand
  g368
  (
    n404,
    n221,
    n147,
    n125,
    n117
  );


  xnor
  g369
  (
    n451,
    n190,
    n17,
    n208,
    n20
  );


  xor
  g370
  (
    n394,
    n183,
    n235,
    n140,
    n244
  );


  or
  g371
  (
    n485,
    n243,
    n260,
    n226,
    n218
  );


  nand
  g372
  (
    n456,
    n187,
    n265,
    n23,
    n143
  );


  or
  g373
  (
    n495,
    n124,
    n219,
    n137,
    n113
  );


  xor
  g374
  (
    n380,
    n233,
    n25,
    n145,
    n224
  );


  nor
  g375
  (
    n334,
    n136,
    n246,
    n252,
    n206
  );


  and
  g376
  (
    n367,
    n104,
    n154,
    n253,
    n147
  );


  nand
  g377
  (
    n406,
    n218,
    n173,
    n23,
    n180
  );


  or
  g378
  (
    n424,
    n245,
    n206,
    n25,
    n116
  );


  nor
  g379
  (
    n312,
    n223,
    n261,
    n229,
    n145
  );


  nor
  g380
  (
    n341,
    n131,
    n189,
    n248,
    n112
  );


  xor
  g381
  (
    KeyWire_0_4,
    n220,
    n228,
    n136,
    n175
  );


  nor
  g382
  (
    n384,
    n24,
    n96,
    n8,
    n233
  );


  xnor
  g383
  (
    n446,
    n234,
    n229,
    n195,
    n154
  );


  nor
  g384
  (
    n274,
    n204,
    n186,
    n209,
    n169
  );


  nand
  g385
  (
    n489,
    n187,
    n196,
    n186,
    n116
  );


  xnor
  g386
  (
    n349,
    n7,
    n151,
    n192,
    n114
  );


  and
  g387
  (
    n477,
    n130,
    n212,
    n19,
    n113
  );


  xnor
  g388
  (
    n376,
    n237,
    n172,
    n226,
    n164
  );


  xnor
  g389
  (
    n350,
    n142,
    n179,
    n7,
    n133
  );


  and
  g390
  (
    n370,
    n138,
    n267,
    n106,
    n133
  );


  xnor
  g391
  (
    n458,
    n159,
    n222,
    n265,
    n204
  );


  nand
  g392
  (
    n357,
    n200,
    n247,
    n199,
    n12
  );


  and
  g393
  (
    n504,
    n13,
    n245,
    n137,
    n102
  );


  or
  g394
  (
    n281,
    n13,
    n157,
    n110,
    n117
  );


  and
  g395
  (
    n345,
    n198,
    n100,
    n248,
    n21
  );


  nor
  g396
  (
    n310,
    n134,
    n191,
    n159,
    n221
  );


  nand
  g397
  (
    n469,
    n138,
    n187,
    n249,
    n131
  );


  xor
  g398
  (
    n343,
    n160,
    n225,
    n212,
    n132
  );


  xnor
  g399
  (
    n426,
    n190,
    n134,
    n197,
    n93
  );


  and
  g400
  (
    n493,
    n269,
    n13,
    n106,
    n8
  );


  nor
  g401
  (
    n438,
    n222,
    n140,
    n258,
    n203
  );


  or
  g402
  (
    n338,
    n24,
    n182,
    n121,
    n201
  );


  nand
  g403
  (
    n428,
    n186,
    n184,
    n120,
    n107
  );


  or
  g404
  (
    n417,
    n157,
    n151,
    n161,
    n185
  );


  xnor
  g405
  (
    n502,
    n258,
    n153,
    n6,
    n251
  );


  or
  g406
  (
    n398,
    n12,
    n129,
    n157,
    n202
  );


  xnor
  g407
  (
    n307,
    n249,
    n221,
    n237,
    n150
  );


  nor
  g408
  (
    n491,
    n161,
    n24,
    n235,
    n129
  );


  xor
  g409
  (
    n483,
    n218,
    n255,
    n8,
    n117
  );


  nand
  g410
  (
    n286,
    n17,
    n24,
    n99,
    n257
  );


  xor
  g411
  (
    n330,
    n206,
    n210,
    n180,
    n183
  );


  nand
  g412
  (
    n315,
    n206,
    n233,
    n121,
    n243
  );


  xor
  g413
  (
    n272,
    n165,
    n101,
    n112,
    n102
  );


  xnor
  g414
  (
    n422,
    n130,
    n267,
    n140,
    n216
  );


  xnor
  g415
  (
    n280,
    n6,
    n104,
    n160,
    n237
  );


  and
  g416
  (
    n347,
    n96,
    n19,
    n179,
    n139
  );


  xnor
  g417
  (
    n420,
    n103,
    n247,
    n148,
    n240
  );


  nand
  g418
  (
    n388,
    n261,
    n197,
    n123,
    n236
  );


  xnor
  g419
  (
    n303,
    n148,
    n14,
    n212,
    n256
  );


  xnor
  g420
  (
    n481,
    n168,
    n200,
    n183,
    n169
  );


  nand
  g421
  (
    n298,
    n177,
    n120,
    n232,
    n182
  );


  nand
  g422
  (
    n374,
    n205,
    n175,
    n139,
    n230
  );


  xnor
  g423
  (
    n498,
    n188,
    n94,
    n262,
    n20
  );


  or
  g424
  (
    n337,
    n96,
    n264,
    n160,
    n152
  );


  xor
  g425
  (
    n301,
    n260,
    n22,
    n159,
    n107
  );


  xor
  g426
  (
    KeyWire_0_3,
    n208,
    n246,
    n223,
    n216
  );


  nor
  g427
  (
    n413,
    n184,
    n233,
    n26,
    n18
  );


  xnor
  g428
  (
    n454,
    n121,
    n219,
    n115,
    n162
  );


  and
  g429
  (
    n431,
    n201,
    n114,
    n236,
    n149
  );


  or
  g430
  (
    n299,
    n207,
    n126,
    n220,
    n199
  );


  nand
  g431
  (
    n363,
    n145,
    n178,
    n259,
    n132
  );


  xnor
  g432
  (
    n360,
    n173,
    n177,
    n141,
    n15
  );


  xnor
  g433
  (
    n470,
    n190,
    n167,
    n135,
    n212
  );


  and
  g434
  (
    n289,
    n180,
    n231,
    n260,
    n228
  );


  and
  g435
  (
    n351,
    n97,
    n238,
    n246,
    n261
  );


  xor
  g436
  (
    n460,
    n229,
    n14,
    n115,
    n94
  );


  or
  g437
  (
    n409,
    n197,
    n193,
    n128,
    n239
  );


  nor
  g438
  (
    n509,
    n188,
    n142,
    n192,
    n18
  );


  nor
  g439
  (
    n425,
    n203,
    n192,
    n98,
    n240
  );


  nand
  g440
  (
    n316,
    n8,
    n17,
    n191,
    n244
  );


  xnor
  g441
  (
    n385,
    n225,
    n122,
    n125,
    n193
  );


  and
  g442
  (
    n390,
    n243,
    n146,
    n228
  );


  xnor
  g443
  (
    n392,
    n108,
    n254,
    n213,
    n234
  );


  or
  g444
  (
    n378,
    n256,
    n97,
    n222,
    n133
  );


  and
  g445
  (
    n323,
    n129,
    n224,
    n187,
    n166
  );


  nand
  g446
  (
    n361,
    n162,
    n25,
    n113,
    n151
  );


  xor
  g447
  (
    n444,
    n198,
    n176,
    n132,
    n255
  );


  nand
  g448
  (
    n412,
    n123,
    n194,
    n100,
    n227
  );


  xnor
  g449
  (
    n423,
    n196,
    n159,
    n168,
    n134
  );


  nand
  g450
  (
    n455,
    n238,
    n250,
    n101,
    n98
  );


  xor
  g451
  (
    n473,
    n231,
    n185,
    n93,
    n224
  );


  xor
  g452
  (
    n336,
    n254,
    n105,
    n153,
    n119
  );


  or
  g453
  (
    n393,
    n163,
    n182,
    n174,
    n93
  );


  xor
  g454
  (
    n421,
    n131,
    n263,
    n15,
    n241
  );


  xor
  g455
  (
    n284,
    n117,
    n144,
    n128
  );


  nor
  g456
  (
    n403,
    n152,
    n128,
    n250,
    n108
  );


  or
  g457
  (
    n325,
    n21,
    n170,
    n227,
    n119
  );


  xor
  g458
  (
    n479,
    n201,
    n219,
    n170,
    n95
  );


  xor
  g459
  (
    n442,
    n259,
    n200,
    n163,
    n7
  );


  or
  g460
  (
    n355,
    n98,
    n199,
    n238,
    n197
  );


  nor
  g461
  (
    n283,
    n217,
    n268,
    n143,
    n104
  );


  nand
  g462
  (
    n366,
    n168,
    n165,
    n95,
    n11
  );


  and
  g463
  (
    n490,
    n155,
    n20,
    n108,
    n171
  );


  xor
  g464
  (
    n467,
    n207,
    n166,
    n150,
    n215
  );


  and
  g465
  (
    n273,
    n194,
    n250,
    n228,
    n244
  );


  and
  g466
  (
    n434,
    n128,
    n194,
    n122,
    n10
  );


  or
  g467
  (
    n466,
    n216,
    n188,
    n145,
    n175
  );


  nand
  g468
  (
    n368,
    n138,
    n137,
    n112,
    n186
  );


  xnor
  g469
  (
    n293,
    n103,
    n266,
    n239,
    n164
  );


  nor
  g470
  (
    n371,
    n239,
    n193,
    n126,
    n152
  );


  and
  g471
  (
    n306,
    n215,
    n263,
    n209,
    n156
  );


  xor
  g472
  (
    n389,
    n227,
    n138,
    n191,
    n171
  );


  xor
  g473
  (
    n319,
    n257,
    n158,
    n154,
    n10
  );


  nand
  g474
  (
    n395,
    n118,
    n122,
    n93,
    n167
  );


  or
  g475
  (
    n447,
    n202,
    n269,
    n101,
    n140
  );


  xor
  g476
  (
    n475,
    n189,
    n116,
    n6,
    n232
  );


  xor
  g477
  (
    n326,
    n121,
    n26,
    n9,
    n109
  );


  xor
  g478
  (
    n531,
    n300,
    n309,
    n282
  );


  or
  g479
  (
    n522,
    n315,
    n307,
    n301,
    n293
  );


  nand
  g480
  (
    n533,
    n281,
    n284,
    n295,
    n291
  );


  xnor
  g481
  (
    n530,
    n305,
    n312,
    n282,
    n278
  );


  nor
  g482
  (
    n521,
    n283,
    n311,
    n290,
    n280
  );


  or
  g483
  (
    n551,
    n278,
    n292,
    n315,
    n306
  );


  or
  g484
  (
    n525,
    n293,
    n306,
    n280,
    n287
  );


  or
  g485
  (
    n539,
    n279,
    n278,
    n283,
    n310
  );


  or
  g486
  (
    n549,
    n298,
    n275,
    n281,
    n312
  );


  nor
  g487
  (
    n512,
    n313,
    n304,
    n311,
    n293
  );


  xor
  g488
  (
    n537,
    n303,
    n276,
    n302,
    n286
  );


  xor
  g489
  (
    n527,
    n312,
    n297,
    n291,
    n280
  );


  nor
  g490
  (
    KeyWire_0_19,
    n290,
    n300,
    n287,
    n280
  );


  and
  g491
  (
    n546,
    n314,
    n290,
    n288,
    n305
  );


  and
  g492
  (
    n524,
    n277,
    n274,
    n315,
    n289
  );


  or
  g493
  (
    n538,
    n294,
    n294,
    n300,
    n285
  );


  nand
  g494
  (
    n552,
    n301,
    n274,
    n311,
    n296
  );


  nand
  g495
  (
    n513,
    n288,
    n308,
    n275
  );


  and
  g496
  (
    n514,
    n314,
    n296,
    n299,
    n291
  );


  xnor
  g497
  (
    n554,
    n310,
    n304,
    n273,
    n286
  );


  and
  g498
  (
    n550,
    n274,
    n287,
    n286,
    n307
  );


  xor
  g499
  (
    n547,
    n308,
    n309,
    n298,
    n299
  );


  xnor
  g500
  (
    n528,
    n289,
    n277,
    n284,
    n285
  );


  xnor
  g501
  (
    n541,
    n283,
    n313,
    n307,
    n279
  );


  nor
  g502
  (
    n542,
    n313,
    n275,
    n304,
    n272
  );


  nand
  g503
  (
    n544,
    n291,
    n282,
    n308,
    n299
  );


  or
  g504
  (
    n532,
    n295,
    n277,
    n300,
    n292
  );


  nand
  g505
  (
    n523,
    n301,
    n296,
    n312,
    n294
  );


  or
  g506
  (
    n520,
    n310,
    n305,
    n298,
    n285
  );


  and
  g507
  (
    n518,
    n311,
    n289,
    n273,
    n310
  );


  nor
  g508
  (
    n540,
    n284,
    n298,
    n292,
    n297
  );


  or
  g509
  (
    n543,
    n283,
    n305,
    n303,
    n297
  );


  xnor
  g510
  (
    n519,
    n287,
    n292,
    n279,
    n304
  );


  nand
  g511
  (
    n545,
    n314,
    n306,
    n273,
    n274
  );


  and
  g512
  (
    n517,
    n284,
    n313,
    n293,
    n289
  );


  and
  g513
  (
    n536,
    n276,
    n281,
    n302,
    n273
  );


  and
  g514
  (
    n515,
    n302,
    n282,
    n297,
    n272
  );


  or
  g515
  (
    n553,
    n272,
    n288,
    n281,
    n295
  );


  nor
  g516
  (
    n516,
    n294,
    n272,
    n302,
    n303
  );


  or
  g517
  (
    n548,
    n290,
    n308,
    n296,
    n276
  );


  or
  g518
  (
    n529,
    n299,
    n303,
    n277,
    n314
  );


  xnor
  g519
  (
    n511,
    n309,
    n286,
    n288,
    n285
  );


  and
  g520
  (
    n534,
    n278,
    n309,
    n307,
    n306
  );


  xor
  g521
  (
    n535,
    n295,
    n301,
    n276,
    n279
  );


  and
  g522
  (
    n589,
    n394,
    n521,
    n382,
    n518
  );


  nor
  g523
  (
    n655,
    n317,
    n526,
    n391,
    n384
  );


  xnor
  g524
  (
    n608,
    n524,
    n355,
    n330,
    n358
  );


  nor
  g525
  (
    n625,
    n374,
    n390,
    n359,
    n539
  );


  xnor
  g526
  (
    n563,
    n395,
    n333,
    n349,
    n354
  );


  nand
  g527
  (
    n664,
    n398,
    n537,
    n393,
    n364
  );


  or
  g528
  (
    n577,
    n524,
    n319,
    n359,
    n364
  );


  xor
  g529
  (
    n627,
    n354,
    n342,
    n319
  );


  and
  g530
  (
    n660,
    n318,
    n530,
    n322,
    n386
  );


  nand
  g531
  (
    n644,
    n383,
    n384,
    n348,
    n529
  );


  nor
  g532
  (
    n636,
    n340,
    n316,
    n370,
    n390
  );


  nor
  g533
  (
    n630,
    n374,
    n353,
    n398,
    n390
  );


  xnor
  g534
  (
    n657,
    n341,
    n380,
    n367,
    n368
  );


  nor
  g535
  (
    n624,
    n363,
    n347,
    n373,
    n376
  );


  nor
  g536
  (
    n574,
    n320,
    n334,
    n318,
    n359
  );


  or
  g537
  (
    n623,
    n326,
    n347,
    n333,
    n368
  );


  xnor
  g538
  (
    n641,
    n514,
    n349,
    n365,
    n322
  );


  and
  g539
  (
    n610,
    n386,
    n532,
    n520,
    n357
  );


  or
  g540
  (
    n666,
    n387,
    n329,
    n396,
    n534
  );


  nand
  g541
  (
    KeyWire_0_9,
    n528,
    n536,
    n512,
    n385
  );


  or
  g542
  (
    n569,
    n317,
    n353,
    n380,
    n381
  );


  nor
  g543
  (
    n628,
    n519,
    n380,
    n320,
    n512
  );


  or
  g544
  (
    n611,
    n335,
    n373,
    n371,
    n535
  );


  xor
  g545
  (
    n586,
    n518,
    n385,
    n323,
    n529
  );


  nand
  g546
  (
    n648,
    n336,
    n536,
    n349,
    n522
  );


  xor
  g547
  (
    n562,
    n387,
    n391,
    n323,
    n397
  );


  nand
  g548
  (
    n639,
    n379,
    n389,
    n339,
    n374
  );


  xnor
  g549
  (
    n622,
    n533,
    n386,
    n538,
    n513
  );


  nand
  g550
  (
    n556,
    n345,
    n324,
    n377
  );


  or
  g551
  (
    n612,
    n365,
    n521,
    n394,
    n373
  );


  xor
  g552
  (
    n651,
    n513,
    n344,
    n346,
    n352
  );


  nor
  g553
  (
    n659,
    n331,
    n331,
    n364,
    n332
  );


  xnor
  g554
  (
    n580,
    n354,
    n324,
    n394,
    n517
  );


  xor
  g555
  (
    n652,
    n330,
    n392,
    n367,
    n535
  );


  and
  g556
  (
    n558,
    n351,
    n518,
    n358,
    n356
  );


  and
  g557
  (
    n619,
    n383,
    n515,
    n372,
    n392
  );


  or
  g558
  (
    n578,
    n317,
    n537,
    n351,
    n527
  );


  nand
  g559
  (
    n640,
    n327,
    n339,
    n366,
    n337
  );


  and
  g560
  (
    n598,
    n322,
    n332,
    n363,
    n520
  );


  and
  g561
  (
    n599,
    n376,
    n514,
    n388,
    n378
  );


  and
  g562
  (
    n601,
    n321,
    n522,
    n334,
    n532
  );


  xnor
  g563
  (
    n616,
    n515,
    n538,
    n388,
    n343
  );


  xnor
  g564
  (
    n603,
    n529,
    n348,
    n391,
    n346
  );


  xnor
  g565
  (
    n587,
    n321,
    n399,
    n527,
    n355
  );


  xnor
  g566
  (
    n646,
    n393,
    n517,
    n327,
    n516
  );


  xor
  g567
  (
    n594,
    n316,
    n333,
    n517,
    n382
  );


  xnor
  g568
  (
    n663,
    n361,
    n352,
    n357,
    n350
  );


  xor
  g569
  (
    n658,
    n331,
    n357,
    n375,
    n345
  );


  and
  g570
  (
    n576,
    n513,
    n382,
    n354,
    n328
  );


  nand
  g571
  (
    n596,
    n325,
    n525,
    n398,
    n329
  );


  nand
  g572
  (
    n635,
    n523,
    n373,
    n341,
    n352
  );


  nor
  g573
  (
    n575,
    n351,
    n387,
    n530,
    n342
  );


  nand
  g574
  (
    n632,
    n335,
    n539,
    n318,
    n532
  );


  nor
  g575
  (
    n633,
    n357,
    n379,
    n332,
    n366
  );


  nor
  g576
  (
    n606,
    n385,
    n384,
    n531,
    n530
  );


  xnor
  g577
  (
    n662,
    n319,
    n533,
    n346,
    n337
  );


  or
  g578
  (
    n665,
    n353,
    n525,
    n372,
    n514
  );


  nand
  g579
  (
    n602,
    n380,
    n398,
    n348,
    n349
  );


  xor
  g580
  (
    n572,
    n338,
    n339,
    n530,
    n337
  );


  or
  g581
  (
    n593,
    n343,
    n395,
    n332,
    n340
  );


  xor
  g582
  (
    n650,
    n396,
    n326,
    n369,
    n523
  );


  xor
  g583
  (
    n637,
    n512,
    n329,
    n374,
    n370
  );


  and
  g584
  (
    n621,
    n386,
    n327,
    n383,
    n528
  );


  nand
  g585
  (
    n604,
    n329,
    n519,
    n534,
    n514
  );


  xor
  g586
  (
    n579,
    n360,
    n325,
    n519,
    n322
  );


  xnor
  g587
  (
    n561,
    n396,
    n534,
    n323,
    n393
  );


  or
  g588
  (
    n661,
    n388,
    n319,
    n317,
    n359
  );


  xor
  g589
  (
    n600,
    n326,
    n353,
    n336,
    n360
  );


  and
  g590
  (
    n617,
    n360,
    n526,
    n397,
    n350
  );


  nor
  g591
  (
    n656,
    n516,
    n531,
    n347,
    n536
  );


  or
  g592
  (
    n573,
    n335,
    n399,
    n361,
    n538
  );


  nor
  g593
  (
    n560,
    n372,
    n383,
    n345,
    n362
  );


  xor
  g594
  (
    n638,
    n529,
    n367,
    n324,
    n369
  );


  xor
  g595
  (
    n581,
    n523,
    n344,
    n392,
    n331
  );


  nand
  g596
  (
    n645,
    n370,
    n368,
    n318,
    n365
  );


  nor
  g597
  (
    n597,
    n528,
    n377,
    n356,
    n376
  );


  or
  g598
  (
    n642,
    n511,
    n390,
    n355
  );


  nor
  g599
  (
    n605,
    n327,
    n361,
    n342,
    n525
  );


  and
  g600
  (
    n559,
    n521,
    n356,
    n351,
    n335
  );


  nor
  g601
  (
    n582,
    n372,
    n341,
    n536,
    n334
  );


  nor
  g602
  (
    n607,
    n340,
    n316,
    n320,
    n511
  );


  nor
  g603
  (
    n584,
    n375,
    n369,
    n330,
    n325
  );


  and
  g604
  (
    n634,
    n364,
    n517,
    n328,
    n382
  );


  nand
  g605
  (
    n571,
    n388,
    n371,
    n350,
    n352
  );


  or
  g606
  (
    n555,
    n328,
    n520,
    n527,
    n397
  );


  xor
  g607
  (
    n654,
    n397,
    n344,
    n391,
    n358
  );


  xor
  g608
  (
    n620,
    n315,
    n358,
    n338,
    n381
  );


  nand
  g609
  (
    n557,
    n533,
    n343,
    n392,
    n340
  );


  nor
  g610
  (
    n629,
    n393,
    n535,
    n323,
    n343
  );


  nand
  g611
  (
    n570,
    n522,
    n375,
    n316,
    n516
  );


  xor
  g612
  (
    n585,
    n338,
    n345,
    n389
  );


  xor
  g613
  (
    n592,
    n378,
    n521,
    n330,
    n368
  );


  or
  g614
  (
    n583,
    n367,
    n523,
    n365,
    n363
  );


  nand
  g615
  (
    n591,
    n378,
    n337,
    n321,
    n538
  );


  nor
  g616
  (
    n566,
    n384,
    n396,
    n375,
    n518
  );


  or
  g617
  (
    n614,
    n362,
    n515,
    n341,
    n370
  );


  nand
  g618
  (
    n631,
    n362,
    n381,
    n526,
    n369
  );


  or
  g619
  (
    n626,
    n519,
    n339,
    n366,
    n532
  );


  and
  g620
  (
    n567,
    n320,
    n344,
    n378,
    n527
  );


  or
  g621
  (
    n647,
    n371,
    n513,
    n511,
    n389
  );


  and
  g622
  (
    n618,
    n360,
    n524,
    n334,
    n537
  );


  xnor
  g623
  (
    n565,
    n377,
    n524,
    n531,
    n533
  );


  and
  g624
  (
    n609,
    n528,
    n350,
    n395,
    n535
  );


  xor
  g625
  (
    n595,
    n381,
    n526,
    n362,
    n385
  );


  xor
  g626
  (
    n568,
    n394,
    n363,
    n346,
    n377
  );


  xnor
  g627
  (
    n588,
    n347,
    n516,
    n537,
    n515
  );


  and
  g628
  (
    n615,
    n348,
    n522,
    n520,
    n325
  );


  and
  g629
  (
    n564,
    n379,
    n376,
    n326,
    n534
  );


  and
  g630
  (
    n649,
    n336,
    n395,
    n525,
    n333
  );


  nand
  g631
  (
    n613,
    n371,
    n328,
    n361,
    n336
  );


  nand
  g632
  (
    n590,
    n379,
    n321,
    n366,
    n531
  );


  xor
  g633
  (
    n643,
    n338,
    n512,
    n387,
    n356
  );


  nand
  g634
  (
    KeyWire_0_1,
    n569,
    n570,
    n578,
    n576
  );


  nor
  g635
  (
    n689,
    n576,
    n561
  );


  nand
  g636
  (
    n678,
    n581,
    n578,
    n555,
    n557
  );


  nand
  g637
  (
    n692,
    n557,
    n571,
    n576,
    n580
  );


  nor
  g638
  (
    n686,
    n563,
    n555,
    n559,
    n573
  );


  nand
  g639
  (
    n676,
    n565,
    n563,
    n575,
    n580
  );


  and
  g640
  (
    n677,
    n560,
    n557,
    n564,
    n567
  );


  or
  g641
  (
    n681,
    n566,
    n559,
    n569,
    n580
  );


  xor
  g642
  (
    n690,
    n580,
    n579,
    n566,
    n562
  );


  nand
  g643
  (
    n684,
    n564,
    n572,
    n566,
    n568
  );


  nor
  g644
  (
    n693,
    n570,
    n559,
    n567,
    n581
  );


  nand
  g645
  (
    n683,
    n562,
    n570,
    n557,
    n578
  );


  nand
  g646
  (
    n670,
    n563,
    n579,
    n556
  );


  nand
  g647
  (
    n673,
    n555,
    n574,
    n556,
    n575
  );


  xor
  g648
  (
    n680,
    n570,
    n569,
    n558,
    n565
  );


  xor
  g649
  (
    n682,
    n566,
    n564,
    n577,
    n575
  );


  xnor
  g650
  (
    n668,
    n571,
    n556,
    n567,
    n573
  );


  and
  g651
  (
    n675,
    n572,
    n568,
    n561,
    n560
  );


  xor
  g652
  (
    n672,
    n565,
    n571,
    n558,
    n572
  );


  nand
  g653
  (
    n679,
    n573,
    n577,
    n563,
    n568
  );


  nor
  g654
  (
    n685,
    n560,
    n558,
    n574
  );


  xor
  g655
  (
    n687,
    n581,
    n556,
    n562,
    n574
  );


  or
  g656
  (
    n667,
    n578,
    n559,
    n560,
    n555
  );


  nor
  g657
  (
    n674,
    n576,
    n562,
    n571,
    n574
  );


  xnor
  g658
  (
    n671,
    n569,
    n568,
    n567,
    n564
  );


  xor
  g659
  (
    n688,
    n565,
    n572,
    n577,
    n579
  );


  nor
  g660
  (
    n691,
    n581,
    n575,
    n577,
    n573
  );


  not
  g661
  (
    n704,
    n674
  );


  xnor
  g662
  (
    n719,
    n602,
    n671,
    n668
  );


  nand
  g663
  (
    n706,
    n582,
    n598,
    n592,
    n668
  );


  and
  g664
  (
    n711,
    n597,
    n593,
    n598
  );


  nand
  g665
  (
    n724,
    n588,
    n589,
    n584,
    n593
  );


  or
  g666
  (
    n716,
    n596,
    n667,
    n598,
    n602
  );


  nor
  g667
  (
    n712,
    n595,
    n593,
    n602,
    n584
  );


  or
  g668
  (
    n708,
    n601,
    n671,
    n584,
    n591
  );


  nor
  g669
  (
    n714,
    n598,
    n600,
    n601,
    n673
  );


  or
  g670
  (
    n696,
    n667,
    n582,
    n672
  );


  or
  g671
  (
    n703,
    n599,
    n592,
    n589,
    n600
  );


  xor
  g672
  (
    n695,
    n669,
    n670,
    n592,
    n600
  );


  xor
  g673
  (
    n722,
    n597,
    n672,
    n670,
    n587
  );


  xnor
  g674
  (
    n700,
    n595,
    n603,
    n586,
    n670
  );


  and
  g675
  (
    n701,
    n674,
    n586,
    n667,
    n599
  );


  and
  g676
  (
    n717,
    n592,
    n600,
    n583,
    n587
  );


  xor
  g677
  (
    n698,
    n603,
    n599,
    n601,
    n582
  );


  xor
  g678
  (
    n702,
    n583,
    n596,
    n588,
    n591
  );


  nor
  g679
  (
    n707,
    n601,
    n594,
    n599,
    n673
  );


  or
  g680
  (
    n709,
    n590,
    n589,
    n603,
    n587
  );


  or
  g681
  (
    n699,
    n595,
    n585,
    n584
  );


  nand
  g682
  (
    n697,
    n669,
    n604,
    n591,
    n588
  );


  or
  g683
  (
    n713,
    n670,
    n596,
    n586,
    n590
  );


  xor
  g684
  (
    n718,
    n603,
    n597,
    n590
  );


  xnor
  g685
  (
    n705,
    n590,
    n673,
    n596,
    n602
  );


  and
  g686
  (
    n723,
    n668,
    n668,
    n669,
    n591
  );


  and
  g687
  (
    n710,
    n672,
    n671,
    n586,
    n583
  );


  nand
  g688
  (
    n720,
    n583,
    n594,
    n673,
    n667
  );


  xnor
  g689
  (
    n715,
    n594,
    n587,
    n595,
    n588
  );


  xnor
  g690
  (
    n721,
    n674,
    n585,
    n594,
    n671
  );


  and
  g691
  (
    n694,
    n669,
    n585,
    n672,
    n589
  );


  nand
  g692
  (
    n725,
    n695,
    n676,
    n675
  );


  nor
  g693
  (
    n727,
    n27,
    n674,
    n678
  );


  or
  g694
  (
    n730,
    n676,
    n694,
    n678,
    n675
  );


  xor
  g695
  (
    n728,
    n27,
    n694,
    n677
  );


  nor
  g696
  (
    n729,
    n696,
    n696,
    n695,
    n694
  );


  nor
  g697
  (
    n726,
    n676,
    n695,
    n677
  );


  and
  g698
  (
    n731,
    n27,
    n675,
    n678
  );


  xor
  g699
  (
    n732,
    n679,
    n677
  );


  xor
  g700
  (
    n751,
    n620,
    n620,
    n616,
    n614
  );


  and
  g701
  (
    n745,
    n725,
    n609,
    n605,
    n619
  );


  xnor
  g702
  (
    n755,
    n609,
    n610,
    n617,
    n731
  );


  xnor
  g703
  (
    n758,
    n618,
    n732,
    n613,
    n726
  );


  or
  g704
  (
    n742,
    n607,
    n605,
    n728,
    n45
  );


  nand
  g705
  (
    n757,
    n613,
    n619,
    n45,
    n614
  );


  nand
  g706
  (
    n741,
    n620,
    n618,
    n696
  );


  xor
  g707
  (
    n736,
    n611,
    n607,
    n618,
    n610
  );


  or
  g708
  (
    n739,
    n612,
    n727,
    n614,
    n731
  );


  nand
  g709
  (
    n734,
    n726,
    n611,
    n697,
    n607
  );


  nor
  g710
  (
    n743,
    n608,
    n697,
    n613,
    n725
  );


  xnor
  g711
  (
    n750,
    n729,
    n610,
    n606,
    n730
  );


  or
  g712
  (
    n738,
    n613,
    n697,
    n619,
    n609
  );


  xnor
  g713
  (
    n752,
    n618,
    n45,
    n610,
    n617
  );


  xnor
  g714
  (
    n746,
    n615,
    n612,
    n605,
    n727
  );


  and
  g715
  (
    n744,
    n730,
    n606,
    n609,
    n614
  );


  nand
  g716
  (
    n756,
    n615,
    n732,
    n617,
    n612
  );


  or
  g717
  (
    n754,
    n605,
    n729,
    n732
  );


  nor
  g718
  (
    n748,
    n616,
    n725,
    n615,
    n620
  );


  and
  g719
  (
    n740,
    n46,
    n45,
    n611,
    n726
  );


  nand
  g720
  (
    n749,
    n728,
    n727,
    n616,
    n607
  );


  and
  g721
  (
    n733,
    n697,
    n606,
    n612,
    n604
  );


  nand
  g722
  (
    n753,
    n731,
    n604,
    n608,
    n606
  );


  or
  g723
  (
    n747,
    n729,
    n616,
    n608,
    n619
  );


  nor
  g724
  (
    n737,
    n611,
    n604,
    n730,
    n617
  );


  xor
  g725
  (
    n735,
    n615,
    n608,
    n731,
    n728
  );


  xor
  g726
  (
    n763,
    n623,
    n621,
    n733,
    n734
  );


  nand
  g727
  (
    n764,
    n624,
    n622
  );


  or
  g728
  (
    n759,
    n621,
    n624,
    n625,
    n622
  );


  nand
  g729
  (
    n761,
    n621,
    n733,
    n623
  );


  or
  g730
  (
    n762,
    n624,
    n734,
    n621
  );


  xor
  g731
  (
    n760,
    n625,
    n623,
    n622
  );


  nand
  g732
  (
    n770,
    n628,
    n401
  );


  xnor
  g733
  (
    n765,
    n761,
    n629,
    n400,
    n626
  );


  xor
  g734
  (
    n773,
    n400,
    n759,
    n628,
    n762
  );


  and
  g735
  (
    n771,
    n762,
    n762,
    n628,
    n627
  );


  xor
  g736
  (
    n774,
    n399,
    n626,
    n625,
    n628
  );


  xnor
  g737
  (
    n769,
    n626,
    n401,
    n400
  );


  xnor
  g738
  (
    n768,
    n625,
    n760,
    n679,
    n399
  );


  or
  g739
  (
    n772,
    n679,
    n627,
    n761,
    n763
  );


  xnor
  g740
  (
    n767,
    n680,
    n760,
    n761,
    n627
  );


  xor
  g741
  (
    n766,
    n759,
    n626,
    n627,
    n629
  );


  not
  g742
  (
    n775,
    n629
  );


  not
  g743
  (
    n777,
    n630
  );


  nand
  g744
  (
    n776,
    n770,
    n768
  );


  and
  g745
  (
    n778,
    n629,
    n767,
    n769,
    n401
  );


  nand
  g746
  (
    n784,
    n632,
    n632,
    n633,
    n637
  );


  nor
  g747
  (
    n779,
    n634,
    n638,
    n636
  );


  and
  g748
  (
    n787,
    n634,
    n776,
    n635,
    n631
  );


  or
  g749
  (
    n788,
    n775,
    n776,
    n632
  );


  nor
  g750
  (
    n790,
    n630,
    n637,
    n631
  );


  xor
  g751
  (
    n785,
    n777,
    n778,
    n631,
    n630
  );


  or
  g752
  (
    n783,
    n635,
    n777,
    n633,
    n637
  );


  xnor
  g753
  (
    n780,
    n633,
    n634,
    n639
  );


  xor
  g754
  (
    n782,
    n777,
    n635,
    n630,
    n636
  );


  or
  g755
  (
    n786,
    n632,
    n638,
    n775
  );


  xnor
  g756
  (
    n781,
    n776,
    n633,
    n637,
    n635
  );


  and
  g757
  (
    n789,
    n777,
    n636,
    n638
  );


  xnor
  g758
  (
    n792,
    n681,
    n680
  );


  or
  g759
  (
    n791,
    n680,
    n779,
    n681
  );


  and
  g760
  (
    n794,
    n682,
    n29
  );


  xnor
  g761
  (
    n795,
    n29,
    n28
  );


  or
  g762
  (
    KeyWire_0_17,
    n792,
    n28,
    n791
  );


  or
  g763
  (
    n793,
    n791,
    n681,
    n29,
    n28
  );


  xor
  g764
  (
    n797,
    n698,
    n699
  );


  nor
  g765
  (
    n801,
    n792,
    n698,
    n639,
    n699
  );


  or
  g766
  (
    n800,
    n698,
    n794,
    n793,
    n699
  );


  or
  g767
  (
    n799,
    n794,
    n639,
    n792,
    n699
  );


  nor
  g768
  (
    n798,
    n792,
    n698,
    n793
  );


  xnor
  g769
  (
    n806,
    n764,
    n763,
    n407,
    n801
  );


  nand
  g770
  (
    n815,
    n404,
    n404,
    n403,
    n778
  );


  or
  g771
  (
    n809,
    n797,
    n800,
    n408,
    n781
  );


  nand
  g772
  (
    n807,
    n798,
    n779,
    n405,
    n407
  );


  xnor
  g773
  (
    n812,
    n404,
    n779,
    n92,
    n778
  );


  or
  g774
  (
    n810,
    n682,
    n403,
    n640,
    n405
  );


  and
  g775
  (
    n804,
    n402,
    n780,
    n403,
    n407
  );


  nor
  g776
  (
    n814,
    n799,
    n801,
    n406,
    n800
  );


  xnor
  g777
  (
    n803,
    n408,
    n797,
    n406,
    n640
  );


  xor
  g778
  (
    n808,
    n406,
    n801,
    n764,
    n408
  );


  or
  g779
  (
    n816,
    n799,
    n402,
    n405,
    n763
  );


  xnor
  g780
  (
    n802,
    n780,
    n408,
    n402,
    n640
  );


  nor
  g781
  (
    n817,
    n402,
    n800,
    n405,
    n407
  );


  nand
  g782
  (
    n805,
    n639,
    n406,
    n798,
    n797
  );


  and
  g783
  (
    n813,
    n799,
    n780,
    n403,
    n640
  );


  or
  g784
  (
    n811,
    n780,
    n404,
    n800,
    n798
  );


  and
  g785
  (
    n825,
    n805,
    n784,
    n788
  );


  nor
  g786
  (
    n820,
    n788,
    n805,
    n785,
    n787
  );


  xor
  g787
  (
    n832,
    n803,
    n790,
    n642,
    n789
  );


  nor
  g788
  (
    n823,
    n789,
    n804,
    n784,
    n802
  );


  nor
  g789
  (
    n819,
    n783,
    n786,
    n642,
    n788
  );


  xor
  g790
  (
    n828,
    n782,
    n785,
    n641,
    n788
  );


  nand
  g791
  (
    n821,
    n782,
    n802,
    n641,
    n784
  );


  or
  g792
  (
    n827,
    n787,
    n802,
    n804,
    n642
  );


  or
  g793
  (
    n831,
    n803,
    n802,
    n804,
    n782
  );


  or
  g794
  (
    n818,
    n783,
    n783,
    n804,
    n803
  );


  xnor
  g795
  (
    n824,
    n787,
    n805,
    n789,
    n782
  );


  nor
  g796
  (
    n829,
    n643,
    n783,
    n786,
    n781
  );


  xor
  g797
  (
    n830,
    n781,
    n803,
    n786,
    n785
  );


  or
  g798
  (
    n822,
    n787,
    n642,
    n641
  );


  or
  g799
  (
    n826,
    n789,
    n786,
    n785,
    n781
  );


  buf
  g800
  (
    n833,
    n825
  );


  buf
  g801
  (
    n834,
    n826
  );


  nor
  g802
  (
    n837,
    n30,
    n834,
    n645,
    n644
  );


  nor
  g803
  (
    n838,
    n834,
    n834,
    n645,
    n833
  );


  and
  g804
  (
    n835,
    n645,
    n643,
    n833
  );


  nor
  g805
  (
    n839,
    n790,
    n644,
    n643
  );


  nand
  g806
  (
    n836,
    n645,
    n790,
    n644
  );


  xnor
  g807
  (
    n846,
    n652,
    n836,
    n649,
    n660
  );


  xor
  g808
  (
    n845,
    n648,
    n649,
    n837,
    n654
  );


  xor
  g809
  (
    n853,
    n647,
    n650,
    n659,
    n652
  );


  xor
  g810
  (
    n840,
    n655,
    n653,
    n649,
    n657
  );


  nand
  g811
  (
    n850,
    n839,
    n837,
    n657,
    n653
  );


  nand
  g812
  (
    n844,
    n836,
    n657,
    n654,
    n655
  );


  xnor
  g813
  (
    n854,
    n838,
    n656,
    n659,
    n837
  );


  xor
  g814
  (
    n851,
    n651,
    n649,
    n652,
    n653
  );


  xnor
  g815
  (
    n859,
    n659,
    n655,
    n651,
    n835
  );


  nor
  g816
  (
    n858,
    n656,
    n838,
    n837
  );


  nand
  g817
  (
    n841,
    n835,
    n646,
    n656,
    n654
  );


  nand
  g818
  (
    n855,
    n646,
    n647,
    n836,
    n656
  );


  and
  g819
  (
    n847,
    n650,
    n646,
    n839,
    n658
  );


  xor
  g820
  (
    n842,
    n836,
    n839,
    n660,
    n646
  );


  or
  g821
  (
    n857,
    n651,
    n658,
    n648
  );


  nand
  g822
  (
    n852,
    n647,
    n653,
    n835,
    n651
  );


  xor
  g823
  (
    n848,
    n652,
    n660,
    n839,
    n838
  );


  nor
  g824
  (
    n843,
    n650,
    n655,
    n659,
    n648
  );


  nand
  g825
  (
    n856,
    n647,
    n654,
    n648,
    n658
  );


  nand
  g826
  (
    n849,
    n660,
    n657,
    n835,
    n650
  );


  and
  g827
  (
    n863,
    n684,
    n683,
    n687
  );


  xnor
  g828
  (
    n860,
    n661,
    n841,
    n687,
    n840
  );


  xor
  g829
  (
    n866,
    n682,
    n685,
    n842
  );


  nor
  g830
  (
    n861,
    n688,
    n686,
    n842,
    n661
  );


  nand
  g831
  (
    n864,
    n841,
    n842,
    n688,
    n685
  );


  or
  g832
  (
    n867,
    n843,
    n686,
    n842,
    n683
  );


  or
  g833
  (
    n868,
    n685,
    n686,
    n840,
    n687
  );


  xor
  g834
  (
    n869,
    n840,
    n684,
    n682
  );


  nand
  g835
  (
    n862,
    n683,
    n687,
    n841,
    n684
  );


  nand
  g836
  (
    n865,
    n686,
    n840,
    n661,
    n841
  );


  or
  g837
  (
    n891,
    n717,
    n717,
    n861,
    n712
  );


  or
  g838
  (
    n885,
    n702,
    n708,
    n710,
    n865
  );


  and
  g839
  (
    n897,
    n869,
    n715,
    n714,
    n705
  );


  nand
  g840
  (
    n880,
    n707,
    n31,
    n706,
    n690
  );


  xor
  g841
  (
    n903,
    n719,
    n710,
    n705,
    n715
  );


  xnor
  g842
  (
    n887,
    n865,
    n705,
    n690,
    n718
  );


  xnor
  g843
  (
    n879,
    n866,
    n689,
    n867,
    n702
  );


  nand
  g844
  (
    n878,
    n703,
    n703,
    n710,
    n720
  );


  or
  g845
  (
    n890,
    n867,
    n721,
    n700
  );


  and
  g846
  (
    n909,
    n709,
    n864,
    n661,
    n707
  );


  nor
  g847
  (
    n884,
    n691,
    n701,
    n713,
    n689
  );


  nor
  g848
  (
    n906,
    n688,
    n704,
    n710,
    n707
  );


  or
  g849
  (
    n881,
    n711,
    n712,
    n868,
    n716
  );


  nor
  g850
  (
    n871,
    n702,
    n719,
    n706,
    n711
  );


  nor
  g851
  (
    n876,
    n700,
    n867,
    n30,
    n704
  );


  nor
  g852
  (
    n889,
    n861,
    n717,
    n711,
    n869
  );


  and
  g853
  (
    n892,
    n720,
    n716,
    n701,
    n860
  );


  xor
  g854
  (
    KeyWire_0_26,
    n719,
    n689,
    n716,
    n709
  );


  or
  g855
  (
    n905,
    n715,
    n862,
    n868,
    n720
  );


  xor
  g856
  (
    n907,
    n864,
    n721,
    n30,
    n714
  );


  nor
  g857
  (
    n902,
    n716,
    n31,
    n702,
    n864
  );


  and
  g858
  (
    n874,
    n862,
    n861,
    n689,
    n796
  );


  and
  g859
  (
    n888,
    n843,
    n864,
    n718,
    n713
  );


  or
  g860
  (
    n908,
    n705,
    n794,
    n862,
    n796
  );


  and
  g861
  (
    n896,
    n704,
    n703,
    n700,
    n861
  );


  xnor
  g862
  (
    n898,
    n707,
    n863,
    n865
  );


  nand
  g863
  (
    n873,
    n863,
    n866,
    n712,
    n708
  );


  and
  g864
  (
    n899,
    n708,
    n30,
    n795,
    n706
  );


  xor
  g865
  (
    n900,
    n715,
    n795,
    n796,
    n701
  );


  nor
  g866
  (
    n894,
    n795,
    n721,
    n796,
    n868
  );


  nor
  g867
  (
    n886,
    n706,
    n778,
    n662,
    n714
  );


  and
  g868
  (
    n882,
    n708,
    n869,
    n795,
    n688
  );


  or
  g869
  (
    n893,
    n866,
    n701,
    n719,
    n717
  );


  nor
  g870
  (
    n875,
    n843,
    n794,
    n713,
    n718
  );


  xnor
  g871
  (
    n870,
    n690,
    n860,
    n868
  );


  xnor
  g872
  (
    n895,
    n862,
    n691,
    n712,
    n690
  );


  and
  g873
  (
    n901,
    n714,
    n709,
    n869,
    n860
  );


  and
  g874
  (
    n904,
    n867,
    n863,
    n711,
    n866
  );


  or
  g875
  (
    n883,
    n720,
    n713,
    n718,
    n703
  );


  or
  g876
  (
    n872,
    n709,
    n865,
    n704,
    n700
  );


  xor
  g877
  (
    n1007,
    n905,
    n878,
    n476,
    n497
  );


  and
  g878
  (
    n1020,
    n434,
    n416,
    n411,
    n454
  );


  xnor
  g879
  (
    n920,
    n422,
    n876,
    n502,
    n440
  );


  xor
  g880
  (
    n951,
    n418,
    n850,
    n501,
    n853
  );


  or
  g881
  (
    n979,
    n908,
    n418,
    n852,
    n450
  );


  xnor
  g882
  (
    n1037,
    n900,
    n896,
    n428,
    n853
  );


  nor
  g883
  (
    n960,
    n461,
    n898,
    n479,
    n471
  );


  nand
  g884
  (
    n939,
    n473,
    n895,
    n851,
    n852
  );


  and
  g885
  (
    n962,
    n663,
    n496,
    n463,
    n447
  );


  and
  g886
  (
    n929,
    n909,
    n449,
    n901,
    n444
  );


  nand
  g887
  (
    n961,
    n881,
    n448,
    n442,
    n439
  );


  xor
  g888
  (
    n1005,
    n434,
    n482,
    n500,
    n488
  );


  xor
  g889
  (
    n1029,
    n903,
    n429,
    n508,
    n451
  );


  or
  g890
  (
    n975,
    n472,
    n724,
    n451,
    n894
  );


  nor
  g891
  (
    n1003,
    n440,
    n470,
    n846
  );


  nor
  g892
  (
    n1053,
    n433,
    n494,
    n846,
    n412
  );


  xor
  g893
  (
    n984,
    n877,
    n462,
    n891,
    n410
  );


  and
  g894
  (
    n996,
    n416,
    n452,
    n492,
    n887
  );


  nor
  g895
  (
    n1054,
    n421,
    n457,
    n884,
    n444
  );


  xor
  g896
  (
    n972,
    n465,
    n882,
    n467,
    n450
  );


  xnor
  g897
  (
    n968,
    n485,
    n723,
    n509,
    n491
  );


  or
  g898
  (
    n1002,
    n448,
    n871,
    n478,
    n510
  );


  or
  g899
  (
    n986,
    n893,
    n905,
    n488,
    n436
  );


  xnor
  g900
  (
    n954,
    n848,
    n906,
    n898,
    n503
  );


  and
  g901
  (
    n1028,
    n424,
    n723,
    n896,
    n724
  );


  nand
  g902
  (
    n949,
    n903,
    n459,
    n441,
    n414
  );


  xor
  g903
  (
    n1009,
    n492,
    n692,
    n875,
    n489
  );


  xor
  g904
  (
    n980,
    n468,
    n885,
    n447,
    n425
  );


  or
  g905
  (
    n1069,
    n692,
    n888,
    n479,
    n433
  );


  xnor
  g906
  (
    n917,
    n479,
    n495,
    n886,
    n874
  );


  xnor
  g907
  (
    n1049,
    n411,
    n449,
    n420,
    n419
  );


  xnor
  g908
  (
    n998,
    n462,
    n435,
    n410,
    n409
  );


  or
  g909
  (
    n989,
    n894,
    n904,
    n491,
    n902
  );


  or
  g910
  (
    n1059,
    n850,
    n907,
    n506,
    n874
  );


  nand
  g911
  (
    n1045,
    n452,
    n430,
    n875,
    n872
  );


  nor
  g912
  (
    n963,
    n878,
    n438,
    n884,
    n413
  );


  nor
  g913
  (
    n1061,
    n489,
    n415,
    n890,
    n427
  );


  xnor
  g914
  (
    n1019,
    n472,
    n461,
    n412,
    n415
  );


  nand
  g915
  (
    n947,
    n844,
    n471,
    n902,
    n453
  );


  nor
  g916
  (
    n942,
    n878,
    n502,
    n889,
    n478
  );


  nor
  g917
  (
    n910,
    n422,
    n844,
    n457,
    n851
  );


  xnor
  g918
  (
    n1012,
    n472,
    n416,
    n871,
    n427
  );


  and
  g919
  (
    n967,
    n879,
    n848,
    n410,
    n466
  );


  xnor
  g920
  (
    n992,
    n471,
    n482,
    n446,
    n451
  );


  and
  g921
  (
    n918,
    n435,
    n440,
    n846,
    n426
  );


  xor
  g922
  (
    n927,
    n481,
    n897,
    n457,
    n466
  );


  or
  g923
  (
    n983,
    n909,
    n445,
    n885,
    n432
  );


  and
  g924
  (
    n988,
    n458,
    n426,
    n874,
    n434
  );


  and
  g925
  (
    n1021,
    n846,
    n505,
    n890,
    n454
  );


  xnor
  g926
  (
    n916,
    n844,
    n853,
    n499,
    n849
  );


  xnor
  g927
  (
    n1040,
    n464,
    n490,
    n907,
    n845
  );


  and
  g928
  (
    n1026,
    n430,
    n722,
    n421,
    n903
  );


  and
  g929
  (
    n1031,
    n909,
    n899,
    n883,
    n481
  );


  nor
  g930
  (
    n971,
    n469,
    n445,
    n419,
    n886
  );


  nor
  g931
  (
    n946,
    n899,
    n409,
    n475,
    n461
  );


  xor
  g932
  (
    n1055,
    n500,
    n847,
    n415
  );


  xnor
  g933
  (
    n941,
    n439,
    n499,
    n417,
    n435
  );


  nor
  g934
  (
    n931,
    n893,
    n724,
    n446,
    n480
  );


  xor
  g935
  (
    n1063,
    n413,
    n480,
    n446,
    n723
  );


  nand
  g936
  (
    n1060,
    n443,
    n452,
    n437,
    n496
  );


  xor
  g937
  (
    n990,
    n852,
    n480,
    n850,
    n458
  );


  and
  g938
  (
    n936,
    n904,
    n500,
    n456,
    n505
  );


  xnor
  g939
  (
    n1051,
    n425,
    n476,
    n872,
    n504
  );


  xnor
  g940
  (
    n959,
    n888,
    n881,
    n847,
    n474
  );


  xor
  g941
  (
    n1033,
    n447,
    n487,
    n480
  );


  xor
  g942
  (
    n1016,
    n498,
    n493,
    n872,
    n457
  );


  or
  g943
  (
    n993,
    n413,
    n467,
    n468,
    n444
  );


  and
  g944
  (
    n1057,
    n508,
    n906,
    n894,
    n886
  );


  and
  g945
  (
    n914,
    n882,
    n426,
    n424,
    n473
  );


  xor
  g946
  (
    n1052,
    n494,
    n896,
    n426,
    n468
  );


  xnor
  g947
  (
    n926,
    n433,
    n507,
    n463,
    n458
  );


  nor
  g948
  (
    n1062,
    n891,
    n502,
    n443,
    n504
  );


  nor
  g949
  (
    n1030,
    n443,
    n418,
    n446,
    n497
  );


  or
  g950
  (
    n925,
    n423,
    n508,
    n852,
    n456
  );


  and
  g951
  (
    n945,
    n849,
    n439,
    n462,
    n893
  );


  xor
  g952
  (
    n976,
    n498,
    n901,
    n432,
    n471
  );


  nand
  g953
  (
    n981,
    n431,
    n871,
    n897,
    n455
  );


  xor
  g954
  (
    n1032,
    n486,
    n479,
    n722,
    n444
  );


  or
  g955
  (
    n911,
    n420,
    n509,
    n899,
    n414
  );


  or
  g956
  (
    n1058,
    n491,
    n895,
    n908,
    n452
  );


  xor
  g957
  (
    n997,
    n892,
    n424,
    n474,
    n508
  );


  xor
  g958
  (
    n1034,
    n412,
    n430,
    n900
  );


  xor
  g959
  (
    n1050,
    n888,
    n468,
    n902,
    n432
  );


  xnor
  g960
  (
    n995,
    n510,
    n441,
    n490,
    n875
  );


  nand
  g961
  (
    n965,
    n903,
    n871,
    n880,
    n463
  );


  nand
  g962
  (
    n991,
    n427,
    n448,
    n507,
    n899
  );


  xnor
  g963
  (
    n974,
    n507,
    n484,
    n879,
    n904
  );


  nand
  g964
  (
    n937,
    n882,
    n491,
    n419,
    n662
  );


  nand
  g965
  (
    n923,
    n844,
    n467,
    n907,
    n484
  );


  xnor
  g966
  (
    n1046,
    n411,
    n412,
    n472,
    n443
  );


  and
  g967
  (
    n978,
    n848,
    n453,
    n475,
    n486
  );


  nor
  g968
  (
    KeyWire_0_21,
    n478,
    n431,
    n460
  );


  or
  g969
  (
    n1038,
    n433,
    n898,
    n693,
    n845
  );


  nand
  g970
  (
    n1064,
    n873,
    n455,
    n881,
    n889
  );


  xnor
  g971
  (
    n932,
    n506,
    n476,
    n442
  );


  nor
  g972
  (
    n969,
    n416,
    n503,
    n483,
    n448
  );


  and
  g973
  (
    n1035,
    n469,
    n909,
    n450,
    n423
  );


  nand
  g974
  (
    n1041,
    n889,
    n483,
    n485,
    n419
  );


  nand
  g975
  (
    n1022,
    n892,
    n438,
    n456,
    n889
  );


  xnor
  g976
  (
    n1004,
    n473,
    n434,
    n885,
    n883
  );


  nor
  g977
  (
    n966,
    n693,
    n879,
    n475,
    n465
  );


  xnor
  g978
  (
    n994,
    n428,
    n454,
    n906,
    n880
  );


  or
  g979
  (
    n1024,
    n415,
    n890,
    n463,
    n459
  );


  or
  g980
  (
    n1042,
    n487,
    n411,
    n440,
    n488
  );


  and
  g981
  (
    n1000,
    n485,
    n429,
    n474,
    n436
  );


  xnor
  g982
  (
    n921,
    n449,
    n431,
    n464,
    n481
  );


  xnor
  g983
  (
    n1001,
    n873,
    n501,
    n878,
    n425
  );


  and
  g984
  (
    n1008,
    n410,
    n467,
    n882,
    n486
  );


  nand
  g985
  (
    n1010,
    n498,
    n504,
    n500,
    n474
  );


  or
  g986
  (
    n1013,
    n874,
    n496,
    n870,
    n454
  );


  nand
  g987
  (
    n1018,
    n908,
    n876,
    n881,
    n897
  );


  xnor
  g988
  (
    n934,
    n494,
    n887,
    n417,
    n896
  );


  xor
  g989
  (
    n933,
    n425,
    n493,
    n905,
    n870
  );


  nor
  g990
  (
    n1017,
    n422,
    n428,
    n875,
    n873
  );


  xor
  g991
  (
    n940,
    n877,
    n438,
    n873,
    n900
  );


  nor
  g992
  (
    n1011,
    n503,
    n843,
    n905,
    n722
  );


  xor
  g993
  (
    n985,
    n465,
    n459,
    n879,
    n895
  );


  nand
  g994
  (
    n943,
    n895,
    n499,
    n724,
    n464
  );


  and
  g995
  (
    n1056,
    n477,
    n494,
    n461,
    n418
  );


  xnor
  g996
  (
    n913,
    n447,
    n499,
    n442,
    n420
  );


  and
  g997
  (
    n1006,
    n484,
    n477,
    n663
  );


  xor
  g998
  (
    n919,
    n483,
    n466,
    n487,
    n884
  );


  xnor
  g999
  (
    n970,
    n904,
    n501,
    n482,
    n429
  );


  nand
  g1000
  (
    n950,
    n432,
    n764,
    n880,
    n851
  );


  nor
  g1001
  (
    n928,
    n506,
    n885,
    n847,
    n492
  );


  or
  g1002
  (
    n955,
    n692,
    n506,
    n428,
    n901
  );


  xor
  g1003
  (
    n930,
    n877,
    n884,
    n430,
    n486
  );


  or
  g1004
  (
    n1015,
    n484,
    n489,
    n436,
    n507
  );


  and
  g1005
  (
    n953,
    n876,
    n850,
    n851,
    n505
  );


  or
  g1006
  (
    n912,
    n883,
    n664,
    n504,
    n483
  );


  and
  g1007
  (
    n982,
    n691,
    n436,
    n880,
    n427
  );


  nor
  g1008
  (
    n964,
    n470,
    n723,
    n887,
    n877
  );


  nand
  g1009
  (
    n1068,
    n663,
    n509,
    n453,
    n441
  );


  or
  g1010
  (
    n935,
    n872,
    n481,
    n423,
    n501
  );


  nand
  g1011
  (
    n999,
    n496,
    n435,
    n495,
    n451
  );


  xnor
  g1012
  (
    KeyWire_0_20,
    n493,
    n876,
    n476,
    n886
  );


  or
  g1013
  (
    n1048,
    n485,
    n849,
    n438,
    n478
  );


  xor
  g1014
  (
    KeyWire_0_6,
    n849,
    n439,
    n908,
    n455
  );


  or
  g1015
  (
    n1043,
    n470,
    n466,
    n891,
    n464
  );


  or
  g1016
  (
    n1047,
    n662,
    n437,
    n414,
    n460
  );


  or
  g1017
  (
    n1065,
    n898,
    n449,
    n892,
    n490
  );


  nand
  g1018
  (
    KeyWire_0_18,
    n456,
    n662,
    n663,
    n475
  );


  nor
  g1019
  (
    n938,
    n414,
    n489,
    n469,
    n495
  );


  xor
  g1020
  (
    n915,
    n482,
    n906,
    n509,
    n888
  );


  or
  g1021
  (
    n1025,
    n887,
    n870,
    n445
  );


  xor
  g1022
  (
    KeyWire_0_5,
    n421,
    n510,
    n420,
    n473
  );


  and
  g1023
  (
    n924,
    n502,
    n664,
    n460,
    n492
  );


  or
  g1024
  (
    n1023,
    n891,
    n901,
    n505,
    n465
  );


  or
  g1025
  (
    n956,
    n429,
    n497,
    n897,
    n892
  );


  and
  g1026
  (
    n987,
    n883,
    n445,
    n488,
    n469
  );


  or
  g1027
  (
    n977,
    n417,
    n437,
    n455
  );


  xor
  g1028
  (
    n952,
    n894,
    n490,
    n890,
    n853
  );


  xor
  g1029
  (
    n1067,
    n462,
    n664,
    n692,
    n498
  );


  nor
  g1030
  (
    n1036,
    n477,
    n722,
    n503,
    n423
  );


  and
  g1031
  (
    n944,
    n497,
    n845,
    n453,
    n458
  );


  and
  g1032
  (
    n957,
    n510,
    n424,
    n893,
    n459
  );


  xnor
  g1033
  (
    n973,
    n493,
    n495,
    n417,
    n409
  );


  nor
  g1034
  (
    n958,
    n409,
    n413,
    n431,
    n902
  );


  or
  g1035
  (
    n1039,
    n848,
    n422,
    n450,
    n845
  );


  nor
  g1036
  (
    n948,
    n907,
    n691,
    n441,
    n421
  );


  xnor
  g1037
  (
    n1262,
    n270,
    n1028,
    n553,
    n1015
  );


  nand
  g1038
  (
    n1083,
    n737,
    n808,
    n1012,
    n1023
  );


  nand
  g1039
  (
    KeyWire_0_11,
    n1061,
    n773,
    n1063,
    n1008
  );


  nor
  g1040
  (
    n1150,
    n994,
    n951,
    n552,
    n1050
  );


  xor
  g1041
  (
    n1257,
    n919,
    n986,
    n961,
    n978
  );


  nand
  g1042
  (
    n1291,
    n1003,
    n935,
    n930,
    n926
  );


  and
  g1043
  (
    n1140,
    n982,
    n910,
    n937,
    n1020
  );


  xnor
  g1044
  (
    n1287,
    n922,
    n753,
    n978,
    n911
  );


  nand
  g1045
  (
    n1085,
    n918,
    n541,
    n856,
    n953
  );


  or
  g1046
  (
    n1202,
    n270,
    n1066,
    n744,
    n939
  );


  xnor
  g1047
  (
    n1211,
    n937,
    n975,
    n1005,
    n1041
  );


  and
  g1048
  (
    n1204,
    n546,
    n1011,
    n46,
    n953
  );


  nor
  g1049
  (
    n1112,
    n960,
    n944,
    n926,
    n950
  );


  nand
  g1050
  (
    n1170,
    n923,
    n970,
    n911,
    n543
  );


  xnor
  g1051
  (
    n1159,
    n1014,
    n1006,
    n859,
    n1029
  );


  xnor
  g1052
  (
    n1217,
    n808,
    n945,
    n854,
    n1047
  );


  or
  g1053
  (
    n1205,
    n551,
    n986,
    n936,
    n928
  );


  xnor
  g1054
  (
    n1116,
    n1042,
    n991,
    n1045,
    n1064
  );


  and
  g1055
  (
    n1186,
    n1069,
    n740,
    n1062,
    n978
  );


  xor
  g1056
  (
    n1244,
    n965,
    n554,
    n928,
    n985
  );


  xor
  g1057
  (
    n1279,
    n923,
    n736,
    n966,
    n985
  );


  nor
  g1058
  (
    n1142,
    n982,
    n971,
    n985,
    n954
  );


  xnor
  g1059
  (
    n1254,
    n1050,
    n954,
    n1056,
    n992
  );


  nand
  g1060
  (
    n1160,
    n550,
    n1019,
    n1020,
    n1033
  );


  nand
  g1061
  (
    n1195,
    n981,
    n1022,
    n937,
    n1049
  );


  xor
  g1062
  (
    n1268,
    n1028,
    n1053,
    n1027,
    n755
  );


  xnor
  g1063
  (
    n1245,
    n952,
    n811,
    n924,
    n550
  );


  nand
  g1064
  (
    n1075,
    n998,
    n926,
    n1006,
    n549
  );


  xnor
  g1065
  (
    n1175,
    n934,
    n995,
    n988,
    n807
  );


  nor
  g1066
  (
    n1234,
    n746,
    n978,
    n949,
    n552
  );


  xnor
  g1067
  (
    n1249,
    n1060,
    n1008,
    n1018,
    n755
  );


  nor
  g1068
  (
    n1225,
    n757,
    n942,
    n1016,
    n918
  );


  nand
  g1069
  (
    n1276,
    n976,
    n930,
    n856,
    n1044
  );


  and
  g1070
  (
    n1221,
    n1009,
    n1037,
    n735,
    n541
  );


  and
  g1071
  (
    n1110,
    n748,
    n972,
    n749,
    n1068
  );


  or
  g1072
  (
    n1207,
    n949,
    n979,
    n1062,
    n664
  );


  nand
  g1073
  (
    n1278,
    n1007,
    n747,
    n944,
    n989
  );


  nor
  g1074
  (
    n1267,
    n960,
    n547,
    n553,
    n807
  );


  nor
  g1075
  (
    n1168,
    n809,
    n1044,
    n737,
    n1056
  );


  xor
  g1076
  (
    n1220,
    n1014,
    n547,
    n743,
    n1019
  );


  nand
  g1077
  (
    n1098,
    n547,
    n999,
    n968,
    n1057
  );


  or
  g1078
  (
    n1117,
    n1048,
    n758,
    n746,
    n1027
  );


  and
  g1079
  (
    n1103,
    n814,
    n812,
    n973,
    n996
  );


  nand
  g1080
  (
    n1105,
    n940,
    n736,
    n963,
    n932
  );


  nand
  g1081
  (
    n1269,
    n1031,
    n1043,
    n743,
    n736
  );


  nand
  g1082
  (
    n1199,
    n953,
    n1013,
    n950,
    n974
  );


  nor
  g1083
  (
    n1164,
    n1031,
    n957,
    n1000,
    n940
  );


  xnor
  g1084
  (
    n1184,
    n919,
    n1036,
    n970,
    n1009
  );


  xnor
  g1085
  (
    n1078,
    n1024,
    n815,
    n984,
    n46
  );


  and
  g1086
  (
    n1072,
    n1040,
    n912,
    n972,
    n539
  );


  nor
  g1087
  (
    n1143,
    n1000,
    n813,
    n950,
    n956
  );


  nor
  g1088
  (
    n1090,
    n915,
    n933,
    n1054,
    n857
  );


  xnor
  g1089
  (
    n1077,
    n554,
    n922,
    n983,
    n915
  );


  or
  g1090
  (
    n1114,
    n545,
    n1061,
    n962,
    n1052
  );


  xnor
  g1091
  (
    n1206,
    n747,
    n754,
    n739,
    n947
  );


  and
  g1092
  (
    n1136,
    n929,
    n938,
    n969,
    n983
  );


  or
  g1093
  (
    n1104,
    n813,
    n1034,
    n992,
    n972
  );


  nor
  g1094
  (
    n1224,
    n1067,
    n831,
    n47,
    n960
  );


  nor
  g1095
  (
    n1208,
    n927,
    n1040,
    n855,
    n924
  );


  nor
  g1096
  (
    n1274,
    n1052,
    n1059,
    n1056,
    n913
  );


  nand
  g1097
  (
    n1281,
    n749,
    n548,
    n816,
    n806
  );


  and
  g1098
  (
    n1091,
    n929,
    n927,
    n996,
    n1055
  );


  nor
  g1099
  (
    n1179,
    n1047,
    n975,
    n923,
    n1068
  );


  xor
  g1100
  (
    n1139,
    n757,
    n939,
    n977,
    n548
  );


  xnor
  g1101
  (
    n1174,
    n1023,
    n990,
    n807,
    n957
  );


  and
  g1102
  (
    n1129,
    n928,
    n981,
    n1044,
    n970
  );


  xnor
  g1103
  (
    n1203,
    n956,
    n1015,
    n542,
    n746
  );


  xor
  g1104
  (
    n1189,
    n999,
    n543,
    n1046,
    n1016
  );


  nand
  g1105
  (
    n1280,
    n1045,
    n1035,
    n980,
    n1025
  );


  xnor
  g1106
  (
    n1126,
    n1055,
    n815,
    n1002,
    n955
  );


  nand
  g1107
  (
    n1289,
    n1029,
    n975,
    n927,
    n982
  );


  nand
  g1108
  (
    n1149,
    n1030,
    n747,
    n817,
    n946
  );


  xor
  g1109
  (
    n1277,
    n548,
    n1021,
    n755,
    n973
  );


  nand
  g1110
  (
    n1188,
    n994,
    n1017,
    n1007,
    n997
  );


  nand
  g1111
  (
    n1080,
    n740,
    n1000,
    n1066,
    n976
  );


  nand
  g1112
  (
    n1183,
    n1030,
    n913,
    n933,
    n1013
  );


  nand
  g1113
  (
    n1232,
    n940,
    n944,
    n1039,
    n910
  );


  or
  g1114
  (
    n1194,
    n758,
    n989,
    n1034,
    n984
  );


  or
  g1115
  (
    n1210,
    n1041,
    n968,
    n753,
    n1018
  );


  nor
  g1116
  (
    KeyWire_0_31,
    n1038,
    n984,
    n271,
    n543
  );


  and
  g1117
  (
    n1215,
    n1052,
    n929,
    n771,
    n974
  );


  xor
  g1118
  (
    n1130,
    n540,
    n1057,
    n944,
    n917
  );


  and
  g1119
  (
    n1138,
    n965,
    n1065,
    n857,
    n983
  );


  or
  g1120
  (
    n1285,
    n1007,
    n748,
    n551,
    n1033
  );


  xor
  g1121
  (
    n1109,
    n741,
    n1040,
    n753,
    n993
  );


  or
  g1122
  (
    n1084,
    n811,
    n946,
    n990,
    n544
  );


  nor
  g1123
  (
    n1167,
    n1031,
    n1013,
    n810,
    n932
  );


  nand
  g1124
  (
    n1165,
    n1014,
    n749,
    n962,
    n974
  );


  and
  g1125
  (
    n1192,
    n973,
    n913,
    n946,
    n1025
  );


  nand
  g1126
  (
    n1171,
    n914,
    n1058,
    n958,
    n856
  );


  xnor
  g1127
  (
    n1230,
    n1028,
    n553,
    n1059,
    n1062
  );


  nor
  g1128
  (
    n1256,
    n1039,
    n1048,
    n740,
    n742
  );


  xnor
  g1129
  (
    n1227,
    n1065,
    n1048,
    n1002,
    n1024
  );


  xnor
  g1130
  (
    n1239,
    n942,
    n989,
    n827,
    n1038
  );


  xor
  g1131
  (
    n1082,
    n947,
    n1049,
    n1034,
    n1022
  );


  xor
  g1132
  (
    n1137,
    n977,
    n1021,
    n1064,
    n939
  );


  xnor
  g1133
  (
    n1190,
    n1020,
    n949,
    n751,
    n928
  );


  xor
  g1134
  (
    n1071,
    n936,
    n1042,
    n947,
    n801
  );


  and
  g1135
  (
    n1148,
    n810,
    n1003,
    n1057,
    n933
  );


  xnor
  g1136
  (
    n1162,
    n1054,
    n1009,
    n817,
    n1032
  );


  xnor
  g1137
  (
    n1182,
    n830,
    n808,
    n1006,
    n922
  );


  nor
  g1138
  (
    n1201,
    n813,
    n921,
    n992,
    n914
  );


  nand
  g1139
  (
    KeyWire_0_24,
    n752,
    n1016,
    n1038,
    n1023
  );


  xnor
  g1140
  (
    n1163,
    n1049,
    n1029,
    n969,
    n1000
  );


  xor
  g1141
  (
    n1158,
    n955,
    n999,
    n931,
    n745
  );


  or
  g1142
  (
    n1213,
    n921,
    n815,
    n1051,
    n922
  );


  nand
  g1143
  (
    n1151,
    n945,
    n965,
    n934,
    n693
  );


  nor
  g1144
  (
    n1156,
    n665,
    n1035,
    n986,
    n933
  );


  nor
  g1145
  (
    n1236,
    n805,
    n960,
    n918,
    n935
  );


  xnor
  g1146
  (
    n1197,
    n539,
    n957,
    n988,
    n807
  );


  nor
  g1147
  (
    n1096,
    n1065,
    n1055,
    n919,
    n859
  );


  nor
  g1148
  (
    n1264,
    n925,
    n993,
    n980,
    n754
  );


  nand
  g1149
  (
    n1284,
    n545,
    n1053,
    n949,
    n938
  );


  nand
  g1150
  (
    n1226,
    n1057,
    n919,
    n1026,
    n743
  );


  or
  g1151
  (
    n1176,
    n756,
    n923,
    n757,
    n1005
  );


  xor
  g1152
  (
    n1185,
    n1037,
    n929,
    n917,
    n991
  );


  and
  g1153
  (
    n1108,
    n1063,
    n1044,
    n971,
    n817
  );


  nand
  g1154
  (
    n1222,
    n951,
    n977,
    n829,
    n915
  );


  and
  g1155
  (
    n1122,
    n1043,
    n1064,
    n985,
    n917
  );


  or
  g1156
  (
    n1177,
    n549,
    n958,
    n981,
    n938
  );


  xnor
  g1157
  (
    n1273,
    n981,
    n948,
    n752,
    n910
  );


  xnor
  g1158
  (
    n1092,
    n806,
    n47,
    n271,
    n961
  );


  and
  g1159
  (
    n1219,
    n1049,
    n1031,
    n939,
    n920
  );


  nand
  g1160
  (
    n1248,
    n937,
    n1037,
    n735,
    n1042
  );


  or
  g1161
  (
    n1125,
    n756,
    n742,
    n1032,
    n987
  );


  xnor
  g1162
  (
    n1235,
    n745,
    n952,
    n270,
    n554
  );


  and
  g1163
  (
    n1266,
    n955,
    n930,
    n995,
    n815
  );


  or
  g1164
  (
    n1231,
    n912,
    n991,
    n921,
    n551
  );


  nor
  g1165
  (
    n1229,
    n751,
    n857,
    n977,
    n542
  );


  xnor
  g1166
  (
    n1087,
    n756,
    n914,
    n828,
    n1014
  );


  and
  g1167
  (
    n1134,
    n1001,
    n1040,
    n1060,
    n1018
  );


  or
  g1168
  (
    n1209,
    n1024,
    n1048,
    n1042,
    n855
  );


  xor
  g1169
  (
    n1118,
    n806,
    n941,
    n956,
    n774
  );


  and
  g1170
  (
    n1193,
    n1043,
    n1065,
    n1059,
    n854
  );


  nor
  g1171
  (
    n1181,
    n816,
    n967,
    n924,
    n1012
  );


  and
  g1172
  (
    n1153,
    n987,
    n735,
    n941
  );


  nor
  g1173
  (
    n1133,
    n959,
    n1061,
    n992
  );


  xnor
  g1174
  (
    n1146,
    n832,
    n744,
    n1018,
    n993
  );


  xnor
  g1175
  (
    n1074,
    n545,
    n809,
    n1017,
    n858
  );


  xnor
  g1176
  (
    n1272,
    n912,
    n996,
    n859,
    n271
  );


  xnor
  g1177
  (
    n1233,
    n936,
    n916,
    n747,
    n546
  );


  or
  g1178
  (
    n1144,
    n997,
    n756,
    n955,
    n920
  );


  and
  g1179
  (
    n1161,
    n754,
    n963,
    n855,
    n752
  );


  xor
  g1180
  (
    n1218,
    n1012,
    n924,
    n1053,
    n546
  );


  nand
  g1181
  (
    n1079,
    n995,
    n1026,
    n746,
    n967
  );


  nand
  g1182
  (
    n1107,
    n932,
    n757,
    n1060,
    n550
  );


  or
  g1183
  (
    n1094,
    n1041,
    n1035,
    n1025,
    n758
  );


  xnor
  g1184
  (
    n1157,
    n751,
    n1010,
    n1051,
    n1053
  );


  or
  g1185
  (
    n1251,
    n1005,
    n1050,
    n1041,
    n1021
  );


  xnor
  g1186
  (
    n1240,
    n968,
    n814,
    n809,
    n1004
  );


  nor
  g1187
  (
    n1070,
    n1068,
    n936,
    n1001,
    n1034
  );


  xor
  g1188
  (
    n1086,
    n858,
    n1036,
    n1033,
    n1038
  );


  nor
  g1189
  (
    n1252,
    n991,
    n1054,
    n1046,
    n542
  );


  xor
  g1190
  (
    n1120,
    n911,
    n854,
    n750,
    n1011
  );


  xor
  g1191
  (
    n1106,
    n1051,
    n814,
    n994,
    n988
  );


  nor
  g1192
  (
    n1246,
    n943,
    n665,
    n811,
    n1063
  );


  nor
  g1193
  (
    n1293,
    n1069,
    n1020,
    n943,
    n739
  );


  and
  g1194
  (
    n1088,
    n916,
    n951,
    n964,
    n1010
  );


  xnor
  g1195
  (
    n1076,
    n916,
    n810,
    n1047,
    n931
  );


  and
  g1196
  (
    n1154,
    n1007,
    n952,
    n665,
    n806
  );


  nand
  g1197
  (
    n1187,
    n1004,
    n966,
    n547,
    n753
  );


  and
  g1198
  (
    n1255,
    n814,
    n46,
    n1023,
    n976
  );


  nand
  g1199
  (
    n1200,
    n1008,
    n1003,
    n921,
    n1017
  );


  nand
  g1200
  (
    n1123,
    n545,
    n1010,
    n958,
    n966
  );


  xor
  g1201
  (
    n1212,
    n752,
    n745,
    n541,
    n974
  );


  and
  g1202
  (
    n1119,
    n1019,
    n979,
    n1067,
    n854
  );


  xor
  g1203
  (
    n1198,
    n1011,
    n541,
    n934,
    n1009
  );


  nand
  g1204
  (
    n1178,
    n926,
    n1026,
    n963,
    n748
  );


  xor
  g1205
  (
    n1228,
    n979,
    n542,
    n540,
    n956
  );


  xor
  g1206
  (
    n1135,
    n1013,
    n1046,
    n816,
    n979
  );


  nand
  g1207
  (
    n1131,
    n739,
    n693,
    n946,
    n930
  );


  or
  g1208
  (
    n1173,
    n665,
    n554,
    n975,
    n914
  );


  nor
  g1209
  (
    n1152,
    n927,
    n961,
    n1069,
    n931
  );


  xor
  g1210
  (
    n1124,
    n1055,
    n1060,
    n971,
    n1008
  );


  and
  g1211
  (
    n1095,
    n812,
    n925,
    n858,
    n1016
  );


  or
  g1212
  (
    n1270,
    n998,
    n947,
    n989,
    n47
  );


  nor
  g1213
  (
    n1100,
    n751,
    n1022,
    n1032,
    n1058
  );


  xnor
  g1214
  (
    n1238,
    n549,
    n269,
    n741,
    n952
  );


  nor
  g1215
  (
    n1113,
    n1012,
    n550,
    n742,
    n976
  );


  xnor
  g1216
  (
    n1166,
    n1001,
    n553,
    n971,
    n1036
  );


  nor
  g1217
  (
    n1259,
    n931,
    n962,
    n920,
    n857
  );


  or
  g1218
  (
    n1115,
    n858,
    n738,
    n1005,
    n964
  );


  and
  g1219
  (
    n1275,
    n750,
    n987,
    n738,
    n1054
  );


  xnor
  g1220
  (
    n1271,
    n962,
    n812,
    n940,
    n749
  );


  nand
  g1221
  (
    n1145,
    n998,
    n1029,
    n1033,
    n549
  );


  nor
  g1222
  (
    n1102,
    n915,
    n918,
    n910,
    n758
  );


  nand
  g1223
  (
    n1101,
    n953,
    n744,
    n997,
    n1050
  );


  and
  g1224
  (
    n1243,
    n988,
    n948,
    n1024,
    n540
  );


  nor
  g1225
  (
    n1258,
    n1045,
    n816,
    n1003,
    n935
  );


  xnor
  g1226
  (
    n1263,
    n271,
    n809,
    n913,
    n942
  );


  nor
  g1227
  (
    n1196,
    n738,
    n1046,
    n808,
    n995
  );


  nor
  g1228
  (
    n1260,
    n1039,
    n743,
    n1066
  );


  or
  g1229
  (
    n1180,
    n959,
    n813,
    n1037,
    n958
  );


  or
  g1230
  (
    n1250,
    n980,
    n1019,
    n741,
    n1001
  );


  nand
  g1231
  (
    n1214,
    n1021,
    n959,
    n1067,
    n982
  );


  or
  g1232
  (
    n1121,
    n945,
    n969,
    n1004,
    n993
  );


  xor
  g1233
  (
    n1253,
    n856,
    n999,
    n540,
    n943
  );


  and
  g1234
  (
    n1216,
    n1010,
    n1002,
    n954,
    n544
  );


  xor
  g1235
  (
    n1097,
    n1032,
    n1067,
    n1004,
    n1045
  );


  nand
  g1236
  (
    KeyWire_0_7,
    n1035,
    n942,
    n1002,
    n964
  );


  xnor
  g1237
  (
    n1241,
    n980,
    n772,
    n1062,
    n1022
  );


  xnor
  g1238
  (
    n1290,
    n750,
    n925,
    n1006,
    n544
  );


  xnor
  g1239
  (
    n1242,
    n1047,
    n1058,
    n954,
    n552
  );


  xor
  g1240
  (
    n1169,
    n748,
    n810,
    n750,
    n1052
  );


  xor
  g1241
  (
    n1292,
    n935,
    n970,
    n967,
    n986
  );


  nand
  g1242
  (
    n1099,
    n812,
    n1063,
    n1039,
    n1030
  );


  or
  g1243
  (
    n1141,
    n943,
    n941,
    n938,
    n543
  );


  nand
  g1244
  (
    n1127,
    n817,
    n551,
    n1068,
    n997
  );


  nor
  g1245
  (
    KeyWire_0_8,
    n754,
    n911,
    n965,
    n972
  );


  nand
  g1246
  (
    n1155,
    n969,
    n1064,
    n1043,
    n859
  );


  xor
  g1247
  (
    n1081,
    n948,
    n920,
    n1017,
    n1058
  );


  nand
  g1248
  (
    n1283,
    n964,
    n990,
    n1026,
    n917
  );


  or
  g1249
  (
    n1132,
    n1027,
    n737,
    n546,
    n996
  );


  nand
  g1250
  (
    n1282,
    n755,
    n1030,
    n987,
    n963
  );


  xor
  g1251
  (
    n1073,
    n990,
    n544,
    n1069,
    n916
  );


  xnor
  g1252
  (
    n1111,
    n998,
    n1056,
    n1051,
    n1015
  );


  and
  g1253
  (
    n1089,
    n951,
    n945,
    n811,
    n932
  );


  xor
  g1254
  (
    n1128,
    n1011,
    n1015,
    n1028,
    n745
  );


  or
  g1255
  (
    n1093,
    n548,
    n983,
    n270,
    n984
  );


  nand
  g1256
  (
    n1261,
    n968,
    n973,
    n957,
    n967
  );


  nand
  g1257
  (
    n1147,
    n948,
    n855,
    n1036,
    n1025
  );


  nor
  g1258
  (
    n1265,
    n961,
    n934,
    n744,
    n959
  );


  xnor
  g1259
  (
    n1172,
    n1027,
    n966,
    n552,
    n1059
  );


  and
  g1260
  (
    n1223,
    n925,
    n950,
    n912,
    n994
  );


  and
  g1261
  (
    n1425,
    n1128,
    n1151,
    n1123,
    n1236
  );


  xnor
  g1262
  (
    n1346,
    n1240,
    n1276,
    n1110,
    n1213
  );


  xnor
  g1263
  (
    n1307,
    n1190,
    n1085,
    n1116,
    n1133
  );


  or
  g1264
  (
    n1389,
    n1190,
    n1143,
    n1288,
    n1076
  );


  and
  g1265
  (
    n1374,
    n1072,
    n1091,
    n1104,
    n1233
  );


  or
  g1266
  (
    n1420,
    n1080,
    n1255,
    n1097,
    n1213
  );


  xor
  g1267
  (
    n1312,
    n1093,
    n1101,
    n1231,
    n1266
  );


  xnor
  g1268
  (
    n1490,
    n1269,
    n1282,
    n1141,
    n1281
  );


  xnor
  g1269
  (
    n1449,
    n1102,
    n1229,
    n1182,
    n1185
  );


  or
  g1270
  (
    n1495,
    n1149,
    n1211,
    n1125,
    n1235
  );


  nor
  g1271
  (
    n1394,
    n1132,
    n1258,
    n1205,
    n1087
  );


  xnor
  g1272
  (
    n1304,
    n1129,
    n1277,
    n1097,
    n1071
  );


  and
  g1273
  (
    n1470,
    n1131,
    n1114,
    n1126,
    n1107
  );


  xor
  g1274
  (
    n1403,
    n1282,
    n1152,
    n1256,
    n1181
  );


  xnor
  g1275
  (
    n1507,
    n1124,
    n1108,
    n1277,
    n1249
  );


  or
  g1276
  (
    n1356,
    n1160,
    n1242,
    n1282,
    n1094
  );


  xor
  g1277
  (
    n1428,
    n1115,
    n1148,
    n1177,
    n1090
  );


  xor
  g1278
  (
    n1376,
    n1140,
    n1291,
    n1212,
    n1257
  );


  and
  g1279
  (
    n1362,
    n1196,
    n1175,
    n1290,
    n1074
  );


  xnor
  g1280
  (
    n1316,
    n1167,
    n1155,
    n1246,
    n1267
  );


  and
  g1281
  (
    n1416,
    n1212,
    n1195,
    n1272,
    n1293
  );


  nor
  g1282
  (
    n1370,
    n1139,
    n1189,
    n1247,
    n1237
  );


  nand
  g1283
  (
    n1462,
    n1110,
    n1139,
    n1119,
    n1093
  );


  xnor
  g1284
  (
    n1322,
    n1156,
    n1283,
    n1292,
    n1163
  );


  xnor
  g1285
  (
    n1471,
    n1178,
    n1264,
    n1164,
    n1130
  );


  xor
  g1286
  (
    n1421,
    n1165,
    n1109,
    n1282,
    n1142
  );


  xnor
  g1287
  (
    n1438,
    n1289,
    n1079,
    n1179,
    n1105
  );


  nor
  g1288
  (
    n1415,
    n1188,
    n1241,
    n1131,
    n1115
  );


  xnor
  g1289
  (
    n1318,
    n1237,
    n1120,
    n1285,
    n1082
  );


  or
  g1290
  (
    n1332,
    n1177,
    n1113,
    n1143,
    n1110
  );


  xnor
  g1291
  (
    n1436,
    n1127,
    n1108,
    n1238,
    n1286
  );


  nor
  g1292
  (
    n1483,
    n1089,
    n1097,
    n1075,
    n1160
  );


  xnor
  g1293
  (
    n1479,
    n1221,
    n1105,
    n1126,
    n1186
  );


  or
  g1294
  (
    n1301,
    n1179,
    n1279,
    n1103,
    n1235
  );


  xor
  g1295
  (
    KeyWire_0_16,
    n1116,
    n1167,
    n1177,
    n1179
  );


  xor
  g1296
  (
    n1382,
    n1248,
    n1142,
    n1161,
    n1140
  );


  or
  g1297
  (
    n1377,
    n1157,
    n1100,
    n1225,
    n1143
  );


  xnor
  g1298
  (
    n1311,
    n1269,
    n666,
    n1160,
    n1208
  );


  nand
  g1299
  (
    n1514,
    n1267,
    n1121,
    n1172,
    n1236
  );


  nand
  g1300
  (
    n1313,
    n1252,
    n1119,
    n1258,
    n1235
  );


  nor
  g1301
  (
    n1342,
    n1089,
    n1073,
    n1117,
    n1072
  );


  xnor
  g1302
  (
    n1481,
    n1289,
    n1162,
    n666,
    n1200
  );


  xnor
  g1303
  (
    n1472,
    n1209,
    n1287,
    n1268,
    n1215
  );


  nand
  g1304
  (
    n1446,
    n1124,
    n1083,
    n1131,
    n1217
  );


  xor
  g1305
  (
    n1460,
    n1187,
    n1192,
    n1262,
    n1141
  );


  xnor
  g1306
  (
    n1482,
    n1266,
    n1274,
    n1194,
    n1228
  );


  xor
  g1307
  (
    n1417,
    n1222,
    n1198,
    n1226,
    n1103
  );


  xor
  g1308
  (
    n1489,
    n1170,
    n1146,
    n1149,
    n1259
  );


  or
  g1309
  (
    n1303,
    n1221,
    n1272,
    n1080,
    n1152
  );


  nor
  g1310
  (
    n1361,
    n1151,
    n1226,
    n1191,
    n1216
  );


  and
  g1311
  (
    n1458,
    n1088,
    n1177,
    n1191,
    n1225
  );


  or
  g1312
  (
    n1378,
    n1142,
    n1223,
    n1112,
    n1269
  );


  and
  g1313
  (
    n1320,
    n1241,
    n1291,
    n1111,
    n1092
  );


  or
  g1314
  (
    n1338,
    n1215,
    n1238,
    n1190,
    n1231
  );


  nor
  g1315
  (
    n1411,
    n1127,
    n1092,
    n1194
  );


  and
  g1316
  (
    n1372,
    n1217,
    n1186,
    n1117,
    n1261
  );


  nor
  g1317
  (
    n1328,
    n1073,
    n1271,
    n1285,
    n1292
  );


  or
  g1318
  (
    n1516,
    n1228,
    n1251,
    n1165,
    n1288
  );


  and
  g1319
  (
    n1352,
    n1211,
    n1226,
    n1196,
    n1085
  );


  nor
  g1320
  (
    n1430,
    n1183,
    n1237,
    n1113,
    n1293
  );


  and
  g1321
  (
    n1488,
    n1156,
    n1175,
    n1158,
    n1153
  );


  nand
  g1322
  (
    n1496,
    n1095,
    n1273,
    n1206,
    n1232
  );


  nand
  g1323
  (
    n1498,
    n1086,
    n1213,
    n1211,
    n1104
  );


  and
  g1324
  (
    n1401,
    n1140,
    n1144,
    n1170,
    n1287
  );


  nor
  g1325
  (
    n1456,
    n1247,
    n1108,
    n1261,
    n1226
  );


  and
  g1326
  (
    n1511,
    n1090,
    n1246,
    n1283,
    n1102
  );


  nand
  g1327
  (
    n1353,
    n1173,
    n1270,
    n1154,
    n1148
  );


  xnor
  g1328
  (
    n1497,
    n1180,
    n1133,
    n1184,
    n1250
  );


  nand
  g1329
  (
    n1339,
    n1223,
    n1133,
    n1122,
    n1183
  );


  or
  g1330
  (
    KeyWire_0_0,
    n1165,
    n1071,
    n1248,
    n1281
  );


  or
  g1331
  (
    n1494,
    n1206,
    n1170,
    n1214,
    n1227
  );


  nor
  g1332
  (
    n1468,
    n1174,
    n1124,
    n1199,
    n1201
  );


  nand
  g1333
  (
    n1418,
    n1091,
    n1189,
    n1086,
    n1252
  );


  and
  g1334
  (
    n1358,
    n1174,
    n1141,
    n1216,
    n1268
  );


  nand
  g1335
  (
    n1398,
    n1125,
    n1169,
    n1159,
    n1216
  );


  and
  g1336
  (
    n1347,
    n1160,
    n1247,
    n1252,
    n1081
  );


  or
  g1337
  (
    n1407,
    n1280,
    n1212,
    n1186,
    n1240
  );


  xor
  g1338
  (
    n1400,
    n1279,
    n1154,
    n1280,
    n1147
  );


  or
  g1339
  (
    n1331,
    n1122,
    n1080,
    n1287,
    n1152
  );


  or
  g1340
  (
    n1386,
    n1083,
    n1099,
    n1121,
    n1081
  );


  nand
  g1341
  (
    n1396,
    n1136,
    n1202,
    n1099,
    n1092
  );


  and
  g1342
  (
    n1393,
    n1227,
    n1240,
    n1210,
    n1112
  );


  nor
  g1343
  (
    n1310,
    n1135,
    n1222,
    n1279,
    n1229
  );


  nor
  g1344
  (
    n1329,
    n1206,
    n1252,
    n1253,
    n1203
  );


  nand
  g1345
  (
    n1493,
    n1225,
    n1070,
    n1090,
    n1157
  );


  and
  g1346
  (
    n1503,
    n1166,
    n1173,
    n1250,
    n1165
  );


  and
  g1347
  (
    n1423,
    n1098,
    n1185,
    n1288,
    n1265
  );


  nor
  g1348
  (
    n1431,
    n1104,
    n1260,
    n1076,
    n1263
  );


  nand
  g1349
  (
    KeyWire_0_13,
    n1171,
    n1083,
    n1145,
    n1166
  );


  nand
  g1350
  (
    n1379,
    n1121,
    n1107,
    n1284,
    n1197
  );


  xor
  g1351
  (
    n1445,
    n1264,
    n1256,
    n1275,
    n1118
  );


  xnor
  g1352
  (
    n1433,
    n1223,
    n1134,
    n1178,
    n1187
  );


  xor
  g1353
  (
    n1383,
    n1230,
    n1290,
    n1157,
    n1265
  );


  and
  g1354
  (
    n1515,
    n1119,
    n1146,
    n1192,
    n1246
  );


  or
  g1355
  (
    n1487,
    n1136,
    n1278,
    n1145,
    n1250
  );


  xor
  g1356
  (
    n1333,
    n1230,
    n1094,
    n1228,
    n1209
  );


  nand
  g1357
  (
    n1439,
    n1229,
    n1077,
    n1136,
    n1073
  );


  nor
  g1358
  (
    n1442,
    n1215,
    n1202,
    n1150,
    n1070
  );


  xnor
  g1359
  (
    n1505,
    n1258,
    n1205,
    n1173,
    n1267
  );


  or
  g1360
  (
    n1302,
    n1175,
    n1154,
    n1208,
    n1085
  );


  or
  g1361
  (
    n1457,
    n1269,
    n1258,
    n1137,
    n1130
  );


  nand
  g1362
  (
    n1512,
    n1163,
    n1162,
    n1142,
    n1147
  );


  xor
  g1363
  (
    n1300,
    n1134,
    n1166,
    n1169,
    n1164
  );


  nand
  g1364
  (
    n1484,
    n1107,
    n1285,
    n1135,
    n1224
  );


  or
  g1365
  (
    n1380,
    n1137,
    n1283,
    n1271,
    n1144
  );


  xor
  g1366
  (
    n1409,
    n1176,
    n1250,
    n1106,
    n1169
  );


  nor
  g1367
  (
    n1408,
    n1168,
    n1095,
    n1263,
    n1085
  );


  and
  g1368
  (
    n1478,
    n1260,
    n1265,
    n1243,
    n1233
  );


  nand
  g1369
  (
    n1381,
    n1217,
    n1257,
    n1204,
    n1273
  );


  nand
  g1370
  (
    n1508,
    n1193,
    n1150,
    n1245,
    n1232
  );


  xor
  g1371
  (
    n1467,
    n1126,
    n1234,
    n1111
  );


  xor
  g1372
  (
    n1350,
    n1260,
    n1219,
    n1277,
    n1171
  );


  or
  g1373
  (
    n1392,
    n1219,
    n1168,
    n1109,
    n1214
  );


  xor
  g1374
  (
    n1359,
    n1074,
    n1127,
    n1202,
    n1207
  );


  nor
  g1375
  (
    n1317,
    n1265,
    n1274,
    n1096,
    n1242
  );


  and
  g1376
  (
    n1469,
    n1147,
    n1276,
    n1271,
    n1267
  );


  xnor
  g1377
  (
    n1475,
    n1236,
    n1211,
    n1239,
    n1182
  );


  or
  g1378
  (
    n1360,
    n1170,
    n1194,
    n1159,
    n1144
  );


  xnor
  g1379
  (
    n1314,
    n1110,
    n1193,
    n1113,
    n1131
  );


  nor
  g1380
  (
    n1294,
    n1077,
    n1129,
    n1238,
    n1214
  );


  nor
  g1381
  (
    n1355,
    n1182,
    n1164,
    n1122,
    n1293
  );


  xor
  g1382
  (
    n1473,
    n1082,
    n1230,
    n1104,
    n1151
  );


  or
  g1383
  (
    n1345,
    n1161,
    n1158,
    n1219,
    n1138
  );


  and
  g1384
  (
    n1499,
    n1078,
    n1243,
    n1188,
    n1091
  );


  and
  g1385
  (
    n1435,
    n1123,
    n1158,
    n1183,
    n1257
  );


  and
  g1386
  (
    n1367,
    n1262,
    n1243,
    n1182,
    n1097
  );


  and
  g1387
  (
    n1506,
    n1120,
    n1126,
    n1163,
    n1286
  );


  xnor
  g1388
  (
    n1402,
    n1187,
    n1087,
    n1239,
    n1141
  );


  or
  g1389
  (
    n1452,
    n1236,
    n1289,
    n1204,
    n1183
  );


  xnor
  g1390
  (
    n1297,
    n1080,
    n1101,
    n1168,
    n1158
  );


  nand
  g1391
  (
    n1330,
    n1109,
    n1199,
    n1101,
    n1248
  );


  nor
  g1392
  (
    n1429,
    n1209,
    n1199,
    n1277,
    n1278
  );


  nor
  g1393
  (
    n1419,
    n1242,
    n1199,
    n1181,
    n1255
  );


  nand
  g1394
  (
    n1334,
    n1272,
    n1153,
    n1112,
    n1084
  );


  xor
  g1395
  (
    n1485,
    n1125,
    n1201,
    n1149,
    n1143
  );


  xnor
  g1396
  (
    n1455,
    n1145,
    n1118,
    n1254,
    n1233
  );


  nand
  g1397
  (
    n1413,
    n1087,
    n1244,
    n1280,
    n1275
  );


  xor
  g1398
  (
    n1369,
    n1168,
    n1224,
    n1113,
    n1253
  );


  xor
  g1399
  (
    n1405,
    n1195,
    n1218,
    n1230,
    n1118
  );


  nand
  g1400
  (
    n1465,
    n1161,
    n1292,
    n1208,
    n1102
  );


  or
  g1401
  (
    n1357,
    n1089,
    n1188,
    n1244,
    n1288
  );


  nor
  g1402
  (
    n1364,
    n1109,
    n1227,
    n1191,
    n1161
  );


  nand
  g1403
  (
    n1502,
    n1095,
    n1139,
    n1082,
    n1100
  );


  nand
  g1404
  (
    n1399,
    n1100,
    n1291,
    n1220,
    n1150
  );


  nor
  g1405
  (
    n1373,
    n1216,
    n1120,
    n1098,
    n1249
  );


  xor
  g1406
  (
    n1298,
    n1078,
    n1271,
    n1128,
    n1233
  );


  nand
  g1407
  (
    n1295,
    n1255,
    n1125,
    n1166,
    n1108
  );


  nand
  g1408
  (
    n1365,
    n1189,
    n1075,
    n1153,
    n1174
  );


  xor
  g1409
  (
    n1344,
    n1263,
    n1152,
    n1185,
    n1077
  );


  or
  g1410
  (
    n1513,
    n1086,
    n1087,
    n1175,
    n1195
  );


  or
  g1411
  (
    n1395,
    n1078,
    n1284,
    n1207,
    n1231
  );


  xor
  g1412
  (
    n1412,
    n1150,
    n1259,
    n1124,
    n1198
  );


  xnor
  g1413
  (
    n1349,
    n1246,
    n1074,
    n1094,
    n1244
  );


  nor
  g1414
  (
    n1406,
    n1137,
    n1209,
    n1180,
    n1286
  );


  xnor
  g1415
  (
    n1385,
    n1148,
    n1138,
    n1128,
    n1096
  );


  or
  g1416
  (
    n1480,
    n1088,
    n1270,
    n1192,
    n1190
  );


  or
  g1417
  (
    n1404,
    n1192,
    n1146,
    n1262,
    n1117
  );


  or
  g1418
  (
    n1422,
    n1093,
    n1210,
    n1203,
    n1201
  );


  nand
  g1419
  (
    n1444,
    n1284,
    n1254,
    n1147,
    n1081
  );


  or
  g1420
  (
    n1461,
    n1099,
    n1076,
    n1198,
    n1249
  );


  and
  g1421
  (
    n1424,
    n1207,
    n1291,
    n1204,
    n1084
  );


  nand
  g1422
  (
    n1440,
    n1081,
    n1188,
    n1220,
    n1195
  );


  xor
  g1423
  (
    n1437,
    n1123,
    n1268,
    n1134,
    n1263
  );


  nand
  g1424
  (
    n1391,
    n1116,
    n1272,
    n1082,
    n1171
  );


  nor
  g1425
  (
    n1340,
    n1084,
    n1249,
    n1244,
    n1114
  );


  nand
  g1426
  (
    n1348,
    n1121,
    n1135,
    n1273,
    n1218
  );


  xnor
  g1427
  (
    n1500,
    n1171,
    n1266,
    n1197,
    n1098
  );


  or
  g1428
  (
    n1375,
    n1245,
    n1293,
    n1106,
    n1207
  );


  nand
  g1429
  (
    n1459,
    n1203,
    n1278,
    n1130,
    n1210
  );


  or
  g1430
  (
    n1343,
    n1154,
    n1105,
    n1218,
    n1254
  );


  and
  g1431
  (
    n1326,
    n1107,
    n1260,
    n1248,
    n1231
  );


  xnor
  g1432
  (
    n1327,
    n1264,
    n1132,
    n1083,
    n1155
  );


  xnor
  g1433
  (
    n1309,
    n1079,
    n1114,
    n1202,
    n1187
  );


  nand
  g1434
  (
    n1341,
    n1157,
    n1096,
    n1163,
    n1219
  );


  nand
  g1435
  (
    n1363,
    n1281,
    n1071,
    n1111,
    n1144
  );


  xnor
  g1436
  (
    n1387,
    n1213,
    n1235,
    n1290,
    n1227
  );


  xor
  g1437
  (
    n1432,
    n1111,
    n1247,
    n1132,
    n1137
  );


  or
  g1438
  (
    n1368,
    n1253,
    n1120,
    n1234,
    n1224
  );


  xnor
  g1439
  (
    n1501,
    n1242,
    n1098,
    n1115,
    n1178
  );


  nand
  g1440
  (
    n1451,
    n1266,
    n1262,
    n1256,
    n1089
  );


  nor
  g1441
  (
    n1414,
    n1127,
    n1200,
    n1196,
    n1133
  );


  xnor
  g1442
  (
    n1476,
    n1243,
    n1217,
    n1279,
    n1123
  );


  or
  g1443
  (
    n1305,
    n1201,
    n1106,
    n1159,
    n1176
  );


  nand
  g1444
  (
    n1426,
    n1072,
    n1078,
    n1256,
    n1273
  );


  nand
  g1445
  (
    n1463,
    n1212,
    n1088,
    n1220,
    n1185
  );


  and
  g1446
  (
    n1325,
    n1178,
    n1220,
    n1117,
    n1118
  );


  nor
  g1447
  (
    n1443,
    n1241,
    n1270,
    n1181,
    n1180
  );


  nor
  g1448
  (
    n1371,
    n1134,
    n1251,
    n1114,
    n1156
  );


  xor
  g1449
  (
    n1454,
    n1283,
    n31,
    n1128,
    n1238
  );


  xnor
  g1450
  (
    n1474,
    n1254,
    n1139,
    n1261,
    n1289
  );


  xor
  g1451
  (
    n1308,
    n1136,
    n1234,
    n1162,
    n1261
  );


  or
  g1452
  (
    n1510,
    n1200,
    n1156,
    n1179,
    n1290
  );


  nor
  g1453
  (
    n1315,
    n1274,
    n1138,
    n1200,
    n1197
  );


  xor
  g1454
  (
    n1509,
    n1151,
    n1180,
    n1162,
    n1284
  );


  nor
  g1455
  (
    n1397,
    n1172,
    n1075,
    n1095,
    n1119
  );


  xor
  g1456
  (
    n1491,
    n1239,
    n1245,
    n1169,
    n1225
  );


  xor
  g1457
  (
    n1299,
    n1174,
    n1122,
    n1223,
    n1135
  );


  xnor
  g1458
  (
    n1337,
    n1155,
    n1264,
    n1091,
    n1206
  );


  nand
  g1459
  (
    n1450,
    n1218,
    n1112,
    n1251,
    n1132
  );


  nand
  g1460
  (
    n1354,
    n1079,
    n1245,
    n1129,
    n1203
  );


  nand
  g1461
  (
    n1466,
    n1255,
    n1176,
    n1205,
    n1099
  );


  nor
  g1462
  (
    n1427,
    n1197,
    n1224,
    n1285,
    n1094
  );


  xor
  g1463
  (
    n1464,
    n1159,
    n1155,
    n1240,
    n1259
  );


  and
  g1464
  (
    n1336,
    n1253,
    n1106,
    n1221,
    n1079
  );


  or
  g1465
  (
    n1296,
    n1093,
    n1268,
    n1232,
    n1222
  );


  xor
  g1466
  (
    n1492,
    n1205,
    n1101,
    n1086,
    n1130
  );


  and
  g1467
  (
    n1453,
    n1286,
    n1275,
    n1232,
    n1292
  );


  nand
  g1468
  (
    KeyWire_0_15,
    n1092,
    n1145,
    n1077,
    n1239
  );


  and
  g1469
  (
    n1486,
    n1184,
    n1193,
    n1275,
    n1090
  );


  or
  g1470
  (
    n1366,
    n1251,
    n1172,
    n1088,
    n1167
  );


  nand
  g1471
  (
    n1323,
    n1241,
    n1257,
    n1208,
    n1215
  );


  nor
  g1472
  (
    KeyWire_0_30,
    n1181,
    n1186,
    n1196,
    n1222
  );


  nor
  g1473
  (
    n1504,
    n1259,
    n1229,
    n1105,
    n1167
  );


  nand
  g1474
  (
    n1477,
    n1070,
    n1103,
    n1129,
    n1096
  );


  nor
  g1475
  (
    n1306,
    n1149,
    n1184,
    n1153,
    n1138
  );


  nand
  g1476
  (
    n1410,
    n1115,
    n1221,
    n1210,
    n1164
  );


  xnor
  g1477
  (
    n1441,
    n1278,
    n1148,
    n1146,
    n1184
  );


  and
  g1478
  (
    n1324,
    n1281,
    n1176,
    n1102,
    n1287
  );


  nor
  g1479
  (
    n1447,
    n1116,
    n1191,
    n1193,
    n1140
  );


  and
  g1480
  (
    n1319,
    n1280,
    n1172,
    n1084,
    n1204
  );


  or
  g1481
  (
    n1448,
    n1237,
    n1103,
    n1276,
    n1274
  );


  or
  g1482
  (
    n1388,
    n1100,
    n1276,
    n1270,
    n1228
  );


  nor
  g1483
  (
    n1321,
    n1198,
    n1214,
    n1173,
    n1189
  );


  xnor
  g1484
  (
    n1579,
    n1428,
    n1350,
    n1438,
    n1450
  );


  or
  g1485
  (
    n1554,
    n1364,
    n1348,
    n1314,
    n1473
  );


  xor
  g1486
  (
    n1544,
    n1512,
    n1353,
    n1401,
    n1514
  );


  nand
  g1487
  (
    n1677,
    n1388,
    n1502,
    n1317,
    n1498
  );


  xor
  g1488
  (
    n1662,
    n1459,
    n1341,
    n1452,
    n1368
  );


  and
  g1489
  (
    n1734,
    n1444,
    n1352,
    n1475,
    n1324
  );


  xor
  g1490
  (
    n1625,
    n1466,
    n1512,
    n1417,
    n1508
  );


  and
  g1491
  (
    n1732,
    n1488,
    n1347,
    n1316
  );


  or
  g1492
  (
    n1571,
    n1332,
    n1391,
    n1364,
    n1507
  );


  nand
  g1493
  (
    n1581,
    n1423,
    n1504,
    n1306,
    n1363
  );


  xnor
  g1494
  (
    n1519,
    n1328,
    n1362,
    n1485,
    n1513
  );


  nand
  g1495
  (
    n1576,
    n1392,
    n1472,
    n1511,
    n1407
  );


  xor
  g1496
  (
    n1657,
    n1409,
    n1369,
    n1489,
    n1346
  );


  xor
  g1497
  (
    n1574,
    n1441,
    n1328,
    n1395,
    n1458
  );


  and
  g1498
  (
    n1634,
    n1398,
    n1490,
    n1424,
    n1515
  );


  nor
  g1499
  (
    n1666,
    n1430,
    n1310,
    n1456,
    n1302
  );


  and
  g1500
  (
    n1523,
    n1451,
    n1403,
    n1463,
    n1322
  );


  or
  g1501
  (
    n1700,
    n1374,
    n1333,
    n1382,
    n1312
  );


  xnor
  g1502
  (
    n1702,
    n1315,
    n1379,
    n1354,
    n1394
  );


  xnor
  g1503
  (
    n1558,
    n1313,
    n1412,
    n1433,
    n1436
  );


  xnor
  g1504
  (
    n1578,
    n1422,
    n1453,
    n1472,
    n1326
  );


  xnor
  g1505
  (
    n1575,
    n1459,
    n1477,
    n1471,
    n1427
  );


  and
  g1506
  (
    n1589,
    n1407,
    n1372,
    n1363,
    n1305
  );


  and
  g1507
  (
    n1524,
    n1456,
    n1429,
    n1451,
    n1442
  );


  xor
  g1508
  (
    n1577,
    n1456,
    n1388,
    n1303,
    n1435
  );


  nor
  g1509
  (
    n1641,
    n1371,
    n1510,
    n1478,
    n1339
  );


  nor
  g1510
  (
    n1650,
    n1361,
    n1419,
    n1418,
    n1415
  );


  xor
  g1511
  (
    n1737,
    n1460,
    n1508,
    n1400,
    n1326
  );


  xnor
  g1512
  (
    n1729,
    n1389,
    n1373,
    n1329,
    n1372
  );


  or
  g1513
  (
    n1614,
    n1321,
    n1428,
    n1431,
    n1492
  );


  nand
  g1514
  (
    n1553,
    n1509,
    n1481,
    n1338,
    n1300
  );


  xor
  g1515
  (
    n1550,
    n1416,
    n1346,
    n1495,
    n1499
  );


  or
  g1516
  (
    n1704,
    n1306,
    n1435,
    n1438,
    n1479
  );


  or
  g1517
  (
    n1613,
    n1387,
    n1358,
    n1337
  );


  nand
  g1518
  (
    n1727,
    n1303,
    n1439,
    n1404,
    n1340
  );


  nand
  g1519
  (
    n1527,
    n1419,
    n1358,
    n1462,
    n1496
  );


  xnor
  g1520
  (
    n1628,
    n1431,
    n1407,
    n1414,
    n1297
  );


  nand
  g1521
  (
    n1537,
    n1383,
    n1308,
    n1353,
    n1349
  );


  xor
  g1522
  (
    n1563,
    n1323,
    n1326,
    n1456,
    n1385
  );


  nor
  g1523
  (
    KeyWire_0_10,
    n1366,
    n1496,
    n1498,
    n1304
  );


  or
  g1524
  (
    n1556,
    n1480,
    n1309,
    n1365,
    n1345
  );


  nor
  g1525
  (
    n1646,
    n1318,
    n47,
    n1379,
    n1311
  );


  nand
  g1526
  (
    n1719,
    n1473,
    n1303,
    n1379,
    n1338
  );


  xnor
  g1527
  (
    n1633,
    n1322,
    n1408,
    n1357,
    n1487
  );


  and
  g1528
  (
    n1687,
    n1372,
    n1373,
    n1465,
    n1403
  );


  xor
  g1529
  (
    n1659,
    n1450,
    n1437,
    n1365,
    n1487
  );


  or
  g1530
  (
    n1663,
    n1304,
    n1457,
    n1445
  );


  xor
  g1531
  (
    n1543,
    n1437,
    n1481,
    n1446,
    n1324
  );


  nor
  g1532
  (
    n1683,
    n1464,
    n1384,
    n1310,
    n1496
  );


  or
  g1533
  (
    n1540,
    n1493,
    n1318,
    n1407,
    n1400
  );


  nand
  g1534
  (
    n1552,
    n1306,
    n1497,
    n1422,
    n1516
  );


  nor
  g1535
  (
    n1522,
    n1406,
    n1307,
    n1327,
    n1437
  );


  or
  g1536
  (
    n1671,
    n1393,
    n1447,
    n1478,
    n1469
  );


  or
  g1537
  (
    n1642,
    n1420,
    n1512,
    n1354,
    n1460
  );


  and
  g1538
  (
    n1603,
    n1350,
    n1304,
    n1502,
    n1334
  );


  xnor
  g1539
  (
    n1602,
    n1314,
    n1402,
    n1370,
    n1498
  );


  nand
  g1540
  (
    n1626,
    n1444,
    n1365,
    n1449,
    n1468
  );


  nor
  g1541
  (
    n1736,
    n1321,
    n1415,
    n1381,
    n1302
  );


  and
  g1542
  (
    n1730,
    n1359,
    n1441,
    n1454,
    n1450
  );


  nor
  g1543
  (
    n1731,
    n1387,
    n1339,
    n1467,
    n1470
  );


  xnor
  g1544
  (
    n1681,
    n1434,
    n1463,
    n1457,
    n1360
  );


  or
  g1545
  (
    n1692,
    n1313,
    n1340,
    n1367,
    n1493
  );


  nor
  g1546
  (
    n1528,
    n1469,
    n1497,
    n1355,
    n1433
  );


  xnor
  g1547
  (
    n1584,
    n1486,
    n1461,
    n1506,
    n1323
  );


  xnor
  g1548
  (
    n1653,
    n1413,
    n1376,
    n1446,
    n1425
  );


  and
  g1549
  (
    n1706,
    n1380,
    n1497,
    n1342,
    n1317
  );


  nand
  g1550
  (
    n1620,
    n1300,
    n1447,
    n1296,
    n1377
  );


  nand
  g1551
  (
    n1604,
    n1362,
    n1398,
    n1417,
    n1485
  );


  nand
  g1552
  (
    n1612,
    n1435,
    n1455,
    n1308,
    n1454
  );


  nor
  g1553
  (
    n1708,
    n1514,
    n1496,
    n1470,
    n1392
  );


  nor
  g1554
  (
    n1643,
    n1467,
    n1477,
    n1413,
    n1451
  );


  nor
  g1555
  (
    n1517,
    n1416,
    n1322,
    n1373,
    n1406
  );


  xor
  g1556
  (
    n1638,
    n1409,
    n1509,
    n1368,
    n1396
  );


  xor
  g1557
  (
    n1649,
    n1472,
    n1411,
    n1310,
    n1403
  );


  nor
  g1558
  (
    n1593,
    n1452,
    n1421,
    n1408,
    n1454
  );


  and
  g1559
  (
    n1722,
    n1381,
    n1360,
    n1462,
    n1463
  );


  xor
  g1560
  (
    n1618,
    n1475,
    n1423,
    n1354
  );


  xor
  g1561
  (
    n1733,
    n1301,
    n1395,
    n1346,
    n1446
  );


  xnor
  g1562
  (
    n1712,
    n1458,
    n1367,
    n1507,
    n1359
  );


  or
  g1563
  (
    n1627,
    n1396,
    n1361,
    n1431,
    n1339
  );


  xor
  g1564
  (
    KeyWire_0_25,
    n1302,
    n1331,
    n1439,
    n1457
  );


  or
  g1565
  (
    n1601,
    n1468,
    n1351,
    n1367,
    n1412
  );


  nand
  g1566
  (
    n1640,
    n1390,
    n1405,
    n1343,
    n1329
  );


  or
  g1567
  (
    n1565,
    n1486,
    n1316,
    n1452,
    n1345
  );


  and
  g1568
  (
    n1559,
    n1397,
    n1298,
    n1402,
    n1384
  );


  xor
  g1569
  (
    n1717,
    n1482,
    n1330,
    n1448,
    n1465
  );


  or
  g1570
  (
    n1645,
    n1307,
    n1479,
    n1378,
    n1320
  );


  nor
  g1571
  (
    n1606,
    n1370,
    n1373,
    n1458,
    n1414
  );


  nand
  g1572
  (
    n1549,
    n1342,
    n1419,
    n1320,
    n1481
  );


  nor
  g1573
  (
    n1548,
    n1384,
    n1336,
    n1495,
    n1399
  );


  xor
  g1574
  (
    n1639,
    n1434,
    n1442,
    n1483,
    n1443
  );


  nand
  g1575
  (
    n1592,
    n1461,
    n1349,
    n1318,
    n1431
  );


  xnor
  g1576
  (
    n1623,
    n1389,
    n1503,
    n1467,
    n1433
  );


  nor
  g1577
  (
    n1699,
    n1347,
    n1424,
    n1502,
    n1506
  );


  nor
  g1578
  (
    n1680,
    n1472,
    n1341,
    n1444,
    n1342
  );


  or
  g1579
  (
    n1674,
    n1386,
    n1358,
    n1355,
    n1463
  );


  xnor
  g1580
  (
    n1595,
    n1515,
    n1320,
    n1343,
    n1351
  );


  xnor
  g1581
  (
    n1709,
    n1347,
    n1468,
    n1328,
    n1491
  );


  xor
  g1582
  (
    n1580,
    n1480,
    n1363,
    n1402,
    n1484
  );


  nor
  g1583
  (
    n1648,
    n1466,
    n1379,
    n1438,
    n1313
  );


  nand
  g1584
  (
    n1529,
    n1511,
    n1410,
    n1397,
    n1386
  );


  nor
  g1585
  (
    n1518,
    n1319,
    n1396,
    n1478,
    n1349
  );


  xor
  g1586
  (
    n1624,
    n1304,
    n1490,
    n1505,
    n1514
  );


  xor
  g1587
  (
    n1694,
    n1418,
    n1338,
    n1447,
    n1422
  );


  nor
  g1588
  (
    n1570,
    n1412,
    n1387,
    n1417,
    n1388
  );


  nand
  g1589
  (
    n1534,
    n1455,
    n1315,
    n1305,
    n1399
  );


  nor
  g1590
  (
    n1586,
    n1475,
    n1476,
    n1482,
    n1294
  );


  xor
  g1591
  (
    n1698,
    n1360,
    n1438,
    n1459,
    n1488
  );


  nor
  g1592
  (
    n1555,
    n1399,
    n1426,
    n1479,
    n1323
  );


  or
  g1593
  (
    n1567,
    n1508,
    n1516,
    n1426,
    n1483
  );


  and
  g1594
  (
    n1545,
    n1321,
    n1377,
    n1420,
    n1471
  );


  xnor
  g1595
  (
    n1568,
    n1380,
    n1375,
    n1345,
    n1348
  );


  xor
  g1596
  (
    n1686,
    n1376,
    n1454,
    n1491,
    n1295
  );


  xnor
  g1597
  (
    n1661,
    n1421,
    n1319,
    n1366,
    n1329
  );


  nand
  g1598
  (
    n1693,
    n1513,
    n1503,
    n1380,
    n1448
  );


  and
  g1599
  (
    n1521,
    n1381,
    n1432,
    n1352,
    n1404
  );


  xor
  g1600
  (
    n1689,
    n1319,
    n1308,
    n1474,
    n1306
  );


  xnor
  g1601
  (
    n1738,
    n1412,
    n1404,
    n1411,
    n1318
  );


  nor
  g1602
  (
    n1608,
    n1299,
    n1500,
    n1473,
    n1295
  );


  xnor
  g1603
  (
    n1673,
    n1443,
    n1389,
    n1416,
    n1405
  );


  and
  g1604
  (
    n1696,
    n1444,
    n1436,
    n1411,
    n1465
  );


  and
  g1605
  (
    n1611,
    n1339,
    n1359,
    n1426,
    n1303
  );


  xor
  g1606
  (
    n1536,
    n1333,
    n1425,
    n1474,
    n1351
  );


  and
  g1607
  (
    KeyWire_0_29,
    n1309,
    n1314,
    n1455,
    n1377
  );


  nand
  g1608
  (
    n1551,
    n1485,
    n1294,
    n1374,
    n1361
  );


  xor
  g1609
  (
    n1609,
    n1432,
    n1393,
    n1415,
    n1335
  );


  and
  g1610
  (
    n1658,
    n1374,
    n1500,
    n1473,
    n1395
  );


  nor
  g1611
  (
    n1530,
    n1500,
    n1462,
    n1507,
    n1427
  );


  xnor
  g1612
  (
    n1591,
    n1301,
    n1360,
    n1428,
    n32
  );


  nand
  g1613
  (
    n1560,
    n1425,
    n1322,
    n1397,
    n1419
  );


  xor
  g1614
  (
    n1675,
    n1376,
    n1371,
    n1418,
    n1448
  );


  xnor
  g1615
  (
    n1590,
    n1488,
    n1466,
    n1350,
    n1391
  );


  nor
  g1616
  (
    n1587,
    n1354,
    n1482,
    n1387,
    n1461
  );


  and
  g1617
  (
    n1678,
    n1483,
    n1507,
    n1409,
    n1505
  );


  and
  g1618
  (
    n1619,
    n1491,
    n1296,
    n1501,
    n1510
  );


  xor
  g1619
  (
    n1520,
    n1470,
    n1491,
    n1469,
    n1493
  );


  nor
  g1620
  (
    n1665,
    n1352,
    n1316,
    n1357,
    n1446
  );


  xor
  g1621
  (
    n1713,
    n1404,
    n1340,
    n1332,
    n1486
  );


  and
  g1622
  (
    n1573,
    n1406,
    n1490,
    n1474,
    n1460
  );


  nand
  g1623
  (
    n1644,
    n1380,
    n1504,
    n1309,
    n1297
  );


  nand
  g1624
  (
    n1716,
    n1516,
    n1401,
    n1329,
    n1324
  );


  xnor
  g1625
  (
    n1541,
    n1350,
    n1362,
    n1297,
    n1390
  );


  or
  g1626
  (
    n1637,
    n1504,
    n1341,
    n1410,
    n1513
  );


  nor
  g1627
  (
    n1724,
    n1461,
    n1345,
    n1443,
    n1457
  );


  xnor
  g1628
  (
    n1564,
    n1364,
    n1436,
    n1386,
    n1335
  );


  nor
  g1629
  (
    n1651,
    n1343,
    n1489,
    n1482,
    n1475
  );


  or
  g1630
  (
    n1703,
    n1343,
    n1492,
    n1390,
    n1501
  );


  xnor
  g1631
  (
    n1685,
    n1384,
    n1476,
    n1432,
    n1366
  );


  xor
  g1632
  (
    n1533,
    n1503,
    n1331,
    n1296,
    n1405
  );


  or
  g1633
  (
    n1664,
    n1369,
    n1374,
    n1477,
    n1357
  );


  nor
  g1634
  (
    n1654,
    n1426,
    n1479,
    n1401
  );


  nor
  g1635
  (
    n1631,
    n1487,
    n1316,
    n1489,
    n1506
  );


  nor
  g1636
  (
    n1667,
    n1344,
    n1311,
    n1376,
    n1395
  );


  or
  g1637
  (
    n1594,
    n1307,
    n1390,
    n1312,
    n1497
  );


  xnor
  g1638
  (
    n1688,
    n1480,
    n1427,
    n1369,
    n1414
  );


  and
  g1639
  (
    n1726,
    n1483,
    n1301,
    n1305,
    n1372
  );


  and
  g1640
  (
    n1635,
    n1295,
    n1314,
    n1476,
    n1338
  );


  nor
  g1641
  (
    n1598,
    n1417,
    n1335,
    n1448,
    n1405
  );


  xnor
  g1642
  (
    n1632,
    n1326,
    n1484,
    n1394,
    n1381
  );


  nor
  g1643
  (
    n1690,
    n1508,
    n1359,
    n1495,
    n1308
  );


  and
  g1644
  (
    n1630,
    n1367,
    n1356,
    n1363,
    n1319
  );


  xor
  g1645
  (
    n1582,
    n1436,
    n1383,
    n1453,
    n1349
  );


  xnor
  g1646
  (
    n1526,
    n1348,
    n1481,
    n1300,
    n1382
  );


  xnor
  g1647
  (
    n1636,
    n1435,
    n1433,
    n1499,
    n1430
  );


  nor
  g1648
  (
    n1656,
    n1298,
    n1449,
    n1311,
    n1414
  );


  or
  g1649
  (
    n1629,
    n1310,
    n1332,
    n1430,
    n1327
  );


  and
  g1650
  (
    n1622,
    n1492,
    n1471,
    n1515,
    n1452
  );


  nor
  g1651
  (
    n1714,
    n1368,
    n1309,
    n1447,
    n1490
  );


  xnor
  g1652
  (
    n1705,
    n1382,
    n1351,
    n1385,
    n1509
  );


  nand
  g1653
  (
    n1672,
    n1403,
    n1429,
    n1512,
    n1396
  );


  or
  g1654
  (
    n1605,
    n1346,
    n1440,
    n1474,
    n1406
  );


  xor
  g1655
  (
    n1615,
    n1334,
    n1420,
    n1353,
    n1429
  );


  xnor
  g1656
  (
    n1588,
    n1495,
    n1441,
    n1344,
    n1402
  );


  and
  g1657
  (
    n1691,
    n1332,
    n1453,
    n1356,
    n1352
  );


  and
  g1658
  (
    n1676,
    n1325,
    n1468,
    n1398,
    n1477
  );


  and
  g1659
  (
    n1621,
    n1410,
    n1509,
    n1388,
    n1383
  );


  xor
  g1660
  (
    n1728,
    n1315,
    n1439,
    n1421,
    n1370
  );


  xor
  g1661
  (
    n1600,
    n1321,
    n1445,
    n1498,
    n1333
  );


  or
  g1662
  (
    n1569,
    n1335,
    n1485,
    n1328,
    n1399
  );


  nand
  g1663
  (
    n1725,
    n1442,
    n1421,
    n1408,
    n1334
  );


  and
  g1664
  (
    n1670,
    n1441,
    n1443,
    n1458,
    n1440
  );


  or
  g1665
  (
    n1585,
    n1501,
    n1302,
    n1344,
    n1331
  );


  xor
  g1666
  (
    n1596,
    n1451,
    n1364,
    n1356,
    n1400
  );


  nand
  g1667
  (
    n1715,
    n1449,
    n1400,
    n1392,
    n1434
  );


  or
  g1668
  (
    n1599,
    n1409,
    n1410,
    n1299,
    n1393
  );


  xnor
  g1669
  (
    n1542,
    n1506,
    n1511,
    n1317,
    n1486
  );


  xnor
  g1670
  (
    n1707,
    n1348,
    n1413,
    n1375,
    n1337
  );


  xor
  g1671
  (
    n1647,
    n1429,
    n1355,
    n1386,
    n1342
  );


  and
  g1672
  (
    n1597,
    n1470,
    n1325,
    n1418,
    n1385
  );


  or
  g1673
  (
    n1735,
    n1434,
    n1305,
    n1413,
    n1313
  );


  xnor
  g1674
  (
    n1557,
    n1355,
    n1510,
    n1377,
    n1462
  );


  xor
  g1675
  (
    n1669,
    n1378,
    n1391,
    n1494,
    n1424
  );


  nor
  g1676
  (
    n1525,
    n1484,
    n1516,
    n31,
    n1450
  );


  and
  g1677
  (
    n1547,
    n1340,
    n1437,
    n1432,
    n1370
  );


  nor
  g1678
  (
    n1607,
    n1453,
    n1424,
    n1389,
    n1385
  );


  and
  g1679
  (
    n1610,
    n1411,
    n1362,
    n1330,
    n1478
  );


  nor
  g1680
  (
    n1679,
    n1459,
    n1449,
    n1476,
    n1333
  );


  xor
  g1681
  (
    n1684,
    n1294,
    n1327,
    n1492,
    n1422
  );


  nor
  g1682
  (
    n1566,
    n1331,
    n1330,
    n1398,
    n1430
  );


  nand
  g1683
  (
    n1616,
    n1442,
    n1341,
    n1510,
    n1505
  );


  nand
  g1684
  (
    n1697,
    n1466,
    n1336,
    n1501,
    n1369
  );


  xnor
  g1685
  (
    n1583,
    n1325,
    n1488,
    n1336,
    n1358
  );


  or
  g1686
  (
    n1695,
    n1503,
    n1356,
    n1494,
    n1392
  );


  or
  g1687
  (
    n1711,
    n1511,
    n1325,
    n1312,
    n1315
  );


  or
  g1688
  (
    n1546,
    n1502,
    n1440,
    n1471,
    n1365
  );


  and
  g1689
  (
    n1701,
    n1375,
    n1378,
    n1494,
    n1330
  );


  nor
  g1690
  (
    n1538,
    n1337,
    n1464,
    n1383,
    n1371
  );


  nor
  g1691
  (
    n1539,
    n1375,
    n1327,
    n1324,
    n1361
  );


  nor
  g1692
  (
    n1562,
    n1420,
    n1500,
    n1425,
    n1489
  );


  xor
  g1693
  (
    n1572,
    n1484,
    n1394,
    n1323,
    n1336
  );


  nor
  g1694
  (
    n1682,
    n1494,
    n1334,
    n1415,
    n1312
  );


  nand
  g1695
  (
    n1668,
    n1480,
    n1467,
    n1504,
    n1493
  );


  and
  g1696
  (
    n1532,
    n1393,
    n1499,
    n1469,
    n1439
  );


  xnor
  g1697
  (
    n1710,
    n1487,
    n1465,
    n1394,
    n1317
  );


  xnor
  g1698
  (
    n1721,
    n1357,
    n1460,
    n1499,
    n1391
  );


  nor
  g1699
  (
    n1660,
    n1344,
    n1416,
    n1298,
    n1382
  );


  nor
  g1700
  (
    n1561,
    n1378,
    n1366,
    n1397,
    n1455
  );


  xnor
  g1701
  (
    n1535,
    n1445,
    n1299,
    n1371,
    n1427
  );


  nor
  g1702
  (
    n1652,
    n1464,
    n1428,
    n1423,
    n1368
  );


  xnor
  g1703
  (
    n1531,
    n1307,
    n1301,
    n1505,
    n1311
  );


  or
  g1704
  (
    n1718,
    n1513,
    n1464,
    n1514,
    n1353
  );


  nor
  g1705
  (
    n1655,
    n1515,
    n1440,
    n1408,
    n1320
  );


  and
  g1706
  (
    n1884,
    n1621,
    n1563,
    n1567,
    n1541
  );


  xnor
  g1707
  (
    n1896,
    n1565,
    n1727,
    n1606,
    n1613
  );


  nand
  g1708
  (
    n1793,
    n1728,
    n1645,
    n1671,
    n1578
  );


  xnor
  g1709
  (
    n1849,
    n1711,
    n1517,
    n1717,
    n1703
  );


  and
  g1710
  (
    n1876,
    n1625,
    n1531,
    n1551,
    n1605
  );


  nand
  g1711
  (
    n1914,
    n1585,
    n1737,
    n1658,
    n1642
  );


  or
  g1712
  (
    n1819,
    n1632,
    n1648,
    n1699,
    n1573
  );


  or
  g1713
  (
    n1838,
    n1596,
    n1704,
    n1627,
    n1593
  );


  xnor
  g1714
  (
    n1773,
    n1543,
    n1706,
    n1704,
    n1617
  );


  nor
  g1715
  (
    n1790,
    n1689,
    n1641,
    n1732,
    n1547
  );


  xor
  g1716
  (
    n1753,
    n1638,
    n1636,
    n1732,
    n1551
  );


  xor
  g1717
  (
    n1829,
    n1654,
    n1630,
    n1575,
    n1722
  );


  nand
  g1718
  (
    n1833,
    n1637,
    n1614,
    n1710,
    n1576
  );


  and
  g1719
  (
    n1780,
    n1640,
    n1705,
    n1582,
    n1583
  );


  xnor
  g1720
  (
    n1824,
    n1655,
    n1648,
    n1571,
    n1595
  );


  xor
  g1721
  (
    n1840,
    n1565,
    n1578,
    n1686,
    n1643
  );


  and
  g1722
  (
    n1902,
    n1602,
    n1667,
    n1646,
    n1556
  );


  nand
  g1723
  (
    n1885,
    n1611,
    n1644,
    n1642,
    n1656
  );


  xor
  g1724
  (
    n1888,
    n1699,
    n1560,
    n1738,
    n1656
  );


  nor
  g1725
  (
    n1825,
    n1675,
    n1702,
    n1691,
    n1733
  );


  xnor
  g1726
  (
    n1889,
    n1635,
    n1629,
    n1518,
    n1553
  );


  nand
  g1727
  (
    n1760,
    n1583,
    n1591,
    n1521,
    n1604
  );


  and
  g1728
  (
    n1918,
    n1631,
    n1597,
    n1560,
    n1737
  );


  nand
  g1729
  (
    n1774,
    n1639,
    n1718,
    n1727,
    n1553
  );


  or
  g1730
  (
    n1746,
    n1634,
    n1583,
    n1563,
    n1690
  );


  nand
  g1731
  (
    n1750,
    n1707,
    n1733,
    n1584,
    n1628
  );


  xnor
  g1732
  (
    n1766,
    n1560,
    n1729,
    n1718,
    n1534
  );


  nor
  g1733
  (
    n1878,
    n1629,
    n1536,
    n1685,
    n1535
  );


  nand
  g1734
  (
    n1910,
    n1655,
    n1543,
    n1602,
    n1552
  );


  nand
  g1735
  (
    n1768,
    n1547,
    n1604,
    n1586,
    n1700
  );


  nor
  g1736
  (
    n1795,
    n1558,
    n1719,
    n1595,
    n1628
  );


  xnor
  g1737
  (
    n1908,
    n1708,
    n1546,
    n1698,
    n1662
  );


  nor
  g1738
  (
    n1786,
    n1540,
    n1712,
    n1681,
    n1710
  );


  nand
  g1739
  (
    n1743,
    n1697,
    n1681,
    n32,
    n1565
  );


  xor
  g1740
  (
    n1839,
    n1556,
    n1532,
    n1685,
    n1581
  );


  xnor
  g1741
  (
    n1769,
    n1555,
    n1637,
    n1620,
    n1575
  );


  or
  g1742
  (
    n1777,
    n1725,
    n1570,
    n1724,
    n1630
  );


  and
  g1743
  (
    n1813,
    n1728,
    n1725,
    n1549,
    n1685
  );


  or
  g1744
  (
    n1894,
    n1605,
    n1559,
    n1611,
    n1648
  );


  or
  g1745
  (
    n1844,
    n1537,
    n1532,
    n1678,
    n1732
  );


  xnor
  g1746
  (
    n1756,
    n1712,
    n1693,
    n1719,
    n1603
  );


  nor
  g1747
  (
    n1807,
    n1536,
    n1536,
    n1598,
    n1518
  );


  nor
  g1748
  (
    n1905,
    n1607,
    n1550,
    n1653,
    n1641
  );


  nor
  g1749
  (
    n1848,
    n1652,
    n1608,
    n1654,
    n1730
  );


  xnor
  g1750
  (
    n1763,
    n1723,
    n1692,
    n1524,
    n1531
  );


  nor
  g1751
  (
    n1801,
    n1725,
    n1541,
    n1531,
    n1523
  );


  and
  g1752
  (
    n1752,
    n1567,
    n1568,
    n1607,
    n1594
  );


  nor
  g1753
  (
    n1855,
    n1656,
    n1635,
    n32,
    n1724
  );


  nor
  g1754
  (
    n1827,
    n1591,
    n1564,
    n1538,
    n1610
  );


  xor
  g1755
  (
    n1822,
    n1628,
    n1603,
    n1663,
    n1666
  );


  xnor
  g1756
  (
    n1808,
    n1526,
    n1694,
    n1543,
    n1572
  );


  xnor
  g1757
  (
    n1867,
    n1627,
    n1713,
    n1568,
    n1714
  );


  nor
  g1758
  (
    n1803,
    n1567,
    n1663,
    n1735,
    n1723
  );


  or
  g1759
  (
    n1846,
    n1638,
    n1704,
    n1730,
    n1688
  );


  xor
  g1760
  (
    n1797,
    n1602,
    n1714,
    n1606,
    n1658
  );


  nor
  g1761
  (
    n1791,
    n1717,
    n1674,
    n1542,
    n1654
  );


  and
  g1762
  (
    n1764,
    n1696,
    n1597,
    n1612,
    n1578
  );


  nand
  g1763
  (
    n1890,
    n1540,
    n1710,
    n1675,
    n1706
  );


  nand
  g1764
  (
    n1765,
    n1705,
    n1660,
    n1665,
    n1714
  );


  nand
  g1765
  (
    n1870,
    n1572,
    n1517,
    n1708,
    n1727
  );


  or
  g1766
  (
    n1882,
    n1573,
    n1657,
    n1598,
    n1736
  );


  xor
  g1767
  (
    n1864,
    n1720,
    n1716,
    n1694,
    n1612
  );


  xnor
  g1768
  (
    n1776,
    n1528,
    n1698,
    n1678,
    n1636
  );


  and
  g1769
  (
    n1879,
    n1676,
    n1722,
    n1564,
    n1601
  );


  or
  g1770
  (
    n1815,
    n1668,
    n1712,
    n1559,
    n1673
  );


  xor
  g1771
  (
    n1861,
    n1710,
    n1644,
    n1690,
    n1662
  );


  nand
  g1772
  (
    n1904,
    n1626,
    n1614,
    n1727,
    n1530
  );


  or
  g1773
  (
    n1796,
    n1708,
    n1626,
    n1693,
    n1737
  );


  xor
  g1774
  (
    n1912,
    n1695,
    n1610,
    n1576,
    n1689
  );


  xnor
  g1775
  (
    n1775,
    n1529,
    n1525,
    n1707,
    n1695
  );


  nand
  g1776
  (
    n1881,
    n1700,
    n1561,
    n1680,
    n1706
  );


  nand
  g1777
  (
    n1812,
    n1574,
    n1632,
    n1718,
    n1699
  );


  xor
  g1778
  (
    n1831,
    n1642,
    n1527,
    n1577,
    n1666
  );


  nor
  g1779
  (
    n1913,
    n1736,
    n1692,
    n1647,
    n1726
  );


  or
  g1780
  (
    n1830,
    n1571,
    n1686,
    n1621,
    n1657
  );


  or
  g1781
  (
    n1740,
    n1729,
    n1683,
    n1624,
    n1549
  );


  nor
  g1782
  (
    n1886,
    n1577,
    n1624,
    n1592,
    n1702
  );


  nor
  g1783
  (
    n1853,
    n1557,
    n1608,
    n1738,
    n1577
  );


  nor
  g1784
  (
    n1883,
    n1715,
    n1725,
    n1704,
    n1635
  );


  or
  g1785
  (
    n1850,
    n1631,
    n1679,
    n1644,
    n1524
  );


  nor
  g1786
  (
    n1832,
    n1700,
    n1616,
    n1527,
    n1574
  );


  xor
  g1787
  (
    n1747,
    n1659,
    n1590,
    n1700,
    n1697
  );


  or
  g1788
  (
    n1814,
    n1542,
    n1579,
    n1534,
    n1698
  );


  xor
  g1789
  (
    n1804,
    n1588,
    n1707,
    n1528,
    n1636
  );


  xnor
  g1790
  (
    n1906,
    n1616,
    n1529,
    n1556
  );


  nand
  g1791
  (
    n1860,
    n1569,
    n1614,
    n1588,
    n1736
  );


  or
  g1792
  (
    n1866,
    n1713,
    n1533,
    n1689,
    n1678
  );


  xnor
  g1793
  (
    n1772,
    n1574,
    n1709,
    n1653,
    n1544
  );


  or
  g1794
  (
    n1744,
    n1713,
    n1677,
    n1554,
    n1521
  );


  xor
  g1795
  (
    n1845,
    n1623,
    n1552,
    n1606,
    n1651
  );


  and
  g1796
  (
    n1758,
    n1687,
    n1657,
    n1713,
    n1691
  );


  nor
  g1797
  (
    n1847,
    n1538,
    n1672,
    n1613,
    n1634
  );


  xor
  g1798
  (
    n1739,
    n1664,
    n1666,
    n1630,
    n1615
  );


  nand
  g1799
  (
    n1778,
    n1730,
    n1724,
    n1616,
    n1625
  );


  nand
  g1800
  (
    n1903,
    n1734,
    n1555,
    n1721,
    n1660
  );


  nor
  g1801
  (
    n1900,
    n1570,
    n1605,
    n1677,
    n1696
  );


  and
  g1802
  (
    n1745,
    n1649,
    n1669,
    n1691,
    n1548
  );


  or
  g1803
  (
    n1854,
    n1610,
    n1544,
    n1554,
    n1575
  );


  or
  g1804
  (
    n1781,
    n1676,
    n1591,
    n1692,
    n1629
  );


  xor
  g1805
  (
    n1761,
    n1557,
    n1520,
    n1545,
    n1715
  );


  or
  g1806
  (
    n1857,
    n1609,
    n1672,
    n1661,
    n1716
  );


  nand
  g1807
  (
    n1856,
    n1600,
    n1715,
    n1609,
    n1733
  );


  nor
  g1808
  (
    n1821,
    n1647,
    n1535,
    n1723,
    n1522
  );


  and
  g1809
  (
    n1800,
    n1545,
    n1733,
    n1594,
    n1524
  );


  xor
  g1810
  (
    n1782,
    n1547,
    n1582,
    n1735,
    n1566
  );


  xnor
  g1811
  (
    n1741,
    n1596,
    n1566,
    n1562,
    n1533
  );


  xnor
  g1812
  (
    n1810,
    n1581,
    n1623,
    n1597,
    n1603
  );


  or
  g1813
  (
    n1893,
    n1729,
    n1696,
    n1687,
    n1706
  );


  nor
  g1814
  (
    n1907,
    n1599,
    n1589,
    n1639,
    n1549
  );


  xnor
  g1815
  (
    n1868,
    n1617,
    n1736,
    n1701,
    n1723
  );


  xor
  g1816
  (
    n1794,
    n1622,
    n1582,
    n1729,
    n1633
  );


  xnor
  g1817
  (
    n1767,
    n1589,
    n1674,
    n1622,
    n1716
  );


  and
  g1818
  (
    n1852,
    n1579,
    n1612,
    n1592,
    n1590
  );


  xor
  g1819
  (
    n1836,
    n1738,
    n1558,
    n1586,
    n1673
  );


  or
  g1820
  (
    n1841,
    n1525,
    n1569,
    n1584,
    n1650
  );


  nor
  g1821
  (
    n1859,
    n1632,
    n1665,
    n1563,
    n1734
  );


  xnor
  g1822
  (
    n1887,
    n1535,
    n1548,
    n1546,
    n1718
  );


  or
  g1823
  (
    n1835,
    n1522,
    n1677,
    n1711,
    n1592
  );


  nor
  g1824
  (
    n1759,
    n1519,
    n1722,
    n1737,
    n1633
  );


  xor
  g1825
  (
    n1891,
    n1717,
    n1638,
    n1720,
    n1683
  );


  or
  g1826
  (
    n1783,
    n1611,
    n1588,
    n1694,
    n1731
  );


  or
  g1827
  (
    n1798,
    n1684,
    n1728,
    n1711,
    n1585
  );


  nor
  g1828
  (
    n1834,
    n1695,
    n1683,
    n1601,
    n1593
  );


  nand
  g1829
  (
    n1792,
    n1695,
    n1561,
    n1662,
    n1580
  );


  and
  g1830
  (
    n1820,
    n1682,
    n1696,
    n1618,
    n1681
  );


  xor
  g1831
  (
    n1811,
    n1714,
    n1555,
    n1680,
    n1523
  );


  nand
  g1832
  (
    n1909,
    n1552,
    n1688,
    n1671,
    n1674
  );


  nand
  g1833
  (
    n1901,
    n1595,
    n1554,
    n1641,
    n1655
  );


  or
  g1834
  (
    n1874,
    n1735,
    n1680,
    n1728,
    n1671
  );


  nor
  g1835
  (
    n1757,
    n1569,
    n1544,
    n1703,
    n1599
  );


  and
  g1836
  (
    n1751,
    n1692,
    n1622,
    n1679,
    n1600
  );


  and
  g1837
  (
    n1911,
    n1619,
    n1608,
    n1645,
    n1719
  );


  or
  g1838
  (
    n1809,
    n1540,
    n1701,
    n1566,
    n1625
  );


  xor
  g1839
  (
    n1789,
    n1542,
    n1651,
    n1587,
    n1617
  );


  and
  g1840
  (
    n1754,
    n1703,
    n1716,
    n1663,
    n1546
  );


  xnor
  g1841
  (
    n1871,
    n1613,
    n1719,
    n1731,
    n1518
  );


  xor
  g1842
  (
    n1875,
    n1559,
    n1545,
    n1698,
    n1517
  );


  xor
  g1843
  (
    n1837,
    n1585,
    n1550,
    n1633,
    n1652
  );


  nor
  g1844
  (
    n1748,
    n1551,
    n1587,
    n1580,
    n1526
  );


  xor
  g1845
  (
    n1895,
    n1639,
    n1684,
    n1701,
    n1726
  );


  and
  g1846
  (
    n1858,
    n1721,
    n1609,
    n1553,
    n1707
  );


  nand
  g1847
  (
    n1877,
    n1539,
    n1580,
    n1658,
    n1521
  );


  xor
  g1848
  (
    n1817,
    n1615,
    n1581,
    n1537,
    n1624
  );


  xor
  g1849
  (
    n1843,
    n1615,
    n1703,
    n1686,
    n1584
  );


  nor
  g1850
  (
    n1784,
    n1732,
    n1573,
    n1664,
    n1731
  );


  nor
  g1851
  (
    n1770,
    n1646,
    n1717,
    n1634,
    n1720
  );


  nand
  g1852
  (
    n1805,
    n1623,
    n1619,
    n1653,
    n1596
  );


  xor
  g1853
  (
    n1872,
    n1670,
    n1726,
    n1572
  );


  nor
  g1854
  (
    n1917,
    n1709,
    n1534,
    n1579,
    n1618
  );


  or
  g1855
  (
    n1816,
    n1626,
    n1643,
    n1519,
    n1676
  );


  and
  g1856
  (
    n1755,
    n1586,
    n1587,
    n1712,
    n1557
  );


  nor
  g1857
  (
    n1749,
    n1541,
    n1711,
    n1734
  );


  xor
  g1858
  (
    n1826,
    n1689,
    n1607,
    n1530,
    n1562
  );


  and
  g1859
  (
    n1873,
    n1593,
    n1649,
    n1721,
    n1619
  );


  xnor
  g1860
  (
    n1863,
    n1550,
    n1598,
    n1735,
    n1690
  );


  and
  g1861
  (
    n1869,
    n1640,
    n1589,
    n1669,
    n1664
  );


  xor
  g1862
  (
    n1779,
    n1576,
    n1522,
    n1643,
    n1523
  );


  nor
  g1863
  (
    n1762,
    n1721,
    n1665,
    n1673,
    n1533
  );


  xor
  g1864
  (
    n1806,
    n1532,
    n1646,
    n1561,
    n1539
  );


  and
  g1865
  (
    n1799,
    n1670,
    n1730,
    n1649,
    n1705
  );


  nand
  g1866
  (
    n1788,
    n1709,
    n1675,
    n1682,
    n1618
  );


  xor
  g1867
  (
    n1898,
    n1620,
    n1690,
    n1650,
    n1548
  );


  or
  g1868
  (
    n1742,
    n1693,
    n1647,
    n1527,
    n1620
  );


  xnor
  g1869
  (
    n1880,
    n1520,
    n1526,
    n1568,
    n1637
  );


  nor
  g1870
  (
    n1787,
    n1645,
    n1702,
    n1724,
    n1682
  );


  and
  g1871
  (
    n1771,
    n1697,
    n1667,
    n1684,
    n1659
  );


  and
  g1872
  (
    n1851,
    n1640,
    n1590,
    n1661,
    n1687
  );


  nor
  g1873
  (
    n1842,
    n1538,
    n1699,
    n1686,
    n1691
  );


  xnor
  g1874
  (
    n1785,
    n1599,
    n1709,
    n1571,
    n1520
  );


  nor
  g1875
  (
    n1892,
    n1537,
    n1604,
    n1688,
    n1668
  );


  and
  g1876
  (
    KeyWire_0_27,
    n1701,
    n1650,
    n1594,
    n1668
  );


  xnor
  g1877
  (
    n1916,
    n1669,
    n1702,
    n1539,
    n1601
  );


  and
  g1878
  (
    n1865,
    n1687,
    n1519,
    n1564,
    n1679
  );


  nor
  g1879
  (
    n1828,
    n1558,
    n1651,
    n1528,
    n1525
  );


  nand
  g1880
  (
    n1818,
    n1660,
    n1600,
    n1670,
    n1693
  );


  xnor
  g1881
  (
    n1802,
    n1659,
    n1722,
    n1731,
    n1667
  );


  xnor
  g1882
  (
    n1862,
    n1530,
    n1697,
    n1672,
    n1562
  );


  xor
  g1883
  (
    n1915,
    n1688,
    n1715,
    n1621,
    n1705
  );


  xnor
  g1884
  (
    n1897,
    n1652,
    n1661,
    n1627,
    n1570
  );


  xnor
  g1885
  (
    n1899,
    n1708,
    n1694,
    n1720,
    n1631
  );


  or
  g1886
  (
    n1944,
    n1910,
    n1905,
    n1764,
    n1867
  );


  nor
  g1887
  (
    n1996,
    n1879,
    n1760,
    n1765,
    n1873
  );


  xnor
  g1888
  (
    n1927,
    n1841,
    n1844,
    n1776,
    n1751
  );


  or
  g1889
  (
    n2007,
    n1845,
    n1758,
    n1849,
    n1848
  );


  nor
  g1890
  (
    n1984,
    n1771,
    n1854,
    n1813,
    n1892
  );


  or
  g1891
  (
    n1985,
    n1818,
    n1915,
    n1865,
    n1741
  );


  xnor
  g1892
  (
    n1951,
    n1828,
    n1861,
    n1888,
    n1791
  );


  xor
  g1893
  (
    n1991,
    n1741,
    n1846,
    n1797,
    n1871
  );


  nand
  g1894
  (
    n1987,
    n1861,
    n1800,
    n1899,
    n1804
  );


  xor
  g1895
  (
    n1940,
    n1868,
    n1880,
    n1883,
    n1850
  );


  nand
  g1896
  (
    n1989,
    n1864,
    n1756,
    n1793,
    n1832
  );


  nand
  g1897
  (
    n1925,
    n1754,
    n1896,
    n1799,
    n1916
  );


  nor
  g1898
  (
    n1950,
    n1858,
    n1773,
    n1868,
    n1916
  );


  nand
  g1899
  (
    n1986,
    n1876,
    n1775,
    n1766,
    n1902
  );


  nor
  g1900
  (
    n1935,
    n1742,
    n1763,
    n1852,
    n1847
  );


  nor
  g1901
  (
    n1941,
    n1837,
    n1830,
    n1866,
    n1807
  );


  nor
  g1902
  (
    n2009,
    n1886,
    n1779,
    n1794,
    n1859
  );


  and
  g1903
  (
    n1963,
    n1823,
    n1914,
    n1905,
    n1878
  );


  and
  g1904
  (
    n1966,
    n1752,
    n1766,
    n1789,
    n1888
  );


  and
  g1905
  (
    n1946,
    n1812,
    n1761,
    n1904,
    n1906
  );


  nor
  g1906
  (
    n1938,
    n1854,
    n1821,
    n1827,
    n1885
  );


  xor
  g1907
  (
    n1921,
    n1910,
    n1756,
    n1767,
    n1798
  );


  and
  g1908
  (
    n1945,
    n1839,
    n1829,
    n1915,
    n1739
  );


  and
  g1909
  (
    n1932,
    n1802,
    n1743,
    n1799,
    n1820
  );


  nand
  g1910
  (
    n1976,
    n1884,
    n1911,
    n1909,
    n1897
  );


  and
  g1911
  (
    n1937,
    n1805,
    n1836,
    n1893,
    n1807
  );


  and
  g1912
  (
    n1952,
    n1809,
    n1844,
    n1862,
    n1832
  );


  and
  g1913
  (
    n2004,
    n1740,
    n1872,
    n1790,
    n1900
  );


  and
  g1914
  (
    n1919,
    n1787,
    n1822,
    n1745,
    n1917
  );


  xor
  g1915
  (
    n1942,
    n1853,
    n1803,
    n1810,
    n1891
  );


  nor
  g1916
  (
    n2008,
    n1863,
    n1780,
    n1826,
    n1753
  );


  nor
  g1917
  (
    n1965,
    n1852,
    n1745,
    n1814,
    n1819
  );


  xnor
  g1918
  (
    n2000,
    n1770,
    n1901,
    n1902,
    n1914
  );


  xnor
  g1919
  (
    n1920,
    n1869,
    n1906,
    n1863,
    n1774
  );


  xor
  g1920
  (
    n1956,
    n1813,
    n1793,
    n1739,
    n1758
  );


  and
  g1921
  (
    n1968,
    n1816,
    n1893,
    n1903,
    n1878
  );


  or
  g1922
  (
    n1982,
    n1841,
    n1786,
    n1797,
    n1772
  );


  xnor
  g1923
  (
    n1936,
    n1817,
    n1743,
    n1894,
    n1840
  );


  nand
  g1924
  (
    n1978,
    n1783,
    n1875,
    n1819,
    n1749
  );


  nand
  g1925
  (
    n1961,
    n666,
    n1855,
    n1846,
    n1777
  );


  and
  g1926
  (
    n1949,
    n1779,
    n1877,
    n1757,
    n1912
  );


  and
  g1927
  (
    n1933,
    n1847,
    n1887,
    n1808,
    n1907
  );


  xor
  g1928
  (
    n2006,
    n1763,
    n1864,
    n1865,
    n1907
  );


  xnor
  g1929
  (
    n2001,
    n1757,
    n1781,
    n1909,
    n1785
  );


  xor
  g1930
  (
    n2005,
    n1761,
    n1857,
    n1897,
    n1856
  );


  or
  g1931
  (
    n1964,
    n1746,
    n1747,
    n1778,
    n1900
  );


  xnor
  g1932
  (
    n2003,
    n1826,
    n1838,
    n1801,
    n1744
  );


  xnor
  g1933
  (
    n1929,
    n1825,
    n1804,
    n1859,
    n1881
  );


  nand
  g1934
  (
    n2002,
    n1843,
    n1855,
    n1784,
    n1874
  );


  xor
  g1935
  (
    n1995,
    n1769,
    n1814,
    n1751,
    n1795
  );


  or
  g1936
  (
    n1947,
    n1913,
    n1898,
    n1834,
    n1838
  );


  xnor
  g1937
  (
    n1962,
    n1875,
    n1824,
    n1802,
    n1781
  );


  xnor
  g1938
  (
    n1924,
    n1809,
    n1783,
    n1890,
    n1885
  );


  xor
  g1939
  (
    n1977,
    n1744,
    n1768,
    n1774,
    n1831
  );


  nand
  g1940
  (
    n1975,
    n1790,
    n1773,
    n1842,
    n1778
  );


  and
  g1941
  (
    n1969,
    n1874,
    n1901,
    n1886,
    n1908
  );


  xnor
  g1942
  (
    n1988,
    n1917,
    n1803,
    n1835,
    n1780
  );


  xor
  g1943
  (
    n1922,
    n1828,
    n1831,
    n1858,
    n1871
  );


  or
  g1944
  (
    n1958,
    n1750,
    n1752,
    n1851,
    n1908
  );


  nand
  g1945
  (
    n1979,
    n1795,
    n1918,
    n1788,
    n1823
  );


  nor
  g1946
  (
    n1960,
    n1764,
    n1880,
    n1800,
    n1881
  );


  and
  g1947
  (
    n1954,
    n1777,
    n1873,
    n1860,
    n1866
  );


  xor
  g1948
  (
    n1973,
    n1782,
    n1827,
    n1850,
    n1869
  );


  xnor
  g1949
  (
    n1994,
    n1747,
    n1839,
    n1788,
    n1768
  );


  nand
  g1950
  (
    n1980,
    n1887,
    n1815,
    n1753,
    n1785
  );


  nand
  g1951
  (
    n1993,
    n1833,
    n1767,
    n1771,
    n1749
  );


  or
  g1952
  (
    n1970,
    n1830,
    n1811,
    n1889,
    n1876
  );


  and
  g1953
  (
    n1971,
    n1842,
    n1834,
    n1759,
    n1870
  );


  or
  g1954
  (
    n1930,
    n1884,
    n1818,
    n1862,
    n1824
  );


  xnor
  g1955
  (
    n1926,
    n1765,
    n1810,
    n1792,
    n1740
  );


  nor
  g1956
  (
    n1934,
    n1817,
    n1829,
    n1913,
    n1746
  );


  xnor
  g1957
  (
    n1939,
    n1755,
    n1860,
    n1835,
    n1801
  );


  xor
  g1958
  (
    n1931,
    n1879,
    n1848,
    n1892,
    n1796
  );


  xnor
  g1959
  (
    n1997,
    n1849,
    n1918,
    n1891,
    n1883
  );


  and
  g1960
  (
    n1923,
    n1833,
    n1769,
    n1816,
    n1845
  );


  and
  g1961
  (
    n1953,
    n1775,
    n1811,
    n1895,
    n666
  );


  nor
  g1962
  (
    n1957,
    n1748,
    n1843,
    n1898,
    n1770
  );


  and
  g1963
  (
    n1998,
    n1853,
    n1890,
    n1872,
    n1812
  );


  nor
  g1964
  (
    n1983,
    n1762,
    n1856,
    n1760,
    n1857
  );


  nand
  g1965
  (
    n1972,
    n1754,
    n1784,
    n1911,
    n1755
  );


  or
  g1966
  (
    n1928,
    n1808,
    n1806,
    n1748,
    n1805
  );


  nor
  g1967
  (
    n1992,
    n1867,
    n1792,
    n1759,
    n1750
  );


  or
  g1968
  (
    n1999,
    n1742,
    n1787,
    n1762,
    n1882
  );


  xnor
  g1969
  (
    n1955,
    n1821,
    n1786,
    n1904,
    n1820
  );


  and
  g1970
  (
    n1990,
    n1806,
    n1851,
    n1776,
    n1895
  );


  xnor
  g1971
  (
    n1974,
    n1896,
    n1889,
    n1772,
    n1840
  );


  xor
  g1972
  (
    n1981,
    n1789,
    n1825,
    n1738,
    n1794
  );


  xor
  g1973
  (
    n1967,
    n1837,
    n1877,
    n1870,
    n1882
  );


  nor
  g1974
  (
    n1943,
    n1822,
    n1815,
    n32,
    n1836
  );


  xor
  g1975
  (
    n1959,
    n1796,
    n1791,
    n1912,
    n1903
  );


  nand
  g1976
  (
    n1948,
    n1782,
    n1894,
    n1798,
    n1899
  );


  and
  g1977
  (
    n2026,
    n1980,
    n1952,
    n1919,
    n1935
  );


  or
  g1978
  (
    n2013,
    n1928,
    n1925,
    n1953,
    n1978
  );


  nand
  g1979
  (
    n2018,
    n1943,
    n1934,
    n1964,
    n1926
  );


  nor
  g1980
  (
    n2023,
    n1997,
    n1955,
    n1962,
    n1960
  );


  and
  g1981
  (
    n2011,
    n1981,
    n1940,
    n1987,
    n1992
  );


  xor
  g1982
  (
    n2010,
    n1929,
    n1963,
    n1923,
    n1979
  );


  xnor
  g1983
  (
    n2028,
    n1947,
    n1946,
    n1973,
    n1969
  );


  and
  g1984
  (
    n2022,
    n1939,
    n2001,
    n1933,
    n1937
  );


  or
  g1985
  (
    n2014,
    n1949,
    n2000,
    n1983,
    n2008
  );


  xor
  g1986
  (
    n2030,
    n1971,
    n2007,
    n1936,
    n1927
  );


  or
  g1987
  (
    n2025,
    n1985,
    n1958,
    n1938,
    n1988
  );


  nor
  g1988
  (
    n2015,
    n1991,
    n1944,
    n1999,
    n1990
  );


  xnor
  g1989
  (
    n2031,
    n1976,
    n1970,
    n2002,
    n1994
  );


  and
  g1990
  (
    n2024,
    n1957,
    n1948,
    n1945,
    n1982
  );


  and
  g1991
  (
    n2027,
    n1975,
    n1922,
    n1993,
    n1942
  );


  and
  g1992
  (
    n2029,
    n1950,
    n1959,
    n1967,
    n1968
  );


  nor
  g1993
  (
    n2021,
    n1954,
    n1921,
    n1965,
    n2003
  );


  xnor
  g1994
  (
    n2017,
    n1986,
    n1966,
    n1931,
    n1972
  );


  nand
  g1995
  (
    n2032,
    n1977,
    n1974,
    n1998,
    n1995
  );


  and
  g1996
  (
    n2019,
    n1930,
    n1984,
    n1932,
    n1956
  );


  xor
  g1997
  (
    n2016,
    n1989,
    n2009,
    n1961,
    n1996
  );


  nor
  g1998
  (
    n2020,
    n1941,
    n2009,
    n1920,
    n1951
  );


  or
  g1999
  (
    n2012,
    n2006,
    n2005,
    n2004,
    n1924
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1384,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n669,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n118,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n382,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n348,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1014,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1027,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1237,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1286,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n653,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n1617,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1191,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n41,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1390,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n457,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1434,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n1335,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n796,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1044,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n526,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1066,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n922,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n36,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n222,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n1288,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n1723,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n877,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1823,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n235,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1720,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n1351,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1247,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

