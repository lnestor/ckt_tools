

module Stat_221_421
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n231,
  n212,
  n208,
  n238,
  n207,
  n226,
  n218,
  n214,
  n220,
  n227,
  n234,
  n235,
  n228,
  n222,
  n223,
  n209,
  n230,
  n224,
  n221,
  n210,
  n233,
  n216,
  n219,
  n237,
  n236,
  n232,
  n217,
  n213,
  n229,
  n215,
  n211,
  n225
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n231;output n212;output n208;output n238;output n207;output n226;output n218;output n214;output n220;output n227;output n234;output n235;output n228;output n222;output n223;output n209;output n230;output n224;output n221;output n210;output n233;output n216;output n219;output n237;output n236;output n232;output n217;output n213;output n229;output n215;output n211;output n225;
  wire n18;wire n19;wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n28,
    n2
  );


  buf
  g1
  (
    n18,
    n3
  );


  not
  g2
  (
    n26,
    n3
  );


  not
  g3
  (
    n32,
    n1
  );


  buf
  g4
  (
    n22,
    n5
  );


  buf
  g5
  (
    n30,
    n1
  );


  buf
  g6
  (
    n23,
    n3
  );


  not
  g7
  (
    KeyWire_0_9,
    n5
  );


  buf
  g8
  (
    n19,
    n2
  );


  not
  g9
  (
    n21,
    n5
  );


  not
  g10
  (
    n20,
    n1
  );


  buf
  g11
  (
    n29,
    n4
  );


  buf
  g12
  (
    KeyWire_0_1,
    n2
  );


  buf
  g13
  (
    n27,
    n4
  );


  not
  g14
  (
    n24,
    n4
  );


  buf
  g15
  (
    n78,
    n23
  );


  not
  g16
  (
    n58,
    n21
  );


  not
  g17
  (
    n53,
    n22
  );


  not
  g18
  (
    n62,
    n32
  );


  not
  g19
  (
    KeyWire_0_22,
    n22
  );


  buf
  g20
  (
    n59,
    n24
  );


  buf
  g21
  (
    n48,
    n21
  );


  buf
  g22
  (
    n61,
    n20
  );


  not
  g23
  (
    n67,
    n26
  );


  not
  g24
  (
    n65,
    n18
  );


  not
  g25
  (
    n52,
    n30
  );


  buf
  g26
  (
    KeyWire_0_6,
    n32
  );


  not
  g27
  (
    n73,
    n28
  );


  not
  g28
  (
    n40,
    n31
  );


  not
  g29
  (
    n50,
    n20
  );


  buf
  g30
  (
    n43,
    n23
  );


  not
  g31
  (
    n44,
    n19
  );


  not
  g32
  (
    n34,
    n18
  );


  buf
  g33
  (
    n37,
    n29
  );


  buf
  g34
  (
    n42,
    n25
  );


  not
  g35
  (
    KeyWire_0_2,
    n28
  );


  not
  g36
  (
    n70,
    n18
  );


  not
  g37
  (
    n41,
    n27
  );


  not
  g38
  (
    n47,
    n29
  );


  not
  g39
  (
    KeyWire_0_29,
    n24
  );


  buf
  g40
  (
    n55,
    n30
  );


  not
  g41
  (
    n68,
    n22
  );


  buf
  g42
  (
    n38,
    n20
  );


  buf
  g43
  (
    n64,
    n28
  );


  buf
  g44
  (
    n72,
    n24
  );


  not
  g45
  (
    n33,
    n27
  );


  buf
  g46
  (
    n39,
    n26
  );


  buf
  g47
  (
    n51,
    n19
  );


  buf
  g48
  (
    n54,
    n30
  );


  not
  g49
  (
    n63,
    n26
  );


  not
  g50
  (
    n45,
    n21
  );


  buf
  g51
  (
    n60,
    n27
  );


  buf
  g52
  (
    n75,
    n32
  );


  buf
  g53
  (
    n36,
    n19
  );


  buf
  g54
  (
    n71,
    n25
  );


  buf
  g55
  (
    KeyWire_0_8,
    n31
  );


  buf
  g56
  (
    KeyWire_0_30,
    n23
  );


  not
  g57
  (
    n66,
    n32
  );


  not
  g58
  (
    KeyWire_0_0,
    n29
  );


  not
  g59
  (
    n76,
    n31
  );


  buf
  g60
  (
    n56,
    n25
  );


  buf
  g61
  (
    n174,
    n33
  );


  buf
  g62
  (
    n101,
    n60
  );


  not
  g63
  (
    n94,
    n45
  );


  buf
  g64
  (
    KeyWire_0_26,
    n77
  );


  buf
  g65
  (
    n104,
    n48
  );


  not
  g66
  (
    n155,
    n52
  );


  not
  g67
  (
    n201,
    n9
  );


  buf
  g68
  (
    n143,
    n76
  );


  not
  g69
  (
    n91,
    n71
  );


  buf
  g70
  (
    n165,
    n34
  );


  buf
  g71
  (
    KeyWire_0_20,
    n35
  );


  not
  g72
  (
    n199,
    n65
  );


  not
  g73
  (
    n106,
    n77
  );


  not
  g74
  (
    KeyWire_0_16,
    n57
  );


  buf
  g75
  (
    n176,
    n53
  );


  buf
  g76
  (
    n178,
    n75
  );


  not
  g77
  (
    n108,
    n17
  );


  not
  g78
  (
    n141,
    n59
  );


  buf
  g79
  (
    n150,
    n45
  );


  not
  g80
  (
    KeyWire_0_3,
    n41
  );


  buf
  g81
  (
    n203,
    n77
  );


  not
  g82
  (
    n128,
    n69
  );


  not
  g83
  (
    KeyWire_0_28,
    n39
  );


  not
  g84
  (
    n102,
    n67
  );


  buf
  g85
  (
    n156,
    n46
  );


  buf
  g86
  (
    n139,
    n41
  );


  buf
  g87
  (
    n205,
    n78
  );


  buf
  g88
  (
    n132,
    n47
  );


  not
  g89
  (
    n127,
    n50
  );


  not
  g90
  (
    n133,
    n61
  );


  buf
  g91
  (
    n197,
    n60
  );


  buf
  g92
  (
    n84,
    n69
  );


  not
  g93
  (
    n136,
    n78
  );


  buf
  g94
  (
    n80,
    n65
  );


  buf
  g95
  (
    n125,
    n38
  );


  not
  g96
  (
    n182,
    n14
  );


  buf
  g97
  (
    n81,
    n41
  );


  buf
  g98
  (
    KeyWire_0_21,
    n7
  );


  buf
  g99
  (
    n123,
    n66
  );


  not
  g100
  (
    n160,
    n14
  );


  buf
  g101
  (
    n87,
    n65
  );


  buf
  g102
  (
    n118,
    n55
  );


  buf
  g103
  (
    n138,
    n36
  );


  not
  g104
  (
    n170,
    n8
  );


  not
  g105
  (
    n154,
    n72
  );


  not
  g106
  (
    n188,
    n70
  );


  not
  g107
  (
    n145,
    n54
  );


  buf
  g108
  (
    KeyWire_0_14,
    n44
  );


  not
  g109
  (
    n130,
    n76
  );


  buf
  g110
  (
    n206,
    n73
  );


  buf
  g111
  (
    n149,
    n52
  );


  buf
  g112
  (
    n90,
    n35
  );


  not
  g113
  (
    KeyWire_0_17,
    n42
  );


  not
  g114
  (
    n192,
    n8
  );


  not
  g115
  (
    n111,
    n74
  );


  buf
  g116
  (
    n117,
    n74
  );


  buf
  g117
  (
    n129,
    n7
  );


  not
  g118
  (
    n202,
    n15
  );


  not
  g119
  (
    n166,
    n49
  );


  buf
  g120
  (
    n114,
    n6
  );


  buf
  g121
  (
    KeyWire_0_27,
    n47
  );


  not
  g122
  (
    n142,
    n59
  );


  not
  g123
  (
    n96,
    n33
  );


  buf
  g124
  (
    n147,
    n15
  );


  buf
  g125
  (
    n157,
    n53
  );


  not
  g126
  (
    KeyWire_0_7,
    n34
  );


  buf
  g127
  (
    n151,
    n58
  );


  not
  g128
  (
    n183,
    n10
  );


  not
  g129
  (
    KeyWire_0_10,
    n66
  );


  buf
  g130
  (
    n169,
    n64
  );


  buf
  g131
  (
    KeyWire_0_23,
    n45
  );


  not
  g132
  (
    n92,
    n73
  );


  not
  g133
  (
    n109,
    n40
  );


  not
  g134
  (
    n93,
    n59
  );


  buf
  g135
  (
    n85,
    n9
  );


  buf
  g136
  (
    n131,
    n74
  );


  not
  g137
  (
    n122,
    n71
  );


  not
  g138
  (
    n163,
    n51
  );


  buf
  g139
  (
    n88,
    n62
  );


  not
  g140
  (
    n82,
    n43
  );


  buf
  g141
  (
    n146,
    n75
  );


  buf
  g142
  (
    n193,
    n40
  );


  buf
  g143
  (
    n158,
    n37
  );


  not
  g144
  (
    KeyWire_0_5,
    n50
  );


  buf
  g145
  (
    n100,
    n49
  );


  not
  g146
  (
    n140,
    n71
  );


  buf
  g147
  (
    n110,
    n49
  );


  buf
  g148
  (
    n186,
    n38
  );


  buf
  g149
  (
    n191,
    n57
  );


  not
  g150
  (
    n119,
    n43
  );


  not
  g151
  (
    n198,
    n37
  );


  not
  g152
  (
    n194,
    n37
  );


  not
  g153
  (
    n180,
    n46
  );


  buf
  g154
  (
    n162,
    n48
  );


  buf
  g155
  (
    n83,
    n48
  );


  not
  g156
  (
    n148,
    n66
  );


  buf
  g157
  (
    n195,
    n13
  );


  not
  g158
  (
    n95,
    n54
  );


  not
  g159
  (
    n204,
    n10
  );


  buf
  g160
  (
    n86,
    n14
  );


  buf
  g161
  (
    KeyWire_0_18,
    n75
  );


  buf
  g162
  (
    KeyWire_0_19,
    n55
  );


  not
  g163
  (
    KeyWire_0_31,
    n39
  );


  buf
  g164
  (
    n200,
    n35
  );


  buf
  g165
  (
    n168,
    n73
  );


  not
  g166
  (
    KeyWire_0_15,
    n34
  );


  not
  g167
  (
    n190,
    n53
  );


  buf
  g168
  (
    n171,
    n72
  );


  not
  g169
  (
    n115,
    n68
  );


  not
  g170
  (
    n79,
    n61
  );


  buf
  g171
  (
    KeyWire_0_13,
    n15
  );


  not
  g172
  (
    n153,
    n33
  );


  nor
  g173
  (
    n144,
    n16,
    n17
  );


  xor
  g174
  (
    n105,
    n57,
    n6,
    n38,
    n36
  );


  or
  g175
  (
    n164,
    n70,
    n56,
    n11,
    n50
  );


  xor
  g176
  (
    n107,
    n70,
    n9,
    n12,
    n56
  );


  and
  g177
  (
    KeyWire_0_11,
    n17,
    n55,
    n68,
    n46
  );


  nand
  g178
  (
    n179,
    n10,
    n78,
    n6,
    n16
  );


  nand
  g179
  (
    n116,
    n13,
    n44,
    n64,
    n42
  );


  and
  g180
  (
    n121,
    n7,
    n51,
    n64,
    n72
  );


  and
  g181
  (
    n184,
    n39,
    n44,
    n8,
    n47
  );


  and
  g182
  (
    n159,
    n68,
    n67,
    n54,
    n61
  );


  xor
  g183
  (
    n173,
    n60,
    n16,
    n58,
    n52
  );


  xor
  g184
  (
    n167,
    n76,
    n12,
    n63,
    n67
  );


  or
  g185
  (
    n134,
    n62,
    n63,
    n69
  );


  xor
  g186
  (
    n113,
    n56,
    n36,
    n12,
    n51
  );


  nor
  g187
  (
    n135,
    n43,
    n11,
    n62,
    n58
  );


  xnor
  g188
  (
    n89,
    n13,
    n40,
    n11,
    n42
  );


  xnor
  g189
  (
    n220,
    n121,
    n135,
    n101,
    n184
  );


  and
  g190
  (
    n222,
    n204,
    n199,
    n196,
    n119
  );


  nand
  g191
  (
    n213,
    n87,
    n126,
    n206,
    n194
  );


  or
  g192
  (
    n208,
    n139,
    n120,
    n92,
    n183
  );


  and
  g193
  (
    n219,
    n154,
    n198,
    n202,
    n163
  );


  and
  g194
  (
    n232,
    n109,
    n107,
    n96,
    n146
  );


  and
  g195
  (
    n225,
    n178,
    n158,
    n160,
    n102
  );


  xnor
  g196
  (
    n227,
    n179,
    n157,
    n145,
    n192
  );


  nand
  g197
  (
    n210,
    n83,
    n85,
    n193,
    n190
  );


  and
  g198
  (
    n218,
    n86,
    n182,
    n156,
    n148
  );


  xnor
  g199
  (
    n231,
    n99,
    n162,
    n128,
    n147
  );


  xor
  g200
  (
    n214,
    n169,
    n116,
    n88,
    n165
  );


  and
  g201
  (
    n224,
    n98,
    n79,
    n123,
    n143
  );


  and
  g202
  (
    n238,
    n104,
    n134,
    n132,
    n108
  );


  nand
  g203
  (
    n237,
    n136,
    n131,
    n176,
    n172
  );


  or
  g204
  (
    n223,
    n170,
    n175,
    n106,
    n140
  );


  or
  g205
  (
    n216,
    n186,
    n166,
    n168,
    n82
  );


  and
  g206
  (
    n209,
    n110,
    n94,
    n173,
    n124
  );


  and
  g207
  (
    n211,
    n115,
    n138,
    n153,
    n149
  );


  and
  g208
  (
    n215,
    n195,
    n111,
    n137,
    n100
  );


  nand
  g209
  (
    n229,
    n129,
    n197,
    n114,
    n95
  );


  xnor
  g210
  (
    n234,
    n151,
    n122,
    n91,
    n81
  );


  nand
  g211
  (
    n212,
    n167,
    n150,
    n185,
    n171
  );


  xnor
  g212
  (
    KeyWire_0_4,
    n187,
    n103,
    n152,
    n203
  );


  and
  g213
  (
    n235,
    n177,
    n105,
    n181,
    n113
  );


  and
  g214
  (
    KeyWire_0_24,
    n84,
    n130,
    n191,
    n141
  );


  and
  g215
  (
    KeyWire_0_12,
    n188,
    n161,
    n200,
    n180
  );


  or
  g216
  (
    n236,
    n144,
    n89,
    n118,
    n142
  );


  xnor
  g217
  (
    n226,
    n112,
    n125,
    n97,
    n164
  );


  nor
  g218
  (
    KeyWire_0_25,
    n90,
    n127,
    n189,
    n93
  );


  xor
  g219
  (
    n207,
    n159,
    n117,
    n80,
    n174
  );


  and
  g220
  (
    n228,
    n201,
    n133,
    n155,
    n205
  );


  xor
  KeyGate_0_0
  (
    n46,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n31,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n74,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n124,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n217,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n152,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n57,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n97,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n77,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n25,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n185,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n103,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n230,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n177,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n137,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n172,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n98,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n120,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n189,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n175,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n99,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n112,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n69,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n161,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n221,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n233,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n181,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n126,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n196,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n49,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n35,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n187,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


