

module Stat_1399_20_5
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n1392,
  n1401,
  n1373,
  n1375,
  n1359,
  n1376,
  n1353,
  n1391,
  n1403,
  n1363,
  n1367,
  n1366,
  n1381,
  n1397,
  n1380,
  n1386,
  n1371,
  n1354,
  n1378,
  n1384,
  n1358,
  n1356,
  n1393,
  n1398,
  n1355,
  n1370,
  n1389,
  n1421,
  n1419,
  n1418,
  n1420
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1392;output n1401;output n1373;output n1375;output n1359;output n1376;output n1353;output n1391;output n1403;output n1363;output n1367;output n1366;output n1381;output n1397;output n1380;output n1386;output n1371;output n1354;output n1378;output n1384;output n1358;output n1356;output n1393;output n1398;output n1355;output n1370;output n1389;output n1421;output n1419;output n1418;output n1420;
  wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1357;wire n1360;wire n1361;wire n1362;wire n1364;wire n1365;wire n1368;wire n1369;wire n1372;wire n1374;wire n1377;wire n1379;wire n1382;wire n1383;wire n1385;wire n1387;wire n1388;wire n1390;wire n1394;wire n1395;wire n1396;wire n1399;wire n1400;wire n1402;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n103,
    n18
  );


  buf
  g1
  (
    n87,
    n10
  );


  not
  g2
  (
    n31,
    n2
  );


  buf
  g3
  (
    n42,
    n21
  );


  not
  g4
  (
    n78,
    n18
  );


  buf
  g5
  (
    n67,
    n19
  );


  not
  g6
  (
    n106,
    n13
  );


  not
  g7
  (
    n40,
    n11
  );


  buf
  g8
  (
    KeyWire_0_28,
    n5
  );


  not
  g9
  (
    n58,
    n19
  );


  not
  g10
  (
    n37,
    n20
  );


  not
  g11
  (
    n39,
    n5
  );


  buf
  g12
  (
    n55,
    n4
  );


  buf
  g13
  (
    n36,
    n21
  );


  not
  g14
  (
    n47,
    n22
  );


  not
  g15
  (
    n64,
    n10
  );


  buf
  g16
  (
    n80,
    n9
  );


  not
  g17
  (
    n28,
    n20
  );


  not
  g18
  (
    n29,
    n18
  );


  not
  g19
  (
    n49,
    n6
  );


  not
  g20
  (
    n91,
    n19
  );


  buf
  g21
  (
    n104,
    n3
  );


  buf
  g22
  (
    n34,
    n13
  );


  buf
  g23
  (
    n92,
    n12
  );


  not
  g24
  (
    n60,
    n16
  );


  not
  g25
  (
    n25,
    n13
  );


  not
  g26
  (
    n23,
    n6
  );


  buf
  g27
  (
    n102,
    n19
  );


  buf
  g28
  (
    n56,
    n22
  );


  not
  g29
  (
    n35,
    n2
  );


  not
  g30
  (
    n54,
    n14
  );


  buf
  g31
  (
    n43,
    n10
  );


  not
  g32
  (
    n46,
    n4
  );


  not
  g33
  (
    n66,
    n15
  );


  buf
  g34
  (
    n33,
    n12
  );


  buf
  g35
  (
    n27,
    n12
  );


  not
  g36
  (
    n89,
    n8
  );


  not
  g37
  (
    n68,
    n12
  );


  buf
  g38
  (
    n65,
    n21
  );


  not
  g39
  (
    n96,
    n17
  );


  buf
  g40
  (
    n41,
    n17
  );


  buf
  g41
  (
    n83,
    n9
  );


  buf
  g42
  (
    n107,
    n13
  );


  buf
  g43
  (
    n71,
    n22
  );


  not
  g44
  (
    n52,
    n1
  );


  buf
  g45
  (
    n82,
    n11
  );


  buf
  g46
  (
    n94,
    n9
  );


  buf
  g47
  (
    n85,
    n8
  );


  not
  g48
  (
    n98,
    n8
  );


  not
  g49
  (
    n30,
    n10
  );


  not
  g50
  (
    n53,
    n2
  );


  buf
  g51
  (
    n70,
    n7
  );


  not
  g52
  (
    n63,
    n3
  );


  buf
  g53
  (
    n61,
    n3
  );


  not
  g54
  (
    n38,
    n6
  );


  not
  g55
  (
    n77,
    n7
  );


  buf
  g56
  (
    n74,
    n5
  );


  buf
  g57
  (
    n24,
    n5
  );


  not
  g58
  (
    n44,
    n17
  );


  buf
  g59
  (
    n101,
    n22
  );


  buf
  g60
  (
    n73,
    n6
  );


  not
  g61
  (
    n100,
    n15
  );


  not
  g62
  (
    n26,
    n14
  );


  not
  g63
  (
    n57,
    n2
  );


  buf
  g64
  (
    n97,
    n7
  );


  not
  g65
  (
    n79,
    n7
  );


  not
  g66
  (
    n48,
    n14
  );


  buf
  g67
  (
    n32,
    n15
  );


  buf
  g68
  (
    n76,
    n15
  );


  buf
  g69
  (
    n105,
    n17
  );


  buf
  g70
  (
    n69,
    n8
  );


  not
  g71
  (
    n45,
    n16
  );


  buf
  g72
  (
    n93,
    n21
  );


  buf
  g73
  (
    n84,
    n11
  );


  buf
  g74
  (
    n81,
    n20
  );


  not
  g75
  (
    n72,
    n18
  );


  buf
  g76
  (
    n51,
    n9
  );


  buf
  g77
  (
    n59,
    n16
  );


  not
  g78
  (
    n88,
    n16
  );


  buf
  g79
  (
    n99,
    n20
  );


  not
  g80
  (
    n62,
    n4
  );


  buf
  g81
  (
    n90,
    n11
  );


  not
  g82
  (
    n86,
    n3
  );


  not
  g83
  (
    n95,
    n4
  );


  buf
  g84
  (
    n75,
    n14
  );


  not
  g85
  (
    n285,
    n81
  );


  buf
  g86
  (
    n182,
    n93
  );


  buf
  g87
  (
    n208,
    n107
  );


  not
  g88
  (
    n232,
    n23
  );


  buf
  g89
  (
    n345,
    n70
  );


  buf
  g90
  (
    n197,
    n61
  );


  buf
  g91
  (
    n164,
    n74
  );


  buf
  g92
  (
    n184,
    n86
  );


  buf
  g93
  (
    n429,
    n74
  );


  buf
  g94
  (
    n262,
    n56
  );


  not
  g95
  (
    n322,
    n94
  );


  not
  g96
  (
    n296,
    n72
  );


  buf
  g97
  (
    n223,
    n45
  );


  not
  g98
  (
    n123,
    n87
  );


  buf
  g99
  (
    n245,
    n105
  );


  buf
  g100
  (
    n313,
    n39
  );


  buf
  g101
  (
    n238,
    n24
  );


  not
  g102
  (
    n174,
    n28
  );


  buf
  g103
  (
    n441,
    n35
  );


  buf
  g104
  (
    n240,
    n78
  );


  not
  g105
  (
    n196,
    n84
  );


  not
  g106
  (
    n124,
    n37
  );


  not
  g107
  (
    KeyWire_0_19,
    n23
  );


  buf
  g108
  (
    n403,
    n41
  );


  buf
  g109
  (
    n374,
    n66
  );


  buf
  g110
  (
    n417,
    n41
  );


  not
  g111
  (
    n171,
    n100
  );


  not
  g112
  (
    KeyWire_0_23,
    n107
  );


  buf
  g113
  (
    n279,
    n71
  );


  buf
  g114
  (
    n377,
    n35
  );


  buf
  g115
  (
    n408,
    n87
  );


  not
  g116
  (
    n192,
    n102
  );


  not
  g117
  (
    n433,
    n24
  );


  buf
  g118
  (
    n227,
    n85
  );


  not
  g119
  (
    n442,
    n30
  );


  not
  g120
  (
    n235,
    n65
  );


  buf
  g121
  (
    n388,
    n76
  );


  buf
  g122
  (
    n126,
    n72
  );


  not
  g123
  (
    n439,
    n103
  );


  not
  g124
  (
    n294,
    n48
  );


  buf
  g125
  (
    n340,
    n65
  );


  buf
  g126
  (
    n405,
    n94
  );


  buf
  g127
  (
    n390,
    n81
  );


  not
  g128
  (
    n136,
    n69
  );


  not
  g129
  (
    n187,
    n58
  );


  buf
  g130
  (
    n329,
    n31
  );


  not
  g131
  (
    n287,
    n76
  );


  buf
  g132
  (
    n331,
    n74
  );


  not
  g133
  (
    n148,
    n80
  );


  not
  g134
  (
    n256,
    n87
  );


  buf
  g135
  (
    n193,
    n68
  );


  buf
  g136
  (
    n229,
    n25
  );


  buf
  g137
  (
    n423,
    n62
  );


  not
  g138
  (
    n250,
    n41
  );


  buf
  g139
  (
    n407,
    n29
  );


  buf
  g140
  (
    n225,
    n89
  );


  buf
  g141
  (
    n114,
    n91
  );


  not
  g142
  (
    n145,
    n51
  );


  buf
  g143
  (
    n258,
    n56
  );


  not
  g144
  (
    n209,
    n66
  );


  buf
  g145
  (
    n257,
    n77
  );


  not
  g146
  (
    n353,
    n91
  );


  not
  g147
  (
    n202,
    n104
  );


  not
  g148
  (
    n143,
    n93
  );


  buf
  g149
  (
    n363,
    n83
  );


  not
  g150
  (
    n302,
    n55
  );


  not
  g151
  (
    n432,
    n105
  );


  buf
  g152
  (
    n266,
    n60
  );


  buf
  g153
  (
    n418,
    n61
  );


  buf
  g154
  (
    n409,
    n99
  );


  buf
  g155
  (
    n204,
    n101
  );


  buf
  g156
  (
    n275,
    n37
  );


  buf
  g157
  (
    n168,
    n35
  );


  buf
  g158
  (
    n295,
    n38
  );


  not
  g159
  (
    n416,
    n67
  );


  buf
  g160
  (
    n370,
    n41
  );


  buf
  g161
  (
    n419,
    n71
  );


  not
  g162
  (
    n344,
    n33
  );


  buf
  g163
  (
    n214,
    n48
  );


  not
  g164
  (
    n198,
    n95
  );


  not
  g165
  (
    n216,
    n82
  );


  buf
  g166
  (
    n312,
    n77
  );


  buf
  g167
  (
    n365,
    n53
  );


  not
  g168
  (
    n281,
    n106
  );


  not
  g169
  (
    n436,
    n63
  );


  buf
  g170
  (
    n203,
    n59
  );


  buf
  g171
  (
    n355,
    n83
  );


  buf
  g172
  (
    n254,
    n61
  );


  buf
  g173
  (
    n146,
    n74
  );


  not
  g174
  (
    n375,
    n36
  );


  not
  g175
  (
    n396,
    n50
  );


  not
  g176
  (
    n165,
    n97
  );


  not
  g177
  (
    n149,
    n60
  );


  not
  g178
  (
    n133,
    n82
  );


  buf
  g179
  (
    n166,
    n102
  );


  not
  g180
  (
    n414,
    n48
  );


  not
  g181
  (
    n243,
    n81
  );


  not
  g182
  (
    n383,
    n34
  );


  buf
  g183
  (
    n267,
    n27
  );


  not
  g184
  (
    n205,
    n82
  );


  not
  g185
  (
    n154,
    n43
  );


  not
  g186
  (
    n137,
    n87
  );


  not
  g187
  (
    n241,
    n98
  );


  not
  g188
  (
    n277,
    n95
  );


  not
  g189
  (
    n354,
    n72
  );


  not
  g190
  (
    n270,
    n98
  );


  buf
  g191
  (
    n406,
    n26
  );


  buf
  g192
  (
    n330,
    n95
  );


  not
  g193
  (
    n399,
    n64
  );


  not
  g194
  (
    n430,
    n52
  );


  not
  g195
  (
    n237,
    n57
  );


  not
  g196
  (
    n152,
    n83
  );


  buf
  g197
  (
    n108,
    n55
  );


  not
  g198
  (
    n230,
    n39
  );


  not
  g199
  (
    n303,
    n66
  );


  not
  g200
  (
    n392,
    n63
  );


  buf
  g201
  (
    n309,
    n31
  );


  buf
  g202
  (
    n239,
    n45
  );


  buf
  g203
  (
    n304,
    n61
  );


  buf
  g204
  (
    n253,
    n27
  );


  not
  g205
  (
    n420,
    n100
  );


  buf
  g206
  (
    n368,
    n58
  );


  not
  g207
  (
    n177,
    n57
  );


  buf
  g208
  (
    n321,
    n82
  );


  not
  g209
  (
    n425,
    n100
  );


  buf
  g210
  (
    n162,
    n38
  );


  buf
  g211
  (
    n350,
    n84
  );


  buf
  g212
  (
    n335,
    n67
  );


  buf
  g213
  (
    n131,
    n88
  );


  not
  g214
  (
    n226,
    n33
  );


  buf
  g215
  (
    n194,
    n52
  );


  not
  g216
  (
    n181,
    n97
  );


  not
  g217
  (
    n178,
    n60
  );


  not
  g218
  (
    n269,
    n29
  );


  buf
  g219
  (
    n129,
    n73
  );


  buf
  g220
  (
    n122,
    n44
  );


  buf
  g221
  (
    n112,
    n89
  );


  not
  g222
  (
    n380,
    n55
  );


  buf
  g223
  (
    n426,
    n27
  );


  buf
  g224
  (
    n385,
    n39
  );


  not
  g225
  (
    n215,
    n53
  );


  buf
  g226
  (
    n282,
    n40
  );


  not
  g227
  (
    n127,
    n71
  );


  not
  g228
  (
    n342,
    n92
  );


  not
  g229
  (
    n411,
    n75
  );


  not
  g230
  (
    n263,
    n42
  );


  buf
  g231
  (
    n273,
    n54
  );


  not
  g232
  (
    n283,
    n96
  );


  not
  g233
  (
    n116,
    n83
  );


  buf
  g234
  (
    n111,
    n91
  );


  buf
  g235
  (
    n185,
    n106
  );


  not
  g236
  (
    n156,
    n50
  );


  not
  g237
  (
    n291,
    n35
  );


  buf
  g238
  (
    n120,
    n45
  );


  buf
  g239
  (
    n395,
    n62
  );


  not
  g240
  (
    n348,
    n73
  );


  not
  g241
  (
    n412,
    n90
  );


  buf
  g242
  (
    n186,
    n77
  );


  buf
  g243
  (
    n190,
    n62
  );


  not
  g244
  (
    n228,
    n40
  );


  not
  g245
  (
    n337,
    n49
  );


  not
  g246
  (
    n332,
    n65
  );


  not
  g247
  (
    n132,
    n78
  );


  buf
  g248
  (
    n328,
    n78
  );


  not
  g249
  (
    n158,
    n70
  );


  not
  g250
  (
    n341,
    n55
  );


  not
  g251
  (
    n402,
    n47
  );


  buf
  g252
  (
    n347,
    n37
  );


  buf
  g253
  (
    n361,
    n36
  );


  not
  g254
  (
    n371,
    n49
  );


  not
  g255
  (
    n440,
    n104
  );


  buf
  g256
  (
    n400,
    n47
  );


  not
  g257
  (
    n289,
    n49
  );


  buf
  g258
  (
    n224,
    n96
  );


  buf
  g259
  (
    n339,
    n95
  );


  not
  g260
  (
    n138,
    n38
  );


  buf
  g261
  (
    n338,
    n43
  );


  buf
  g262
  (
    n118,
    n76
  );


  not
  g263
  (
    n125,
    n45
  );


  not
  g264
  (
    n259,
    n37
  );


  not
  g265
  (
    n221,
    n54
  );


  buf
  g266
  (
    n346,
    n75
  );


  not
  g267
  (
    n176,
    n80
  );


  not
  g268
  (
    n244,
    n88
  );


  not
  g269
  (
    n128,
    n93
  );


  not
  g270
  (
    n382,
    n51
  );


  buf
  g271
  (
    n318,
    n43
  );


  not
  g272
  (
    n415,
    n31
  );


  not
  g273
  (
    n364,
    n56
  );


  buf
  g274
  (
    n274,
    n33
  );


  not
  g275
  (
    n424,
    n102
  );


  not
  g276
  (
    n113,
    n69
  );


  not
  g277
  (
    n173,
    n103
  );


  not
  g278
  (
    n233,
    n70
  );


  not
  g279
  (
    n366,
    n101
  );


  buf
  g280
  (
    n410,
    n86
  );


  not
  g281
  (
    n255,
    n93
  );


  buf
  g282
  (
    n300,
    n28
  );


  buf
  g283
  (
    n160,
    n75
  );


  not
  g284
  (
    n220,
    n92
  );


  buf
  g285
  (
    n115,
    n99
  );


  not
  g286
  (
    n140,
    n59
  );


  buf
  g287
  (
    n247,
    n63
  );


  buf
  g288
  (
    n298,
    n97
  );


  buf
  g289
  (
    KeyWire_0_14,
    n27
  );


  not
  g290
  (
    n376,
    n107
  );


  not
  g291
  (
    n144,
    n101
  );


  not
  g292
  (
    n169,
    n105
  );


  not
  g293
  (
    n401,
    n49
  );


  buf
  g294
  (
    n437,
    n106
  );


  not
  g295
  (
    n170,
    n53
  );


  not
  g296
  (
    n308,
    n32
  );


  buf
  g297
  (
    n443,
    n79
  );


  not
  g298
  (
    n362,
    n26
  );


  buf
  g299
  (
    n384,
    n44
  );


  buf
  g300
  (
    n280,
    n42
  );


  buf
  g301
  (
    n157,
    n46
  );


  not
  g302
  (
    n435,
    n33
  );


  buf
  g303
  (
    n147,
    n48
  );


  buf
  g304
  (
    n387,
    n70
  );


  not
  g305
  (
    n119,
    n104
  );


  not
  g306
  (
    n301,
    n65
  );


  buf
  g307
  (
    n325,
    n80
  );


  buf
  g308
  (
    n427,
    n99
  );


  buf
  g309
  (
    KeyWire_0_6,
    n58
  );


  buf
  g310
  (
    n189,
    n38
  );


  buf
  g311
  (
    n293,
    n54
  );


  buf
  g312
  (
    n317,
    n63
  );


  buf
  g313
  (
    n422,
    n60
  );


  not
  g314
  (
    n324,
    n103
  );


  not
  g315
  (
    n333,
    n78
  );


  not
  g316
  (
    n207,
    n51
  );


  not
  g317
  (
    n284,
    n53
  );


  buf
  g318
  (
    n314,
    n62
  );


  not
  g319
  (
    n394,
    n40
  );


  not
  g320
  (
    n159,
    n90
  );


  buf
  g321
  (
    n315,
    n76
  );


  not
  g322
  (
    n288,
    n89
  );


  not
  g323
  (
    n367,
    n30
  );


  buf
  g324
  (
    n305,
    n81
  );


  not
  g325
  (
    n217,
    n29
  );


  buf
  g326
  (
    n445,
    n59
  );


  not
  g327
  (
    n150,
    n40
  );


  not
  g328
  (
    n213,
    n94
  );


  buf
  g329
  (
    n195,
    n36
  );


  buf
  g330
  (
    n246,
    n25
  );


  not
  g331
  (
    n431,
    n73
  );


  buf
  g332
  (
    KeyWire_0_27,
    n29
  );


  not
  g333
  (
    n334,
    n46
  );


  not
  g334
  (
    n188,
    n91
  );


  buf
  g335
  (
    n110,
    n31
  );


  buf
  g336
  (
    n234,
    n73
  );


  buf
  g337
  (
    n434,
    n56
  );


  buf
  g338
  (
    n299,
    n30
  );


  not
  g339
  (
    n326,
    n69
  );


  buf
  g340
  (
    n381,
    n43
  );


  not
  g341
  (
    n373,
    n50
  );


  not
  g342
  (
    n180,
    n106
  );


  not
  g343
  (
    n121,
    n85
  );


  buf
  g344
  (
    n210,
    n97
  );


  not
  g345
  (
    n252,
    n47
  );


  not
  g346
  (
    n167,
    n26
  );


  buf
  g347
  (
    n212,
    n25
  );


  not
  g348
  (
    n379,
    n34
  );


  not
  g349
  (
    n179,
    n28
  );


  not
  g350
  (
    KeyWire_0_3,
    n68
  );


  not
  g351
  (
    n261,
    n77
  );


  buf
  g352
  (
    n260,
    n24
  );


  not
  g353
  (
    n201,
    n30
  );


  buf
  g354
  (
    n271,
    n42
  );


  not
  g355
  (
    n219,
    n98
  );


  not
  g356
  (
    n316,
    n85
  );


  not
  g357
  (
    n428,
    n52
  );


  buf
  g358
  (
    n183,
    n52
  );


  buf
  g359
  (
    n378,
    n50
  );


  buf
  g360
  (
    n264,
    n90
  );


  not
  g361
  (
    n421,
    n59
  );


  not
  g362
  (
    n141,
    n32
  );


  not
  g363
  (
    n397,
    n104
  );


  not
  g364
  (
    n231,
    n32
  );


  buf
  g365
  (
    n135,
    n68
  );


  not
  g366
  (
    n398,
    n80
  );


  not
  g367
  (
    n323,
    n100
  );


  not
  g368
  (
    n206,
    n90
  );


  buf
  g369
  (
    n286,
    n28
  );


  not
  g370
  (
    n265,
    n86
  );


  not
  g371
  (
    n297,
    n57
  );


  buf
  g372
  (
    n310,
    n54
  );


  not
  g373
  (
    n117,
    n105
  );


  buf
  g374
  (
    n151,
    n67
  );


  not
  g375
  (
    n327,
    n47
  );


  buf
  g376
  (
    n336,
    n32
  );


  buf
  g377
  (
    n236,
    n92
  );


  buf
  g378
  (
    n161,
    n42
  );


  not
  g379
  (
    n290,
    n64
  );


  not
  g380
  (
    n438,
    n58
  );


  not
  g381
  (
    n251,
    n25
  );


  buf
  g382
  (
    n139,
    n103
  );


  not
  g383
  (
    n349,
    n84
  );


  buf
  g384
  (
    n249,
    n64
  );


  buf
  g385
  (
    n272,
    n24
  );


  not
  g386
  (
    n163,
    n44
  );


  buf
  g387
  (
    n134,
    n51
  );


  buf
  g388
  (
    n199,
    n79
  );


  not
  g389
  (
    n109,
    n88
  );


  buf
  g390
  (
    n292,
    n44
  );


  buf
  g391
  (
    n444,
    n92
  );


  not
  g392
  (
    n404,
    n96
  );


  buf
  g393
  (
    n319,
    n75
  );


  buf
  g394
  (
    n172,
    n98
  );


  buf
  g395
  (
    n393,
    n34
  );


  not
  g396
  (
    n218,
    n46
  );


  not
  g397
  (
    n191,
    n89
  );


  not
  g398
  (
    n386,
    n84
  );


  not
  g399
  (
    n276,
    n67
  );


  not
  g400
  (
    n352,
    n46
  );


  buf
  g401
  (
    n413,
    n39
  );


  not
  g402
  (
    n142,
    n36
  );


  buf
  g403
  (
    n351,
    n94
  );


  buf
  g404
  (
    n268,
    n96
  );


  not
  g405
  (
    n356,
    n23
  );


  buf
  g406
  (
    n358,
    n66
  );


  buf
  g407
  (
    KeyWire_0_25,
    n88
  );


  buf
  g408
  (
    n391,
    n79
  );


  buf
  g409
  (
    n278,
    n72
  );


  not
  g410
  (
    n343,
    n26
  );


  not
  g411
  (
    n155,
    n102
  );


  not
  g412
  (
    n357,
    n79
  );


  not
  g413
  (
    n200,
    n86
  );


  buf
  g414
  (
    n369,
    n99
  );


  buf
  g415
  (
    n372,
    n101
  );


  not
  g416
  (
    n311,
    n68
  );


  not
  g417
  (
    n306,
    n71
  );


  buf
  g418
  (
    n307,
    n23
  );


  buf
  g419
  (
    n130,
    n69
  );


  buf
  g420
  (
    n211,
    n64
  );


  not
  g421
  (
    n175,
    n34
  );


  nand
  g422
  (
    n222,
    n85,
    n57
  );


  xor
  g423
  (
    n518,
    n329,
    n431,
    n223,
    n347
  );


  and
  g424
  (
    n515,
    n422,
    n307,
    n279,
    n256
  );


  xor
  g425
  (
    n460,
    n311,
    n232,
    n319,
    n159
  );


  nor
  g426
  (
    n521,
    n239,
    n368,
    n391,
    n421
  );


  and
  g427
  (
    n483,
    n276,
    n167,
    n419,
    n369
  );


  nand
  g428
  (
    n475,
    n379,
    n300,
    n380,
    n386
  );


  nor
  g429
  (
    n466,
    n289,
    n250,
    n406,
    n154
  );


  nor
  g430
  (
    n454,
    n199,
    n402,
    n149,
    n242
  );


  or
  g431
  (
    n465,
    n194,
    n230,
    n225,
    n176
  );


  xnor
  g432
  (
    n476,
    n203,
    n352,
    n326,
    n346
  );


  xnor
  g433
  (
    n497,
    n165,
    n383,
    n127,
    n152
  );


  xor
  g434
  (
    n494,
    n410,
    n309,
    n443,
    n192
  );


  or
  g435
  (
    n486,
    n171,
    n136,
    n417,
    n375
  );


  xor
  g436
  (
    KeyWire_0_0,
    n111,
    n268,
    n144,
    n312
  );


  and
  g437
  (
    n482,
    n313,
    n376,
    n292,
    n328
  );


  nor
  g438
  (
    KeyWire_0_26,
    n384,
    n186,
    n443,
    n116
  );


  xnor
  g439
  (
    n484,
    n290,
    n374,
    n148,
    n295
  );


  xnor
  g440
  (
    n471,
    n187,
    n273,
    n207,
    n299
  );


  nor
  g441
  (
    n523,
    n353,
    n424,
    n126,
    n170
  );


  xnor
  g442
  (
    n495,
    n291,
    n286,
    n206,
    n153
  );


  nand
  g443
  (
    n457,
    n243,
    n177,
    n120,
    n444
  );


  nand
  g444
  (
    n458,
    n123,
    n244,
    n293,
    n172
  );


  and
  g445
  (
    n508,
    n110,
    n215,
    n414,
    n443
  );


  nand
  g446
  (
    n499,
    n335,
    n420,
    n394,
    n388
  );


  xnor
  g447
  (
    n459,
    n261,
    n363,
    n124,
    n109
  );


  and
  g448
  (
    n489,
    n235,
    n316,
    n409,
    n141
  );


  nor
  g449
  (
    KeyWire_0_5,
    n439,
    n341,
    n218,
    n357
  );


  and
  g450
  (
    n479,
    n125,
    n282,
    n366,
    n285
  );


  nand
  g451
  (
    n488,
    n331,
    n284,
    n224,
    n164
  );


  xnor
  g452
  (
    n447,
    n178,
    n301,
    n430,
    n382
  );


  nand
  g453
  (
    n502,
    n270,
    n150,
    n168,
    n441
  );


  or
  g454
  (
    n487,
    n401,
    n405,
    n404,
    n355
  );


  and
  g455
  (
    n450,
    n433,
    n189,
    n156,
    n343
  );


  and
  g456
  (
    n462,
    n275,
    n135,
    n181,
    n137
  );


  xor
  g457
  (
    n520,
    n184,
    n333,
    n130,
    n255
  );


  nor
  g458
  (
    n503,
    n332,
    n348,
    n188,
    n241
  );


  nand
  g459
  (
    n464,
    n396,
    n119,
    n226,
    n336
  );


  and
  g460
  (
    n524,
    n408,
    n434,
    n272,
    n305
  );


  or
  g461
  (
    n485,
    n129,
    n107,
    n280,
    n392
  );


  xnor
  g462
  (
    n511,
    n211,
    n412,
    n365,
    n323
  );


  and
  g463
  (
    n455,
    n163,
    n358,
    n415,
    n399
  );


  and
  g464
  (
    n519,
    n246,
    n183,
    n443,
    n370
  );


  nor
  g465
  (
    n473,
    n429,
    n271,
    n373,
    n200
  );


  nor
  g466
  (
    n463,
    n147,
    n281,
    n354,
    n303
  );


  xnor
  g467
  (
    n478,
    n321,
    n214,
    n330,
    n205
  );


  xor
  g468
  (
    n468,
    n212,
    n428,
    n361,
    n185
  );


  nor
  g469
  (
    n480,
    n425,
    n390,
    n155,
    n423
  );


  xnor
  g470
  (
    n501,
    n108,
    n315,
    n400,
    n233
  );


  xnor
  g471
  (
    n449,
    n296,
    n175,
    n160,
    n283
  );


  and
  g472
  (
    n504,
    n302,
    n442,
    n432,
    n362
  );


  xor
  g473
  (
    n530,
    n360,
    n310,
    n139,
    n437
  );


  and
  g474
  (
    n506,
    n314,
    n146,
    n413,
    n356
  );


  xnor
  g475
  (
    n531,
    n217,
    n198,
    n134,
    n371
  );


  xor
  g476
  (
    n500,
    n377,
    n440,
    n351,
    n201
  );


  or
  g477
  (
    n514,
    n121,
    n253,
    n131,
    n228
  );


  xor
  g478
  (
    n491,
    n277,
    n444,
    n143,
    n287
  );


  nand
  g479
  (
    n512,
    n173,
    n113,
    n387,
    n267
  );


  nand
  g480
  (
    n516,
    n389,
    n248,
    n344,
    n133
  );


  nor
  g481
  (
    n517,
    n247,
    n325,
    n210,
    n237
  );


  xor
  g482
  (
    n522,
    n385,
    n367,
    n234,
    n158
  );


  and
  g483
  (
    n448,
    n162,
    n249,
    n259,
    n138
  );


  xor
  g484
  (
    n472,
    n298,
    n180,
    n118,
    n245
  );


  or
  g485
  (
    n498,
    n145,
    n213,
    n112,
    n438
  );


  nor
  g486
  (
    n509,
    n320,
    n381,
    n208,
    n339
  );


  xnor
  g487
  (
    n510,
    n266,
    n403,
    n182,
    n342
  );


  or
  g488
  (
    n453,
    n350,
    n322,
    n436,
    n142
  );


  xor
  g489
  (
    n474,
    n209,
    n398,
    n338,
    n169
  );


  nand
  g490
  (
    n513,
    n257,
    n364,
    n324,
    n397
  );


  nor
  g491
  (
    n467,
    n337,
    n318,
    n227,
    n190
  );


  xor
  g492
  (
    n469,
    n304,
    n260,
    n238,
    n327
  );


  nand
  g493
  (
    n493,
    n222,
    n115,
    n426,
    n294
  );


  xor
  g494
  (
    n452,
    n288,
    n197,
    n306,
    n308
  );


  nand
  g495
  (
    n490,
    n411,
    n254,
    n252,
    n258
  );


  nand
  g496
  (
    n492,
    n221,
    n345,
    n264,
    n418
  );


  and
  g497
  (
    n529,
    n349,
    n117,
    n435,
    n193
  );


  xnor
  g498
  (
    n481,
    n372,
    n262,
    n204,
    n297
  );


  xor
  g499
  (
    n525,
    n219,
    n265,
    n278,
    n416
  );


  nor
  g500
  (
    n496,
    n166,
    n395,
    n191,
    n114
  );


  xnor
  g501
  (
    n526,
    n140,
    n269,
    n157,
    n128
  );


  or
  g502
  (
    n528,
    n340,
    n334,
    n122,
    n359
  );


  nor
  g503
  (
    n461,
    n196,
    n179,
    n174,
    n263
  );


  nor
  g504
  (
    n507,
    n378,
    n274,
    n151,
    n317
  );


  and
  g505
  (
    n505,
    n231,
    n220,
    n444,
    n229
  );


  or
  g506
  (
    n451,
    n161,
    n427,
    n251,
    n407
  );


  nor
  g507
  (
    n446,
    n195,
    n132,
    n202,
    n240
  );


  xor
  g508
  (
    n477,
    n444,
    n216,
    n236,
    n393
  );


  buf
  g509
  (
    n550,
    n469
  );


  buf
  g510
  (
    n552,
    n452
  );


  buf
  g511
  (
    n547,
    n457
  );


  not
  g512
  (
    n533,
    n467
  );


  buf
  g513
  (
    n554,
    n462
  );


  buf
  g514
  (
    n546,
    n460
  );


  buf
  g515
  (
    n548,
    n450
  );


  buf
  g516
  (
    n551,
    n453
  );


  buf
  g517
  (
    n539,
    n454
  );


  buf
  g518
  (
    n543,
    n451
  );


  buf
  g519
  (
    n535,
    n456
  );


  not
  g520
  (
    n538,
    n447
  );


  buf
  g521
  (
    n553,
    n471
  );


  not
  g522
  (
    n542,
    n472
  );


  not
  g523
  (
    n537,
    n465
  );


  buf
  g524
  (
    n540,
    n468
  );


  not
  g525
  (
    n534,
    n455
  );


  not
  g526
  (
    n555,
    n466
  );


  buf
  g527
  (
    n544,
    n448
  );


  buf
  g528
  (
    n536,
    n446
  );


  not
  g529
  (
    n541,
    n464
  );


  not
  g530
  (
    n557,
    n458
  );


  buf
  g531
  (
    n549,
    n463
  );


  buf
  g532
  (
    n532,
    n470
  );


  buf
  g533
  (
    n545,
    n473
  );


  buf
  g534
  (
    KeyWire_0_7,
    n449
  );


  not
  g535
  (
    KeyWire_0_29,
    n461
  );


  not
  g536
  (
    n556,
    n459
  );


  not
  g537
  (
    n560,
    n532
  );


  not
  g538
  (
    n561,
    n532
  );


  nand
  g539
  (
    n564,
    n475,
    n482,
    n483,
    n476
  );


  or
  g540
  (
    n563,
    n490,
    n496,
    n561,
    n474
  );


  and
  g541
  (
    n567,
    n486,
    n560,
    n481,
    n478
  );


  nand
  g542
  (
    n566,
    n497,
    n561,
    n489,
    n487
  );


  and
  g543
  (
    n565,
    n560,
    n480,
    n484,
    n495
  );


  and
  g544
  (
    n569,
    n561,
    n560,
    n488,
    n479
  );


  xnor
  g545
  (
    n568,
    n561,
    n491,
    n560,
    n477
  );


  xnor
  g546
  (
    n562,
    n492,
    n494,
    n493,
    n485
  );


  not
  g547
  (
    n576,
    n563
  );


  buf
  g548
  (
    n572,
    n565
  );


  not
  g549
  (
    n570,
    n563
  );


  buf
  g550
  (
    n575,
    n565
  );


  buf
  g551
  (
    n586,
    n566
  );


  buf
  g552
  (
    n584,
    n564
  );


  not
  g553
  (
    n573,
    n564
  );


  not
  g554
  (
    n589,
    n565
  );


  not
  g555
  (
    n585,
    n562
  );


  buf
  g556
  (
    n583,
    n563
  );


  buf
  g557
  (
    n580,
    n564
  );


  buf
  g558
  (
    n578,
    n565
  );


  buf
  g559
  (
    n579,
    n562
  );


  buf
  g560
  (
    n582,
    n562
  );


  buf
  g561
  (
    n577,
    n566
  );


  buf
  g562
  (
    n571,
    n562
  );


  not
  g563
  (
    n581,
    n564
  );


  buf
  g564
  (
    n587,
    n563
  );


  not
  g565
  (
    n588,
    n566
  );


  not
  g566
  (
    n574,
    n566
  );


  buf
  g567
  (
    n665,
    n577
  );


  not
  g568
  (
    n625,
    n577
  );


  buf
  g569
  (
    n654,
    n582
  );


  buf
  g570
  (
    n601,
    n588
  );


  not
  g571
  (
    n618,
    n577
  );


  buf
  g572
  (
    n648,
    n573
  );


  buf
  g573
  (
    n590,
    n580
  );


  buf
  g574
  (
    n614,
    n575
  );


  not
  g575
  (
    n652,
    n588
  );


  buf
  g576
  (
    n593,
    n581
  );


  buf
  g577
  (
    n612,
    n574
  );


  buf
  g578
  (
    n637,
    n575
  );


  buf
  g579
  (
    n632,
    n584
  );


  buf
  g580
  (
    n649,
    n571
  );


  not
  g581
  (
    n658,
    n570
  );


  buf
  g582
  (
    n596,
    n582
  );


  not
  g583
  (
    n595,
    n577
  );


  not
  g584
  (
    n608,
    n570
  );


  not
  g585
  (
    n634,
    n583
  );


  not
  g586
  (
    n653,
    n572
  );


  buf
  g587
  (
    n663,
    n584
  );


  not
  g588
  (
    n646,
    n587
  );


  buf
  g589
  (
    n667,
    n579
  );


  buf
  g590
  (
    n597,
    n580
  );


  not
  g591
  (
    n604,
    n579
  );


  buf
  g592
  (
    n621,
    n571
  );


  not
  g593
  (
    n599,
    n576
  );


  buf
  g594
  (
    n605,
    n578
  );


  buf
  g595
  (
    n615,
    n572
  );


  not
  g596
  (
    n633,
    n573
  );


  buf
  g597
  (
    n617,
    n583
  );


  not
  g598
  (
    n610,
    n587
  );


  buf
  g599
  (
    n609,
    n575
  );


  not
  g600
  (
    n600,
    n585
  );


  buf
  g601
  (
    n657,
    n589
  );


  buf
  g602
  (
    KeyWire_0_8,
    n588
  );


  not
  g603
  (
    n643,
    n573
  );


  buf
  g604
  (
    n656,
    n589
  );


  buf
  g605
  (
    n603,
    n581
  );


  not
  g606
  (
    n602,
    n570
  );


  buf
  g607
  (
    n591,
    n578
  );


  buf
  g608
  (
    n661,
    n576
  );


  buf
  g609
  (
    n647,
    n583
  );


  buf
  g610
  (
    n640,
    n587
  );


  not
  g611
  (
    n636,
    n579
  );


  not
  g612
  (
    n629,
    n589
  );


  not
  g613
  (
    n613,
    n576
  );


  buf
  g614
  (
    n624,
    n584
  );


  not
  g615
  (
    n662,
    n571
  );


  buf
  g616
  (
    n594,
    n574
  );


  not
  g617
  (
    n635,
    n574
  );


  buf
  g618
  (
    n645,
    n586
  );


  buf
  g619
  (
    n606,
    n585
  );


  not
  g620
  (
    n622,
    n585
  );


  not
  g621
  (
    n660,
    n589
  );


  buf
  g622
  (
    n620,
    n579
  );


  buf
  g623
  (
    n607,
    n578
  );


  buf
  g624
  (
    n628,
    n581
  );


  not
  g625
  (
    n669,
    n586
  );


  not
  g626
  (
    n631,
    n575
  );


  not
  g627
  (
    n616,
    n585
  );


  buf
  g628
  (
    n619,
    n587
  );


  buf
  g629
  (
    n639,
    n584
  );


  not
  g630
  (
    n664,
    n571
  );


  not
  g631
  (
    n630,
    n578
  );


  buf
  g632
  (
    n666,
    n586
  );


  not
  g633
  (
    n651,
    n580
  );


  buf
  g634
  (
    n638,
    n583
  );


  buf
  g635
  (
    n659,
    n573
  );


  not
  g636
  (
    n592,
    n574
  );


  buf
  g637
  (
    n641,
    n588
  );


  buf
  g638
  (
    n627,
    n572
  );


  buf
  g639
  (
    n626,
    n582
  );


  not
  g640
  (
    n650,
    n586
  );


  not
  g641
  (
    n644,
    n576
  );


  buf
  g642
  (
    n623,
    n572
  );


  buf
  g643
  (
    n642,
    n582
  );


  buf
  g644
  (
    n598,
    n580
  );


  not
  g645
  (
    n655,
    n570
  );


  buf
  g646
  (
    n668,
    n581
  );


  not
  g647
  (
    n865,
    n612
  );


  buf
  g648
  (
    n963,
    n594
  );


  not
  g649
  (
    n863,
    n647
  );


  not
  g650
  (
    n955,
    n590
  );


  not
  g651
  (
    n915,
    n598
  );


  not
  g652
  (
    n796,
    n543
  );


  buf
  g653
  (
    n827,
    n663
  );


  not
  g654
  (
    n705,
    n621
  );


  buf
  g655
  (
    n779,
    n639
  );


  buf
  g656
  (
    n821,
    n614
  );


  buf
  g657
  (
    n899,
    n598
  );


  not
  g658
  (
    n730,
    n556
  );


  not
  g659
  (
    n789,
    n534
  );


  not
  g660
  (
    n761,
    n626
  );


  buf
  g661
  (
    n770,
    n655
  );


  not
  g662
  (
    n856,
    n619
  );


  not
  g663
  (
    n776,
    n596
  );


  buf
  g664
  (
    n867,
    n595
  );


  not
  g665
  (
    n976,
    n637
  );


  not
  g666
  (
    n842,
    n623
  );


  buf
  g667
  (
    n743,
    n640
  );


  buf
  g668
  (
    n787,
    n593
  );


  not
  g669
  (
    n670,
    n622
  );


  not
  g670
  (
    n788,
    n593
  );


  not
  g671
  (
    n913,
    n595
  );


  not
  g672
  (
    n782,
    n591
  );


  buf
  g673
  (
    n837,
    n606
  );


  not
  g674
  (
    n971,
    n568
  );


  not
  g675
  (
    n859,
    n591
  );


  not
  g676
  (
    n783,
    n535
  );


  not
  g677
  (
    n984,
    n615
  );


  buf
  g678
  (
    n681,
    n533
  );


  buf
  g679
  (
    n876,
    n627
  );


  buf
  g680
  (
    n895,
    n602
  );


  buf
  g681
  (
    n759,
    n603
  );


  not
  g682
  (
    n718,
    n636
  );


  buf
  g683
  (
    n957,
    n612
  );


  buf
  g684
  (
    n711,
    n618
  );


  buf
  g685
  (
    n757,
    n649
  );


  not
  g686
  (
    n801,
    n607
  );


  not
  g687
  (
    n846,
    n627
  );


  buf
  g688
  (
    n910,
    n639
  );


  not
  g689
  (
    n838,
    n659
  );


  not
  g690
  (
    n869,
    n646
  );


  not
  g691
  (
    n708,
    n538
  );


  not
  g692
  (
    n852,
    n646
  );


  not
  g693
  (
    n735,
    n629
  );


  not
  g694
  (
    n841,
    n557
  );


  buf
  g695
  (
    n857,
    n557
  );


  buf
  g696
  (
    n786,
    n596
  );


  not
  g697
  (
    n832,
    n662
  );


  not
  g698
  (
    n715,
    n535
  );


  buf
  g699
  (
    n900,
    n559
  );


  buf
  g700
  (
    n695,
    n603
  );


  not
  g701
  (
    n673,
    n559
  );


  not
  g702
  (
    n820,
    n550
  );


  buf
  g703
  (
    n977,
    n617
  );


  buf
  g704
  (
    n890,
    n541
  );


  buf
  g705
  (
    KeyWire_0_11,
    n623
  );


  buf
  g706
  (
    n974,
    n602
  );


  buf
  g707
  (
    KeyWire_0_1,
    n648
  );


  not
  g708
  (
    n817,
    n539
  );


  not
  g709
  (
    n721,
    n633
  );


  buf
  g710
  (
    n960,
    n593
  );


  buf
  g711
  (
    n729,
    n603
  );


  not
  g712
  (
    n725,
    n549
  );


  not
  g713
  (
    n868,
    n643
  );


  buf
  g714
  (
    n753,
    n610
  );


  buf
  g715
  (
    n843,
    n534
  );


  buf
  g716
  (
    n970,
    n594
  );


  not
  g717
  (
    n983,
    n504
  );


  buf
  g718
  (
    n747,
    n541
  );


  buf
  g719
  (
    n936,
    n622
  );


  buf
  g720
  (
    n862,
    n632
  );


  buf
  g721
  (
    n826,
    n633
  );


  buf
  g722
  (
    n798,
    n556
  );


  buf
  g723
  (
    n961,
    n533
  );


  not
  g724
  (
    n964,
    n660
  );


  buf
  g725
  (
    n917,
    n549
  );


  buf
  g726
  (
    n851,
    n642
  );


  buf
  g727
  (
    n741,
    n594
  );


  buf
  g728
  (
    n864,
    n538
  );


  not
  g729
  (
    n968,
    n547
  );


  not
  g730
  (
    n750,
    n643
  );


  not
  g731
  (
    n985,
    n665
  );


  buf
  g732
  (
    n671,
    n611
  );


  not
  g733
  (
    n703,
    n666
  );


  not
  g734
  (
    n896,
    n556
  );


  not
  g735
  (
    n815,
    n647
  );


  not
  g736
  (
    n745,
    n608
  );


  not
  g737
  (
    n953,
    n552
  );


  not
  g738
  (
    n720,
    n656
  );


  buf
  g739
  (
    n736,
    n631
  );


  not
  g740
  (
    n797,
    n551
  );


  not
  g741
  (
    n941,
    n667
  );


  not
  g742
  (
    n847,
    n668
  );


  buf
  g743
  (
    n793,
    n533
  );


  not
  g744
  (
    n946,
    n642
  );


  buf
  g745
  (
    n914,
    n610
  );


  buf
  g746
  (
    n828,
    n536
  );


  buf
  g747
  (
    n849,
    n555
  );


  buf
  g748
  (
    n774,
    n620
  );


  buf
  g749
  (
    n756,
    n669
  );


  not
  g750
  (
    n965,
    n599
  );


  not
  g751
  (
    n922,
    n658
  );


  not
  g752
  (
    n824,
    n619
  );


  buf
  g753
  (
    n902,
    n550
  );


  buf
  g754
  (
    n702,
    n656
  );


  buf
  g755
  (
    n688,
    n600
  );


  not
  g756
  (
    n950,
    n591
  );


  not
  g757
  (
    n923,
    n643
  );


  buf
  g758
  (
    KeyWire_0_30,
    n626
  );


  not
  g759
  (
    n903,
    n636
  );


  buf
  g760
  (
    n680,
    n655
  );


  buf
  g761
  (
    n858,
    n597
  );


  not
  g762
  (
    n755,
    n618
  );


  not
  g763
  (
    n933,
    n604
  );


  not
  g764
  (
    n700,
    n625
  );


  buf
  g765
  (
    n879,
    n666
  );


  not
  g766
  (
    n898,
    n606
  );


  buf
  g767
  (
    n959,
    n639
  );


  not
  g768
  (
    n816,
    n646
  );


  not
  g769
  (
    n905,
    n661
  );


  buf
  g770
  (
    n945,
    n544
  );


  buf
  g771
  (
    n752,
    n599
  );


  not
  g772
  (
    n784,
    n659
  );


  buf
  g773
  (
    n728,
    n543
  );


  buf
  g774
  (
    n931,
    n664
  );


  buf
  g775
  (
    n758,
    n599
  );


  buf
  g776
  (
    n763,
    n621
  );


  buf
  g777
  (
    KeyWire_0_20,
    n554
  );


  not
  g778
  (
    n714,
    n595
  );


  buf
  g779
  (
    n944,
    n534
  );


  not
  g780
  (
    n981,
    n630
  );


  buf
  g781
  (
    n701,
    n567
  );


  not
  g782
  (
    n830,
    n548
  );


  buf
  g783
  (
    n834,
    n545
  );


  buf
  g784
  (
    n699,
    n542
  );


  buf
  g785
  (
    n823,
    n629
  );


  buf
  g786
  (
    n691,
    n623
  );


  buf
  g787
  (
    n911,
    n661
  );


  not
  g788
  (
    n948,
    n662
  );


  buf
  g789
  (
    n717,
    n644
  );


  buf
  g790
  (
    n966,
    n630
  );


  not
  g791
  (
    n860,
    n622
  );


  not
  g792
  (
    n805,
    n652
  );


  not
  g793
  (
    n930,
    n649
  );


  not
  g794
  (
    n937,
    n636
  );


  not
  g795
  (
    n986,
    n628
  );


  buf
  g796
  (
    n762,
    n541
  );


  not
  g797
  (
    n727,
    n546
  );


  not
  g798
  (
    n881,
    n643
  );


  buf
  g799
  (
    n871,
    n627
  );


  buf
  g800
  (
    n769,
    n537
  );


  not
  g801
  (
    n952,
    n546
  );


  not
  g802
  (
    n694,
    n663
  );


  not
  g803
  (
    n891,
    n615
  );


  not
  g804
  (
    n811,
    n609
  );


  not
  g805
  (
    n853,
    n568
  );


  not
  g806
  (
    n818,
    n657
  );


  buf
  g807
  (
    n822,
    n650
  );


  not
  g808
  (
    n771,
    n659
  );


  not
  g809
  (
    KeyWire_0_4,
    n609
  );


  not
  g810
  (
    n794,
    n548
  );


  buf
  g811
  (
    n795,
    n658
  );


  not
  g812
  (
    n684,
    n617
  );


  buf
  g813
  (
    KeyWire_0_24,
    n631
  );


  buf
  g814
  (
    n696,
    n655
  );


  buf
  g815
  (
    n848,
    n567
  );


  buf
  g816
  (
    n825,
    n647
  );


  not
  g817
  (
    n829,
    n558
  );


  not
  g818
  (
    n975,
    n660
  );


  not
  g819
  (
    n781,
    n625
  );


  not
  g820
  (
    n740,
    n645
  );


  not
  g821
  (
    n766,
    n615
  );


  buf
  g822
  (
    n693,
    n537
  );


  not
  g823
  (
    n835,
    n650
  );


  buf
  g824
  (
    n768,
    n543
  );


  not
  g825
  (
    n926,
    n606
  );


  not
  g826
  (
    n958,
    n546
  );


  not
  g827
  (
    n935,
    n601
  );


  buf
  g828
  (
    n760,
    n592
  );


  not
  g829
  (
    n775,
    n548
  );


  not
  g830
  (
    n932,
    n568
  );


  buf
  g831
  (
    n676,
    n552
  );


  not
  g832
  (
    n790,
    n605
  );


  not
  g833
  (
    n887,
    n553
  );


  not
  g834
  (
    n908,
    n547
  );


  not
  g835
  (
    n894,
    n568
  );


  not
  g836
  (
    n919,
    n611
  );


  buf
  g837
  (
    n912,
    n638
  );


  buf
  g838
  (
    n866,
    n536
  );


  not
  g839
  (
    n722,
    n613
  );


  not
  g840
  (
    n850,
    n595
  );


  not
  g841
  (
    n901,
    n644
  );


  not
  g842
  (
    n672,
    n616
  );


  not
  g843
  (
    n839,
    n506
  );


  buf
  g844
  (
    n765,
    n598
  );


  buf
  g845
  (
    n878,
    n545
  );


  not
  g846
  (
    n954,
    n632
  );


  buf
  g847
  (
    n803,
    n624
  );


  buf
  g848
  (
    n880,
    n665
  );


  not
  g849
  (
    n943,
    n555
  );


  buf
  g850
  (
    n973,
    n604
  );


  not
  g851
  (
    n812,
    n614
  );


  not
  g852
  (
    n738,
    n548
  );


  buf
  g853
  (
    n893,
    n621
  );


  not
  g854
  (
    n921,
    n554
  );


  buf
  g855
  (
    n810,
    n609
  );


  not
  g856
  (
    n686,
    n559
  );


  buf
  g857
  (
    n883,
    n535
  );


  not
  g858
  (
    n814,
    n537
  );


  not
  g859
  (
    n710,
    n598
  );


  not
  g860
  (
    n892,
    n601
  );


  not
  g861
  (
    n939,
    n597
  );


  buf
  g862
  (
    n928,
    n542
  );


  buf
  g863
  (
    n833,
    n668
  );


  not
  g864
  (
    n692,
    n637
  );


  not
  g865
  (
    n697,
    n638
  );


  not
  g866
  (
    n877,
    n550
  );


  not
  g867
  (
    n873,
    n535
  );


  not
  g868
  (
    n861,
    n556
  );


  not
  g869
  (
    n929,
    n590
  );


  buf
  g870
  (
    n713,
    n552
  );


  not
  g871
  (
    n683,
    n540
  );


  not
  g872
  (
    n791,
    n594
  );


  not
  g873
  (
    n716,
    n634
  );


  buf
  g874
  (
    n967,
    n649
  );


  not
  g875
  (
    n704,
    n635
  );


  not
  g876
  (
    n978,
    n635
  );


  not
  g877
  (
    n739,
    n538
  );


  not
  g878
  (
    n800,
    n622
  );


  not
  g879
  (
    n927,
    n604
  );


  not
  g880
  (
    n792,
    n608
  );


  not
  g881
  (
    n916,
    n616
  );


  not
  g882
  (
    n742,
    n646
  );


  buf
  g883
  (
    n882,
    n559
  );


  buf
  g884
  (
    n987,
    n632
  );


  not
  g885
  (
    KeyWire_0_2,
    n547
  );


  not
  g886
  (
    n773,
    n593
  );


  buf
  g887
  (
    n726,
    n591
  );


  buf
  g888
  (
    n886,
    n607
  );


  buf
  g889
  (
    n685,
    n558
  );


  not
  g890
  (
    n840,
    n638
  );


  buf
  g891
  (
    n956,
    n540
  );


  buf
  g892
  (
    n844,
    n657
  );


  not
  g893
  (
    n689,
    n654
  );


  buf
  g894
  (
    n819,
    n553
  );


  not
  g895
  (
    n778,
    n549
  );


  not
  g896
  (
    n724,
    n661
  );


  not
  g897
  (
    n972,
    n500
  );


  not
  g898
  (
    n764,
    n605
  );


  not
  g899
  (
    n907,
    n637
  );


  not
  g900
  (
    n872,
    n636
  );


  not
  g901
  (
    n813,
    n553
  );


  not
  g902
  (
    n884,
    n624
  );


  buf
  g903
  (
    n888,
    n607
  );


  not
  g904
  (
    n942,
    n650
  );


  buf
  g905
  (
    n807,
    n659
  );


  not
  g906
  (
    n874,
    n540
  );


  not
  g907
  (
    n675,
    n653
  );


  buf
  g908
  (
    n870,
    n657
  );


  not
  g909
  (
    n909,
    n551
  );


  not
  g910
  (
    n924,
    n641
  );


  buf
  g911
  (
    n906,
    n545
  );


  buf
  g912
  (
    n749,
    n549
  );


  not
  g913
  (
    n875,
    n625
  );


  buf
  g914
  (
    n734,
    n645
  );


  buf
  g915
  (
    n918,
    n628
  );


  not
  g916
  (
    n706,
    n645
  );


  not
  g917
  (
    n674,
    n620
  );


  buf
  g918
  (
    n980,
    n532
  );


  not
  g919
  (
    n885,
    n536
  );


  not
  g920
  (
    n951,
    n599
  );


  nand
  g921
  (
    n751,
    n651,
    n614
  );


  xor
  g922
  (
    n934,
    n644,
    n616,
    n619,
    n640
  );


  nor
  g923
  (
    n709,
    n603,
    n613,
    n547,
    n658
  );


  and
  g924
  (
    n969,
    n542,
    n658,
    n654,
    n633
  );


  xnor
  g925
  (
    n831,
    n601,
    n557,
    n617,
    n652
  );


  xor
  g926
  (
    n731,
    n610,
    n502,
    n650,
    n536
  );


  nor
  g927
  (
    n719,
    n567,
    n567,
    n654,
    n532
  );


  nand
  g928
  (
    n712,
    n669,
    n639,
    n626,
    n645
  );


  or
  g929
  (
    n947,
    n628,
    n498,
    n669,
    n554
  );


  nand
  g930
  (
    n809,
    n661,
    n641,
    n544
  );


  xor
  g931
  (
    n679,
    n629,
    n499,
    n543,
    n551
  );


  xor
  g932
  (
    n737,
    n606,
    n602,
    n613,
    n539
  );


  nand
  g933
  (
    n982,
    n539,
    n653,
    n545,
    n637
  );


  xor
  g934
  (
    n698,
    n665,
    n663,
    n619,
    n601
  );


  xnor
  g935
  (
    n682,
    n505,
    n609,
    n592,
    n644
  );


  xnor
  g936
  (
    n845,
    n602,
    n596,
    n634,
    n592
  );


  or
  g937
  (
    n767,
    n546,
    n642,
    n608,
    n631
  );


  xnor
  g938
  (
    n746,
    n608,
    n663,
    n539,
    n503
  );


  nor
  g939
  (
    n772,
    n640,
    n630,
    n652,
    n553
  );


  or
  g940
  (
    n777,
    n669,
    n610,
    n533,
    n600
  );


  nand
  g941
  (
    n979,
    n640,
    n540,
    n612,
    n635
  );


  xnor
  g942
  (
    n785,
    n633,
    n666,
    n550,
    n656
  );


  nand
  g943
  (
    n754,
    n534,
    n635,
    n654,
    n631
  );


  xnor
  g944
  (
    n690,
    n605,
    n618,
    n668,
    n667
  );


  nor
  g945
  (
    n925,
    n596,
    n615,
    n648,
    n651
  );


  xnor
  g946
  (
    n938,
    n501,
    n665,
    n551,
    n648
  );


  or
  g947
  (
    n904,
    n620,
    n660,
    n664,
    n507
  );


  nand
  g948
  (
    n962,
    n624,
    n612,
    n604,
    n607
  );


  nor
  g949
  (
    n780,
    n537,
    n611,
    n600,
    n653
  );


  xor
  g950
  (
    n802,
    n620,
    n555,
    n634
  );


  and
  g951
  (
    n732,
    n557,
    n624,
    n621,
    n653
  );


  nand
  g952
  (
    n744,
    n664,
    n667,
    n558,
    n634
  );


  xor
  g953
  (
    n855,
    n641,
    n651,
    n648,
    n542
  );


  xor
  g954
  (
    n799,
    n592,
    n618,
    n656,
    n628
  );


  xnor
  g955
  (
    n806,
    n541,
    n666,
    n600,
    n558
  );


  xnor
  g956
  (
    n897,
    n662,
    n652,
    n617,
    n605
  );


  nor
  g957
  (
    n920,
    n597,
    n544,
    n667
  );


  xor
  g958
  (
    n678,
    n625,
    n538,
    n660,
    n623
  );


  xor
  g959
  (
    n677,
    n657,
    n611,
    n627,
    n651
  );


  nor
  g960
  (
    n949,
    n647,
    n629,
    n554,
    n664
  );


  nand
  g961
  (
    n889,
    n642,
    n638,
    n616,
    n630
  );


  and
  g962
  (
    n804,
    n649,
    n597,
    n626,
    n655
  );


  xnor
  g963
  (
    n854,
    n614,
    n613,
    n668,
    n590
  );


  xnor
  g964
  (
    n940,
    n662,
    n632,
    n552,
    n590
  );


  buf
  g965
  (
    n996,
    n682
  );


  not
  g966
  (
    n993,
    n679
  );


  not
  g967
  (
    n995,
    n678
  );


  not
  g968
  (
    n989,
    n671
  );


  not
  g969
  (
    n997,
    n677
  );


  buf
  g970
  (
    n994,
    n683
  );


  not
  g971
  (
    n1000,
    n684
  );


  buf
  g972
  (
    n1002,
    n681
  );


  buf
  g973
  (
    n1001,
    n674
  );


  buf
  g974
  (
    n999,
    n675
  );


  not
  g975
  (
    n988,
    n670
  );


  buf
  g976
  (
    n991,
    n672
  );


  buf
  g977
  (
    n992,
    n685
  );


  buf
  g978
  (
    n990,
    n676
  );


  and
  g979
  (
    n998,
    n680,
    n673
  );


  not
  g980
  (
    n1011,
    n994
  );


  buf
  g981
  (
    n1019,
    n990
  );


  not
  g982
  (
    n1021,
    n998
  );


  buf
  g983
  (
    n1005,
    n989
  );


  not
  g984
  (
    n1009,
    n995
  );


  not
  g985
  (
    n1008,
    n999
  );


  not
  g986
  (
    n1013,
    n1001
  );


  buf
  g987
  (
    n1016,
    n1000
  );


  buf
  g988
  (
    n1020,
    n992
  );


  not
  g989
  (
    n1004,
    n1000
  );


  buf
  g990
  (
    n1017,
    n1002
  );


  not
  g991
  (
    n1012,
    n991
  );


  buf
  g992
  (
    n1003,
    n993
  );


  not
  g993
  (
    n1015,
    n1001
  );


  buf
  g994
  (
    n1018,
    n1000
  );


  buf
  g995
  (
    n1022,
    n997
  );


  not
  g996
  (
    n1007,
    n1002
  );


  not
  g997
  (
    n1006,
    n1000
  );


  not
  g998
  (
    n1024,
    n988
  );


  not
  g999
  (
    n1014,
    n1001
  );


  not
  g1000
  (
    n1023,
    n996
  );


  buf
  g1001
  (
    n1010,
    n1001
  );


  nand
  g1002
  (
    n1085,
    n792,
    n902,
    n940,
    n853
  );


  nand
  g1003
  (
    n1066,
    n701,
    n919,
    n915,
    n1013
  );


  and
  g1004
  (
    n1101,
    n1009,
    n748,
    n1011,
    n769
  );


  xor
  g1005
  (
    n1091,
    n717,
    n780,
    n820,
    n897
  );


  and
  g1006
  (
    n1078,
    n749,
    n754,
    n931,
    n850
  );


  xor
  g1007
  (
    n1054,
    n927,
    n788,
    n1005,
    n1010
  );


  nand
  g1008
  (
    n1048,
    n943,
    n880,
    n844,
    n1013
  );


  or
  g1009
  (
    n1032,
    n904,
    n819,
    n921,
    n822
  );


  xor
  g1010
  (
    n1029,
    n884,
    n727,
    n705,
    n874
  );


  and
  g1011
  (
    n1072,
    n756,
    n941,
    n703,
    n1022
  );


  xor
  g1012
  (
    n1074,
    n737,
    n872,
    n768,
    n901
  );


  xnor
  g1013
  (
    n1071,
    n707,
    n1011,
    n716,
    n799
  );


  and
  g1014
  (
    n1058,
    n1008,
    n752,
    n761,
    n755
  );


  nor
  g1015
  (
    n1031,
    n895,
    n690,
    n827,
    n1013
  );


  and
  g1016
  (
    n1088,
    n1012,
    n686,
    n777,
    n917
  );


  xnor
  g1017
  (
    n1070,
    n936,
    n1015,
    n813,
    n841
  );


  nor
  g1018
  (
    n1104,
    n702,
    n1014,
    n1015,
    n886
  );


  nor
  g1019
  (
    n1065,
    n1010,
    n858,
    n775,
    n1004
  );


  xor
  g1020
  (
    n1075,
    n876,
    n713,
    n857,
    n773
  );


  nor
  g1021
  (
    n1097,
    n866,
    n803,
    n818,
    n729
  );


  nor
  g1022
  (
    n1092,
    n738,
    n719,
    n861,
    n770
  );


  xnor
  g1023
  (
    n1025,
    n1012,
    n1018,
    n1007
  );


  nor
  g1024
  (
    KeyWire_0_9,
    n1019,
    n753,
    n691,
    n945
  );


  xor
  g1025
  (
    n1052,
    n694,
    n782,
    n1004,
    n767
  );


  and
  g1026
  (
    n1044,
    n837,
    n787,
    n843,
    n948
  );


  xor
  g1027
  (
    n1053,
    n860,
    n877,
    n845,
    n720
  );


  nand
  g1028
  (
    n1034,
    n706,
    n1016,
    n1019,
    n898
  );


  and
  g1029
  (
    n1036,
    n781,
    n854,
    n825,
    n789
  );


  and
  g1030
  (
    n1045,
    n928,
    n784,
    n846,
    n747
  );


  and
  g1031
  (
    n1067,
    n771,
    n1003,
    n757,
    n772
  );


  nand
  g1032
  (
    n1076,
    n839,
    n1006,
    n791,
    n1003
  );


  xor
  g1033
  (
    n1079,
    n920,
    n712,
    n923,
    n1021
  );


  and
  g1034
  (
    n1086,
    n865,
    n912,
    n842,
    n1006
  );


  xor
  g1035
  (
    n1042,
    n811,
    n726,
    n736,
    n1022
  );


  or
  g1036
  (
    n1105,
    n743,
    n750,
    n700,
    n933
  );


  xnor
  g1037
  (
    n1055,
    n746,
    n758,
    n1007,
    n1005
  );


  and
  g1038
  (
    n1041,
    n1022,
    n821,
    n1009,
    n1016
  );


  xnor
  g1039
  (
    n1033,
    n833,
    n693,
    n1008,
    n869
  );


  or
  g1040
  (
    n1087,
    n1014,
    n1006,
    n835
  );


  or
  g1041
  (
    n1111,
    n689,
    n1021,
    n1004,
    n910
  );


  and
  g1042
  (
    n1028,
    n1019,
    n724,
    n805,
    n826
  );


  and
  g1043
  (
    n1051,
    n812,
    n836,
    n734,
    n739
  );


  nand
  g1044
  (
    n1039,
    n938,
    n1017,
    n742,
    n1015
  );


  or
  g1045
  (
    n1068,
    n864,
    n744,
    n778,
    n889
  );


  and
  g1046
  (
    KeyWire_0_12,
    n1017,
    n763,
    n890,
    n715
  );


  and
  g1047
  (
    n1069,
    n900,
    n862,
    n1016,
    n882
  );


  nand
  g1048
  (
    n1110,
    n793,
    n859,
    n883,
    n1008
  );


  xnor
  g1049
  (
    n1057,
    n1015,
    n1018,
    n944,
    n937
  );


  xor
  g1050
  (
    n1046,
    n856,
    n1017,
    n765,
    n1010
  );


  and
  g1051
  (
    n1099,
    n1009,
    n908,
    n688,
    n696
  );


  nor
  g1052
  (
    n1060,
    n830,
    n1022,
    n831,
    n1003
  );


  or
  g1053
  (
    n1026,
    n1024,
    n714,
    n1023,
    n774
  );


  xor
  g1054
  (
    n1077,
    n732,
    n722,
    n1020
  );


  and
  g1055
  (
    n1062,
    n815,
    n802,
    n1014,
    n741
  );


  xor
  g1056
  (
    n1100,
    n1021,
    n1004,
    n847,
    n709
  );


  nand
  g1057
  (
    n1103,
    n867,
    n949,
    n785,
    n786
  );


  xor
  g1058
  (
    n1096,
    n916,
    n711,
    n906,
    n779
  );


  nor
  g1059
  (
    KeyWire_0_15,
    n733,
    n922,
    n929,
    n888
  );


  or
  g1060
  (
    n1030,
    n878,
    n695,
    n834,
    n848
  );


  or
  g1061
  (
    n1059,
    n925,
    n790,
    n704,
    n764
  );


  or
  g1062
  (
    n1106,
    n699,
    n816,
    n728,
    n698
  );


  nor
  g1063
  (
    n1084,
    n1012,
    n725,
    n794,
    n766
  );


  and
  g1064
  (
    n1050,
    n1011,
    n838,
    n817,
    n855
  );


  nand
  g1065
  (
    n1040,
    n934,
    n849,
    n804,
    n801
  );


  and
  g1066
  (
    n1112,
    n891,
    n808,
    n932,
    n926
  );


  or
  g1067
  (
    n1089,
    n851,
    n896,
    n730,
    n751
  );


  xor
  g1068
  (
    n1095,
    n824,
    n913,
    n731,
    n776
  );


  xnor
  g1069
  (
    n1037,
    n907,
    n759,
    n795,
    n1023
  );


  nor
  g1070
  (
    n1064,
    n797,
    n1024,
    n723,
    n809
  );


  nor
  g1071
  (
    n1035,
    n914,
    n1018,
    n1024,
    n1005
  );


  xor
  g1072
  (
    n1098,
    n708,
    n823,
    n721,
    n762
  );


  nor
  g1073
  (
    n1080,
    n939,
    n905,
    n1017,
    n1011
  );


  nor
  g1074
  (
    KeyWire_0_21,
    n893,
    n875,
    n863,
    n918
  );


  xor
  g1075
  (
    n1056,
    n930,
    n873,
    n1016,
    n894
  );


  or
  g1076
  (
    n1090,
    n885,
    n1009,
    n807,
    n1024
  );


  and
  g1077
  (
    n1038,
    n692,
    n798,
    n832,
    n1020
  );


  and
  g1078
  (
    n1109,
    n829,
    n810,
    n892,
    n1005
  );


  nor
  g1079
  (
    n1082,
    n946,
    n697,
    n814,
    n1012
  );


  nor
  g1080
  (
    n1108,
    n800,
    n911,
    n879,
    n1003
  );


  nor
  g1081
  (
    n1081,
    n1007,
    n1020,
    n710,
    n871
  );


  xnor
  g1082
  (
    n1043,
    n881,
    n935,
    n1021,
    n796
  );


  nor
  g1083
  (
    n1049,
    n852,
    n947,
    n870,
    n1007
  );


  and
  g1084
  (
    n1093,
    n840,
    n899,
    n806,
    n868
  );


  xnor
  g1085
  (
    n1027,
    n1013,
    n1014,
    n760,
    n718
  );


  xor
  g1086
  (
    n1073,
    n828,
    n942,
    n1023,
    n909
  );


  nor
  g1087
  (
    n1063,
    n745,
    n1023,
    n903,
    n1010
  );


  nand
  g1088
  (
    n1102,
    n687,
    n1019,
    n1008,
    n740
  );


  and
  g1089
  (
    n1047,
    n783,
    n887,
    n735,
    n924
  );


  buf
  g1090
  (
    n1113,
    n1034
  );


  buf
  g1091
  (
    n1128,
    n1043
  );


  not
  g1092
  (
    n1126,
    n445
  );


  not
  g1093
  (
    n1124,
    n1044
  );


  not
  g1094
  (
    n1131,
    n1046
  );


  not
  g1095
  (
    n1115,
    n1031
  );


  buf
  g1096
  (
    n1117,
    n445
  );


  buf
  g1097
  (
    n1133,
    n1040
  );


  not
  g1098
  (
    n1132,
    n1039
  );


  not
  g1099
  (
    n1119,
    n1041
  );


  not
  g1100
  (
    n1130,
    n1032
  );


  not
  g1101
  (
    n1116,
    n1042
  );


  buf
  g1102
  (
    KeyWire_0_16,
    n1047
  );


  not
  g1103
  (
    n1134,
    n1037
  );


  buf
  g1104
  (
    n1129,
    n1036
  );


  not
  g1105
  (
    n1135,
    n1025
  );


  buf
  g1106
  (
    n1118,
    n1030
  );


  not
  g1107
  (
    n1127,
    n1027
  );


  buf
  g1108
  (
    n1121,
    n1048
  );


  buf
  g1109
  (
    n1120,
    n1045
  );


  not
  g1110
  (
    n1125,
    n1038
  );


  not
  g1111
  (
    n1114,
    n1029
  );


  buf
  g1112
  (
    n1123,
    n1035
  );


  nand
  g1113
  (
    n1122,
    n1028,
    n1033,
    n1026
  );


  nand
  g1114
  (
    n1146,
    n520,
    n955,
    n967,
    n980
  );


  xor
  g1115
  (
    n1139,
    n978,
    n979,
    n1113
  );


  and
  g1116
  (
    n1143,
    n1116,
    n1113,
    n952,
    n521
  );


  and
  g1117
  (
    n1153,
    n1118,
    n980,
    n954,
    n976
  );


  xnor
  g1118
  (
    n1140,
    n961,
    n1116,
    n510,
    n1119
  );


  or
  g1119
  (
    n1150,
    n519,
    n970,
    n516,
    n1114
  );


  xor
  g1120
  (
    n1152,
    n974,
    n1115,
    n1117
  );


  nand
  g1121
  (
    n1137,
    n968,
    n508,
    n512,
    n964
  );


  and
  g1122
  (
    n1159,
    n977,
    n960,
    n980,
    n972
  );


  xnor
  g1123
  (
    n1145,
    n957,
    n968,
    n1115,
    n1117
  );


  xnor
  g1124
  (
    n1161,
    n1119,
    n969,
    n1114,
    n976
  );


  nand
  g1125
  (
    n1157,
    n958,
    n975,
    n977
  );


  xor
  g1126
  (
    n1151,
    n1115,
    n1118,
    n966,
    n979
  );


  nand
  g1127
  (
    n1156,
    n977,
    n978,
    n515,
    n968
  );


  xor
  g1128
  (
    n1148,
    n965,
    n509,
    n1114,
    n1117
  );


  xnor
  g1129
  (
    n1141,
    n980,
    n970,
    n1113,
    n1116
  );


  nand
  g1130
  (
    n1147,
    n518,
    n976,
    n978,
    n1118
  );


  and
  g1131
  (
    n1158,
    n517,
    n1114,
    n977,
    n511
  );


  xnor
  g1132
  (
    n1163,
    n976,
    n969,
    n973,
    n971
  );


  nand
  g1133
  (
    n1164,
    n975,
    n974,
    n1115
  );


  xnor
  g1134
  (
    n1142,
    n978,
    n971,
    n951,
    n1119
  );


  nand
  g1135
  (
    n1162,
    n513,
    n962,
    n1118,
    n979
  );


  nor
  g1136
  (
    n1144,
    n514,
    n973,
    n959,
    n970
  );


  nor
  g1137
  (
    n1155,
    n953,
    n973,
    n1119,
    n972
  );


  or
  g1138
  (
    n1160,
    n970,
    n972,
    n975,
    n969
  );


  or
  g1139
  (
    n1149,
    n968,
    n950,
    n963,
    n971
  );


  nor
  g1140
  (
    n1154,
    n974,
    n1116,
    n971,
    n956
  );


  xor
  g1141
  (
    n1138,
    n969,
    n973,
    n972,
    n1113
  );


  or
  g1142
  (
    n1188,
    n1085,
    n1086,
    n1061,
    n1074
  );


  or
  g1143
  (
    KeyWire_0_18,
    n1091,
    n1073,
    n1002,
    n1050
  );


  and
  g1144
  (
    n1181,
    n1095,
    n1053,
    n1072,
    n1148
  );


  xnor
  g1145
  (
    n1186,
    n1081,
    n1054,
    n1073,
    n1163
  );


  nor
  g1146
  (
    n1192,
    n1083,
    n1083,
    n1094,
    n1086
  );


  nand
  g1147
  (
    n1167,
    n1075,
    n1159,
    n1162,
    n1083
  );


  and
  g1148
  (
    n1169,
    n1162,
    n1089,
    n1002,
    n1090
  );


  xor
  g1149
  (
    n1196,
    n1052,
    n1162,
    n1082,
    n1079
  );


  nor
  g1150
  (
    n1202,
    n1071,
    n1153,
    n1094,
    n1143
  );


  or
  g1151
  (
    n1168,
    n1068,
    n1090,
    n1088,
    n1146
  );


  and
  g1152
  (
    n1182,
    n1161,
    n1079,
    n1075,
    n1076
  );


  and
  g1153
  (
    n1184,
    n1163,
    n1092,
    n1088,
    n1154
  );


  or
  g1154
  (
    n1189,
    n1084,
    n1080,
    n1091,
    n1074
  );


  and
  g1155
  (
    n1203,
    n1083,
    n1089,
    n1075,
    n1085
  );


  nor
  g1156
  (
    n1165,
    n1093,
    n1152,
    n1086,
    n1078
  );


  xor
  g1157
  (
    n1170,
    n1087,
    n1164,
    n1049,
    n1090
  );


  or
  g1158
  (
    n1174,
    n1092,
    n1056,
    n1082,
    n1077
  );


  and
  g1159
  (
    n1185,
    n1057,
    n1138,
    n1065,
    n1072
  );


  nor
  g1160
  (
    n1179,
    n1139,
    n1095,
    n1164,
    n1079
  );


  and
  g1161
  (
    n1176,
    n1089,
    n1094,
    n1091,
    n1081
  );


  or
  g1162
  (
    n1177,
    n1055,
    n1164,
    n1081,
    n1078
  );


  or
  g1163
  (
    n1187,
    n1088,
    n1087,
    n1149,
    n1161
  );


  xor
  g1164
  (
    n1195,
    n1077,
    n1076,
    n1058,
    n1092
  );


  and
  g1165
  (
    n1178,
    n1059,
    n1089,
    n1093,
    n1147
  );


  xor
  g1166
  (
    n1171,
    n1085,
    n1162,
    n1064,
    n1137
  );


  nand
  g1167
  (
    n1166,
    n1073,
    n1076,
    n1092,
    n1144
  );


  nor
  g1168
  (
    n1180,
    n1096,
    n1158,
    n1074,
    n1163
  );


  xor
  g1169
  (
    n1198,
    n1164,
    n1140,
    n1087,
    n1145
  );


  nand
  g1170
  (
    n1175,
    n1076,
    n1093,
    n1160,
    n1063
  );


  and
  g1171
  (
    n1199,
    n1051,
    n1062,
    n1163,
    n1078
  );


  or
  g1172
  (
    n1191,
    n1060,
    n1077,
    n1080,
    n1090
  );


  nand
  g1173
  (
    n1197,
    n1075,
    n1080,
    n1094,
    n1066
  );


  xnor
  g1174
  (
    n1193,
    n1069,
    n1074,
    n1088,
    n1080
  );


  nor
  g1175
  (
    n1204,
    n1079,
    n1141,
    n1070,
    n1084
  );


  nand
  g1176
  (
    n1200,
    n1077,
    n1087,
    n1095,
    n1091
  );


  nand
  g1177
  (
    n1201,
    n1078,
    n1082,
    n1156,
    n1067
  );


  xor
  g1178
  (
    n1183,
    n1142,
    n1071,
    n1161,
    n1151
  );


  nand
  g1179
  (
    n1190,
    n1085,
    n1095,
    n1157,
    n1081
  );


  and
  g1180
  (
    n1172,
    n1086,
    n1084,
    n1082,
    n1150
  );


  xor
  g1181
  (
    n1173,
    n1155,
    n1161,
    n1084,
    n1093
  );


  not
  g1182
  (
    n1297,
    n1124
  );


  not
  g1183
  (
    n1262,
    n1197
  );


  not
  g1184
  (
    n1242,
    n1178
  );


  not
  g1185
  (
    n1299,
    n1196
  );


  buf
  g1186
  (
    n1295,
    n982
  );


  not
  g1187
  (
    n1350,
    n1171
  );


  not
  g1188
  (
    n1346,
    n1121
  );


  not
  g1189
  (
    n1215,
    n1128
  );


  not
  g1190
  (
    n1244,
    n981
  );


  not
  g1191
  (
    n1222,
    n1180
  );


  not
  g1192
  (
    n1287,
    n1123
  );


  buf
  g1193
  (
    n1302,
    n528
  );


  buf
  g1194
  (
    n1334,
    n983
  );


  buf
  g1195
  (
    n1255,
    n1174
  );


  buf
  g1196
  (
    n1260,
    n1131
  );


  not
  g1197
  (
    n1338,
    n1182
  );


  buf
  g1198
  (
    n1293,
    n1191
  );


  not
  g1199
  (
    n1246,
    n1175
  );


  not
  g1200
  (
    n1229,
    n1187
  );


  not
  g1201
  (
    n1335,
    n1181
  );


  not
  g1202
  (
    n1218,
    n1183
  );


  buf
  g1203
  (
    KeyWire_0_13,
    n1193
  );


  not
  g1204
  (
    n1296,
    n1122
  );


  not
  g1205
  (
    n1216,
    n1175
  );


  buf
  g1206
  (
    n1300,
    n1120
  );


  not
  g1207
  (
    n1211,
    n1203
  );


  buf
  g1208
  (
    n1265,
    n1120
  );


  buf
  g1209
  (
    n1236,
    n1167
  );


  buf
  g1210
  (
    n1328,
    n1193
  );


  buf
  g1211
  (
    n1349,
    n1182
  );


  not
  g1212
  (
    n1271,
    n1129
  );


  not
  g1213
  (
    n1304,
    n1123
  );


  buf
  g1214
  (
    n1320,
    n1179
  );


  buf
  g1215
  (
    n1226,
    n1187
  );


  buf
  g1216
  (
    n1212,
    n1180
  );


  buf
  g1217
  (
    n1234,
    n1197
  );


  buf
  g1218
  (
    n1208,
    n1180
  );


  not
  g1219
  (
    n1282,
    n1192
  );


  buf
  g1220
  (
    n1280,
    n1188
  );


  not
  g1221
  (
    n1258,
    n1125
  );


  not
  g1222
  (
    n1309,
    n1185
  );


  buf
  g1223
  (
    n1256,
    n1183
  );


  buf
  g1224
  (
    n1261,
    n1190
  );


  buf
  g1225
  (
    n1321,
    n1191
  );


  not
  g1226
  (
    n1341,
    n1175
  );


  buf
  g1227
  (
    n1301,
    n445
  );


  buf
  g1228
  (
    n1323,
    n1194
  );


  buf
  g1229
  (
    n1257,
    n1191
  );


  not
  g1230
  (
    n1276,
    n982
  );


  not
  g1231
  (
    n1266,
    n1174
  );


  buf
  g1232
  (
    n1288,
    n1124
  );


  buf
  g1233
  (
    n1259,
    n1170
  );


  not
  g1234
  (
    n1223,
    n1176
  );


  buf
  g1235
  (
    n1230,
    n1198
  );


  not
  g1236
  (
    n1241,
    n1190
  );


  not
  g1237
  (
    n1306,
    n1129
  );


  buf
  g1238
  (
    n1289,
    n1176
  );


  buf
  g1239
  (
    n1303,
    n1199
  );


  buf
  g1240
  (
    n1263,
    n984
  );


  not
  g1241
  (
    n1235,
    n1127
  );


  buf
  g1242
  (
    n1205,
    n1183
  );


  not
  g1243
  (
    n1311,
    n1185
  );


  buf
  g1244
  (
    n1278,
    n1133
  );


  not
  g1245
  (
    n1272,
    n1126
  );


  buf
  g1246
  (
    n1247,
    n524
  );


  not
  g1247
  (
    n1342,
    n1124
  );


  not
  g1248
  (
    n1250,
    n1177
  );


  buf
  g1249
  (
    n1264,
    n1184
  );


  not
  g1250
  (
    n1307,
    n1201
  );


  buf
  g1251
  (
    n1348,
    n1200
  );


  not
  g1252
  (
    n1344,
    n1203
  );


  not
  g1253
  (
    n1273,
    n1173
  );


  buf
  g1254
  (
    n1253,
    n1179
  );


  not
  g1255
  (
    n1327,
    n1195
  );


  buf
  g1256
  (
    n1252,
    n1173
  );


  buf
  g1257
  (
    n1240,
    n1188
  );


  buf
  g1258
  (
    n1330,
    n1175
  );


  buf
  g1259
  (
    n1284,
    n1096
  );


  not
  g1260
  (
    n1277,
    n982
  );


  buf
  g1261
  (
    n1217,
    n1197
  );


  buf
  g1262
  (
    n1220,
    n1130
  );


  buf
  g1263
  (
    n1221,
    n1199
  );


  not
  g1264
  (
    n1331,
    n1176
  );


  not
  g1265
  (
    n1322,
    n1176
  );


  buf
  g1266
  (
    n1228,
    n1202
  );


  not
  g1267
  (
    KeyWire_0_10,
    n1131
  );


  buf
  g1268
  (
    n1298,
    n1166
  );


  not
  g1269
  (
    n1270,
    n1126
  );


  not
  g1270
  (
    n1285,
    n1135
  );


  buf
  g1271
  (
    n1206,
    n1189
  );


  not
  g1272
  (
    n1254,
    n1194
  );


  not
  g1273
  (
    n1245,
    n1180
  );


  buf
  g1274
  (
    n1325,
    n1179
  );


  not
  g1275
  (
    n1249,
    n1192
  );


  not
  g1276
  (
    n1231,
    n1133
  );


  not
  g1277
  (
    n1243,
    n1168
  );


  not
  g1278
  (
    n1290,
    n1127
  );


  not
  g1279
  (
    n1308,
    n1121
  );


  buf
  g1280
  (
    n1232,
    n1201
  );


  buf
  g1281
  (
    n1314,
    n983
  );


  not
  g1282
  (
    n1318,
    n1130
  );


  not
  g1283
  (
    n1294,
    n1200
  );


  not
  g1284
  (
    n1210,
    n1123
  );


  buf
  g1285
  (
    n1227,
    n1166
  );


  not
  g1286
  (
    n1269,
    n1193
  );


  buf
  g1287
  (
    n1233,
    n982
  );


  not
  g1288
  (
    n1279,
    n1177
  );


  buf
  g1289
  (
    KeyWire_0_31,
    n522
  );


  buf
  g1290
  (
    n1345,
    n1177
  );


  buf
  g1291
  (
    n1347,
    n1134
  );


  xnor
  g1292
  (
    n1275,
    n1191,
    n981,
    n1203,
    n1178
  );


  and
  g1293
  (
    KeyWire_0_17,
    n523,
    n1197,
    n1182,
    n1199
  );


  nand
  g1294
  (
    n1336,
    n1192,
    n1184,
    n1165,
    n529
  );


  xor
  g1295
  (
    n1333,
    n1171,
    n1185,
    n1134,
    n1128
  );


  and
  g1296
  (
    n1319,
    n1132,
    n1131,
    n1184,
    n1134
  );


  xor
  g1297
  (
    n1339,
    n1184,
    n1187,
    n1129,
    n1169
  );


  xor
  g1298
  (
    n1312,
    n1203,
    n1136,
    n984
  );


  or
  g1299
  (
    n1313,
    n981,
    n983,
    n1168,
    n1186
  );


  xnor
  g1300
  (
    n1337,
    n1186,
    n1177,
    n1122,
    n1173
  );


  or
  g1301
  (
    n1329,
    n1166,
    n1188,
    n527,
    n1198
  );


  xnor
  g1302
  (
    n1316,
    n1169,
    n1172,
    n1201,
    n1125
  );


  and
  g1303
  (
    n1224,
    n1167,
    n1182,
    n1165,
    n1186
  );


  xor
  g1304
  (
    n1274,
    n1189,
    n1133,
    n1169,
    n1204
  );


  xnor
  g1305
  (
    n1332,
    n1171,
    n1194,
    n526,
    n1132
  );


  and
  g1306
  (
    n1248,
    n1202,
    n1128,
    n1195,
    n1196
  );


  xor
  g1307
  (
    n1207,
    n1120,
    n1125,
    n1132,
    n1165
  );


  nand
  g1308
  (
    n1283,
    n1172,
    n1172,
    n1124,
    n1186
  );


  or
  g1309
  (
    n1214,
    n1127,
    n1192,
    n1122,
    n1165
  );


  nand
  g1310
  (
    n1286,
    n1200,
    n981,
    n1181,
    n1129
  );


  nand
  g1311
  (
    n1209,
    n1195,
    n1190,
    n1123,
    n1183
  );


  xnor
  g1312
  (
    n1281,
    n1170,
    n1178,
    n1185,
    n1128
  );


  xnor
  g1313
  (
    n1310,
    n1135,
    n1204,
    n445,
    n1130
  );


  or
  g1314
  (
    n1340,
    n1181,
    n525,
    n1200,
    n1125
  );


  nand
  g1315
  (
    n1326,
    n1187,
    n1189,
    n1130,
    n1170
  );


  or
  g1316
  (
    n1315,
    n1178,
    n1126,
    n1173,
    n1196
  );


  nand
  g1317
  (
    n1219,
    n984,
    n1188,
    n1204,
    n1201
  );


  xnor
  g1318
  (
    n1343,
    n1170,
    n1179,
    n1193,
    n1168
  );


  and
  g1319
  (
    n1267,
    n1171,
    n1126,
    n1122,
    n1167
  );


  xor
  g1320
  (
    n1238,
    n1202,
    n1189,
    n1121,
    n1133
  );


  xor
  g1321
  (
    n1291,
    n1204,
    n1195,
    n1135,
    n1168
  );


  or
  g1322
  (
    n1251,
    n1121,
    n1194,
    n1135,
    n1167
  );


  nand
  g1323
  (
    n1213,
    n1181,
    n1198,
    n984
  );


  and
  g1324
  (
    n1324,
    n1169,
    n1166,
    n1132,
    n1174
  );


  nand
  g1325
  (
    n1268,
    n1190,
    n1127,
    n983,
    n1172
  );


  nand
  g1326
  (
    n1239,
    n1136,
    n1199,
    n1120,
    n1174
  );


  nand
  g1327
  (
    n1292,
    n1131,
    n1136,
    n1202,
    n1196
  );


  nor
  g1328
  (
    n1367,
    n530,
    n1101,
    n1311,
    n1278
  );


  nor
  g1329
  (
    n1396,
    n1239,
    n1244,
    n1110,
    n1243
  );


  xnor
  g1330
  (
    n1353,
    n1328,
    n1096,
    n1305,
    n1217
  );


  xnor
  g1331
  (
    n1404,
    n1108,
    n1102,
    n1346,
    n1240
  );


  xnor
  g1332
  (
    n1369,
    n1106,
    n1299,
    n1111,
    n1286
  );


  xor
  g1333
  (
    n1387,
    n1320,
    n1213,
    n1103,
    n1105
  );


  or
  g1334
  (
    n1352,
    n1097,
    n1234,
    n986,
    n1225
  );


  xnor
  g1335
  (
    n1401,
    n1272,
    n1097,
    n1101,
    n1334
  );


  xor
  g1336
  (
    n1377,
    n1098,
    n1341,
    n1242,
    n1109
  );


  and
  g1337
  (
    n1398,
    n1098,
    n1230,
    n1108,
    n1229
  );


  and
  g1338
  (
    n1403,
    n1099,
    n1262,
    n1104,
    n1325
  );


  xnor
  g1339
  (
    n1363,
    n1316,
    n1107,
    n1218,
    n1326
  );


  and
  g1340
  (
    n1366,
    n1340,
    n1271,
    n1338,
    n1284
  );


  nor
  g1341
  (
    n1397,
    n1312,
    n1261,
    n1281,
    n1327
  );


  xnor
  g1342
  (
    n1374,
    n1303,
    n1101,
    n1246,
    n1291
  );


  nor
  g1343
  (
    n1405,
    n1233,
    n1339,
    n1267,
    n1106
  );


  or
  g1344
  (
    n1400,
    n1105,
    n1307,
    n1097,
    n1283
  );


  and
  g1345
  (
    n1399,
    n1250,
    n1347,
    n1350,
    n1298
  );


  xnor
  g1346
  (
    n1361,
    n1112,
    n1323,
    n1253,
    n1302
  );


  or
  g1347
  (
    KeyWire_0_22,
    n1275,
    n1241,
    n569,
    n1263
  );


  or
  g1348
  (
    n1382,
    n1304,
    n1102,
    n569,
    n1098
  );


  or
  g1349
  (
    n1359,
    n1099,
    n1296,
    n1110,
    n1333
  );


  nor
  g1350
  (
    n1386,
    n1112,
    n1321,
    n1342,
    n1322
  );


  and
  g1351
  (
    n1364,
    n1247,
    n1310,
    n1287,
    n1279
  );


  or
  g1352
  (
    n1380,
    n985,
    n1285,
    n1318,
    n1235
  );


  xnor
  g1353
  (
    n1351,
    n1212,
    n1248,
    n1216,
    n1105
  );


  xnor
  g1354
  (
    n1383,
    n1264,
    n1226,
    n1265,
    n1344
  );


  and
  g1355
  (
    n1375,
    n1345,
    n1236,
    n1103,
    n1096
  );


  xor
  g1356
  (
    n1372,
    n1111,
    n1223,
    n1100,
    n569
  );


  nand
  g1357
  (
    n1371,
    n1300,
    n1269,
    n1105,
    n1343
  );


  nor
  g1358
  (
    n1392,
    n1292,
    n1104,
    n1112,
    n985
  );


  nand
  g1359
  (
    n1391,
    n986,
    n1308,
    n1210,
    n1319
  );


  xnor
  g1360
  (
    n1406,
    n1301,
    n1259,
    n1268,
    n1108
  );


  or
  g1361
  (
    n1402,
    n1219,
    n1324,
    n1335,
    n1112
  );


  xor
  g1362
  (
    n1360,
    n1349,
    n1277,
    n1290,
    n1231
  );


  and
  g1363
  (
    n1393,
    n1315,
    n1109,
    n1222,
    n1276
  );


  and
  g1364
  (
    n1356,
    n1103,
    n1109,
    n1288,
    n1337
  );


  and
  g1365
  (
    n1354,
    n1336,
    n1329,
    n1227,
    n1237
  );


  or
  g1366
  (
    n1355,
    n1251,
    n1228,
    n986,
    n1306
  );


  and
  g1367
  (
    n1385,
    n1348,
    n1256,
    n1104,
    n1273
  );


  and
  g1368
  (
    n1362,
    n1108,
    n1289,
    n985,
    n1098
  );


  nand
  g1369
  (
    n1368,
    n1101,
    n1215,
    n1274,
    n1102
  );


  xor
  g1370
  (
    n1370,
    n1208,
    n1211,
    n1107,
    n1252
  );


  or
  g1371
  (
    n1394,
    n1270,
    n1245,
    n1209,
    n1293
  );


  and
  g1372
  (
    n1395,
    n1255,
    n1100,
    n1295,
    n1297
  );


  xor
  g1373
  (
    n1373,
    n1109,
    n1294,
    n1313,
    n569
  );


  or
  g1374
  (
    n1357,
    n1110,
    n1111,
    n1317,
    n1207
  );


  xor
  g1375
  (
    n1365,
    n1257,
    n1282,
    n1220,
    n1107
  );


  and
  g1376
  (
    n1389,
    n1206,
    n1100,
    n1099,
    n1103
  );


  xor
  g1377
  (
    n1379,
    n1097,
    n1224,
    n1254,
    n1331
  );


  xnor
  g1378
  (
    n1384,
    n1111,
    n1266,
    n1100,
    n1104
  );


  nor
  g1379
  (
    n1358,
    n1205,
    n1106,
    n1258
  );


  nand
  g1380
  (
    n1378,
    n1314,
    n1214,
    n1102,
    n1280
  );


  nor
  g1381
  (
    n1376,
    n1309,
    n1332,
    n1107,
    n1110
  );


  nand
  g1382
  (
    n1390,
    n1221,
    n1249,
    n1330,
    n1232
  );


  xor
  g1383
  (
    n1381,
    n1260,
    n985,
    n1099,
    n1238
  );


  not
  g1384
  (
    n1407,
    n1383
  );


  not
  g1385
  (
    n1410,
    n1378
  );


  buf
  g1386
  (
    n1409,
    n1384
  );


  not
  g1387
  (
    n1408,
    n1386
  );


  and
  g1388
  (
    n1412,
    n1380,
    n1382
  );


  nand
  g1389
  (
    n1411,
    n1385,
    n1387,
    n1379,
    n1381
  );


  nand
  g1390
  (
    n1414,
    n1390,
    n1396,
    n1412,
    n1393
  );


  xnor
  g1391
  (
    n1416,
    n1395,
    n1388,
    n1394,
    n1410
  );


  or
  g1392
  (
    n1413,
    n1400,
    n1398,
    n1392,
    n1401
  );


  nand
  g1393
  (
    n1415,
    n1411,
    n1391,
    n1389,
    n1397
  );


  or
  g1394
  (
    n1417,
    n1408,
    n1409,
    n1407,
    n1399
  );


  nor
  g1395
  (
    n1419,
    n1415,
    n531,
    n987,
    n1413
  );


  nor
  g1396
  (
    n1418,
    n1405,
    n1417,
    n1406,
    n987
  );


  or
  g1397
  (
    n1421,
    n1416,
    n986,
    n1403,
    n1404
  );


  xnor
  g1398
  (
    n1420,
    n1402,
    n1414,
    n987
  );


  xnor
  KeyGate_0_0
  (
    n470,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n836,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n733,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n359,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n748,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n456,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n389,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n559,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n611,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1094,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n1317,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n687,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1061,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1237,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n320,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1107,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1136,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1305,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1194,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n248,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n808,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1083,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1388,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n242,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n707,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n360,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n527,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n153,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n50,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n558,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n723,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1225,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


