

module Stat_2757_36_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n2301,
  n2318,
  n2343,
  n2341,
  n2333,
  n2336,
  n2334,
  n2342,
  n2335,
  n2418,
  n2684,
  n2682,
  n2691,
  n2753,
  n2778,
  n2766,
  n2762,
  n2749,
  n2777,
  n2764,
  n2769,
  n2758,
  n2770,
  n2751,
  n2779,
  n2759,
  n2771,
  n2776,
  n2756,
  n2760,
  n2761,
  n2774,
  n2750,
  n2768,
  n2765,
  n2780,
  n2763,
  n2757,
  n2767,
  n2752,
  n2754,
  n2775,
  n2755,
  n2781,
  n2772,
  n2773
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n2301;output n2318;output n2343;output n2341;output n2333;output n2336;output n2334;output n2342;output n2335;output n2418;output n2684;output n2682;output n2691;output n2753;output n2778;output n2766;output n2762;output n2749;output n2777;output n2764;output n2769;output n2758;output n2770;output n2751;output n2779;output n2759;output n2771;output n2776;output n2756;output n2760;output n2761;output n2774;output n2750;output n2768;output n2765;output n2780;output n2763;output n2757;output n2767;output n2752;output n2754;output n2775;output n2755;output n2781;output n2772;output n2773;
  wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2337;wire n2338;wire n2339;wire n2340;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2683;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;

  buf
  g0
  (
    n110,
    n12
  );


  not
  g1
  (
    n94,
    n19
  );


  not
  g2
  (
    n77,
    n11
  );


  buf
  g3
  (
    n62,
    n13
  );


  buf
  g4
  (
    n87,
    n3
  );


  buf
  g5
  (
    n25,
    n6
  );


  buf
  g6
  (
    n113,
    n15
  );


  not
  g7
  (
    n42,
    n9
  );


  buf
  g8
  (
    n56,
    n7
  );


  buf
  g9
  (
    n82,
    n7
  );


  not
  g10
  (
    n66,
    n3
  );


  buf
  g11
  (
    n57,
    n24
  );


  not
  g12
  (
    n43,
    n18
  );


  buf
  g13
  (
    n102,
    n2
  );


  not
  g14
  (
    n31,
    n16
  );


  not
  g15
  (
    n84,
    n5
  );


  not
  g16
  (
    n92,
    n8
  );


  buf
  g17
  (
    n53,
    n8
  );


  buf
  g18
  (
    n88,
    n13
  );


  buf
  g19
  (
    n65,
    n13
  );


  not
  g20
  (
    n81,
    n5
  );


  buf
  g21
  (
    n91,
    n17
  );


  buf
  g22
  (
    n108,
    n4
  );


  buf
  g23
  (
    n111,
    n10
  );


  not
  g24
  (
    n27,
    n10
  );


  buf
  g25
  (
    n51,
    n1
  );


  buf
  g26
  (
    n39,
    n16
  );


  buf
  g27
  (
    n83,
    n12
  );


  buf
  g28
  (
    n115,
    n22
  );


  not
  g29
  (
    n107,
    n10
  );


  not
  g30
  (
    n26,
    n20
  );


  buf
  g31
  (
    n71,
    n22
  );


  buf
  g32
  (
    n58,
    n21
  );


  buf
  g33
  (
    n109,
    n4
  );


  not
  g34
  (
    n112,
    n6
  );


  buf
  g35
  (
    n75,
    n17
  );


  buf
  g36
  (
    n76,
    n6
  );


  buf
  g37
  (
    n67,
    n8
  );


  buf
  g38
  (
    n68,
    n15
  );


  buf
  g39
  (
    n48,
    n24
  );


  not
  g40
  (
    n49,
    n11
  );


  not
  g41
  (
    n54,
    n9
  );


  not
  g42
  (
    n35,
    n19
  );


  buf
  g43
  (
    n34,
    n18
  );


  buf
  g44
  (
    n73,
    n6
  );


  not
  g45
  (
    n69,
    n5
  );


  not
  g46
  (
    n55,
    n15
  );


  not
  g47
  (
    n96,
    n9
  );


  not
  g48
  (
    n98,
    n20
  );


  not
  g49
  (
    n116,
    n14
  );


  buf
  g50
  (
    n36,
    n19
  );


  buf
  g51
  (
    n64,
    n23
  );


  buf
  g52
  (
    n103,
    n14
  );


  buf
  g53
  (
    n44,
    n22
  );


  not
  g54
  (
    n45,
    n4
  );


  buf
  g55
  (
    n95,
    n21
  );


  buf
  g56
  (
    n50,
    n12
  );


  buf
  g57
  (
    n29,
    n1
  );


  buf
  g58
  (
    n60,
    n15
  );


  not
  g59
  (
    n106,
    n2
  );


  not
  g60
  (
    n59,
    n11
  );


  not
  g61
  (
    n61,
    n18
  );


  not
  g62
  (
    n119,
    n4
  );


  not
  g63
  (
    n41,
    n18
  );


  not
  g64
  (
    n80,
    n23
  );


  not
  g65
  (
    n114,
    n1
  );


  buf
  g66
  (
    n120,
    n17
  );


  not
  g67
  (
    n89,
    n2
  );


  not
  g68
  (
    n97,
    n5
  );


  not
  g69
  (
    n46,
    n20
  );


  buf
  g70
  (
    n47,
    n11
  );


  not
  g71
  (
    n79,
    n24
  );


  not
  g72
  (
    n63,
    n23
  );


  buf
  g73
  (
    n28,
    n2
  );


  buf
  g74
  (
    n70,
    n8
  );


  buf
  g75
  (
    n33,
    n21
  );


  not
  g76
  (
    n85,
    n10
  );


  not
  g77
  (
    n74,
    n17
  );


  not
  g78
  (
    n52,
    n12
  );


  not
  g79
  (
    n104,
    n3
  );


  not
  g80
  (
    n105,
    n7
  );


  buf
  g81
  (
    n90,
    n22
  );


  not
  g82
  (
    n101,
    n9
  );


  buf
  g83
  (
    n100,
    n7
  );


  not
  g84
  (
    n99,
    n1
  );


  buf
  g85
  (
    n117,
    n16
  );


  not
  g86
  (
    n72,
    n24
  );


  buf
  g87
  (
    n93,
    n3
  );


  not
  g88
  (
    n30,
    n19
  );


  not
  g89
  (
    n86,
    n14
  );


  not
  g90
  (
    n118,
    n13
  );


  not
  g91
  (
    n40,
    n20
  );


  not
  g92
  (
    n78,
    n16
  );


  not
  g93
  (
    n32,
    n14
  );


  buf
  g94
  (
    n37,
    n21
  );


  not
  g95
  (
    n38,
    n23
  );


  not
  g96
  (
    n325,
    n38
  );


  not
  g97
  (
    n403,
    n76
  );


  not
  g98
  (
    n341,
    n94
  );


  buf
  g99
  (
    n273,
    n43
  );


  buf
  g100
  (
    n245,
    n28
  );


  buf
  g101
  (
    n329,
    n84
  );


  buf
  g102
  (
    n494,
    n44
  );


  buf
  g103
  (
    n489,
    n112
  );


  not
  g104
  (
    n217,
    n97
  );


  not
  g105
  (
    n306,
    n104
  );


  not
  g106
  (
    n254,
    n103
  );


  not
  g107
  (
    n274,
    n38
  );


  buf
  g108
  (
    n130,
    n111
  );


  buf
  g109
  (
    n263,
    n57
  );


  buf
  g110
  (
    n491,
    n35
  );


  not
  g111
  (
    n169,
    n53
  );


  buf
  g112
  (
    n294,
    n118
  );


  not
  g113
  (
    n474,
    n81
  );


  not
  g114
  (
    n370,
    n109
  );


  buf
  g115
  (
    n173,
    n39
  );


  buf
  g116
  (
    n218,
    n75
  );


  buf
  g117
  (
    n326,
    n75
  );


  not
  g118
  (
    n439,
    n43
  );


  not
  g119
  (
    n487,
    n102
  );


  not
  g120
  (
    n163,
    n116
  );


  buf
  g121
  (
    n456,
    n61
  );


  buf
  g122
  (
    n412,
    n64
  );


  not
  g123
  (
    n414,
    n62
  );


  buf
  g124
  (
    n238,
    n30
  );


  buf
  g125
  (
    n209,
    n74
  );


  not
  g126
  (
    n242,
    n62
  );


  not
  g127
  (
    n480,
    n52
  );


  not
  g128
  (
    n157,
    n26
  );


  not
  g129
  (
    n321,
    n102
  );


  not
  g130
  (
    n335,
    n90
  );


  buf
  g131
  (
    n285,
    n119
  );


  buf
  g132
  (
    n477,
    n81
  );


  not
  g133
  (
    n195,
    n90
  );


  not
  g134
  (
    n388,
    n77
  );


  not
  g135
  (
    n427,
    n70
  );


  not
  g136
  (
    n303,
    n83
  );


  buf
  g137
  (
    n444,
    n95
  );


  buf
  g138
  (
    n164,
    n30
  );


  not
  g139
  (
    n215,
    n104
  );


  not
  g140
  (
    n284,
    n29
  );


  not
  g141
  (
    n255,
    n49
  );


  buf
  g142
  (
    n280,
    n35
  );


  not
  g143
  (
    n183,
    n58
  );


  buf
  g144
  (
    n333,
    n114
  );


  buf
  g145
  (
    n213,
    n25
  );


  not
  g146
  (
    n424,
    n56
  );


  buf
  g147
  (
    n438,
    n113
  );


  buf
  g148
  (
    n385,
    n60
  );


  buf
  g149
  (
    n249,
    n91
  );


  buf
  g150
  (
    n353,
    n116
  );


  not
  g151
  (
    n348,
    n103
  );


  not
  g152
  (
    n181,
    n80
  );


  buf
  g153
  (
    n441,
    n64
  );


  buf
  g154
  (
    n401,
    n55
  );


  buf
  g155
  (
    n208,
    n112
  );


  buf
  g156
  (
    n143,
    n80
  );


  not
  g157
  (
    n283,
    n93
  );


  not
  g158
  (
    n276,
    n40
  );


  not
  g159
  (
    n132,
    n76
  );


  buf
  g160
  (
    n172,
    n28
  );


  buf
  g161
  (
    n257,
    n48
  );


  buf
  g162
  (
    n162,
    n65
  );


  not
  g163
  (
    n498,
    n72
  );


  not
  g164
  (
    n150,
    n90
  );


  buf
  g165
  (
    n449,
    n73
  );


  buf
  g166
  (
    n394,
    n81
  );


  buf
  g167
  (
    n154,
    n55
  );


  not
  g168
  (
    n379,
    n92
  );


  buf
  g169
  (
    n200,
    n73
  );


  buf
  g170
  (
    n368,
    n63
  );


  buf
  g171
  (
    n500,
    n62
  );


  buf
  g172
  (
    n442,
    n76
  );


  not
  g173
  (
    n302,
    n46
  );


  buf
  g174
  (
    n259,
    n93
  );


  not
  g175
  (
    n211,
    n31
  );


  buf
  g176
  (
    n453,
    n94
  );


  not
  g177
  (
    n359,
    n92
  );


  not
  g178
  (
    n278,
    n72
  );


  not
  g179
  (
    n380,
    n45
  );


  buf
  g180
  (
    n387,
    n31
  );


  buf
  g181
  (
    n476,
    n101
  );


  not
  g182
  (
    n247,
    n113
  );


  not
  g183
  (
    n346,
    n85
  );


  buf
  g184
  (
    n457,
    n86
  );


  not
  g185
  (
    n466,
    n71
  );


  buf
  g186
  (
    n133,
    n75
  );


  buf
  g187
  (
    n499,
    n117
  );


  not
  g188
  (
    n275,
    n82
  );


  not
  g189
  (
    n431,
    n119
  );


  not
  g190
  (
    n330,
    n114
  );


  buf
  g191
  (
    n471,
    n76
  );


  buf
  g192
  (
    n377,
    n118
  );


  buf
  g193
  (
    n134,
    n29
  );


  not
  g194
  (
    n309,
    n41
  );


  buf
  g195
  (
    n131,
    n114
  );


  not
  g196
  (
    n482,
    n73
  );


  buf
  g197
  (
    n365,
    n26
  );


  not
  g198
  (
    n324,
    n53
  );


  buf
  g199
  (
    n409,
    n40
  );


  buf
  g200
  (
    n297,
    n42
  );


  not
  g201
  (
    n318,
    n94
  );


  buf
  g202
  (
    n234,
    n66
  );


  buf
  g203
  (
    n479,
    n78
  );


  buf
  g204
  (
    n415,
    n98
  );


  buf
  g205
  (
    n239,
    n27
  );


  buf
  g206
  (
    n354,
    n118
  );


  buf
  g207
  (
    n250,
    n49
  );


  buf
  g208
  (
    n188,
    n65
  );


  buf
  g209
  (
    n372,
    n62
  );


  buf
  g210
  (
    n138,
    n88
  );


  buf
  g211
  (
    n436,
    n44
  );


  buf
  g212
  (
    n216,
    n98
  );


  buf
  g213
  (
    n452,
    n97
  );


  buf
  g214
  (
    n266,
    n106
  );


  not
  g215
  (
    n233,
    n73
  );


  buf
  g216
  (
    n166,
    n116
  );


  not
  g217
  (
    n147,
    n71
  );


  not
  g218
  (
    n224,
    n43
  );


  not
  g219
  (
    n434,
    n47
  );


  buf
  g220
  (
    n139,
    n117
  );


  buf
  g221
  (
    n296,
    n32
  );


  not
  g222
  (
    n363,
    n34
  );


  buf
  g223
  (
    n121,
    n111
  );


  not
  g224
  (
    n458,
    n70
  );


  buf
  g225
  (
    n271,
    n79
  );


  not
  g226
  (
    n504,
    n69
  );


  buf
  g227
  (
    n190,
    n89
  );


  not
  g228
  (
    n417,
    n119
  );


  not
  g229
  (
    n338,
    n86
  );


  not
  g230
  (
    n270,
    n72
  );


  buf
  g231
  (
    n393,
    n105
  );


  buf
  g232
  (
    n300,
    n59
  );


  not
  g233
  (
    n191,
    n104
  );


  not
  g234
  (
    n165,
    n37
  );


  buf
  g235
  (
    n155,
    n59
  );


  buf
  g236
  (
    n290,
    n110
  );


  not
  g237
  (
    n142,
    n79
  );


  not
  g238
  (
    n305,
    n107
  );


  not
  g239
  (
    n397,
    n25
  );


  buf
  g240
  (
    n287,
    n84
  );


  not
  g241
  (
    n194,
    n93
  );


  buf
  g242
  (
    n148,
    n51
  );


  not
  g243
  (
    n376,
    n45
  );


  not
  g244
  (
    n501,
    n110
  );


  buf
  g245
  (
    n136,
    n54
  );


  not
  g246
  (
    n223,
    n50
  );


  not
  g247
  (
    n192,
    n116
  );


  buf
  g248
  (
    n310,
    n91
  );


  not
  g249
  (
    n299,
    n58
  );


  not
  g250
  (
    n327,
    n27
  );


  not
  g251
  (
    n472,
    n39
  );


  not
  g252
  (
    n288,
    n50
  );


  not
  g253
  (
    n177,
    n87
  );


  not
  g254
  (
    n315,
    n78
  );


  buf
  g255
  (
    n492,
    n92
  );


  buf
  g256
  (
    n135,
    n44
  );


  buf
  g257
  (
    KeyWire_0_8,
    n30
  );


  buf
  g258
  (
    n146,
    n102
  );


  not
  g259
  (
    n381,
    n25
  );


  not
  g260
  (
    n448,
    n114
  );


  not
  g261
  (
    n465,
    n78
  );


  not
  g262
  (
    n337,
    n52
  );


  buf
  g263
  (
    n360,
    n42
  );


  not
  g264
  (
    n314,
    n91
  );


  not
  g265
  (
    n352,
    n60
  );


  buf
  g266
  (
    n289,
    n45
  );


  not
  g267
  (
    n202,
    n106
  );


  buf
  g268
  (
    n189,
    n36
  );


  not
  g269
  (
    n214,
    n42
  );


  buf
  g270
  (
    n186,
    n101
  );


  buf
  g271
  (
    n496,
    n49
  );


  not
  g272
  (
    n295,
    n82
  );


  buf
  g273
  (
    n124,
    n34
  );


  buf
  g274
  (
    n356,
    n86
  );


  not
  g275
  (
    n235,
    n115
  );


  buf
  g276
  (
    n272,
    n36
  );


  buf
  g277
  (
    n432,
    n79
  );


  buf
  g278
  (
    n320,
    n67
  );


  not
  g279
  (
    n460,
    n108
  );


  not
  g280
  (
    n367,
    n46
  );


  not
  g281
  (
    n246,
    n98
  );


  buf
  g282
  (
    n405,
    n68
  );


  not
  g283
  (
    n237,
    n58
  );


  buf
  g284
  (
    n170,
    n37
  );


  not
  g285
  (
    n265,
    n55
  );


  not
  g286
  (
    n451,
    n66
  );


  not
  g287
  (
    n248,
    n86
  );


  not
  g288
  (
    KeyWire_0_12,
    n99
  );


  not
  g289
  (
    n470,
    n87
  );


  buf
  g290
  (
    n410,
    n80
  );


  not
  g291
  (
    n229,
    n83
  );


  not
  g292
  (
    n332,
    n56
  );


  not
  g293
  (
    n425,
    n110
  );


  not
  g294
  (
    n362,
    n41
  );


  not
  g295
  (
    n286,
    n44
  );


  buf
  g296
  (
    n334,
    n53
  );


  not
  g297
  (
    n389,
    n94
  );


  buf
  g298
  (
    n343,
    n61
  );


  not
  g299
  (
    n339,
    n31
  );


  buf
  g300
  (
    n316,
    n80
  );


  buf
  g301
  (
    n311,
    n50
  );


  not
  g302
  (
    n323,
    n38
  );


  buf
  g303
  (
    n167,
    n34
  );


  buf
  g304
  (
    n437,
    n77
  );


  not
  g305
  (
    n252,
    n70
  );


  not
  g306
  (
    n407,
    n63
  );


  buf
  g307
  (
    n391,
    n115
  );


  not
  g308
  (
    n502,
    n85
  );


  not
  g309
  (
    n123,
    n112
  );


  not
  g310
  (
    n402,
    n26
  );


  not
  g311
  (
    n301,
    n31
  );


  not
  g312
  (
    n307,
    n45
  );


  buf
  g313
  (
    n404,
    n46
  );


  not
  g314
  (
    n382,
    n104
  );


  buf
  g315
  (
    n198,
    n92
  );


  buf
  g316
  (
    n464,
    n47
  );


  not
  g317
  (
    n225,
    n95
  );


  buf
  g318
  (
    n390,
    n89
  );


  buf
  g319
  (
    n291,
    n60
  );


  buf
  g320
  (
    n406,
    n33
  );


  buf
  g321
  (
    n197,
    n108
  );


  buf
  g322
  (
    n468,
    n110
  );


  buf
  g323
  (
    n473,
    n42
  );


  not
  g324
  (
    n201,
    n60
  );


  not
  g325
  (
    n145,
    n109
  );


  not
  g326
  (
    n293,
    n67
  );


  not
  g327
  (
    n160,
    n95
  );


  buf
  g328
  (
    n171,
    n35
  );


  not
  g329
  (
    n268,
    n65
  );


  not
  g330
  (
    n207,
    n81
  );


  buf
  g331
  (
    n319,
    n35
  );


  buf
  g332
  (
    n433,
    n83
  );


  not
  g333
  (
    n454,
    n47
  );


  not
  g334
  (
    n219,
    n33
  );


  buf
  g335
  (
    n484,
    n27
  );


  not
  g336
  (
    n205,
    n68
  );


  buf
  g337
  (
    n446,
    n106
  );


  not
  g338
  (
    n261,
    n41
  );


  not
  g339
  (
    n440,
    n49
  );


  not
  g340
  (
    n374,
    n59
  );


  not
  g341
  (
    n344,
    n100
  );


  not
  g342
  (
    n149,
    n108
  );


  buf
  g343
  (
    n450,
    n57
  );


  not
  g344
  (
    n351,
    n82
  );


  buf
  g345
  (
    n340,
    n87
  );


  buf
  g346
  (
    n418,
    n37
  );


  buf
  g347
  (
    n408,
    n88
  );


  not
  g348
  (
    n462,
    n120
  );


  not
  g349
  (
    n153,
    n109
  );


  buf
  g350
  (
    n445,
    n61
  );


  buf
  g351
  (
    n336,
    n101
  );


  buf
  g352
  (
    n369,
    n67
  );


  not
  g353
  (
    n262,
    n98
  );


  buf
  g354
  (
    n140,
    n89
  );


  buf
  g355
  (
    n384,
    n105
  );


  buf
  g356
  (
    n258,
    n70
  );


  not
  g357
  (
    n375,
    n43
  );


  buf
  g358
  (
    n308,
    n118
  );


  not
  g359
  (
    n358,
    n39
  );


  not
  g360
  (
    n227,
    n102
  );


  buf
  g361
  (
    n361,
    n96
  );


  not
  g362
  (
    n357,
    n107
  );


  not
  g363
  (
    n331,
    n26
  );


  buf
  g364
  (
    n256,
    n107
  );


  not
  g365
  (
    n159,
    n103
  );


  buf
  g366
  (
    n423,
    n99
  );


  not
  g367
  (
    n490,
    n54
  );


  not
  g368
  (
    n313,
    n32
  );


  buf
  g369
  (
    n222,
    n113
  );


  buf
  g370
  (
    n420,
    n41
  );


  buf
  g371
  (
    n399,
    n100
  );


  buf
  g372
  (
    n503,
    n119
  );


  not
  g373
  (
    n350,
    n112
  );


  buf
  g374
  (
    n126,
    n88
  );


  buf
  g375
  (
    n125,
    n71
  );


  buf
  g376
  (
    n174,
    n74
  );


  buf
  g377
  (
    n364,
    n75
  );


  buf
  g378
  (
    n244,
    n97
  );


  buf
  g379
  (
    n144,
    n99
  );


  not
  g380
  (
    n430,
    n77
  );


  buf
  g381
  (
    n253,
    n95
  );


  not
  g382
  (
    n179,
    n34
  );


  buf
  g383
  (
    n228,
    n83
  );


  buf
  g384
  (
    n241,
    n38
  );


  buf
  g385
  (
    n232,
    n63
  );


  buf
  g386
  (
    n260,
    n117
  );


  not
  g387
  (
    n212,
    n56
  );


  buf
  g388
  (
    n429,
    n48
  );


  buf
  g389
  (
    n282,
    n51
  );


  not
  g390
  (
    n355,
    n66
  );


  buf
  g391
  (
    n467,
    n40
  );


  buf
  g392
  (
    n317,
    n120
  );


  not
  g393
  (
    n196,
    n69
  );


  not
  g394
  (
    n269,
    n107
  );


  buf
  g395
  (
    n137,
    n30
  );


  buf
  g396
  (
    n497,
    n68
  );


  buf
  g397
  (
    n184,
    n111
  );


  not
  g398
  (
    n495,
    n109
  );


  buf
  g399
  (
    n127,
    n36
  );


  not
  g400
  (
    n463,
    n51
  );


  not
  g401
  (
    n396,
    n100
  );


  not
  g402
  (
    n312,
    n57
  );


  not
  g403
  (
    n151,
    n55
  );


  buf
  g404
  (
    n478,
    n33
  );


  not
  g405
  (
    n426,
    n33
  );


  not
  g406
  (
    n230,
    n85
  );


  not
  g407
  (
    n413,
    n93
  );


  not
  g408
  (
    n328,
    n29
  );


  buf
  g409
  (
    n231,
    n66
  );


  not
  g410
  (
    n292,
    n56
  );


  buf
  g411
  (
    n180,
    n48
  );


  not
  g412
  (
    n488,
    n39
  );


  buf
  g413
  (
    n203,
    n89
  );


  buf
  g414
  (
    n243,
    n84
  );


  not
  g415
  (
    n378,
    n105
  );


  not
  g416
  (
    n416,
    n72
  );


  buf
  g417
  (
    n304,
    n54
  );


  buf
  g418
  (
    n371,
    n91
  );


  buf
  g419
  (
    n277,
    n25
  );


  not
  g420
  (
    n267,
    n90
  );


  not
  g421
  (
    n156,
    n36
  );


  buf
  g422
  (
    n141,
    n111
  );


  not
  g423
  (
    n236,
    n46
  );


  buf
  g424
  (
    n193,
    n50
  );


  not
  g425
  (
    n128,
    n52
  );


  not
  g426
  (
    n455,
    n28
  );


  buf
  g427
  (
    n176,
    n40
  );


  not
  g428
  (
    n347,
    n113
  );


  not
  g429
  (
    n373,
    n78
  );


  buf
  g430
  (
    n158,
    n99
  );


  not
  g431
  (
    n168,
    n88
  );


  buf
  g432
  (
    n422,
    n82
  );


  buf
  g433
  (
    n461,
    n67
  );


  buf
  g434
  (
    n383,
    n48
  );


  not
  g435
  (
    n129,
    n87
  );


  not
  g436
  (
    n443,
    n103
  );


  buf
  g437
  (
    n481,
    n96
  );


  not
  g438
  (
    n349,
    n117
  );


  buf
  g439
  (
    n122,
    n47
  );


  not
  g440
  (
    n182,
    n68
  );


  buf
  g441
  (
    n226,
    n61
  );


  not
  g442
  (
    n459,
    n97
  );


  not
  g443
  (
    n322,
    n32
  );


  buf
  g444
  (
    n395,
    n85
  );


  not
  g445
  (
    n221,
    n84
  );


  not
  g446
  (
    n187,
    n69
  );


  buf
  g447
  (
    n486,
    n115
  );


  buf
  g448
  (
    n161,
    n29
  );


  not
  g449
  (
    n342,
    n27
  );


  buf
  g450
  (
    n428,
    n32
  );


  buf
  g451
  (
    n279,
    n96
  );


  buf
  g452
  (
    n152,
    n64
  );


  not
  g453
  (
    n185,
    n54
  );


  not
  g454
  (
    n483,
    n63
  );


  not
  g455
  (
    n493,
    n28
  );


  not
  g456
  (
    n298,
    n79
  );


  not
  g457
  (
    n220,
    n105
  );


  buf
  g458
  (
    n435,
    n115
  );


  buf
  g459
  (
    n485,
    n108
  );


  buf
  g460
  (
    n421,
    n69
  );


  not
  g461
  (
    n264,
    n57
  );


  not
  g462
  (
    n178,
    n96
  );


  buf
  g463
  (
    n366,
    n53
  );


  not
  g464
  (
    n206,
    n74
  );


  not
  g465
  (
    n175,
    n101
  );


  buf
  g466
  (
    n411,
    n65
  );


  not
  g467
  (
    n386,
    n77
  );


  not
  g468
  (
    n281,
    n106
  );


  buf
  g469
  (
    n251,
    n52
  );


  buf
  g470
  (
    n204,
    n74
  );


  buf
  g471
  (
    n199,
    n51
  );


  not
  g472
  (
    n419,
    n100
  );


  not
  g473
  (
    n475,
    n58
  );


  not
  g474
  (
    KeyWire_0_15,
    n71
  );


  buf
  g475
  (
    n398,
    n120
  );


  not
  g476
  (
    n210,
    n64
  );


  not
  g477
  (
    n345,
    n120
  );


  not
  g478
  (
    n400,
    n37
  );


  buf
  g479
  (
    n392,
    n59
  );


  buf
  g480
  (
    n1457,
    n264
  );


  not
  g481
  (
    n752,
    n393
  );


  not
  g482
  (
    n708,
    n494
  );


  not
  g483
  (
    n565,
    n312
  );


  buf
  g484
  (
    n1505,
    n350
  );


  buf
  g485
  (
    n615,
    n301
  );


  buf
  g486
  (
    n1232,
    n259
  );


  not
  g487
  (
    n1157,
    n351
  );


  not
  g488
  (
    n1191,
    n383
  );


  buf
  g489
  (
    n1299,
    n340
  );


  not
  g490
  (
    n748,
    n289
  );


  not
  g491
  (
    n1062,
    n292
  );


  buf
  g492
  (
    n1340,
    n474
  );


  buf
  g493
  (
    n511,
    n488
  );


  not
  g494
  (
    n508,
    n130
  );


  not
  g495
  (
    n843,
    n376
  );


  not
  g496
  (
    n1383,
    n342
  );


  not
  g497
  (
    n869,
    n179
  );


  buf
  g498
  (
    n854,
    n294
  );


  buf
  g499
  (
    n541,
    n333
  );


  buf
  g500
  (
    n1332,
    n467
  );


  not
  g501
  (
    n672,
    n317
  );


  not
  g502
  (
    n1251,
    n128
  );


  not
  g503
  (
    n912,
    n342
  );


  buf
  g504
  (
    n781,
    n381
  );


  not
  g505
  (
    n983,
    n256
  );


  buf
  g506
  (
    n1393,
    n310
  );


  not
  g507
  (
    n1360,
    n465
  );


  buf
  g508
  (
    n936,
    n443
  );


  buf
  g509
  (
    n1248,
    n385
  );


  buf
  g510
  (
    KeyWire_0_11,
    n263
  );


  buf
  g511
  (
    n665,
    n469
  );


  buf
  g512
  (
    n1249,
    n350
  );


  not
  g513
  (
    n522,
    n406
  );


  buf
  g514
  (
    n1305,
    n423
  );


  not
  g515
  (
    n1229,
    n456
  );


  not
  g516
  (
    n1322,
    n151
  );


  not
  g517
  (
    n1485,
    n424
  );


  buf
  g518
  (
    n580,
    n437
  );


  buf
  g519
  (
    n635,
    n466
  );


  not
  g520
  (
    n1370,
    n471
  );


  buf
  g521
  (
    n1483,
    n451
  );


  buf
  g522
  (
    n772,
    n408
  );


  buf
  g523
  (
    n518,
    n275
  );


  not
  g524
  (
    n990,
    n234
  );


  not
  g525
  (
    n825,
    n429
  );


  not
  g526
  (
    n571,
    n364
  );


  buf
  g527
  (
    n1087,
    n209
  );


  buf
  g528
  (
    n1074,
    n354
  );


  buf
  g529
  (
    n584,
    n394
  );


  buf
  g530
  (
    n757,
    n482
  );


  buf
  g531
  (
    n1186,
    n480
  );


  not
  g532
  (
    n1412,
    n482
  );


  not
  g533
  (
    n882,
    n447
  );


  not
  g534
  (
    n1467,
    n446
  );


  not
  g535
  (
    n1306,
    n501
  );


  not
  g536
  (
    n600,
    n319
  );


  not
  g537
  (
    n529,
    n241
  );


  buf
  g538
  (
    n714,
    n460
  );


  buf
  g539
  (
    n850,
    n445
  );


  not
  g540
  (
    n563,
    n399
  );


  buf
  g541
  (
    n1314,
    n377
  );


  buf
  g542
  (
    n634,
    n427
  );


  buf
  g543
  (
    n703,
    n375
  );


  not
  g544
  (
    n1390,
    n353
  );


  buf
  g545
  (
    n1091,
    n408
  );


  not
  g546
  (
    n723,
    n437
  );


  buf
  g547
  (
    n999,
    n329
  );


  not
  g548
  (
    n1446,
    n387
  );


  buf
  g549
  (
    n1101,
    n491
  );


  not
  g550
  (
    n670,
    n387
  );


  buf
  g551
  (
    n1416,
    n281
  );


  not
  g552
  (
    n1280,
    n418
  );


  not
  g553
  (
    n778,
    n325
  );


  buf
  g554
  (
    n1086,
    n481
  );


  buf
  g555
  (
    n728,
    n356
  );


  buf
  g556
  (
    n819,
    n431
  );


  not
  g557
  (
    n1272,
    n321
  );


  buf
  g558
  (
    n606,
    n292
  );


  not
  g559
  (
    n1085,
    n215
  );


  buf
  g560
  (
    n1391,
    n286
  );


  buf
  g561
  (
    n840,
    n395
  );


  buf
  g562
  (
    n1207,
    n377
  );


  not
  g563
  (
    n1313,
    n323
  );


  buf
  g564
  (
    n1113,
    n444
  );


  not
  g565
  (
    n726,
    n383
  );


  not
  g566
  (
    n835,
    n364
  );


  buf
  g567
  (
    n839,
    n392
  );


  not
  g568
  (
    n1481,
    n452
  );


  buf
  g569
  (
    n924,
    n400
  );


  buf
  g570
  (
    n797,
    n478
  );


  buf
  g571
  (
    n1204,
    n419
  );


  buf
  g572
  (
    n1065,
    n263
  );


  buf
  g573
  (
    n1286,
    n492
  );


  not
  g574
  (
    n833,
    n396
  );


  not
  g575
  (
    n521,
    n492
  );


  not
  g576
  (
    n1339,
    n444
  );


  not
  g577
  (
    n675,
    n193
  );


  not
  g578
  (
    n842,
    n489
  );


  buf
  g579
  (
    n881,
    n415
  );


  not
  g580
  (
    n1298,
    n361
  );


  not
  g581
  (
    n964,
    n291
  );


  not
  g582
  (
    n765,
    n423
  );


  not
  g583
  (
    n1169,
    n240
  );


  buf
  g584
  (
    n1119,
    n440
  );


  buf
  g585
  (
    n1364,
    n185
  );


  not
  g586
  (
    n857,
    n317
  );


  not
  g587
  (
    n805,
    n455
  );


  not
  g588
  (
    n785,
    n413
  );


  buf
  g589
  (
    n1459,
    n302
  );


  not
  g590
  (
    n1429,
    n433
  );


  buf
  g591
  (
    n908,
    n479
  );


  not
  g592
  (
    n810,
    n157
  );


  buf
  g593
  (
    n1092,
    n429
  );


  buf
  g594
  (
    n1203,
    n412
  );


  buf
  g595
  (
    n1037,
    n359
  );


  buf
  g596
  (
    n1419,
    n345
  );


  buf
  g597
  (
    n1475,
    n484
  );


  not
  g598
  (
    n760,
    n160
  );


  buf
  g599
  (
    n952,
    n423
  );


  buf
  g600
  (
    n716,
    n334
  );


  not
  g601
  (
    n1441,
    n372
  );


  buf
  g602
  (
    n1294,
    n385
  );


  not
  g603
  (
    n1060,
    n335
  );


  not
  g604
  (
    n1077,
    n388
  );


  not
  g605
  (
    n1123,
    n462
  );


  buf
  g606
  (
    n1316,
    n439
  );


  not
  g607
  (
    n687,
    n404
  );


  not
  g608
  (
    n1010,
    n283
  );


  buf
  g609
  (
    n864,
    n368
  );


  buf
  g610
  (
    n1323,
    n461
  );


  buf
  g611
  (
    n861,
    n483
  );


  buf
  g612
  (
    n662,
    n421
  );


  not
  g613
  (
    n986,
    n330
  );


  not
  g614
  (
    n1342,
    n389
  );


  not
  g615
  (
    n627,
    n475
  );


  buf
  g616
  (
    n533,
    n437
  );


  buf
  g617
  (
    n923,
    n323
  );


  not
  g618
  (
    n1240,
    n259
  );


  buf
  g619
  (
    n866,
    n498
  );


  not
  g620
  (
    n1428,
    n373
  );


  buf
  g621
  (
    n1219,
    n217
  );


  not
  g622
  (
    n1082,
    n453
  );


  buf
  g623
  (
    n1224,
    n224
  );


  not
  g624
  (
    n743,
    n341
  );


  buf
  g625
  (
    n815,
    n370
  );


  buf
  g626
  (
    n622,
    n496
  );


  not
  g627
  (
    n910,
    n322
  );


  buf
  g628
  (
    n1254,
    n330
  );


  not
  g629
  (
    n652,
    n347
  );


  not
  g630
  (
    n595,
    n170
  );


  not
  g631
  (
    n931,
    n353
  );


  not
  g632
  (
    n1255,
    n290
  );


  not
  g633
  (
    n1466,
    n147
  );


  not
  g634
  (
    n1252,
    n421
  );


  not
  g635
  (
    n1501,
    n401
  );


  not
  g636
  (
    n1084,
    n377
  );


  not
  g637
  (
    n1405,
    n142
  );


  buf
  g638
  (
    n1182,
    n296
  );


  buf
  g639
  (
    n1263,
    n322
  );


  buf
  g640
  (
    n664,
    n278
  );


  not
  g641
  (
    n1041,
    n471
  );


  buf
  g642
  (
    n896,
    n307
  );


  not
  g643
  (
    n1433,
    n330
  );


  not
  g644
  (
    n1451,
    n247
  );


  not
  g645
  (
    n1357,
    n267
  );


  buf
  g646
  (
    n871,
    n454
  );


  not
  g647
  (
    n1129,
    n416
  );


  not
  g648
  (
    n1435,
    n417
  );


  buf
  g649
  (
    n526,
    n171
  );


  buf
  g650
  (
    n996,
    n321
  );


  buf
  g651
  (
    n736,
    n484
  );


  not
  g652
  (
    n1490,
    n367
  );


  not
  g653
  (
    n1345,
    n249
  );


  buf
  g654
  (
    n700,
    n479
  );


  buf
  g655
  (
    n1161,
    n406
  );


  buf
  g656
  (
    n1019,
    n500
  );


  not
  g657
  (
    n1328,
    n493
  );


  buf
  g658
  (
    n775,
    n320
  );


  not
  g659
  (
    n527,
    n331
  );


  buf
  g660
  (
    n582,
    n441
  );


  not
  g661
  (
    n1381,
    n260
  );


  buf
  g662
  (
    n1278,
    n149
  );


  not
  g663
  (
    n1126,
    n477
  );


  buf
  g664
  (
    n913,
    n373
  );


  not
  g665
  (
    n1284,
    n355
  );


  not
  g666
  (
    n520,
    n493
  );


  not
  g667
  (
    n1422,
    n267
  );


  buf
  g668
  (
    n1333,
    n424
  );


  not
  g669
  (
    n1190,
    n464
  );


  buf
  g670
  (
    n509,
    n475
  );


  buf
  g671
  (
    n1478,
    n295
  );


  not
  g672
  (
    n786,
    n137
  );


  buf
  g673
  (
    n735,
    n284
  );


  not
  g674
  (
    n940,
    n313
  );


  not
  g675
  (
    n1162,
    n470
  );


  not
  g676
  (
    n570,
    n439
  );


  buf
  g677
  (
    n616,
    n362
  );


  buf
  g678
  (
    n1373,
    n359
  );


  not
  g679
  (
    n1209,
    n140
  );


  not
  g680
  (
    n1355,
    n343
  );


  buf
  g681
  (
    n1424,
    n449
  );


  not
  g682
  (
    n1470,
    n452
  );


  not
  g683
  (
    n1235,
    n308
  );


  buf
  g684
  (
    n771,
    n343
  );


  not
  g685
  (
    n713,
    n262
  );


  not
  g686
  (
    n1035,
    n405
  );


  buf
  g687
  (
    n1138,
    n202
  );


  buf
  g688
  (
    n645,
    n169
  );


  not
  g689
  (
    n588,
    n475
  );


  not
  g690
  (
    n1260,
    n298
  );


  not
  g691
  (
    n1257,
    n333
  );


  not
  g692
  (
    n979,
    n289
  );


  buf
  g693
  (
    n1013,
    n435
  );


  not
  g694
  (
    n1135,
    n354
  );


  not
  g695
  (
    n1301,
    n466
  );


  buf
  g696
  (
    n995,
    n268
  );


  not
  g697
  (
    n1474,
    n474
  );


  buf
  g698
  (
    n1315,
    n488
  );


  not
  g699
  (
    n1011,
    n466
  );


  buf
  g700
  (
    n980,
    n274
  );


  buf
  g701
  (
    n697,
    n253
  );


  buf
  g702
  (
    n558,
    n349
  );


  not
  g703
  (
    n516,
    n332
  );


  buf
  g704
  (
    n614,
    n153
  );


  buf
  g705
  (
    n1137,
    n317
  );


  buf
  g706
  (
    n578,
    n425
  );


  buf
  g707
  (
    n812,
    n428
  );


  not
  g708
  (
    n613,
    n404
  );


  not
  g709
  (
    n653,
    n390
  );


  not
  g710
  (
    n1024,
    n456
  );


  not
  g711
  (
    n639,
    n383
  );


  buf
  g712
  (
    n788,
    n198
  );


  buf
  g713
  (
    n1494,
    n374
  );


  buf
  g714
  (
    n1185,
    n380
  );


  not
  g715
  (
    n911,
    n381
  );


  not
  g716
  (
    n1023,
    n463
  );


  buf
  g717
  (
    n655,
    n338
  );


  buf
  g718
  (
    n970,
    n319
  );


  not
  g719
  (
    n1281,
    n464
  );


  buf
  g720
  (
    n1008,
    n408
  );


  not
  g721
  (
    n566,
    n316
  );


  not
  g722
  (
    n1063,
    n369
  );


  not
  g723
  (
    n814,
    n220
  );


  buf
  g724
  (
    n961,
    n341
  );


  buf
  g725
  (
    n1165,
    n405
  );


  not
  g726
  (
    n1144,
    n489
  );


  not
  g727
  (
    n685,
    n370
  );


  not
  g728
  (
    n965,
    n410
  );


  not
  g729
  (
    n1443,
    n489
  );


  buf
  g730
  (
    n998,
    n490
  );


  buf
  g731
  (
    n1398,
    n348
  );


  not
  g732
  (
    n873,
    n393
  );


  buf
  g733
  (
    n532,
    n380
  );


  not
  g734
  (
    n1052,
    n266
  );


  not
  g735
  (
    n676,
    n456
  );


  not
  g736
  (
    n1308,
    n385
  );


  not
  g737
  (
    n690,
    n189
  );


  buf
  g738
  (
    n804,
    n311
  );


  not
  g739
  (
    n1425,
    n424
  );


  not
  g740
  (
    n1427,
    n148
  );


  buf
  g741
  (
    n702,
    n368
  );


  buf
  g742
  (
    n1468,
    n339
  );


  buf
  g743
  (
    n663,
    n264
  );


  not
  g744
  (
    n1044,
    n452
  );


  not
  g745
  (
    n1034,
    n391
  );


  not
  g746
  (
    n1214,
    n326
  );


  buf
  g747
  (
    n1226,
    n334
  );


  buf
  g748
  (
    n929,
    n458
  );


  not
  g749
  (
    n1335,
    n244
  );


  buf
  g750
  (
    n783,
    n371
  );


  buf
  g751
  (
    n988,
    n428
  );


  buf
  g752
  (
    n954,
    n250
  );


  not
  g753
  (
    n1115,
    n485
  );


  not
  g754
  (
    n1033,
    n312
  );


  buf
  g755
  (
    n901,
    n303
  );


  not
  g756
  (
    n1070,
    n348
  );


  buf
  g757
  (
    n640,
    n360
  );


  buf
  g758
  (
    n773,
    n426
  );


  not
  g759
  (
    n1170,
    n499
  );


  buf
  g760
  (
    n678,
    n392
  );


  not
  g761
  (
    n1385,
    n255
  );


  not
  g762
  (
    n888,
    n407
  );


  buf
  g763
  (
    n811,
    n477
  );


  not
  g764
  (
    n969,
    n144
  );


  buf
  g765
  (
    n1192,
    n164
  );


  not
  g766
  (
    n1120,
    n388
  );


  not
  g767
  (
    n1319,
    n396
  );


  buf
  g768
  (
    n1334,
    n416
  );


  buf
  g769
  (
    n841,
    n486
  );


  buf
  g770
  (
    n691,
    n313
  );


  not
  g771
  (
    n1496,
    n427
  );


  not
  g772
  (
    n1031,
    n456
  );


  buf
  g773
  (
    n1206,
    n460
  );


  not
  g774
  (
    n1145,
    n444
  );


  not
  g775
  (
    n604,
    n440
  );


  buf
  g776
  (
    n682,
    n450
  );


  buf
  g777
  (
    n946,
    n439
  );


  not
  g778
  (
    n1488,
    n399
  );


  not
  g779
  (
    n883,
    n344
  );


  not
  g780
  (
    n801,
    n501
  );


  buf
  g781
  (
    n657,
    n428
  );


  not
  g782
  (
    n724,
    n474
  );


  not
  g783
  (
    n1463,
    n500
  );


  buf
  g784
  (
    n868,
    n361
  );


  not
  g785
  (
    n1358,
    n417
  );


  not
  g786
  (
    n1075,
    n210
  );


  buf
  g787
  (
    n766,
    n469
  );


  buf
  g788
  (
    n1142,
    n488
  );


  not
  g789
  (
    n1495,
    n238
  );


  not
  g790
  (
    n1017,
    n316
  );


  not
  g791
  (
    n1028,
    n192
  );


  buf
  g792
  (
    n1005,
    n411
  );


  not
  g793
  (
    n1230,
    n494
  );


  buf
  g794
  (
    n1406,
    n419
  );


  not
  g795
  (
    n1421,
    n346
  );


  buf
  g796
  (
    n513,
    n398
  );


  buf
  g797
  (
    n560,
    n251
  );


  buf
  g798
  (
    n1061,
    n222
  );


  buf
  g799
  (
    n696,
    n272
  );


  buf
  g800
  (
    n658,
    n419
  );


  not
  g801
  (
    n505,
    n480
  );


  not
  g802
  (
    n770,
    n188
  );


  not
  g803
  (
    n617,
    n434
  );


  buf
  g804
  (
    n1379,
    n254
  );


  buf
  g805
  (
    n802,
    n314
  );


  not
  g806
  (
    n1112,
    n414
  );


  buf
  g807
  (
    n1152,
    n409
  );


  buf
  g808
  (
    n1295,
    n122
  );


  not
  g809
  (
    n568,
    n333
  );


  not
  g810
  (
    n893,
    n334
  );


  not
  g811
  (
    n838,
    n281
  );


  not
  g812
  (
    n506,
    n299
  );


  not
  g813
  (
    n729,
    n257
  );


  not
  g814
  (
    n1050,
    n343
  );


  buf
  g815
  (
    n1304,
    n477
  );


  not
  g816
  (
    n987,
    n384
  );


  buf
  g817
  (
    n1256,
    n407
  );


  buf
  g818
  (
    n960,
    n494
  );


  not
  g819
  (
    n985,
    n366
  );


  not
  g820
  (
    n656,
    n333
  );


  not
  g821
  (
    n1200,
    n432
  );


  buf
  g822
  (
    KeyWire_0_10,
    n427
  );


  not
  g823
  (
    n895,
    n366
  );


  not
  g824
  (
    n1265,
    n325
  );


  not
  g825
  (
    n860,
    n351
  );


  not
  g826
  (
    n879,
    n138
  );


  not
  g827
  (
    n1109,
    n328
  );


  not
  g828
  (
    n1032,
    n290
  );


  not
  g829
  (
    n1016,
    n421
  );


  buf
  g830
  (
    n1154,
    n211
  );


  not
  g831
  (
    n1130,
    n397
  );


  buf
  g832
  (
    n1400,
    n296
  );


  not
  g833
  (
    n791,
    n481
  );


  not
  g834
  (
    n1282,
    n330
  );


  buf
  g835
  (
    n1343,
    n235
  );


  buf
  g836
  (
    n856,
    n465
  );


  not
  g837
  (
    n821,
    n448
  );


  not
  g838
  (
    n605,
    n277
  );


  buf
  g839
  (
    n799,
    n150
  );


  not
  g840
  (
    n972,
    n285
  );


  buf
  g841
  (
    n1139,
    n325
  );


  not
  g842
  (
    n1363,
    n132
  );


  buf
  g843
  (
    n1489,
    n354
  );


  buf
  g844
  (
    n1477,
    n352
  );


  buf
  g845
  (
    n1458,
    n336
  );


  buf
  g846
  (
    n1246,
    n381
  );


  not
  g847
  (
    n603,
    n481
  );


  not
  g848
  (
    n1499,
    n406
  );


  buf
  g849
  (
    n612,
    n435
  );


  buf
  g850
  (
    n1199,
    n305
  );


  buf
  g851
  (
    n978,
    n323
  );


  buf
  g852
  (
    n755,
    n453
  );


  buf
  g853
  (
    n741,
    n390
  );


  buf
  g854
  (
    n1289,
    n177
  );


  not
  g855
  (
    n1197,
    n378
  );


  not
  g856
  (
    n1504,
    n464
  );


  not
  g857
  (
    n623,
    n369
  );


  buf
  g858
  (
    n1238,
    n476
  );


  not
  g859
  (
    n1158,
    n265
  );


  not
  g860
  (
    n1361,
    n339
  );


  buf
  g861
  (
    n1131,
    n125
  );


  not
  g862
  (
    n1059,
    n379
  );


  buf
  g863
  (
    n874,
    n403
  );


  buf
  g864
  (
    n669,
    n363
  );


  not
  g865
  (
    n631,
    n205
  );


  not
  g866
  (
    n1067,
    n360
  );


  not
  g867
  (
    n915,
    n397
  );


  not
  g868
  (
    n686,
    n288
  );


  buf
  g869
  (
    n539,
    n176
  );


  buf
  g870
  (
    n1114,
    n451
  );


  buf
  g871
  (
    n1321,
    n315
  );


  buf
  g872
  (
    n1069,
    n183
  );


  buf
  g873
  (
    n1237,
    n304
  );


  not
  g874
  (
    n547,
    n495
  );


  not
  g875
  (
    n1042,
    n344
  );


  not
  g876
  (
    n1015,
    n375
  );


  not
  g877
  (
    n1047,
    n477
  );


  buf
  g878
  (
    n1106,
    n399
  );


  buf
  g879
  (
    n1049,
    n501
  );


  not
  g880
  (
    n738,
    n450
  );


  not
  g881
  (
    n569,
    n442
  );


  buf
  g882
  (
    n920,
    n459
  );


  buf
  g883
  (
    n1409,
    n395
  );


  not
  g884
  (
    n737,
    n459
  );


  not
  g885
  (
    n1354,
    n214
  );


  not
  g886
  (
    n852,
    n445
  );


  buf
  g887
  (
    n746,
    n435
  );


  not
  g888
  (
    n897,
    n357
  );


  not
  g889
  (
    n1072,
    n458
  );


  buf
  g890
  (
    n1007,
    n390
  );


  not
  g891
  (
    n1057,
    n300
  );


  not
  g892
  (
    n1001,
    n401
  );


  buf
  g893
  (
    n1442,
    n233
  );


  not
  g894
  (
    n1507,
    n418
  );


  not
  g895
  (
    n1465,
    n500
  );


  not
  g896
  (
    n1148,
    n402
  );


  not
  g897
  (
    n646,
    n391
  );


  not
  g898
  (
    n1212,
    n152
  );


  not
  g899
  (
    n1183,
    n496
  );


  buf
  g900
  (
    n1222,
    n434
  );


  not
  g901
  (
    n1450,
    n232
  );


  buf
  g902
  (
    n848,
    n165
  );


  not
  g903
  (
    n902,
    n199
  );


  buf
  g904
  (
    n711,
    n374
  );


  not
  g905
  (
    n1436,
    n204
  );


  not
  g906
  (
    n875,
    n388
  );


  not
  g907
  (
    n1287,
    n316
  );


  buf
  g908
  (
    n894,
    n182
  );


  not
  g909
  (
    n1195,
    n306
  );


  buf
  g910
  (
    n1432,
    n203
  );


  not
  g911
  (
    n1193,
    n186
  );


  buf
  g912
  (
    n878,
    n317
  );


  buf
  g913
  (
    n1160,
    n410
  );


  not
  g914
  (
    n706,
    n314
  );


  not
  g915
  (
    n769,
    n410
  );


  buf
  g916
  (
    n1388,
    n432
  );


  buf
  g917
  (
    n575,
    n390
  );


  buf
  g918
  (
    n628,
    n154
  );


  buf
  g919
  (
    n865,
    n401
  );


  buf
  g920
  (
    n777,
    n353
  );


  not
  g921
  (
    n886,
    n382
  );


  not
  g922
  (
    n948,
    n371
  );


  not
  g923
  (
    n763,
    n499
  );


  buf
  g924
  (
    n1121,
    n328
  );


  not
  g925
  (
    n644,
    n430
  );


  not
  g926
  (
    n794,
    n458
  );


  buf
  g927
  (
    n1125,
    n431
  );


  not
  g928
  (
    n1038,
    n442
  );


  not
  g929
  (
    n1384,
    n197
  );


  not
  g930
  (
    n780,
    n340
  );


  buf
  g931
  (
    n1132,
    n457
  );


  not
  g932
  (
    n1348,
    n380
  );


  buf
  g933
  (
    n1014,
    n467
  );


  not
  g934
  (
    n1320,
    n337
  );


  not
  g935
  (
    n984,
    n270
  );


  buf
  g936
  (
    n567,
    n393
  );


  not
  g937
  (
    n1056,
    n172
  );


  not
  g938
  (
    n1366,
    n268
  );


  not
  g939
  (
    n557,
    n196
  );


  buf
  g940
  (
    n592,
    n218
  );


  not
  g941
  (
    n722,
    n417
  );


  not
  g942
  (
    n1309,
    n438
  );


  not
  g943
  (
    n754,
    n293
  );


  buf
  g944
  (
    n699,
    n483
  );


  not
  g945
  (
    n1239,
    n162
  );


  not
  g946
  (
    n1133,
    n425
  );


  buf
  g947
  (
    n546,
    n369
  );


  buf
  g948
  (
    n884,
    n266
  );


  buf
  g949
  (
    n1410,
    n491
  );


  not
  g950
  (
    n1079,
    n472
  );


  not
  g951
  (
    n636,
    n321
  );


  buf
  g952
  (
    n621,
    n319
  );


  not
  g953
  (
    n930,
    n338
  );


  buf
  g954
  (
    n507,
    n365
  );


  buf
  g955
  (
    n1201,
    n407
  );


  buf
  g956
  (
    n1403,
    n490
  );


  buf
  g957
  (
    n932,
    n318
  );


  not
  g958
  (
    n1508,
    n353
  );


  buf
  g959
  (
    n1180,
    n404
  );


  not
  g960
  (
    n966,
    n363
  );


  not
  g961
  (
    n1434,
    n346
  );


  not
  g962
  (
    n651,
    n395
  );


  buf
  g963
  (
    n1156,
    n422
  );


  not
  g964
  (
    n826,
    n216
  );


  buf
  g965
  (
    n1486,
    n409
  );


  not
  g966
  (
    n1000,
    n256
  );


  not
  g967
  (
    n867,
    n190
  );


  buf
  g968
  (
    n967,
    n335
  );


  buf
  g969
  (
    n827,
    n282
  );


  buf
  g970
  (
    n1476,
    n382
  );


  buf
  g971
  (
    n762,
    n321
  );


  not
  g972
  (
    n750,
    n496
  );


  buf
  g973
  (
    n809,
    n449
  );


  buf
  g974
  (
    n749,
    n480
  );


  buf
  g975
  (
    n1324,
    n373
  );


  not
  g976
  (
    n997,
    n206
  );


  buf
  g977
  (
    n717,
    n476
  );


  not
  g978
  (
    n1150,
    n461
  );


  buf
  g979
  (
    n906,
    n271
  );


  not
  g980
  (
    n597,
    n414
  );


  buf
  g981
  (
    n1022,
    n406
  );


  buf
  g982
  (
    n916,
    n324
  );


  buf
  g983
  (
    n642,
    n397
  );


  not
  g984
  (
    n822,
    n422
  );


  not
  g985
  (
    n1211,
    n421
  );


  not
  g986
  (
    n937,
    n450
  );


  buf
  g987
  (
    n1374,
    n410
  );


  buf
  g988
  (
    n519,
    n404
  );


  buf
  g989
  (
    n1352,
    n426
  );


  not
  g990
  (
    n734,
    n397
  );


  buf
  g991
  (
    n1310,
    n403
  );


  buf
  g992
  (
    n1124,
    n415
  );


  not
  g993
  (
    n1068,
    n331
  );


  not
  g994
  (
    n1236,
    n443
  );


  not
  g995
  (
    n692,
    n229
  );


  not
  g996
  (
    n958,
    n417
  );


  not
  g997
  (
    n1234,
    n379
  );


  buf
  g998
  (
    n740,
    n441
  );


  not
  g999
  (
    n594,
    n207
  );


  buf
  g1000
  (
    n1274,
    n315
  );


  buf
  g1001
  (
    n1071,
    n327
  );


  not
  g1002
  (
    n1118,
    n212
  );


  not
  g1003
  (
    n1325,
    n492
  );


  buf
  g1004
  (
    n715,
    n476
  );


  not
  g1005
  (
    n1163,
    n302
  );


  not
  g1006
  (
    n554,
    n400
  );


  not
  g1007
  (
    n531,
    n258
  );


  not
  g1008
  (
    n514,
    n297
  );


  not
  g1009
  (
    n683,
    n376
  );


  buf
  g1010
  (
    n1009,
    n385
  );


  not
  g1011
  (
    n733,
    n391
  );


  not
  g1012
  (
    n1269,
    n398
  );


  not
  g1013
  (
    n1510,
    n320
  );


  buf
  g1014
  (
    n820,
    n420
  );


  not
  g1015
  (
    n1480,
    n362
  );


  not
  g1016
  (
    n1111,
    n338
  );


  not
  g1017
  (
    n1055,
    n411
  );


  not
  g1018
  (
    n942,
    n359
  );


  not
  g1019
  (
    n1455,
    n484
  );


  not
  g1020
  (
    n1471,
    n454
  );


  buf
  g1021
  (
    n1168,
    n441
  );


  not
  g1022
  (
    n1093,
    n360
  );


  not
  g1023
  (
    n530,
    n184
  );


  not
  g1024
  (
    n1136,
    n161
  );


  not
  g1025
  (
    n1411,
    n490
  );


  buf
  g1026
  (
    n784,
    n457
  );


  not
  g1027
  (
    n807,
    n415
  );


  buf
  g1028
  (
    n862,
    n489
  );


  buf
  g1029
  (
    n1408,
    n334
  );


  not
  g1030
  (
    n808,
    n465
  );


  not
  g1031
  (
    n968,
    n133
  );


  buf
  g1032
  (
    n1213,
    n447
  );


  buf
  g1033
  (
    n585,
    n399
  );


  buf
  g1034
  (
    n625,
    n328
  );


  not
  g1035
  (
    n633,
    n407
  );


  buf
  g1036
  (
    n1347,
    n463
  );


  not
  g1037
  (
    n637,
    n401
  );


  buf
  g1038
  (
    n1003,
    n181
  );


  buf
  g1039
  (
    n1178,
    n358
  );


  buf
  g1040
  (
    n1453,
    n319
  );


  not
  g1041
  (
    n1040,
    n491
  );


  not
  g1042
  (
    n559,
    n315
  );


  buf
  g1043
  (
    n1290,
    n366
  );


  not
  g1044
  (
    n1472,
    n433
  );


  not
  g1045
  (
    n1259,
    n487
  );


  buf
  g1046
  (
    n1297,
    n430
  );


  buf
  g1047
  (
    n1149,
    n343
  );


  buf
  g1048
  (
    n1399,
    n445
  );


  buf
  g1049
  (
    n564,
    n345
  );


  not
  g1050
  (
    n900,
    n371
  );


  not
  g1051
  (
    n553,
    n344
  );


  not
  g1052
  (
    n517,
    n436
  );


  buf
  g1053
  (
    n1300,
    n223
  );


  not
  g1054
  (
    n1155,
    n394
  );


  not
  g1055
  (
    n1261,
    n403
  );


  not
  g1056
  (
    n957,
    n414
  );


  buf
  g1057
  (
    n534,
    n391
  );


  not
  g1058
  (
    n1107,
    n467
  );


  buf
  g1059
  (
    n732,
    n371
  );


  buf
  g1060
  (
    n528,
    n383
  );


  buf
  g1061
  (
    n1271,
    n324
  );


  not
  g1062
  (
    n947,
    n381
  );


  buf
  g1063
  (
    n1258,
    n479
  );


  buf
  g1064
  (
    n1181,
    n326
  );


  buf
  g1065
  (
    n1231,
    n332
  );


  buf
  g1066
  (
    n1205,
    n446
  );


  buf
  g1067
  (
    n548,
    n324
  );


  not
  g1068
  (
    n688,
    n308
  );


  not
  g1069
  (
    n1439,
    n389
  );


  buf
  g1070
  (
    n525,
    n452
  );


  buf
  g1071
  (
    n1445,
    n131
  );


  buf
  g1072
  (
    n742,
    n462
  );


  buf
  g1073
  (
    n1177,
    n332
  );


  buf
  g1074
  (
    n1140,
    n341
  );


  buf
  g1075
  (
    n927,
    n303
  );


  not
  g1076
  (
    n538,
    n367
  );


  buf
  g1077
  (
    n618,
    n345
  );


  buf
  g1078
  (
    n679,
    n485
  );


  not
  g1079
  (
    n693,
    n426
  );


  buf
  g1080
  (
    n1127,
    n329
  );


  not
  g1081
  (
    n1116,
    n427
  );


  not
  g1082
  (
    n552,
    n346
  );


  buf
  g1083
  (
    n1089,
    n449
  );


  not
  g1084
  (
    n976,
    n355
  );


  buf
  g1085
  (
    n1337,
    n443
  );


  buf
  g1086
  (
    n1426,
    n339
  );


  not
  g1087
  (
    n891,
    n482
  );


  buf
  g1088
  (
    n1167,
    n282
  );


  buf
  g1089
  (
    n847,
    n471
  );


  buf
  g1090
  (
    n836,
    n402
  );


  not
  g1091
  (
    n1151,
    n252
  );


  not
  g1092
  (
    n1051,
    n394
  );


  not
  g1093
  (
    n889,
    n438
  );


  not
  g1094
  (
    n1449,
    n285
  );


  buf
  g1095
  (
    n1500,
    n357
  );


  buf
  g1096
  (
    n793,
    n356
  );


  not
  g1097
  (
    n540,
    n451
  );


  not
  g1098
  (
    n523,
    n382
  );


  buf
  g1099
  (
    n1491,
    n428
  );


  buf
  g1100
  (
    n1356,
    n300
  );


  buf
  g1101
  (
    n510,
    n396
  );


  not
  g1102
  (
    n1302,
    n488
  );


  not
  g1103
  (
    n1012,
    n248
  );


  buf
  g1104
  (
    n562,
    n126
  );


  buf
  g1105
  (
    n1389,
    n121
  );


  not
  g1106
  (
    n824,
    n311
  );


  buf
  g1107
  (
    n1228,
    n374
  );


  buf
  g1108
  (
    n545,
    n340
  );


  buf
  g1109
  (
    n1362,
    n464
  );


  not
  g1110
  (
    n1266,
    n470
  );


  not
  g1111
  (
    n1413,
    n476
  );


  not
  g1112
  (
    n992,
    n278
  );


  buf
  g1113
  (
    n1053,
    n440
  );


  not
  g1114
  (
    n1094,
    n168
  );


  buf
  g1115
  (
    n745,
    n139
  );


  buf
  g1116
  (
    n1291,
    n146
  );


  buf
  g1117
  (
    n761,
    n392
  );


  buf
  g1118
  (
    n756,
    n287
  );


  buf
  g1119
  (
    n1448,
    n495
  );


  buf
  g1120
  (
    n1350,
    n335
  );


  not
  g1121
  (
    n1365,
    n322
  );


  buf
  g1122
  (
    n590,
    n341
  );


  buf
  g1123
  (
    n694,
    n457
  );


  not
  g1124
  (
    n1103,
    n123
  );


  not
  g1125
  (
    n973,
    n368
  );


  buf
  g1126
  (
    n829,
    n294
  );


  not
  g1127
  (
    n939,
    n430
  );


  not
  g1128
  (
    n1223,
    n461
  );


  buf
  g1129
  (
    n1394,
    n448
  );


  not
  g1130
  (
    n1351,
    n419
  );


  not
  g1131
  (
    n677,
    n273
  );


  not
  g1132
  (
    n1159,
    n500
  );


  not
  g1133
  (
    n1341,
    n497
  );


  not
  g1134
  (
    n650,
    n398
  );


  buf
  g1135
  (
    n1359,
    n422
  );


  buf
  g1136
  (
    n1108,
    n378
  );


  not
  g1137
  (
    n744,
    n342
  );


  buf
  g1138
  (
    n579,
    n416
  );


  buf
  g1139
  (
    n1493,
    n191
  );


  not
  g1140
  (
    n602,
    n411
  );


  not
  g1141
  (
    n1048,
    n483
  );


  buf
  g1142
  (
    n853,
    n392
  );


  not
  g1143
  (
    n1317,
    n378
  );


  buf
  g1144
  (
    n1039,
    n386
  );


  buf
  g1145
  (
    n877,
    n454
  );


  not
  g1146
  (
    n727,
    n208
  );


  buf
  g1147
  (
    n1245,
    n342
  );


  not
  g1148
  (
    n638,
    n402
  );


  buf
  g1149
  (
    n649,
    n221
  );


  buf
  g1150
  (
    n934,
    n310
  );


  not
  g1151
  (
    n1444,
    n332
  );


  buf
  g1152
  (
    n1452,
    n431
  );


  buf
  g1153
  (
    n1029,
    n475
  );


  buf
  g1154
  (
    n684,
    n301
  );


  buf
  g1155
  (
    n1143,
    n226
  );


  not
  g1156
  (
    n611,
    n457
  );


  not
  g1157
  (
    n1473,
    n444
  );


  not
  g1158
  (
    n1396,
    n328
  );


  buf
  g1159
  (
    n1376,
    n194
  );


  buf
  g1160
  (
    n1164,
    n372
  );


  buf
  g1161
  (
    n1173,
    n340
  );


  not
  g1162
  (
    n721,
    n257
  );


  not
  g1163
  (
    n1283,
    n134
  );


  not
  g1164
  (
    n938,
    n129
  );


  buf
  g1165
  (
    n1081,
    n354
  );


  not
  g1166
  (
    n855,
    n358
  );


  buf
  g1167
  (
    n803,
    n260
  );


  not
  g1168
  (
    n573,
    n433
  );


  buf
  g1169
  (
    n764,
    n357
  );


  not
  g1170
  (
    n800,
    n480
  );


  not
  g1171
  (
    n1312,
    n327
  );


  buf
  g1172
  (
    n747,
    n309
  );


  not
  g1173
  (
    n719,
    n350
  );


  not
  g1174
  (
    n1479,
    n284
  );


  not
  g1175
  (
    n1105,
    n490
  );


  buf
  g1176
  (
    n1100,
    n447
  );


  buf
  g1177
  (
    n922,
    n498
  );


  buf
  g1178
  (
    n1247,
    n402
  );


  not
  g1179
  (
    n1377,
    n323
  );


  not
  g1180
  (
    n837,
    n499
  );


  buf
  g1181
  (
    n831,
    n486
  );


  not
  g1182
  (
    n1285,
    n379
  );


  buf
  g1183
  (
    n1368,
    n324
  );


  not
  g1184
  (
    n1461,
    n493
  );


  buf
  g1185
  (
    n725,
    n497
  );


  buf
  g1186
  (
    n1492,
    n322
  );


  buf
  g1187
  (
    n1367,
    n261
  );


  buf
  g1188
  (
    n1189,
    n384
  );


  buf
  g1189
  (
    n1078,
    n460
  );


  buf
  g1190
  (
    n1386,
    n436
  );


  buf
  g1191
  (
    n977,
    n472
  );


  not
  g1192
  (
    n892,
    n326
  );


  buf
  g1193
  (
    KeyWire_0_14,
    n435
  );


  not
  g1194
  (
    n661,
    n307
  );


  not
  g1195
  (
    n1503,
    n442
  );


  buf
  g1196
  (
    n1349,
    n448
  );


  not
  g1197
  (
    n859,
    n387
  );


  not
  g1198
  (
    n1276,
    n494
  );


  buf
  g1199
  (
    n1369,
    n386
  );


  not
  g1200
  (
    n858,
    n472
  );


  not
  g1201
  (
    n899,
    n348
  );


  not
  g1202
  (
    n904,
    n409
  );


  not
  g1203
  (
    n1395,
    n373
  );


  buf
  g1204
  (
    n1227,
    n436
  );


  buf
  g1205
  (
    n1244,
    n449
  );


  not
  g1206
  (
    n1318,
    n327
  );


  not
  g1207
  (
    n1080,
    n269
  );


  not
  g1208
  (
    n1371,
    n163
  );


  buf
  g1209
  (
    n1392,
    n349
  );


  buf
  g1210
  (
    n751,
    n200
  );


  buf
  g1211
  (
    n659,
    n462
  );


  not
  g1212
  (
    n1122,
    n414
  );


  buf
  g1213
  (
    n885,
    n359
  );


  not
  g1214
  (
    n1498,
    n298
  );


  not
  g1215
  (
    n681,
    n386
  );


  not
  g1216
  (
    n1045,
    n413
  );


  not
  g1217
  (
    n1273,
    n265
  );


  buf
  g1218
  (
    n1117,
    n446
  );


  buf
  g1219
  (
    n730,
    n409
  );


  buf
  g1220
  (
    KeyWire_0_4,
    n413
  );


  not
  g1221
  (
    n1346,
    n305
  );


  buf
  g1222
  (
    n574,
    n350
  );


  not
  g1223
  (
    n1036,
    n497
  );


  buf
  g1224
  (
    n1110,
    n450
  );


  buf
  g1225
  (
    n1330,
    n255
  );


  not
  g1226
  (
    n718,
    n380
  );


  not
  g1227
  (
    n589,
    n355
  );


  not
  g1228
  (
    n1066,
    n365
  );


  not
  g1229
  (
    n1187,
    n379
  );


  not
  g1230
  (
    n880,
    n242
  );


  not
  g1231
  (
    n1292,
    n352
  );


  buf
  g1232
  (
    n561,
    n293
  );


  not
  g1233
  (
    n849,
    n429
  );


  not
  g1234
  (
    n515,
    n472
  );


  buf
  g1235
  (
    n1225,
    n275
  );


  not
  g1236
  (
    n1431,
    n155
  );


  buf
  g1237
  (
    n698,
    n127
  );


  not
  g1238
  (
    n1020,
    n355
  );


  buf
  g1239
  (
    n598,
    n423
  );


  not
  g1240
  (
    n796,
    n413
  );


  buf
  g1241
  (
    n991,
    n344
  );


  not
  g1242
  (
    n1464,
    n485
  );


  buf
  g1243
  (
    n704,
    n451
  );


  not
  g1244
  (
    n712,
    n447
  );


  buf
  g1245
  (
    n1296,
    n318
  );


  not
  g1246
  (
    n876,
    n395
  );


  buf
  g1247
  (
    n907,
    n466
  );


  buf
  g1248
  (
    n1043,
    n346
  );


  not
  g1249
  (
    n1184,
    n478
  );


  buf
  g1250
  (
    n556,
    n440
  );


  buf
  g1251
  (
    n555,
    n276
  );


  buf
  g1252
  (
    n1264,
    n436
  );


  not
  g1253
  (
    n1462,
    n411
  );


  buf
  g1254
  (
    n935,
    n143
  );


  buf
  g1255
  (
    n581,
    n372
  );


  buf
  g1256
  (
    n1241,
    n315
  );


  buf
  g1257
  (
    n971,
    n124
  );


  not
  g1258
  (
    n845,
    n405
  );


  buf
  g1259
  (
    n832,
    n403
  );


  buf
  g1260
  (
    n844,
    n327
  );


  buf
  g1261
  (
    n1025,
    n279
  );


  not
  g1262
  (
    n1174,
    n314
  );


  not
  g1263
  (
    n1076,
    n400
  );


  not
  g1264
  (
    n1176,
    n136
  );


  not
  g1265
  (
    n551,
    n400
  );


  buf
  g1266
  (
    n918,
    n361
  );


  buf
  g1267
  (
    n1415,
    n473
  );


  not
  g1268
  (
    n949,
    n471
  );


  buf
  g1269
  (
    n641,
    n318
  );


  buf
  g1270
  (
    n1220,
    n499
  );


  buf
  g1271
  (
    n1242,
    n367
  );


  buf
  g1272
  (
    n1460,
    n420
  );


  buf
  g1273
  (
    n629,
    n167
  );


  not
  g1274
  (
    n768,
    n426
  );


  buf
  g1275
  (
    n1456,
    n360
  );


  not
  g1276
  (
    n779,
    n306
  );


  buf
  g1277
  (
    n887,
    n318
  );


  buf
  g1278
  (
    n1372,
    n415
  );


  buf
  g1279
  (
    n1375,
    n460
  );


  not
  g1280
  (
    n550,
    n454
  );


  not
  g1281
  (
    n543,
    n434
  );


  buf
  g1282
  (
    n609,
    n175
  );


  not
  g1283
  (
    n1102,
    n237
  );


  buf
  g1284
  (
    n1387,
    n166
  );


  buf
  g1285
  (
    n1171,
    n438
  );


  buf
  g1286
  (
    n1179,
    n174
  );


  buf
  g1287
  (
    n1006,
    n433
  );


  not
  g1288
  (
    n671,
    n351
  );


  not
  g1289
  (
    n1437,
    n372
  );


  buf
  g1290
  (
    n620,
    n368
  );


  not
  g1291
  (
    n813,
    n483
  );


  not
  g1292
  (
    n975,
    n261
  );


  not
  g1293
  (
    KeyWire_0_5,
    n173
  );


  buf
  g1294
  (
    n917,
    n473
  );


  not
  g1295
  (
    n587,
    n387
  );


  not
  g1296
  (
    n535,
    n486
  );


  buf
  g1297
  (
    n919,
    n375
  );


  buf
  g1298
  (
    n593,
    n478
  );


  not
  g1299
  (
    n572,
    n459
  );


  not
  g1300
  (
    n1098,
    n459
  );


  buf
  g1301
  (
    n1380,
    n432
  );


  not
  g1302
  (
    n660,
    n336
  );


  not
  g1303
  (
    n1329,
    n468
  );


  buf
  g1304
  (
    n1215,
    n487
  );


  not
  g1305
  (
    n981,
    n274
  );


  buf
  g1306
  (
    n720,
    n337
  );


  not
  g1307
  (
    n1482,
    n337
  );


  not
  g1308
  (
    n731,
    n201
  );


  buf
  g1309
  (
    n926,
    n465
  );


  not
  g1310
  (
    n1146,
    n339
  );


  not
  g1311
  (
    KeyWire_0_6,
    n363
  );


  not
  g1312
  (
    n816,
    n347
  );


  not
  g1313
  (
    n632,
    n453
  );


  not
  g1314
  (
    n599,
    n145
  );


  buf
  g1315
  (
    n1447,
    n463
  );


  not
  g1316
  (
    n654,
    n420
  );


  not
  g1317
  (
    n925,
    n455
  );


  not
  g1318
  (
    n666,
    n313
  );


  buf
  g1319
  (
    n1401,
    n376
  );


  buf
  g1320
  (
    n1506,
    n277
  );


  not
  g1321
  (
    n1243,
    n467
  );


  not
  g1322
  (
    n1440,
    n366
  );


  not
  g1323
  (
    n914,
    n438
  );


  buf
  g1324
  (
    n608,
    n156
  );


  buf
  g1325
  (
    n1326,
    n320
  );


  buf
  g1326
  (
    n962,
    n349
  );


  buf
  g1327
  (
    n1497,
    n351
  );


  buf
  g1328
  (
    n1438,
    n374
  );


  buf
  g1329
  (
    n1307,
    n304
  );


  buf
  g1330
  (
    n872,
    n279
  );


  not
  g1331
  (
    n610,
    n478
  );


  buf
  g1332
  (
    n759,
    n495
  );


  buf
  g1333
  (
    n1196,
    n462
  );


  buf
  g1334
  (
    n1404,
    n335
  );


  not
  g1335
  (
    n1250,
    n352
  );


  not
  g1336
  (
    n963,
    n498
  );


  buf
  g1337
  (
    n647,
    n326
  );


  buf
  g1338
  (
    n1188,
    n497
  );


  buf
  g1339
  (
    n1418,
    n473
  );


  not
  g1340
  (
    n953,
    n389
  );


  buf
  g1341
  (
    n989,
    n299
  );


  buf
  g1342
  (
    n1275,
    n276
  );


  buf
  g1343
  (
    n1141,
    n470
  );


  not
  g1344
  (
    n549,
    n388
  );


  buf
  g1345
  (
    n1058,
    n443
  );


  buf
  g1346
  (
    n828,
    n329
  );


  not
  g1347
  (
    n701,
    n473
  );


  buf
  g1348
  (
    n834,
    n376
  );


  not
  g1349
  (
    n630,
    n377
  );


  buf
  g1350
  (
    n643,
    n367
  );


  not
  g1351
  (
    n974,
    n365
  );


  buf
  g1352
  (
    n577,
    n239
  );


  buf
  g1353
  (
    n1430,
    n482
  );


  buf
  g1354
  (
    n1397,
    n405
  );


  not
  g1355
  (
    n1509,
    n348
  );


  not
  g1356
  (
    n542,
    n269
  );


  buf
  g1357
  (
    n1454,
    n325
  );


  buf
  g1358
  (
    n798,
    n486
  );


  not
  g1359
  (
    n903,
    n432
  );


  not
  g1360
  (
    n537,
    n492
  );


  buf
  g1361
  (
    n941,
    n246
  );


  buf
  g1362
  (
    n1021,
    n396
  );


  not
  g1363
  (
    n1147,
    n386
  );


  buf
  g1364
  (
    n1469,
    n362
  );


  buf
  g1365
  (
    n601,
    n370
  );


  buf
  g1366
  (
    n1233,
    n412
  );


  not
  g1367
  (
    n767,
    n416
  );


  not
  g1368
  (
    n1270,
    n420
  );


  buf
  g1369
  (
    n944,
    n434
  );


  buf
  g1370
  (
    n823,
    n338
  );


  buf
  g1371
  (
    n619,
    n425
  );


  buf
  g1372
  (
    n1096,
    n329
  );


  buf
  g1373
  (
    n1288,
    n231
  );


  not
  g1374
  (
    n576,
    n481
  );


  buf
  g1375
  (
    n626,
    n393
  );


  not
  g1376
  (
    n695,
    n412
  );


  buf
  g1377
  (
    n674,
    n356
  );


  not
  g1378
  (
    n787,
    n291
  );


  buf
  g1379
  (
    n1353,
    n365
  );


  buf
  g1380
  (
    n624,
    n498
  );


  buf
  g1381
  (
    n1083,
    n382
  );


  not
  g1382
  (
    n1487,
    n352
  );


  buf
  g1383
  (
    n1407,
    n288
  );


  buf
  g1384
  (
    n956,
    n363
  );


  not
  g1385
  (
    n1194,
    n187
  );


  buf
  g1386
  (
    n1502,
    n195
  );


  buf
  g1387
  (
    n1064,
    n458
  );


  buf
  g1388
  (
    n667,
    n431
  );


  buf
  g1389
  (
    n1002,
    n270
  );


  not
  g1390
  (
    n898,
    n422
  );


  buf
  g1391
  (
    n993,
    n358
  );


  buf
  g1392
  (
    n591,
    n453
  );


  buf
  g1393
  (
    n1054,
    n273
  );


  buf
  g1394
  (
    n596,
    n227
  );


  not
  g1395
  (
    n818,
    n331
  );


  not
  g1396
  (
    n583,
    n230
  );


  buf
  g1397
  (
    n668,
    n479
  );


  buf
  g1398
  (
    n1134,
    n418
  );


  buf
  g1399
  (
    n1166,
    n262
  );


  buf
  g1400
  (
    n1104,
    n501
  );


  buf
  g1401
  (
    n994,
    n441
  );


  buf
  g1402
  (
    n1311,
    n309
  );


  not
  g1403
  (
    n1293,
    n295
  );


  not
  g1404
  (
    n790,
    n287
  );


  buf
  g1405
  (
    n1088,
    n445
  );


  buf
  g1406
  (
    n1267,
    n236
  );


  not
  g1407
  (
    n776,
    n484
  );


  not
  g1408
  (
    n586,
    n369
  );


  not
  g1409
  (
    n959,
    n361
  );


  not
  g1410
  (
    n933,
    n455
  );


  not
  g1411
  (
    n739,
    n336
  );


  buf
  g1412
  (
    n1378,
    n225
  );


  buf
  g1413
  (
    n921,
    n271
  );


  buf
  g1414
  (
    n789,
    n468
  );


  buf
  g1415
  (
    n1279,
    n491
  );


  not
  g1416
  (
    n950,
    n135
  );


  not
  g1417
  (
    n1097,
    n455
  );


  not
  g1418
  (
    n955,
    n219
  );


  not
  g1419
  (
    n1253,
    n280
  );


  buf
  g1420
  (
    n1420,
    n398
  );


  not
  g1421
  (
    n1417,
    n389
  );


  buf
  g1422
  (
    n1046,
    n439
  );


  buf
  g1423
  (
    n1030,
    n283
  );


  buf
  g1424
  (
    n536,
    n286
  );


  buf
  g1425
  (
    n1095,
    n493
  );


  buf
  g1426
  (
    n705,
    n331
  );


  buf
  g1427
  (
    n1099,
    n384
  );


  not
  g1428
  (
    n758,
    n463
  );


  not
  g1429
  (
    n524,
    n487
  );


  not
  g1430
  (
    n870,
    n243
  );


  buf
  g1431
  (
    n1128,
    n408
  );


  buf
  g1432
  (
    n1336,
    n141
  );


  not
  g1433
  (
    n928,
    n320
  );


  not
  g1434
  (
    n890,
    n180
  );


  not
  g1435
  (
    n689,
    n158
  );


  not
  g1436
  (
    n1382,
    n228
  );


  buf
  g1437
  (
    n863,
    n468
  );


  buf
  g1438
  (
    n909,
    n446
  );


  not
  g1439
  (
    n817,
    n418
  );


  not
  g1440
  (
    n1018,
    n314
  );


  not
  g1441
  (
    n1414,
    n349
  );


  not
  g1442
  (
    n1073,
    n429
  );


  not
  g1443
  (
    n1262,
    n347
  );


  buf
  g1444
  (
    n1172,
    n272
  );


  not
  g1445
  (
    n1344,
    n362
  );


  not
  g1446
  (
    n1217,
    n469
  );


  buf
  g1447
  (
    n830,
    n213
  );


  not
  g1448
  (
    n709,
    n412
  );


  buf
  g1449
  (
    n648,
    n437
  );


  buf
  g1450
  (
    n1175,
    n485
  );


  buf
  g1451
  (
    n680,
    n336
  );


  buf
  g1452
  (
    n774,
    n394
  );


  not
  g1453
  (
    n607,
    n474
  );


  not
  g1454
  (
    n1210,
    n442
  );


  buf
  g1455
  (
    n792,
    n245
  );


  buf
  g1456
  (
    n1208,
    n496
  );


  buf
  g1457
  (
    n1327,
    n430
  );


  not
  g1458
  (
    n673,
    n495
  );


  not
  g1459
  (
    n1216,
    n364
  );


  not
  g1460
  (
    n951,
    n337
  );


  not
  g1461
  (
    n1303,
    n316
  );


  not
  g1462
  (
    n1004,
    n378
  );


  not
  g1463
  (
    n1218,
    n258
  );


  not
  g1464
  (
    n1090,
    n178
  );


  not
  g1465
  (
    n851,
    n313
  );


  buf
  g1466
  (
    n1277,
    n297
  );


  not
  g1467
  (
    n846,
    n375
  );


  buf
  g1468
  (
    n512,
    n364
  );


  buf
  g1469
  (
    n806,
    n280
  );


  not
  g1470
  (
    n1338,
    n357
  );


  buf
  g1471
  (
    n1027,
    n345
  );


  not
  g1472
  (
    n1026,
    n370
  );


  buf
  g1473
  (
    n1198,
    n358
  );


  not
  g1474
  (
    n1331,
    n469
  );


  not
  g1475
  (
    n795,
    n425
  );


  not
  g1476
  (
    n982,
    n347
  );


  not
  g1477
  (
    n707,
    n159
  );


  buf
  g1478
  (
    n1402,
    n424
  );


  buf
  g1479
  (
    n945,
    n356
  );


  not
  g1480
  (
    n1268,
    n468
  );


  not
  g1481
  (
    n1423,
    n448
  );


  not
  g1482
  (
    n1484,
    n461
  );


  buf
  g1483
  (
    n1221,
    n487
  );


  not
  g1484
  (
    n782,
    n470
  );


  buf
  g1485
  (
    n1202,
    n384
  );


  buf
  g1486
  (
    n1828,
    n570
  );


  not
  g1487
  (
    n2025,
    n527
  );


  buf
  g1488
  (
    n1979,
    n695
  );


  buf
  g1489
  (
    n1571,
    n644
  );


  buf
  g1490
  (
    n1857,
    n726
  );


  buf
  g1491
  (
    n2168,
    n882
  );


  not
  g1492
  (
    n1825,
    n795
  );


  buf
  g1493
  (
    n2070,
    n517
  );


  buf
  g1494
  (
    n2062,
    n1096
  );


  buf
  g1495
  (
    n1656,
    n591
  );


  buf
  g1496
  (
    n1973,
    n996
  );


  not
  g1497
  (
    n1949,
    n939
  );


  buf
  g1498
  (
    n2063,
    n675
  );


  buf
  g1499
  (
    n1525,
    n691
  );


  buf
  g1500
  (
    n2173,
    n817
  );


  buf
  g1501
  (
    n1754,
    n1070
  );


  not
  g1502
  (
    n2175,
    n522
  );


  not
  g1503
  (
    n1850,
    n1042
  );


  not
  g1504
  (
    n1964,
    n770
  );


  not
  g1505
  (
    n2177,
    n1147
  );


  not
  g1506
  (
    n1824,
    n887
  );


  buf
  g1507
  (
    n2163,
    n941
  );


  buf
  g1508
  (
    n2137,
    n938
  );


  buf
  g1509
  (
    n1629,
    n706
  );


  not
  g1510
  (
    n1913,
    n714
  );


  not
  g1511
  (
    n1721,
    n1027
  );


  buf
  g1512
  (
    n1698,
    n1119
  );


  buf
  g1513
  (
    n2127,
    n556
  );


  buf
  g1514
  (
    n1746,
    n1062
  );


  not
  g1515
  (
    n1567,
    n630
  );


  not
  g1516
  (
    n2001,
    n615
  );


  buf
  g1517
  (
    n2012,
    n1142
  );


  buf
  g1518
  (
    n2113,
    n720
  );


  buf
  g1519
  (
    n1546,
    n857
  );


  buf
  g1520
  (
    n1847,
    n1134
  );


  buf
  g1521
  (
    n1579,
    n596
  );


  buf
  g1522
  (
    n1926,
    n509
  );


  buf
  g1523
  (
    n1956,
    n622
  );


  buf
  g1524
  (
    n1758,
    n954
  );


  not
  g1525
  (
    n1699,
    n1004
  );


  buf
  g1526
  (
    n1863,
    n788
  );


  not
  g1527
  (
    n2083,
    n1099
  );


  not
  g1528
  (
    n1787,
    n821
  );


  not
  g1529
  (
    n1788,
    n516
  );


  not
  g1530
  (
    n2105,
    n734
  );


  buf
  g1531
  (
    n1654,
    n761
  );


  buf
  g1532
  (
    n2116,
    n993
  );


  buf
  g1533
  (
    n1748,
    n525
  );


  buf
  g1534
  (
    n1859,
    n530
  );


  buf
  g1535
  (
    n2120,
    n774
  );


  buf
  g1536
  (
    n1659,
    n963
  );


  buf
  g1537
  (
    n2056,
    n666
  );


  not
  g1538
  (
    n2150,
    n1141
  );


  not
  g1539
  (
    n2043,
    n697
  );


  not
  g1540
  (
    n1910,
    n689
  );


  not
  g1541
  (
    n1764,
    n967
  );


  buf
  g1542
  (
    n1635,
    n647
  );


  buf
  g1543
  (
    n1693,
    n785
  );


  not
  g1544
  (
    n1974,
    n1129
  );


  not
  g1545
  (
    n2050,
    n577
  );


  buf
  g1546
  (
    n1705,
    n822
  );


  not
  g1547
  (
    n1584,
    n743
  );


  not
  g1548
  (
    n1763,
    n922
  );


  buf
  g1549
  (
    n2004,
    n755
  );


  buf
  g1550
  (
    n1535,
    n1074
  );


  buf
  g1551
  (
    KeyWire_0_7,
    n747
  );


  buf
  g1552
  (
    n1800,
    n728
  );


  not
  g1553
  (
    n1548,
    n511
  );


  not
  g1554
  (
    n1808,
    n927
  );


  not
  g1555
  (
    n1557,
    n656
  );


  buf
  g1556
  (
    n1793,
    n1148
  );


  buf
  g1557
  (
    n1624,
    n566
  );


  buf
  g1558
  (
    n1823,
    n1082
  );


  not
  g1559
  (
    n1730,
    n1162
  );


  not
  g1560
  (
    n2053,
    n952
  );


  not
  g1561
  (
    n1714,
    n865
  );


  buf
  g1562
  (
    n1917,
    n765
  );


  buf
  g1563
  (
    n1540,
    n864
  );


  not
  g1564
  (
    n1849,
    n624
  );


  buf
  g1565
  (
    n1961,
    n862
  );


  buf
  g1566
  (
    n1615,
    n722
  );


  not
  g1567
  (
    n1835,
    n1126
  );


  buf
  g1568
  (
    n1651,
    n680
  );


  not
  g1569
  (
    n2006,
    n1059
  );


  buf
  g1570
  (
    n1537,
    n972
  );


  buf
  g1571
  (
    n2079,
    n725
  );


  buf
  g1572
  (
    n1600,
    n895
  );


  buf
  g1573
  (
    n1955,
    n554
  );


  buf
  g1574
  (
    n2164,
    n1066
  );


  buf
  g1575
  (
    n1736,
    n645
  );


  buf
  g1576
  (
    n1940,
    n1031
  );


  not
  g1577
  (
    n1619,
    n975
  );


  buf
  g1578
  (
    n1695,
    n589
  );


  buf
  g1579
  (
    n2121,
    n798
  );


  not
  g1580
  (
    n1912,
    n631
  );


  buf
  g1581
  (
    n1986,
    n958
  );


  not
  g1582
  (
    n1761,
    n569
  );


  buf
  g1583
  (
    n1555,
    n555
  );


  not
  g1584
  (
    n1792,
    n1155
  );


  not
  g1585
  (
    n2084,
    n838
  );


  buf
  g1586
  (
    n1728,
    n1045
  );


  not
  g1587
  (
    n2031,
    n940
  );


  not
  g1588
  (
    n1812,
    n721
  );


  buf
  g1589
  (
    n2103,
    n677
  );


  buf
  g1590
  (
    n2059,
    n1006
  );


  buf
  g1591
  (
    n2139,
    n863
  );


  not
  g1592
  (
    n1675,
    n1048
  );


  buf
  g1593
  (
    n2014,
    n611
  );


  not
  g1594
  (
    n2108,
    n617
  );


  buf
  g1595
  (
    n1775,
    n973
  );


  not
  g1596
  (
    n1578,
    n812
  );


  buf
  g1597
  (
    n1549,
    n1079
  );


  not
  g1598
  (
    n1620,
    n1089
  );


  not
  g1599
  (
    n1575,
    n575
  );


  buf
  g1600
  (
    n1603,
    n1158
  );


  buf
  g1601
  (
    n2046,
    n653
  );


  not
  g1602
  (
    n2040,
    n639
  );


  not
  g1603
  (
    n1958,
    n846
  );


  buf
  g1604
  (
    n2058,
    n989
  );


  not
  g1605
  (
    n1708,
    n1157
  );


  buf
  g1606
  (
    n1559,
    n1181
  );


  buf
  g1607
  (
    n1959,
    n1053
  );


  buf
  g1608
  (
    n1687,
    n898
  );


  not
  g1609
  (
    n1737,
    n1047
  );


  buf
  g1610
  (
    n1672,
    n1073
  );


  buf
  g1611
  (
    n2085,
    n943
  );


  not
  g1612
  (
    n2069,
    n955
  );


  buf
  g1613
  (
    n1935,
    n791
  );


  not
  g1614
  (
    n1997,
    n1115
  );


  buf
  g1615
  (
    n1989,
    n815
  );


  buf
  g1616
  (
    n1753,
    n829
  );


  buf
  g1617
  (
    n2090,
    n836
  );


  buf
  g1618
  (
    n1544,
    n1056
  );


  buf
  g1619
  (
    n1563,
    n625
  );


  not
  g1620
  (
    n1783,
    n702
  );


  not
  g1621
  (
    n2019,
    n804
  );


  not
  g1622
  (
    n1796,
    n612
  );


  buf
  g1623
  (
    n1517,
    n813
  );


  buf
  g1624
  (
    n1621,
    n934
  );


  not
  g1625
  (
    n1734,
    n935
  );


  buf
  g1626
  (
    n2179,
    n1130
  );


  buf
  g1627
  (
    n1953,
    n881
  );


  not
  g1628
  (
    n1550,
    n819
  );


  not
  g1629
  (
    n2106,
    n949
  );


  buf
  g1630
  (
    n1671,
    n1109
  );


  buf
  g1631
  (
    n2132,
    n609
  );


  buf
  g1632
  (
    n1894,
    n1022
  );


  not
  g1633
  (
    n1965,
    n637
  );


  buf
  g1634
  (
    n1589,
    n767
  );


  not
  g1635
  (
    n2104,
    n667
  );


  buf
  g1636
  (
    n1626,
    n515
  );


  not
  g1637
  (
    n2071,
    n588
  );


  buf
  g1638
  (
    n1802,
    n1077
  );


  buf
  g1639
  (
    n1583,
    n1098
  );


  not
  g1640
  (
    n1987,
    n541
  );


  buf
  g1641
  (
    n1821,
    n853
  );


  not
  g1642
  (
    n1658,
    n1020
  );


  buf
  g1643
  (
    n1733,
    n605
  );


  not
  g1644
  (
    n1801,
    n969
  );


  buf
  g1645
  (
    n2023,
    n900
  );


  buf
  g1646
  (
    n1545,
    n729
  );


  buf
  g1647
  (
    n2002,
    n1146
  );


  buf
  g1648
  (
    n1627,
    n871
  );


  buf
  g1649
  (
    n2161,
    n1090
  );


  buf
  g1650
  (
    n1511,
    n1012
  );


  buf
  g1651
  (
    n1925,
    n792
  );


  not
  g1652
  (
    n1937,
    n707
  );


  buf
  g1653
  (
    n1891,
    n688
  );


  buf
  g1654
  (
    n1556,
    n1168
  );


  buf
  g1655
  (
    n2123,
    n1005
  );


  buf
  g1656
  (
    n1901,
    n899
  );


  buf
  g1657
  (
    n1868,
    n538
  );


  not
  g1658
  (
    n2181,
    n1072
  );


  buf
  g1659
  (
    n1984,
    n773
  );


  not
  g1660
  (
    n1616,
    n1029
  );


  not
  g1661
  (
    n1916,
    n842
  );


  not
  g1662
  (
    n1981,
    n1075
  );


  buf
  g1663
  (
    n1715,
    n693
  );


  buf
  g1664
  (
    n1757,
    n1061
  );


  not
  g1665
  (
    n2134,
    n565
  );


  buf
  g1666
  (
    n1605,
    n982
  );


  buf
  g1667
  (
    n1780,
    n1033
  );


  buf
  g1668
  (
    n1534,
    n582
  );


  not
  g1669
  (
    n1606,
    n600
  );


  buf
  g1670
  (
    n1885,
    n655
  );


  buf
  g1671
  (
    n1922,
    n867
  );


  not
  g1672
  (
    n2152,
    n928
  );


  buf
  g1673
  (
    n1670,
    n823
  );


  buf
  g1674
  (
    n1558,
    n1177
  );


  buf
  g1675
  (
    n2160,
    n1065
  );


  buf
  g1676
  (
    n1883,
    n1123
  );


  buf
  g1677
  (
    n1843,
    n1064
  );


  not
  g1678
  (
    n1516,
    n586
  );


  not
  g1679
  (
    n1512,
    n930
  );


  not
  g1680
  (
    n2187,
    n884
  );


  buf
  g1681
  (
    n1530,
    n731
  );


  buf
  g1682
  (
    n2169,
    n552
  );


  buf
  g1683
  (
    n1882,
    n851
  );


  not
  g1684
  (
    n1632,
    n810
  );


  buf
  g1685
  (
    n2015,
    n1136
  );


  buf
  g1686
  (
    n1677,
    n602
  );


  buf
  g1687
  (
    n2030,
    n1118
  );


  not
  g1688
  (
    n2124,
    n551
  );


  buf
  g1689
  (
    n1722,
    n910
  );


  not
  g1690
  (
    n1822,
    n550
  );


  not
  g1691
  (
    n2041,
    n710
  );


  not
  g1692
  (
    n2157,
    n1084
  );


  buf
  g1693
  (
    n1688,
    n1037
  );


  buf
  g1694
  (
    n1839,
    n929
  );


  buf
  g1695
  (
    n1751,
    n784
  );


  buf
  g1696
  (
    n1810,
    n531
  );


  buf
  g1697
  (
    n1854,
    n874
  );


  not
  g1698
  (
    n1657,
    n818
  );


  not
  g1699
  (
    n1595,
    n1144
  );


  buf
  g1700
  (
    n1609,
    n966
  );


  not
  g1701
  (
    n1643,
    n713
  );


  buf
  g1702
  (
    n1590,
    n620
  );


  not
  g1703
  (
    n1870,
    n908
  );


  buf
  g1704
  (
    n1554,
    n1091
  );


  buf
  g1705
  (
    n1541,
    n861
  );


  buf
  g1706
  (
    n2129,
    n1114
  );


  buf
  g1707
  (
    n1867,
    n508
  );


  buf
  g1708
  (
    n2141,
    n623
  );


  not
  g1709
  (
    n1815,
    n1107
  );


  buf
  g1710
  (
    n1930,
    n834
  );


  not
  g1711
  (
    n1860,
    n690
  );


  not
  g1712
  (
    n1562,
    n694
  );


  buf
  g1713
  (
    n1879,
    n684
  );


  not
  g1714
  (
    n1637,
    n789
  );


  not
  g1715
  (
    n1648,
    n629
  );


  not
  g1716
  (
    n1856,
    n893
  );


  buf
  g1717
  (
    n1876,
    n660
  );


  not
  g1718
  (
    n2099,
    n643
  );


  buf
  g1719
  (
    n1645,
    n627
  );


  buf
  g1720
  (
    n2143,
    n923
  );


  buf
  g1721
  (
    n1646,
    n584
  );


  not
  g1722
  (
    n1782,
    n636
  );


  not
  g1723
  (
    n2186,
    n1164
  );


  not
  g1724
  (
    n1633,
    n751
  );


  not
  g1725
  (
    n1992,
    n1052
  );


  buf
  g1726
  (
    n2021,
    n1063
  );


  not
  g1727
  (
    n1939,
    n787
  );


  buf
  g1728
  (
    n1875,
    n670
  );


  buf
  g1729
  (
    n2052,
    n580
  );


  buf
  g1730
  (
    n1874,
    n1175
  );


  buf
  g1731
  (
    n2155,
    n1008
  );


  not
  g1732
  (
    n1724,
    n614
  );


  not
  g1733
  (
    n1971,
    n855
  );


  buf
  g1734
  (
    n2008,
    n832
  );


  buf
  g1735
  (
    n1725,
    n753
  );


  buf
  g1736
  (
    n1719,
    n518
  );


  buf
  g1737
  (
    n1694,
    n1182
  );


  not
  g1738
  (
    n2138,
    n587
  );


  buf
  g1739
  (
    n1729,
    n991
  );


  buf
  g1740
  (
    n1899,
    n756
  );


  not
  g1741
  (
    n1934,
    n520
  );


  buf
  g1742
  (
    n1684,
    n793
  );


  not
  g1743
  (
    n1848,
    n914
  );


  not
  g1744
  (
    n1570,
    n965
  );


  buf
  g1745
  (
    n1527,
    n536
  );


  buf
  g1746
  (
    n1878,
    n1117
  );


  not
  g1747
  (
    n1528,
    n711
  );


  not
  g1748
  (
    n2087,
    n891
  );


  buf
  g1749
  (
    n1588,
    n1018
  );


  buf
  g1750
  (
    n1932,
    n745
  );


  buf
  g1751
  (
    n2018,
    n771
  );


  not
  g1752
  (
    n2136,
    n1152
  );


  buf
  g1753
  (
    n1739,
    n843
  );


  buf
  g1754
  (
    n2145,
    n1046
  );


  not
  g1755
  (
    n1975,
    n652
  );


  buf
  g1756
  (
    n2072,
    n529
  );


  buf
  g1757
  (
    n2068,
    n1183
  );


  not
  g1758
  (
    n2098,
    n1120
  );


  not
  g1759
  (
    n1920,
    n796
  );


  not
  g1760
  (
    n2162,
    n1101
  );


  buf
  g1761
  (
    n2096,
    n512
  );


  not
  g1762
  (
    n1832,
    n888
  );


  not
  g1763
  (
    n2057,
    n913
  );


  not
  g1764
  (
    n2081,
    n599
  );


  not
  g1765
  (
    n2077,
    n962
  );


  not
  g1766
  (
    n2028,
    n513
  );


  buf
  g1767
  (
    n1960,
    n1051
  );


  buf
  g1768
  (
    n1759,
    n716
  );


  not
  g1769
  (
    n2170,
    n858
  );


  buf
  g1770
  (
    n1846,
    n749
  );


  buf
  g1771
  (
    n2180,
    n715
  );


  not
  g1772
  (
    n1969,
    n970
  );


  buf
  g1773
  (
    n1702,
    n986
  );


  buf
  g1774
  (
    n1842,
    n1049
  );


  not
  g1775
  (
    n2074,
    n534
  );


  buf
  g1776
  (
    n2118,
    n724
  );


  not
  g1777
  (
    n2158,
    n681
  );


  buf
  g1778
  (
    n1598,
    n1044
  );


  not
  g1779
  (
    n1994,
    n549
  );


  not
  g1780
  (
    n1623,
    n878
  );


  not
  g1781
  (
    n2092,
    n696
  );


  buf
  g1782
  (
    n2003,
    n831
  );


  not
  g1783
  (
    n2067,
    n739
  );


  buf
  g1784
  (
    n1889,
    n1068
  );


  not
  g1785
  (
    n1631,
    n1133
  );


  buf
  g1786
  (
    n1524,
    n760
  );


  buf
  g1787
  (
    n2073,
    n944
  );


  not
  g1788
  (
    n1904,
    n1060
  );


  not
  g1789
  (
    n1902,
    n984
  );


  buf
  g1790
  (
    n1809,
    n1102
  );


  buf
  g1791
  (
    n2010,
    n1087
  );


  not
  g1792
  (
    n1890,
    n1178
  );


  buf
  g1793
  (
    n1682,
    n797
  );


  buf
  g1794
  (
    n1644,
    n856
  );


  not
  g1795
  (
    n1599,
    n754
  );


  buf
  g1796
  (
    n2044,
    n671
  );


  not
  g1797
  (
    n1880,
    n875
  );


  not
  g1798
  (
    KeyWire_0_0,
    n1103
  );


  buf
  g1799
  (
    n1640,
    n769
  );


  not
  g1800
  (
    n1689,
    n561
  );


  not
  g1801
  (
    n1665,
    n1111
  );


  not
  g1802
  (
    n1798,
    n1036
  );


  buf
  g1803
  (
    n1834,
    n1167
  );


  buf
  g1804
  (
    n2114,
    n872
  );


  not
  g1805
  (
    n1946,
    n1067
  );


  not
  g1806
  (
    n1915,
    n839
  );


  not
  g1807
  (
    n1520,
    n869
  );


  buf
  g1808
  (
    n2088,
    n1026
  );


  buf
  g1809
  (
    n2174,
    n676
  );


  buf
  g1810
  (
    n1887,
    n524
  );


  not
  g1811
  (
    n1951,
    n683
  );


  not
  g1812
  (
    n1928,
    n837
  );


  buf
  g1813
  (
    n1864,
    n1016
  );


  buf
  g1814
  (
    n1978,
    n912
  );


  buf
  g1815
  (
    n1752,
    n1093
  );


  buf
  g1816
  (
    n1662,
    n618
  );


  buf
  g1817
  (
    n1741,
    n1150
  );


  not
  g1818
  (
    n1968,
    n1105
  );


  buf
  g1819
  (
    n2037,
    n659
  );


  buf
  g1820
  (
    n2154,
    n889
  );


  buf
  g1821
  (
    n2097,
    n957
  );


  buf
  g1822
  (
    n1536,
    n616
  );


  not
  g1823
  (
    n1976,
    n901
  );


  buf
  g1824
  (
    n2011,
    n805
  );


  buf
  g1825
  (
    n1950,
    n709
  );


  buf
  g1826
  (
    n1948,
    n633
  );


  not
  g1827
  (
    n2016,
    n1161
  );


  buf
  g1828
  (
    n1760,
    n1166
  );


  buf
  g1829
  (
    n1529,
    n1176
  );


  not
  g1830
  (
    n1610,
    n1113
  );


  not
  g1831
  (
    n1970,
    n514
  );


  buf
  g1832
  (
    n2125,
    n946
  );


  not
  g1833
  (
    n1718,
    n906
  );


  buf
  g1834
  (
    n1594,
    n598
  );


  buf
  g1835
  (
    n1749,
    n553
  );


  buf
  g1836
  (
    n2182,
    n879
  );


  not
  g1837
  (
    n1669,
    n947
  );


  buf
  g1838
  (
    n1774,
    n1165
  );


  not
  g1839
  (
    n1582,
    n896
  );


  buf
  g1840
  (
    n1611,
    n662
  );


  not
  g1841
  (
    n2051,
    n945
  );


  buf
  g1842
  (
    n1568,
    n661
  );


  buf
  g1843
  (
    n2005,
    n894
  );


  buf
  g1844
  (
    n1513,
    n758
  );


  buf
  g1845
  (
    n2184,
    n1108
  );


  not
  g1846
  (
    n1710,
    n897
  );


  not
  g1847
  (
    n2142,
    n803
  );


  buf
  g1848
  (
    n1542,
    n1171
  );


  not
  g1849
  (
    n2112,
    n840
  );


  not
  g1850
  (
    n2027,
    n1034
  );


  not
  g1851
  (
    n1663,
    n1071
  );


  not
  g1852
  (
    n1566,
    n1057
  );


  buf
  g1853
  (
    n1586,
    n1035
  );


  not
  g1854
  (
    n1840,
    n808
  );


  not
  g1855
  (
    n2102,
    n1100
  );


  buf
  g1856
  (
    n2045,
    n708
  );


  not
  g1857
  (
    n1519,
    n1041
  );


  buf
  g1858
  (
    n1929,
    n931
  );


  buf
  g1859
  (
    n1933,
    n664
  );


  not
  g1860
  (
    n2007,
    n809
  );


  buf
  g1861
  (
    n1872,
    n1163
  );


  buf
  g1862
  (
    n1704,
    n979
  );


  buf
  g1863
  (
    n1991,
    n951
  );


  buf
  g1864
  (
    n2035,
    n870
  );


  not
  g1865
  (
    n1523,
    n560
  );


  not
  g1866
  (
    n1947,
    n678
  );


  not
  g1867
  (
    n1587,
    n866
  );


  buf
  g1868
  (
    n2078,
    n988
  );


  not
  g1869
  (
    n1660,
    n933
  );


  not
  g1870
  (
    n1884,
    n651
  );


  buf
  g1871
  (
    n1871,
    n506
  );


  buf
  g1872
  (
    n1622,
    n668
  );


  not
  g1873
  (
    n1607,
    n673
  );


  buf
  g1874
  (
    n1830,
    n1145
  );


  not
  g1875
  (
    n1641,
    n1043
  );


  buf
  g1876
  (
    n1766,
    n672
  );


  buf
  g1877
  (
    n2054,
    n703
  );


  not
  g1878
  (
    n2109,
    n916
  );


  not
  g1879
  (
    n2126,
    n768
  );


  not
  g1880
  (
    n1750,
    n1013
  );


  buf
  g1881
  (
    n1638,
    n1179
  );


  not
  g1882
  (
    n1581,
    n920
  );


  not
  g1883
  (
    n1564,
    n1038
  );


  buf
  g1884
  (
    n1685,
    n909
  );


  buf
  g1885
  (
    n1683,
    n987
  );


  buf
  g1886
  (
    n1985,
    n610
  );


  buf
  g1887
  (
    n1845,
    n1154
  );


  not
  g1888
  (
    n1803,
    n1076
  );


  not
  g1889
  (
    n1593,
    n854
  );


  buf
  g1890
  (
    n1995,
    n685
  );


  not
  g1891
  (
    n1522,
    n1180
  );


  buf
  g1892
  (
    n1954,
    n692
  );


  buf
  g1893
  (
    n1877,
    n540
  );


  buf
  g1894
  (
    n1533,
    n669
  );


  not
  g1895
  (
    n1851,
    n521
  );


  buf
  g1896
  (
    n2178,
    n573
  );


  buf
  g1897
  (
    n1941,
    n905
  );


  not
  g1898
  (
    n1608,
    n860
  );


  not
  g1899
  (
    n1565,
    n1092
  );


  buf
  g1900
  (
    n1931,
    n1078
  );


  buf
  g1901
  (
    n2093,
    n604
  );


  buf
  g1902
  (
    n1735,
    n926
  );


  buf
  g1903
  (
    n2135,
    n932
  );


  not
  g1904
  (
    n1649,
    n727
  );


  not
  g1905
  (
    n2042,
    n806
  );


  buf
  g1906
  (
    n1790,
    n632
  );


  buf
  g1907
  (
    n1831,
    n528
  );


  not
  g1908
  (
    n1897,
    n995
  );


  not
  g1909
  (
    n1778,
    n1032
  );


  buf
  g1910
  (
    n1990,
    n519
  );


  buf
  g1911
  (
    n1727,
    n533
  );


  not
  g1912
  (
    n2133,
    n825
  );


  buf
  g1913
  (
    n1613,
    n1019
  );


  buf
  g1914
  (
    n1799,
    n790
  );


  not
  g1915
  (
    n1706,
    n1040
  );


  not
  g1916
  (
    n2147,
    n559
  );


  buf
  g1917
  (
    n2122,
    n876
  );


  not
  g1918
  (
    n1731,
    n999
  );


  not
  g1919
  (
    n1596,
    n1151
  );


  buf
  g1920
  (
    n2095,
    n657
  );


  not
  g1921
  (
    n2020,
    n1080
  );


  not
  g1922
  (
    n2185,
    n835
  );


  not
  g1923
  (
    n2026,
    n748
  );


  buf
  g1924
  (
    n1862,
    n997
  );


  not
  g1925
  (
    n1655,
    n635
  );


  not
  g1926
  (
    n2144,
    n948
  );


  buf
  g1927
  (
    n2082,
    n1083
  );


  not
  g1928
  (
    n1521,
    n1028
  );


  buf
  g1929
  (
    n1786,
    n1153
  );


  buf
  g1930
  (
    n1771,
    n663
  );


  not
  g1931
  (
    n1612,
    n641
  );


  buf
  g1932
  (
    n1826,
    n736
  );


  buf
  g1933
  (
    n1674,
    n595
  );


  not
  g1934
  (
    n1919,
    n543
  );


  not
  g1935
  (
    n1585,
    n903
  );


  buf
  g1936
  (
    n1732,
    n1050
  );


  not
  g1937
  (
    n2065,
    n1140
  );


  not
  g1938
  (
    n2148,
    n1001
  );


  buf
  g1939
  (
    n1844,
    n998
  );


  not
  g1940
  (
    n1818,
    n978
  );


  not
  g1941
  (
    n2076,
    n698
  );


  not
  g1942
  (
    n1813,
    n990
  );


  buf
  g1943
  (
    n1806,
    n1174
  );


  buf
  g1944
  (
    n2101,
    n658
  );


  buf
  g1945
  (
    n1911,
    n699
  );


  not
  g1946
  (
    n2183,
    n1030
  );


  not
  g1947
  (
    n1918,
    n830
  );


  buf
  g1948
  (
    n1690,
    n1160
  );


  buf
  g1949
  (
    n1967,
    n1017
  );


  not
  g1950
  (
    n2094,
    n1094
  );


  buf
  g1951
  (
    n1726,
    n985
  );


  not
  g1952
  (
    n1820,
    n742
  );


  not
  g1953
  (
    n1827,
    n558
  );


  not
  g1954
  (
    n1957,
    n752
  );


  buf
  g1955
  (
    n1944,
    n1121
  );


  buf
  g1956
  (
    n1602,
    n712
  );


  not
  g1957
  (
    n1738,
    n1024
  );


  not
  g1958
  (
    n2107,
    n568
  );


  buf
  g1959
  (
    n1531,
    n780
  );


  not
  g1960
  (
    n1538,
    n764
  );


  not
  g1961
  (
    n1804,
    n907
  );


  buf
  g1962
  (
    n1560,
    n802
  );


  buf
  g1963
  (
    n2171,
    n1097
  );


  not
  g1964
  (
    n2156,
    n640
  );


  buf
  g1965
  (
    n1518,
    n723
  );


  buf
  g1966
  (
    n2036,
    n719
  );


  not
  g1967
  (
    n1680,
    n977
  );


  not
  g1968
  (
    n1707,
    n841
  );


  buf
  g1969
  (
    n1572,
    n807
  );


  buf
  g1970
  (
    n1838,
    n548
  );


  buf
  g1971
  (
    n1601,
    n759
  );


  buf
  g1972
  (
    n1720,
    n919
  );


  buf
  g1973
  (
    n1636,
    n782
  );


  buf
  g1974
  (
    n1762,
    n1172
  );


  not
  g1975
  (
    n2038,
    n890
  );


  buf
  g1976
  (
    n1898,
    n1139
  );


  not
  g1977
  (
    n1896,
    n868
  );


  not
  g1978
  (
    n1988,
    n579
  );


  buf
  g1979
  (
    n2086,
    n735
  );


  buf
  g1980
  (
    n1673,
    n621
  );


  buf
  g1981
  (
    n1966,
    n921
  );


  buf
  g1982
  (
    n1747,
    n892
  );


  not
  g1983
  (
    n1697,
    n778
  );


  buf
  g1984
  (
    n2159,
    n687
  );


  not
  g1985
  (
    n1791,
    n1159
  );


  not
  g1986
  (
    n2013,
    n974
  );


  not
  g1987
  (
    n2009,
    n886
  );


  buf
  g1988
  (
    n2060,
    n1156
  );


  buf
  g1989
  (
    n1865,
    n544
  );


  not
  g1990
  (
    n2146,
    n953
  );


  buf
  g1991
  (
    n1678,
    n1054
  );


  not
  g1992
  (
    n2165,
    n772
  );


  not
  g1993
  (
    n1703,
    n902
  );


  not
  g1994
  (
    n1905,
    n562
  );


  not
  g1995
  (
    n1784,
    n732
  );


  buf
  g1996
  (
    n1700,
    n603
  );


  buf
  g1997
  (
    n1921,
    n1007
  );


  not
  g1998
  (
    n1614,
    n597
  );


  buf
  g1999
  (
    n1652,
    n574
  );


  buf
  g2000
  (
    n1755,
    n950
  );


  buf
  g2001
  (
    n2111,
    n1132
  );


  not
  g2002
  (
    n1852,
    n845
  );


  not
  g2003
  (
    n1881,
    n646
  );


  buf
  g2004
  (
    n2024,
    n859
  );


  not
  g2005
  (
    n1634,
    n571
  );


  buf
  g2006
  (
    n2049,
    n847
  );


  buf
  g2007
  (
    n2151,
    n563
  );


  buf
  g2008
  (
    n1923,
    n701
  );


  not
  g2009
  (
    n2166,
    n844
  );


  buf
  g2010
  (
    n1743,
    n733
  );


  not
  g2011
  (
    n1795,
    n757
  );


  buf
  g2012
  (
    n1841,
    n779
  );


  buf
  g2013
  (
    n2130,
    n799
  );


  buf
  g2014
  (
    n1829,
    n777
  );


  buf
  g2015
  (
    n1630,
    n542
  );


  not
  g2016
  (
    n1900,
    n786
  );


  not
  g2017
  (
    n1716,
    n848
  );


  buf
  g2018
  (
    n1805,
    n826
  );


  buf
  g2019
  (
    n1888,
    n968
  );


  not
  g2020
  (
    n1667,
    n665
  );


  buf
  g2021
  (
    n1908,
    n814
  );


  not
  g2022
  (
    n1963,
    n911
  );


  buf
  g2023
  (
    n1711,
    n1055
  );


  not
  g2024
  (
    n1666,
    n581
  );


  not
  g2025
  (
    n2017,
    n918
  );


  buf
  g2026
  (
    n1797,
    n1015
  );


  not
  g2027
  (
    n2131,
    n983
  );


  not
  g2028
  (
    n1781,
    n781
  );


  not
  g2029
  (
    n1712,
    n654
  );


  buf
  g2030
  (
    n1551,
    n718
  );


  buf
  g2031
  (
    n2032,
    n776
  );


  buf
  g2032
  (
    n1983,
    n873
  );


  not
  g2033
  (
    n1709,
    n545
  );


  buf
  g2034
  (
    n1618,
    n850
  );


  not
  g2035
  (
    n1676,
    n740
  );


  not
  g2036
  (
    n2091,
    n924
  );


  buf
  g2037
  (
    n1914,
    n650
  );


  not
  g2038
  (
    n1886,
    n811
  );


  buf
  g2039
  (
    n1873,
    n578
  );


  not
  g2040
  (
    n1642,
    n992
  );


  buf
  g2041
  (
    n1701,
    n730
  );


  buf
  g2042
  (
    n2176,
    n607
  );


  buf
  g2043
  (
    n1767,
    n981
  );


  not
  g2044
  (
    n1982,
    n532
  );


  buf
  g2045
  (
    n2149,
    n1122
  );


  buf
  g2046
  (
    n1777,
    n1023
  );


  buf
  g2047
  (
    n1661,
    n820
  );


  not
  g2048
  (
    n2100,
    n1069
  );


  not
  g2049
  (
    n1861,
    n1039
  );


  not
  g2050
  (
    n1768,
    n583
  );


  not
  g2051
  (
    n1691,
    n1131
  );


  not
  g2052
  (
    n2048,
    n682
  );


  not
  g2053
  (
    n1972,
    n634
  );


  not
  g2054
  (
    n1742,
    n1124
  );


  buf
  g2055
  (
    n1628,
    n576
  );


  buf
  g2056
  (
    n2066,
    n794
  );


  buf
  g2057
  (
    n1993,
    n1138
  );


  buf
  g2058
  (
    n1713,
    n649
  );


  not
  g2059
  (
    n2061,
    n1112
  );


  not
  g2060
  (
    n1945,
    n679
  );


  buf
  g2061
  (
    n1779,
    n766
  );


  buf
  g2062
  (
    n1604,
    n1127
  );


  buf
  g2063
  (
    n2172,
    n626
  );


  not
  g2064
  (
    n2080,
    n942
  );


  buf
  g2065
  (
    n2115,
    n961
  );


  not
  g2066
  (
    n2075,
    n1125
  );


  buf
  g2067
  (
    n1532,
    n1085
  );


  buf
  g2068
  (
    n1664,
    n1104
  );


  buf
  g2069
  (
    n1927,
    n904
  );


  buf
  g2070
  (
    n1553,
    n976
  );


  buf
  g2071
  (
    n1938,
    n1143
  );


  buf
  g2072
  (
    n1617,
    n704
  );


  not
  g2073
  (
    n2167,
    n852
  );


  not
  g2074
  (
    n1756,
    n956
  );


  buf
  g2075
  (
    n2117,
    n1011
  );


  buf
  g2076
  (
    n1789,
    n741
  );


  buf
  g2077
  (
    n1692,
    n828
  );


  buf
  g2078
  (
    n1569,
    n1010
  );


  not
  g2079
  (
    n1943,
    n608
  );


  buf
  g2080
  (
    n1592,
    n535
  );


  buf
  g2081
  (
    n1765,
    n1000
  );


  not
  g2082
  (
    n1679,
    n705
  );


  buf
  g2083
  (
    n1539,
    n1170
  );


  buf
  g2084
  (
    n1811,
    n547
  );


  buf
  g2085
  (
    n1647,
    n1184
  );


  buf
  g2086
  (
    n1625,
    n936
  );


  buf
  g2087
  (
    n1817,
    n1110
  );


  not
  g2088
  (
    n1769,
    n885
  );


  buf
  g2089
  (
    n1580,
    n737
  );


  buf
  g2090
  (
    n1744,
    n816
  );


  buf
  g2091
  (
    n1936,
    n750
  );


  buf
  g2092
  (
    n1772,
    n883
  );


  not
  g2093
  (
    n1807,
    n686
  );


  not
  g2094
  (
    n1573,
    n606
  );


  not
  g2095
  (
    n1561,
    n1116
  );


  buf
  g2096
  (
    n1686,
    n642
  );


  not
  g2097
  (
    n1998,
    n564
  );


  not
  g2098
  (
    n2064,
    n1095
  );


  buf
  g2099
  (
    n1816,
    n1169
  );


  not
  g2100
  (
    n1794,
    n775
  );


  not
  g2101
  (
    n1653,
    n937
  );


  not
  g2102
  (
    n2022,
    n783
  );


  buf
  g2103
  (
    n1740,
    n801
  );


  not
  g2104
  (
    n2055,
    n567
  );


  buf
  g2105
  (
    n1833,
    n746
  );


  buf
  g2106
  (
    n1576,
    n1135
  );


  not
  g2107
  (
    n1696,
    n505
  );


  not
  g2108
  (
    n1909,
    n738
  );


  buf
  g2109
  (
    n1906,
    n925
  );


  buf
  g2110
  (
    n1924,
    n971
  );


  not
  g2111
  (
    n1526,
    n648
  );


  buf
  g2112
  (
    n1853,
    n619
  );


  not
  g2113
  (
    n1668,
    n510
  );


  buf
  g2114
  (
    n1543,
    n592
  );


  buf
  g2115
  (
    n2140,
    n674
  );


  not
  g2116
  (
    n1547,
    n526
  );


  buf
  g2117
  (
    n1723,
    n964
  );


  buf
  g2118
  (
    n2110,
    n744
  );


  buf
  g2119
  (
    n2128,
    n1128
  );


  buf
  g2120
  (
    n1952,
    n1009
  );


  not
  g2121
  (
    n1942,
    n1003
  );


  buf
  g2122
  (
    n1980,
    n585
  );


  not
  g2123
  (
    n1717,
    n1058
  );


  not
  g2124
  (
    n1681,
    n700
  );


  not
  g2125
  (
    n2029,
    n1088
  );


  not
  g2126
  (
    n1650,
    n994
  );


  not
  g2127
  (
    n2033,
    n1002
  );


  buf
  g2128
  (
    n1745,
    n1081
  );


  buf
  g2129
  (
    n1773,
    n717
  );


  not
  g2130
  (
    n1903,
    n1149
  );


  buf
  g2131
  (
    n1837,
    n1014
  );


  buf
  g2132
  (
    n1814,
    n1106
  );


  buf
  g2133
  (
    n1866,
    n1086
  );


  not
  g2134
  (
    n1639,
    n960
  );


  buf
  g2135
  (
    n1770,
    n537
  );


  buf
  g2136
  (
    n1597,
    n594
  );


  buf
  g2137
  (
    n1855,
    n917
  );


  not
  g2138
  (
    n2000,
    n601
  );


  buf
  g2139
  (
    n2119,
    n959
  );


  not
  g2140
  (
    n1515,
    n915
  );


  buf
  g2141
  (
    n1996,
    n1173
  );


  buf
  g2142
  (
    n1977,
    n572
  );


  not
  g2143
  (
    n1591,
    n546
  );


  buf
  g2144
  (
    n1858,
    n1025
  );


  buf
  g2145
  (
    n1895,
    n827
  );


  buf
  g2146
  (
    n1776,
    n539
  );


  not
  g2147
  (
    n1999,
    n507
  );


  not
  g2148
  (
    n1893,
    n638
  );


  buf
  g2149
  (
    n1785,
    n762
  );


  not
  g2150
  (
    n2089,
    n593
  );


  buf
  g2151
  (
    n1962,
    n877
  );


  not
  g2152
  (
    n2039,
    n833
  );


  buf
  g2153
  (
    n1819,
    n590
  );


  not
  g2154
  (
    n1869,
    n1021
  );


  buf
  g2155
  (
    n1514,
    n628
  );


  buf
  g2156
  (
    n1836,
    n523
  );


  buf
  g2157
  (
    n2047,
    n880
  );


  not
  g2158
  (
    n1574,
    n800
  );


  not
  g2159
  (
    n1577,
    n763
  );


  not
  g2160
  (
    n1907,
    n613
  );


  xnor
  g2161
  (
    n2153,
    n557,
    n824
  );


  xor
  g2162
  (
    n1892,
    n849,
    n980,
    n1137
  );


  nor
  g2163
  (
    n2203,
    n1240,
    n1519,
    n1185,
    n1224
  );


  nand
  g2164
  (
    n2195,
    n1256,
    n1262,
    n1241,
    n1193
  );


  xor
  g2165
  (
    n2206,
    n1242,
    n1189,
    n1192,
    n1206
  );


  xnor
  g2166
  (
    n2193,
    n1217,
    n1536,
    n1253,
    n1235
  );


  nand
  g2167
  (
    n2210,
    n1214,
    n1522,
    n1523,
    n1225
  );


  or
  g2168
  (
    n2191,
    n1228,
    n1520,
    n1254,
    n1209
  );


  xor
  g2169
  (
    n2209,
    n1239,
    n1237,
    n1186,
    n1203
  );


  nand
  g2170
  (
    n2199,
    n1251,
    n1243,
    n1208,
    n1245
  );


  nor
  g2171
  (
    n2211,
    n1516,
    n1215,
    n1238,
    n1533
  );


  and
  g2172
  (
    n2189,
    n1532,
    n1216,
    n1229,
    n1517
  );


  xor
  g2173
  (
    n2204,
    n1223,
    n1202,
    n1227,
    n1236
  );


  nor
  g2174
  (
    n2208,
    n1212,
    n1219,
    n1231,
    n1250
  );


  or
  g2175
  (
    n2192,
    n1201,
    n1518,
    n1515,
    n1257
  );


  or
  g2176
  (
    n2207,
    n1247,
    n1234,
    n1525,
    n1528
  );


  xnor
  g2177
  (
    n2202,
    n1207,
    n1230,
    n1527,
    n1200
  );


  xnor
  g2178
  (
    n2190,
    n1258,
    n1513,
    n1531,
    n1246
  );


  nor
  g2179
  (
    n2188,
    n1260,
    n1511,
    n1226,
    n1220
  );


  or
  g2180
  (
    n2200,
    n1232,
    n1210,
    n1521,
    n1244
  );


  and
  g2181
  (
    n2198,
    n1194,
    n1197,
    n1205,
    n1534
  );


  xnor
  g2182
  (
    n2205,
    n1529,
    n1233,
    n1514,
    n1526
  );


  xor
  g2183
  (
    n2213,
    n1204,
    n1199,
    n1252,
    n1195
  );


  xnor
  g2184
  (
    n2194,
    n1261,
    n1191,
    n1188,
    n1255
  );


  xnor
  g2185
  (
    n2212,
    n1530,
    n1187,
    n1524,
    n1218
  );


  and
  g2186
  (
    n2197,
    n1512,
    n1248,
    n1190,
    n1211
  );


  nand
  g2187
  (
    n2196,
    n1198,
    n1221,
    n1213,
    n1196
  );


  nor
  g2188
  (
    n2201,
    n1535,
    n1222,
    n1259,
    n1249
  );


  not
  g2189
  (
    n2226,
    n1540
  );


  not
  g2190
  (
    n2220,
    n1539
  );


  not
  g2191
  (
    n2224,
    n2191
  );


  not
  g2192
  (
    n2222,
    n1542
  );


  not
  g2193
  (
    n2218,
    n1551
  );


  buf
  g2194
  (
    n2221,
    n1543
  );


  buf
  g2195
  (
    n2217,
    n1549
  );


  not
  g2196
  (
    n2229,
    n2192
  );


  not
  g2197
  (
    n2215,
    n2200
  );


  buf
  g2198
  (
    n2225,
    n2198
  );


  and
  g2199
  (
    n2228,
    n1552,
    n1548
  );


  nand
  g2200
  (
    n2223,
    n1550,
    n2196,
    n1545,
    n2203
  );


  nand
  g2201
  (
    n2219,
    n2195,
    n1547,
    n1546,
    n2199
  );


  nand
  g2202
  (
    n2227,
    n2202,
    n2201,
    n2190,
    n2194
  );


  xnor
  g2203
  (
    n2216,
    n1541,
    n2188,
    n2189,
    n2193
  );


  and
  g2204
  (
    n2214,
    n1544,
    n1537,
    n2197,
    n1538
  );


  and
  g2205
  (
    n2235,
    n1276,
    n1284,
    n1275,
    n1271
  );


  xnor
  g2206
  (
    n2230,
    n1270,
    n1267,
    n1553,
    n1274
  );


  or
  g2207
  (
    n2232,
    n1266,
    n1280,
    n2214,
    n1277
  );


  nand
  g2208
  (
    n2237,
    n1272,
    n1268,
    n1278,
    n1264
  );


  xor
  g2209
  (
    n2234,
    n1282,
    n1281,
    n1263,
    n2215
  );


  or
  g2210
  (
    n2233,
    n1554,
    n2215,
    n1279,
    n2214
  );


  and
  g2211
  (
    n2231,
    n1283,
    n2215,
    n2214,
    n1273
  );


  nand
  g2212
  (
    n2236,
    n2215,
    n1269,
    n1265,
    n2214
  );


  not
  g2213
  (
    n2240,
    n2237
  );


  buf
  g2214
  (
    n2238,
    n1555
  );


  not
  g2215
  (
    n2242,
    n2230
  );


  buf
  g2216
  (
    n2241,
    n1556
  );


  not
  g2217
  (
    n2244,
    n2234
  );


  buf
  g2218
  (
    n2245,
    n2235
  );


  buf
  g2219
  (
    n2239,
    n2231
  );


  xor
  g2220
  (
    n2243,
    n2233,
    n2232,
    n2236
  );


  not
  g2221
  (
    n2247,
    n2238
  );


  not
  g2222
  (
    n2251,
    n2239
  );


  buf
  g2223
  (
    n2249,
    n2239
  );


  buf
  g2224
  (
    n2250,
    n2241
  );


  not
  g2225
  (
    n2246,
    n2240
  );


  buf
  g2226
  (
    n2248,
    n2240
  );


  nor
  g2227
  (
    n2254,
    n2246,
    n2221,
    n2249,
    n2247
  );


  xnor
  g2228
  (
    n2253,
    n2217,
    n2220,
    n1293,
    n2224
  );


  nand
  g2229
  (
    n2274,
    n1559,
    n2223,
    n2221,
    n1289
  );


  nor
  g2230
  (
    n2256,
    n2216,
    n2248,
    n2217,
    n2226
  );


  or
  g2231
  (
    n2267,
    n2224,
    n2246,
    n2216,
    n2218
  );


  nand
  g2232
  (
    n2259,
    n1562,
    n2250,
    n2251
  );


  xnor
  g2233
  (
    n2265,
    n2226,
    n2223,
    n2227,
    n2247
  );


  nor
  g2234
  (
    n2266,
    n2221,
    n1561,
    n2220,
    n2227
  );


  nor
  g2235
  (
    n2258,
    n2216,
    n2224,
    n2249,
    n2251
  );


  and
  g2236
  (
    n2257,
    n2226,
    n1287,
    n2225,
    n2218
  );


  xnor
  g2237
  (
    n2268,
    n2204,
    n2251,
    n1290,
    n2225
  );


  xnor
  g2238
  (
    n2263,
    n2219,
    n2219,
    n2217,
    n2221
  );


  nand
  g2239
  (
    n2273,
    n1560,
    n1285,
    n2208,
    n2248
  );


  nor
  g2240
  (
    n2262,
    n2222,
    n1557,
    n2247,
    n2219
  );


  and
  g2241
  (
    n2260,
    n2216,
    n2222,
    n2223,
    n2250
  );


  xnor
  g2242
  (
    n2272,
    n2248,
    n1563,
    n2207,
    n2222
  );


  xnor
  g2243
  (
    n2271,
    n2219,
    n2227,
    n2223,
    n1566
  );


  nand
  g2244
  (
    n2255,
    n2217,
    n1286,
    n2218,
    n1565
  );


  xor
  g2245
  (
    n2269,
    n2224,
    n1564,
    n2249,
    n2218
  );


  xnor
  g2246
  (
    n2270,
    n2206,
    n1291,
    n2205,
    n2251
  );


  xor
  g2247
  (
    KeyWire_0_1,
    n2250,
    n2249,
    n2247,
    n2209
  );


  nand
  g2248
  (
    n2252,
    n1558,
    n2246,
    n1288,
    n1292
  );


  or
  g2249
  (
    n2275,
    n2222,
    n2246,
    n2248,
    n2225
  );


  nand
  g2250
  (
    n2264,
    n2220,
    n2220,
    n2225,
    n2226
  );


  or
  g2251
  (
    n2276,
    n2252,
    n1567,
    n1568,
    n1569
  );


  or
  g2252
  (
    n2278,
    n1571,
    n2276,
    n1574
  );


  nand
  g2253
  (
    n2277,
    n1575,
    n1572,
    n1573,
    n1570
  );


  buf
  g2254
  (
    n2286,
    n2277
  );


  not
  g2255
  (
    n2283,
    n1297
  );


  not
  g2256
  (
    n2285,
    n1301
  );


  not
  g2257
  (
    n2281,
    n2278
  );


  not
  g2258
  (
    n2284,
    n2278
  );


  or
  g2259
  (
    n2279,
    n1296,
    n2278,
    n1294
  );


  nand
  g2260
  (
    n2282,
    n1300,
    n1295,
    n2277
  );


  and
  g2261
  (
    n2280,
    n1299,
    n2277,
    n1298,
    n2278
  );


  xnor
  g2262
  (
    n2288,
    n1576,
    n1580,
    n1583,
    n1579
  );


  and
  g2263
  (
    n2287,
    n2280,
    n1584,
    n1582,
    n1578
  );


  or
  g2264
  (
    n2289,
    n1581,
    n1577,
    n2279,
    n2281
  );


  not
  g2265
  (
    n2294,
    n2288
  );


  not
  g2266
  (
    n2290,
    n2288
  );


  buf
  g2267
  (
    n2295,
    n2287
  );


  buf
  g2268
  (
    n2292,
    n2288
  );


  buf
  g2269
  (
    n2293,
    n2253
  );


  nor
  g2270
  (
    n2291,
    n2288,
    n1585,
    n2289,
    n1586
  );


  nand
  g2271
  (
    n2296,
    n502,
    n1309,
    n1587,
    n503
  );


  xnor
  g2272
  (
    n2301,
    n2293,
    n2295,
    n503
  );


  and
  g2273
  (
    n2300,
    n502,
    n2292,
    n1306,
    n1307
  );


  nand
  g2274
  (
    n2299,
    n2291,
    n2294,
    n1310,
    n502
  );


  xnor
  g2275
  (
    n2298,
    n1588,
    n502,
    n1304,
    n1308
  );


  xnor
  g2276
  (
    n2297,
    n1305,
    n1302,
    n1303,
    n2290
  );


  buf
  g2277
  (
    n2306,
    n2300
  );


  not
  g2278
  (
    n2310,
    n2299
  );


  buf
  g2279
  (
    n2315,
    n2301
  );


  buf
  g2280
  (
    n2309,
    n2300
  );


  buf
  g2281
  (
    n2316,
    n2299
  );


  buf
  g2282
  (
    n2308,
    n2301
  );


  buf
  g2283
  (
    n2312,
    n2301
  );


  not
  g2284
  (
    n2304,
    n2296
  );


  buf
  g2285
  (
    n2305,
    n2299
  );


  buf
  g2286
  (
    n2314,
    n2300
  );


  buf
  g2287
  (
    n2307,
    n2297
  );


  not
  g2288
  (
    n2313,
    n2299
  );


  buf
  g2289
  (
    n2303,
    n2301
  );


  buf
  g2290
  (
    n2302,
    n1311
  );


  nor
  g2291
  (
    n2311,
    n2300,
    n2298
  );


  buf
  g2292
  (
    n2317,
    n2302
  );


  buf
  g2293
  (
    n2318,
    n2303
  );


  xnor
  g2294
  (
    n2319,
    n1591,
    n1589,
    n2318,
    n1590
  );


  nand
  g2295
  (
    n2323,
    n1602,
    n1594,
    n1598,
    n1593
  );


  xnor
  g2296
  (
    n2320,
    n1595,
    n1600,
    n1601,
    n2319
  );


  xnor
  g2297
  (
    n2321,
    n1592,
    n2319,
    n1597
  );


  xnor
  g2298
  (
    n2322,
    n1599,
    n2319,
    n1596,
    n1603
  );


  buf
  g2299
  (
    KeyWire_0_2,
    n2323
  );


  not
  g2300
  (
    n2325,
    n2323
  );


  not
  g2301
  (
    KeyWire_0_9,
    n2320
  );


  buf
  g2302
  (
    n2328,
    n2323
  );


  buf
  g2303
  (
    n2327,
    n2322
  );


  not
  g2304
  (
    n2331,
    n2321
  );


  not
  g2305
  (
    n2324,
    n2323
  );


  and
  g2306
  (
    n2330,
    n2322,
    n1605,
    n1604
  );


  xor
  g2307
  (
    n2333,
    n2327,
    n2305,
    n2324,
    n2308
  );


  nand
  g2308
  (
    n2344,
    n2309,
    n2311,
    n1614,
    n2325
  );


  and
  g2309
  (
    n2336,
    n2312,
    n1615,
    n2308,
    n2306
  );


  nor
  g2310
  (
    n2346,
    n1616,
    n2310,
    n2307,
    n2326
  );


  xor
  g2311
  (
    n2340,
    n2311,
    n2308,
    n2326
  );


  xor
  g2312
  (
    n2335,
    n2325,
    n2324,
    n1610,
    n1608
  );


  xor
  g2313
  (
    n2339,
    n2327,
    n2309,
    n2310,
    n1612
  );


  or
  g2314
  (
    n2338,
    n2327,
    n1619,
    n2312,
    n2313
  );


  xor
  g2315
  (
    n2342,
    n2306,
    n2310,
    n1620,
    n1618
  );


  xor
  g2316
  (
    n2332,
    n2307,
    n2309,
    n2325,
    n2313
  );


  nor
  g2317
  (
    n2341,
    n2312,
    n2326,
    n1617,
    n2308
  );


  and
  g2318
  (
    n2334,
    n2310,
    n2325,
    n1613,
    n2311
  );


  nand
  g2319
  (
    n2345,
    n2304,
    n2307,
    n1611
  );


  nand
  g2320
  (
    n2343,
    n1606,
    n2309,
    n1609,
    n1607
  );


  nand
  g2321
  (
    n2337,
    n2311,
    n2324,
    n2312
  );


  nor
  g2322
  (
    n2350,
    n1626,
    n1629,
    n2342,
    n1630
  );


  xor
  g2323
  (
    n2348,
    n1621,
    n1624,
    n1627,
    n2341
  );


  and
  g2324
  (
    n2347,
    n1631,
    n2339,
    n2340,
    n1622
  );


  nor
  g2325
  (
    n2349,
    n1623,
    n1632,
    n1625,
    n1628
  );


  buf
  g2326
  (
    n2355,
    n2245
  );


  not
  g2327
  (
    n2360,
    n2289
  );


  nor
  g2328
  (
    n2356,
    n2314,
    n2289
  );


  nor
  g2329
  (
    n2352,
    n1633,
    n1639,
    n2345,
    n2349
  );


  xnor
  g2330
  (
    n2361,
    n2343,
    n2348,
    n2242
  );


  xnor
  g2331
  (
    n2354,
    n2241,
    n2313,
    n1638,
    n1636
  );


  and
  g2332
  (
    n2358,
    n2244,
    n2313,
    n2349,
    n2346
  );


  or
  g2333
  (
    n2351,
    n2347,
    n2243,
    n1637,
    n2348
  );


  xnor
  g2334
  (
    n2359,
    n2347,
    n1634,
    n2350
  );


  nand
  g2335
  (
    n2357,
    n2243,
    n1635,
    n2314,
    n2350
  );


  xnor
  g2336
  (
    n2353,
    n2244,
    n1640,
    n2289,
    n2349
  );


  nand
  g2337
  (
    n2362,
    n2350,
    n2344,
    n2245,
    n2349
  );


  not
  g2338
  (
    n2379,
    n2329
  );


  not
  g2339
  (
    n2389,
    n2360
  );


  not
  g2340
  (
    n2375,
    n2316
  );


  buf
  g2341
  (
    n2401,
    n2329
  );


  buf
  g2342
  (
    n2378,
    n2351
  );


  buf
  g2343
  (
    n2395,
    n2360
  );


  not
  g2344
  (
    n2388,
    n2228
  );


  buf
  g2345
  (
    n2392,
    n2361
  );


  not
  g2346
  (
    n2391,
    n2259
  );


  buf
  g2347
  (
    n2372,
    n2264
  );


  buf
  g2348
  (
    n2364,
    n2331
  );


  not
  g2349
  (
    n2410,
    n2358
  );


  buf
  g2350
  (
    n2405,
    n2354
  );


  not
  g2351
  (
    n2382,
    n1312
  );


  not
  g2352
  (
    n2402,
    n2257
  );


  not
  g2353
  (
    n2376,
    n2357
  );


  not
  g2354
  (
    n2366,
    n2352
  );


  buf
  g2355
  (
    n2371,
    n2331
  );


  buf
  g2356
  (
    n2394,
    n2355
  );


  not
  g2357
  (
    n2365,
    n2265
  );


  not
  g2358
  (
    n2399,
    n2228
  );


  not
  g2359
  (
    n2369,
    n1320
  );


  buf
  g2360
  (
    n2368,
    n2353
  );


  buf
  g2361
  (
    n2404,
    n2355
  );


  not
  g2362
  (
    n2367,
    n2355
  );


  buf
  g2363
  (
    n2400,
    n2356
  );


  buf
  g2364
  (
    n2393,
    n2352
  );


  not
  g2365
  (
    n2387,
    n2358
  );


  not
  g2366
  (
    n2390,
    n2357
  );


  xnor
  g2367
  (
    n2396,
    n2261,
    n2355,
    n1318,
    n2316
  );


  and
  g2368
  (
    n2408,
    n2356,
    n2260,
    n2227,
    n2360
  );


  nand
  g2369
  (
    n2385,
    n2361,
    n2358,
    n1315,
    n2328
  );


  nor
  g2370
  (
    n2407,
    n2360,
    n2330,
    n2315
  );


  xor
  g2371
  (
    n2373,
    n1323,
    n2351,
    n2359,
    n2354
  );


  xnor
  g2372
  (
    n2406,
    n2359,
    n2315,
    n2254,
    n2316
  );


  xnor
  g2373
  (
    n2397,
    n2314,
    n2362,
    n2330
  );


  xor
  g2374
  (
    n2383,
    n2357,
    n2359,
    n2353,
    n2354
  );


  nand
  g2375
  (
    n2398,
    n2330,
    n2327,
    n2263,
    n1314
  );


  nor
  g2376
  (
    n2363,
    n1324,
    n2362,
    n2358,
    n1321
  );


  xor
  g2377
  (
    n2384,
    n2361,
    n2316,
    n2353,
    n2330
  );


  and
  g2378
  (
    n2370,
    n2329,
    n2328,
    n1317
  );


  or
  g2379
  (
    n2409,
    n2328,
    n2351,
    n2352,
    n2353
  );


  xnor
  g2380
  (
    n2374,
    n1316,
    n2331,
    n2228,
    n2356
  );


  and
  g2381
  (
    n2381,
    n2255,
    n2362,
    n2258,
    n2315
  );


  xnor
  g2382
  (
    n2380,
    n2228,
    n1313,
    n2359,
    n2357
  );


  xor
  g2383
  (
    n2377,
    n2361,
    n2262,
    n2314,
    n2329
  );


  and
  g2384
  (
    n2403,
    n2351,
    n2331,
    n2354,
    n1322
  );


  and
  g2385
  (
    n2386,
    n2352,
    n1319,
    n2356,
    n2256
  );


  buf
  g2386
  (
    n2414,
    n1647
  );


  buf
  g2387
  (
    n2416,
    n1643
  );


  not
  g2388
  (
    n2418,
    n2363
  );


  buf
  g2389
  (
    n2413,
    n2364
  );


  buf
  g2390
  (
    n2412,
    n1644
  );


  buf
  g2391
  (
    n2415,
    n2364
  );


  or
  g2392
  (
    n2417,
    n2364,
    n1641
  );


  or
  g2393
  (
    n2419,
    n2365,
    n2364,
    n1646,
    n1645
  );


  xnor
  g2394
  (
    n2411,
    n1642,
    n2363
  );


  nand
  g2395
  (
    n2447,
    n2414,
    n1415,
    n1370,
    n1336
  );


  or
  g2396
  (
    n2448,
    n1426,
    n1423,
    n1382,
    n2416
  );


  nand
  g2397
  (
    n2435,
    n1332,
    n1425,
    n2415,
    n2413
  );


  xor
  g2398
  (
    n2453,
    n1363,
    n1394,
    n1343,
    n1325
  );


  xnor
  g2399
  (
    n2443,
    n1338,
    n1391,
    n1388,
    n2413
  );


  xnor
  g2400
  (
    n2430,
    n1403,
    n2419,
    n1352,
    n1376
  );


  nor
  g2401
  (
    n2445,
    n1422,
    n1354,
    n1371,
    n1372
  );


  xor
  g2402
  (
    n2424,
    n1355,
    n1331,
    n1412,
    n1359
  );


  or
  g2403
  (
    n2454,
    n2412,
    n1353,
    n2411,
    n1367
  );


  and
  g2404
  (
    n2437,
    n2417,
    n1328,
    n1345,
    n1360
  );


  and
  g2405
  (
    n2420,
    n2414,
    n2415,
    n1361,
    n1383
  );


  nand
  g2406
  (
    n2440,
    n2419,
    n1421,
    n1365,
    n1329
  );


  xor
  g2407
  (
    n2432,
    n1402,
    n1396,
    n1347,
    n1387
  );


  nand
  g2408
  (
    n2421,
    n1362,
    n1334,
    n1418,
    n1405
  );


  xnor
  g2409
  (
    n2423,
    n1335,
    n2418,
    n1648,
    n2413
  );


  and
  g2410
  (
    n2442,
    n1397,
    n1420,
    n1377,
    n1404
  );


  xor
  g2411
  (
    n2438,
    n1375,
    n1385,
    n1400,
    n2413
  );


  and
  g2412
  (
    n2439,
    n1411,
    n1340,
    n1337,
    n1374
  );


  nor
  g2413
  (
    n2441,
    n1409,
    n1401,
    n2412,
    n1414
  );


  and
  g2414
  (
    n2451,
    n1390,
    n1379,
    n2412,
    n1330
  );


  or
  g2415
  (
    n2444,
    n1398,
    n1339,
    n1384,
    n1381
  );


  xnor
  g2416
  (
    n2431,
    n1358,
    n1351,
    n1356,
    n1380
  );


  or
  g2417
  (
    n2426,
    n1364,
    n2415,
    n2419
  );


  nand
  g2418
  (
    n2450,
    n1389,
    n1327,
    n2416,
    n1410
  );


  xnor
  g2419
  (
    n2433,
    n2417,
    n2416,
    n1392,
    n2414
  );


  nand
  g2420
  (
    n2452,
    n1393,
    n2419,
    n2418,
    n1357
  );


  or
  g2421
  (
    n2422,
    n1395,
    n1341,
    n1368,
    n1416
  );


  xnor
  g2422
  (
    n2436,
    n1350,
    n1386,
    n1399,
    n1348
  );


  nand
  g2423
  (
    n2446,
    n2417,
    n1373,
    n1333,
    n1424
  );


  xor
  g2424
  (
    n2425,
    n1326,
    n1369,
    n1417,
    n1419
  );


  nand
  g2425
  (
    n2429,
    n1349,
    n1408,
    n1649,
    n2412
  );


  xnor
  g2426
  (
    n2434,
    n1344,
    n2411,
    n2418,
    n1413
  );


  and
  g2427
  (
    n2427,
    n2417,
    n2416,
    n1378,
    n2414
  );


  or
  g2428
  (
    n2428,
    n2418,
    n1407,
    n1346,
    n1366
  );


  and
  g2429
  (
    n2449,
    n1406,
    n1427,
    n1342,
    n2411
  );


  or
  g2430
  (
    n2527,
    n1807,
    n2066,
    n1873,
    n1826
  );


  nor
  g2431
  (
    n2546,
    n1805,
    n2434,
    n2027,
    n1698
  );


  xnor
  g2432
  (
    n2468,
    n1985,
    n2062,
    n1817,
    n1750
  );


  nor
  g2433
  (
    n2551,
    n1997,
    n1990,
    n1661,
    n1762
  );


  or
  g2434
  (
    n2493,
    n1676,
    n2454,
    n2428,
    n1917
  );


  or
  g2435
  (
    n2487,
    n1948,
    n2444,
    n1766,
    n2448
  );


  xnor
  g2436
  (
    n2514,
    n2426,
    n2432,
    n2048,
    n1881
  );


  nor
  g2437
  (
    n2469,
    n1979,
    n1884,
    n1687,
    n2019
  );


  and
  g2438
  (
    n2582,
    n2437,
    n2055,
    n2426,
    n1658
  );


  and
  g2439
  (
    n2566,
    n1895,
    n2449,
    n2441,
    n2049
  );


  xnor
  g2440
  (
    n2494,
    n2449,
    n2030,
    n1671,
    n2025
  );


  nand
  g2441
  (
    n2489,
    n2420,
    n1994,
    n1988,
    n2001
  );


  and
  g2442
  (
    n2565,
    n1885,
    n1823,
    n1670,
    n2008
  );


  nor
  g2443
  (
    n2547,
    n1704,
    n2440,
    n2420,
    n1935
  );


  nand
  g2444
  (
    n2530,
    n1838,
    n1853,
    n2015,
    n1865
  );


  or
  g2445
  (
    n2545,
    n1755,
    n1840,
    n2445,
    n2064
  );


  and
  g2446
  (
    n2492,
    n1953,
    n1975,
    n2431,
    n2043
  );


  nor
  g2447
  (
    n2584,
    n1947,
    n2045,
    n1797,
    n1915
  );


  or
  g2448
  (
    n2539,
    n1996,
    n1950,
    n1713,
    n1850
  );


  xor
  g2449
  (
    n2560,
    n2441,
    n1773,
    n2436,
    n2423
  );


  and
  g2450
  (
    n2553,
    n1705,
    n1856,
    n1841,
    n1673
  );


  nand
  g2451
  (
    n2456,
    n1694,
    n1710,
    n1706,
    n1714
  );


  nand
  g2452
  (
    n2464,
    n1857,
    n2440,
    n1943,
    n1683
  );


  xnor
  g2453
  (
    n2515,
    n1688,
    n2052,
    n1686,
    n1842
  );


  xnor
  g2454
  (
    n2569,
    n1782,
    n2439,
    n1723,
    n1677
  );


  and
  g2455
  (
    n2471,
    n1928,
    n1690,
    n2420,
    n1656
  );


  xor
  g2456
  (
    n2544,
    n2431,
    n1769,
    n1837,
    n2424
  );


  nand
  g2457
  (
    n2571,
    n2446,
    n1811,
    n1911,
    n1794
  );


  nor
  g2458
  (
    n2513,
    n1651,
    n1680,
    n1736,
    n2438
  );


  xnor
  g2459
  (
    n2522,
    n1810,
    n2451,
    n1982,
    n2444
  );


  xor
  g2460
  (
    n2533,
    n1814,
    n2447,
    n1945,
    n1664
  );


  or
  g2461
  (
    n2574,
    n1939,
    n2450,
    n2426,
    n1844
  );


  and
  g2462
  (
    n2506,
    n1920,
    n1708,
    n2421,
    n2423
  );


  and
  g2463
  (
    n2490,
    n1696,
    n1900,
    n2449,
    n2054
  );


  xnor
  g2464
  (
    n2555,
    n1685,
    n1772,
    n1699,
    n1695
  );


  xnor
  g2465
  (
    n2465,
    n2423,
    n1854,
    n1936,
    n2425
  );


  xnor
  g2466
  (
    n2585,
    n2431,
    n2434,
    n1828,
    n2420
  );


  and
  g2467
  (
    n2495,
    n1754,
    n1851,
    n2021,
    n1944
  );


  nor
  g2468
  (
    n2556,
    n2427,
    n1733,
    n2442,
    n2429
  );


  nand
  g2469
  (
    n2531,
    n1940,
    n2447,
    n2453,
    n2005
  );


  nand
  g2470
  (
    n2589,
    n2046,
    n1894,
    n2428,
    n1720
  );


  nor
  g2471
  (
    n2526,
    n2450,
    n1877,
    n2443,
    n1795
  );


  xor
  g2472
  (
    n2519,
    n1995,
    n1784,
    n1816,
    n1801
  );


  and
  g2473
  (
    n2482,
    n2426,
    n2422,
    n1919,
    n2435
  );


  nor
  g2474
  (
    n2557,
    n1971,
    n1959,
    n2429,
    n1702
  );


  nor
  g2475
  (
    n2475,
    n2423,
    n1880,
    n2451,
    n1813
  );


  and
  g2476
  (
    n2525,
    n1672,
    n1740,
    n1675,
    n1764
  );


  and
  g2477
  (
    n2477,
    n2433,
    n2026,
    n2436,
    n2443
  );


  or
  g2478
  (
    n2499,
    n1781,
    n1993,
    n2430,
    n1765
  );


  or
  g2479
  (
    n2587,
    n1727,
    n2439,
    n2437,
    n2452
  );


  xor
  g2480
  (
    n2481,
    n1679,
    n1663,
    n1904,
    n2454
  );


  xnor
  g2481
  (
    n2541,
    n2056,
    n1768,
    n2037,
    n1689
  );


  nand
  g2482
  (
    n2550,
    n2422,
    n1752,
    n1902,
    n1753
  );


  xor
  g2483
  (
    n2516,
    n1961,
    n1745,
    n2443,
    n1822
  );


  nand
  g2484
  (
    n2507,
    n2433,
    n1930,
    n1654,
    n1949
  );


  or
  g2485
  (
    n2488,
    n2042,
    n1725,
    n2442,
    n1785
  );


  nand
  g2486
  (
    n2592,
    n2435,
    n2446,
    n1748,
    n1650
  );


  nor
  g2487
  (
    n2503,
    n1815,
    n1831,
    n2035,
    n2040
  );


  or
  g2488
  (
    n2578,
    n1927,
    n1820,
    n1759,
    n1786
  );


  xor
  g2489
  (
    n2501,
    n1845,
    n1984,
    n1863,
    n1788
  );


  xnor
  g2490
  (
    n2559,
    n2422,
    n2439,
    n2067,
    n1757
  );


  nor
  g2491
  (
    n2542,
    n1825,
    n2029,
    n1747,
    n1843
  );


  xor
  g2492
  (
    n2461,
    n2009,
    n2444,
    n2068,
    n1923
  );


  xnor
  g2493
  (
    n2496,
    n1749,
    n1778,
    n1861,
    n2041
  );


  nor
  g2494
  (
    n2567,
    n2016,
    n2058,
    n1867,
    n1775
  );


  and
  g2495
  (
    n2480,
    n1972,
    n1709,
    n1712,
    n1933
  );


  nand
  g2496
  (
    n2458,
    n1730,
    n1721,
    n1770,
    n1962
  );


  nor
  g2497
  (
    n2534,
    n1887,
    n2428,
    n2440,
    n1839
  );


  or
  g2498
  (
    n2593,
    n1889,
    n2443,
    n2432,
    n1925
  );


  or
  g2499
  (
    n2467,
    n1716,
    n1934,
    n1724,
    n1942
  );


  xor
  g2500
  (
    n2535,
    n2060,
    n1906,
    n1806,
    n2427
  );


  or
  g2501
  (
    n2564,
    n2051,
    n2039,
    n1803,
    n1783
  );


  nand
  g2502
  (
    n2529,
    n1901,
    n2429,
    n2063,
    n2424
  );


  nor
  g2503
  (
    n2504,
    n2454,
    n1715,
    n1876,
    n1976
  );


  xnor
  g2504
  (
    n2581,
    n2424,
    n1666,
    n2447,
    n2453
  );


  xnor
  g2505
  (
    n2479,
    n2448,
    n1946,
    n1913,
    n1978
  );


  or
  g2506
  (
    n2500,
    n1711,
    n1678,
    n1869,
    n1921
  );


  or
  g2507
  (
    n2509,
    n2428,
    n1956,
    n2452,
    n2427
  );


  and
  g2508
  (
    n2491,
    n1732,
    n2448,
    n1892,
    n1868
  );


  and
  g2509
  (
    n2511,
    n1792,
    n2032,
    n1728,
    n1891
  );


  xnor
  g2510
  (
    n2562,
    n1717,
    n2000,
    n2430,
    n1790
  );


  nand
  g2511
  (
    n2497,
    n1722,
    n1860,
    n1726,
    n2431
  );


  nor
  g2512
  (
    n2575,
    n1729,
    n1739,
    n1804,
    n1970
  );


  nand
  g2513
  (
    n2460,
    n2421,
    n1987,
    n2050,
    n1991
  );


  nor
  g2514
  (
    n2548,
    n1776,
    n1818,
    n1693,
    n1875
  );


  nor
  g2515
  (
    n2486,
    n1737,
    n1898,
    n1878,
    n1761
  );


  and
  g2516
  (
    n2517,
    n1703,
    n1893,
    n2441,
    n1924
  );


  xnor
  g2517
  (
    n2466,
    n1809,
    n1779,
    n1829,
    n1660
  );


  xnor
  g2518
  (
    n2576,
    n2028,
    n1771,
    n2444,
    n2449
  );


  nor
  g2519
  (
    KeyWire_0_3,
    n1888,
    n1914,
    n2442,
    n1731
  );


  xor
  g2520
  (
    n2570,
    n2425,
    n1833,
    n1741,
    n2069
  );


  xnor
  g2521
  (
    n2508,
    n2038,
    n2447,
    n2433,
    n1932
  );


  and
  g2522
  (
    n2518,
    n2452,
    n2438,
    n2006,
    n1966
  );


  xnor
  g2523
  (
    n2591,
    n1986,
    n2014,
    n2433,
    n2010
  );


  and
  g2524
  (
    n2577,
    n1981,
    n1789,
    n1952,
    n2013
  );


  xor
  g2525
  (
    n2573,
    n1760,
    n2435,
    n1738,
    n1954
  );


  xor
  g2526
  (
    n2552,
    n1667,
    n1791,
    n1758,
    n1866
  );


  nor
  g2527
  (
    n2470,
    n1998,
    n2020,
    n2017,
    n1964
  );


  nand
  g2528
  (
    n2538,
    n1653,
    n2434,
    n2435,
    n2011
  );


  or
  g2529
  (
    n2561,
    n1903,
    n1969,
    n2429,
    n1707
  );


  xnor
  g2530
  (
    n2590,
    n2427,
    n2434,
    n1787,
    n1659
  );


  nand
  g2531
  (
    n2523,
    n1951,
    n1852,
    n2439,
    n1846
  );


  nand
  g2532
  (
    n2485,
    n2012,
    n1744,
    n2036,
    n1958
  );


  and
  g2533
  (
    n2543,
    n2445,
    n2436,
    n1941,
    n1965
  );


  nor
  g2534
  (
    n2583,
    n2437,
    n2033,
    n1774,
    n1780
  );


  and
  g2535
  (
    n2528,
    n1798,
    n1821,
    n1938,
    n2061
  );


  xnor
  g2536
  (
    n2594,
    n2453,
    n1929,
    n1960,
    n1682
  );


  or
  g2537
  (
    n2502,
    n1871,
    n1834,
    n2450,
    n1872
  );


  xor
  g2538
  (
    n2462,
    n2441,
    n1910,
    n1848,
    n1886
  );


  or
  g2539
  (
    n2512,
    n1973,
    n1692,
    n1691,
    n1669
  );


  xnor
  g2540
  (
    n2588,
    n2057,
    n1908,
    n2421,
    n1808
  );


  or
  g2541
  (
    n2484,
    n1800,
    n2446,
    n1718,
    n1937
  );


  xor
  g2542
  (
    n2457,
    n1796,
    n2432,
    n2422,
    n1684
  );


  or
  g2543
  (
    n2498,
    n2425,
    n2448,
    n2004,
    n1743
  );


  or
  g2544
  (
    n2455,
    n1883,
    n2059,
    n1742,
    n1767
  );


  nor
  g2545
  (
    n2537,
    n1899,
    n1862,
    n1999,
    n2425
  );


  nand
  g2546
  (
    n2521,
    n1916,
    n2432,
    n2430,
    n2454
  );


  and
  g2547
  (
    n2540,
    n1793,
    n1751,
    n2445,
    n2421
  );


  xor
  g2548
  (
    n2520,
    n2442,
    n2024,
    n2445,
    n1652
  );


  xnor
  g2549
  (
    n2558,
    n1897,
    n1734,
    n2023,
    n1858
  );


  and
  g2550
  (
    n2473,
    n2446,
    n1657,
    n1668,
    n1830
  );


  xor
  g2551
  (
    n2474,
    n1701,
    n1827,
    n1980,
    n2453
  );


  xnor
  g2552
  (
    n2580,
    n2451,
    n1746,
    n1922,
    n1662
  );


  nand
  g2553
  (
    n2463,
    n2440,
    n2034,
    n1874,
    n1931
  );


  or
  g2554
  (
    n2536,
    n1864,
    n1957,
    n1879,
    n1674
  );


  nor
  g2555
  (
    n2568,
    n1989,
    n1835,
    n1907,
    n2044
  );


  nand
  g2556
  (
    n2579,
    n1665,
    n2018,
    n1847,
    n1832
  );


  nor
  g2557
  (
    n2483,
    n1909,
    n2438,
    n2002,
    n1890
  );


  xnor
  g2558
  (
    n2532,
    n1849,
    n1812,
    n1992,
    n1926
  );


  xor
  g2559
  (
    n2554,
    n2022,
    n1697,
    n1655,
    n1824
  );


  xor
  g2560
  (
    n2472,
    n2065,
    n1756,
    n2053,
    n2031
  );


  nor
  g2561
  (
    n2510,
    n2436,
    n2437,
    n1977,
    n1870
  );


  or
  g2562
  (
    n2478,
    n1700,
    n1968,
    n1719,
    n1763
  );


  xnor
  g2563
  (
    n2524,
    n2452,
    n1681,
    n1777,
    n1802
  );


  and
  g2564
  (
    n2505,
    n1819,
    n2007,
    n1859,
    n2438
  );


  xnor
  g2565
  (
    n2586,
    n2430,
    n1836,
    n2047,
    n1963
  );


  or
  g2566
  (
    n2476,
    n1974,
    n1896,
    n1918,
    n2450
  );


  nor
  g2567
  (
    n2563,
    n1905,
    n2424,
    n1983,
    n1855
  );


  and
  g2568
  (
    n2572,
    n1882,
    n1735,
    n1799,
    n2451
  );


  nor
  g2569
  (
    n2549,
    n1912,
    n2003,
    n1955,
    n1967
  );


  or
  g2570
  (
    n2673,
    n2408,
    n504,
    n2410,
    n2366
  );


  xnor
  g2571
  (
    n2677,
    n2371,
    n2482,
    n2384,
    n2080
  );


  nor
  g2572
  (
    n2617,
    n2374,
    n504,
    n2286,
    n2409
  );


  or
  g2573
  (
    n2653,
    n2402,
    n2384,
    n2532,
    n2393
  );


  and
  g2574
  (
    n2656,
    n2481,
    n2398,
    n2491,
    n2559
  );


  and
  g2575
  (
    n2663,
    n2388,
    n2211,
    n2373,
    n2528
  );


  or
  g2576
  (
    n2619,
    n2394,
    n2387,
    n2384,
    n2373
  );


  xor
  g2577
  (
    n2675,
    n2377,
    n2383,
    n2370,
    n2561
  );


  nand
  g2578
  (
    n2651,
    n2524,
    n2409,
    n2390,
    n2283
  );


  xnor
  g2579
  (
    n2602,
    n2538,
    n2375,
    n2378,
    n2560
  );


  nor
  g2580
  (
    n2645,
    n2510,
    n2391,
    n2272,
    n2533
  );


  xnor
  g2581
  (
    n2622,
    n2398,
    n2381,
    n2475,
    n2462
  );


  xnor
  g2582
  (
    n2625,
    n2525,
    n2398,
    n2404,
    n2507
  );


  nor
  g2583
  (
    n2638,
    n2271,
    n2368,
    n2083,
    n2549
  );


  xor
  g2584
  (
    n2628,
    n2553,
    n2076,
    n2397,
    n2212
  );


  or
  g2585
  (
    n2642,
    n2275,
    n2485,
    n2390,
    n2499
  );


  and
  g2586
  (
    n2606,
    n2455,
    n2492,
    n2405,
    n2512
  );


  nor
  g2587
  (
    n2652,
    n2391,
    n2405,
    n2369,
    n2410
  );


  xor
  g2588
  (
    n2624,
    n2369,
    n2367,
    n2518,
    n2557
  );


  xnor
  g2589
  (
    n2640,
    n2484,
    n2213,
    n2519,
    n2400
  );


  nand
  g2590
  (
    n2665,
    n2380,
    n2456,
    n2374,
    n2282
  );


  nor
  g2591
  (
    n2639,
    n2269,
    n2408,
    n2526,
    n2078
  );


  xor
  g2592
  (
    n2613,
    n2371,
    n2377,
    n2410,
    n2275
  );


  nand
  g2593
  (
    n2659,
    n2494,
    n2395,
    n2383,
    n2378
  );


  xnor
  g2594
  (
    n2644,
    n2473,
    n2376,
    n2385,
    n2465
  );


  nand
  g2595
  (
    n2603,
    n2464,
    n2477,
    n2389,
    n2368
  );


  xor
  g2596
  (
    KeyWire_0_13,
    n2393,
    n2550,
    n2389,
    n2551
  );


  xnor
  g2597
  (
    n2616,
    n2382,
    n2070,
    n2558,
    n2400
  );


  and
  g2598
  (
    n2671,
    n2367,
    n2389,
    n2071,
    n2383
  );


  xor
  g2599
  (
    n2598,
    n2372,
    n2527,
    n2365,
    n2381
  );


  and
  g2600
  (
    n2608,
    n2394,
    n2377,
    n2268,
    n2483
  );


  xnor
  g2601
  (
    n2636,
    n2390,
    n2081,
    n2505,
    n2509
  );


  xor
  g2602
  (
    n2650,
    n2273,
    n2379,
    n2395
  );


  or
  g2603
  (
    n2662,
    n2409,
    n2471,
    n2404,
    n2385
  );


  nor
  g2604
  (
    n2672,
    n2410,
    n2072,
    n2403,
    n2474
  );


  or
  g2605
  (
    n2655,
    n2391,
    n2365,
    n2370,
    n2385
  );


  nand
  g2606
  (
    n2674,
    n2366,
    n2502,
    n2382,
    n2405
  );


  xnor
  g2607
  (
    n2666,
    n2389,
    n2402,
    n2073,
    n2273
  );


  xnor
  g2608
  (
    n2596,
    n2396,
    n2468,
    n2536,
    n2388
  );


  xor
  g2609
  (
    n2670,
    n2523,
    n2373,
    n2386,
    n2380
  );


  xor
  g2610
  (
    n2629,
    n2496,
    n2392,
    n2396,
    n2394
  );


  xnor
  g2611
  (
    n2634,
    n2531,
    n2461,
    n2387,
    n2403
  );


  nor
  g2612
  (
    n2618,
    n2516,
    n2404,
    n2394,
    n2275
  );


  and
  g2613
  (
    n2654,
    n2386,
    n2401,
    n2480,
    n2388
  );


  nor
  g2614
  (
    n2604,
    n2407,
    n2275,
    n2396,
    n2368
  );


  and
  g2615
  (
    n2630,
    n2368,
    n2386,
    n2369,
    n2514
  );


  nor
  g2616
  (
    n2646,
    n2380,
    n2375,
    n2476,
    n2511
  );


  nand
  g2617
  (
    n2599,
    n2371,
    n2392,
    n2543,
    n2400
  );


  xor
  g2618
  (
    n2632,
    n2529,
    n2521,
    n2397,
    n2466
  );


  and
  g2619
  (
    n2607,
    n2370,
    n2399,
    n2266,
    n2386
  );


  or
  g2620
  (
    n2621,
    n2495,
    n2522,
    n2372,
    n2537
  );


  xor
  g2621
  (
    n2605,
    n2270,
    n2504,
    n2392,
    n2082
  );


  nand
  g2622
  (
    n2649,
    n2285,
    n2398,
    n2486,
    n2397
  );


  and
  g2623
  (
    n2660,
    n2369,
    n2379,
    n2406,
    n2501
  );


  xor
  g2624
  (
    n2610,
    n2397,
    n503,
    n2375,
    n2373
  );


  nand
  g2625
  (
    n2633,
    n2267,
    n2388,
    n2402,
    n2403
  );


  nand
  g2626
  (
    n2678,
    n2520,
    n2407,
    n2075,
    n2513
  );


  or
  g2627
  (
    n2664,
    n2545,
    n2404,
    n2367,
    n2399
  );


  xor
  g2628
  (
    n2643,
    n2463,
    n2400,
    n2377,
    n2503
  );


  xor
  g2629
  (
    n2611,
    n2379,
    n2381,
    n2470,
    n2274
  );


  and
  g2630
  (
    n2612,
    n2372,
    n2376,
    n2544,
    n2079
  );


  xnor
  g2631
  (
    n2631,
    n2546,
    n2469,
    n2493,
    n2542
  );


  xnor
  g2632
  (
    n2601,
    n2402,
    n2382,
    n2274,
    n2460
  );


  nor
  g2633
  (
    n2627,
    n2376,
    n2458,
    n2406,
    n2396
  );


  xnor
  g2634
  (
    n2658,
    n2374,
    n2472,
    n2554,
    n2366
  );


  nand
  g2635
  (
    n2614,
    n2380,
    n2374,
    n504,
    n2500
  );


  or
  g2636
  (
    n2661,
    n2478,
    n2530,
    n2367,
    n2366
  );


  nor
  g2637
  (
    n2609,
    n2408,
    n2375,
    n2457,
    n2407
  );


  xor
  g2638
  (
    n2648,
    n2401,
    n2403,
    n2399,
    n2085
  );


  nand
  g2639
  (
    n2597,
    n2407,
    n2409,
    n2459,
    n2534
  );


  and
  g2640
  (
    n2668,
    n2284,
    n2540,
    n2074,
    n2515
  );


  nor
  g2641
  (
    n2600,
    n2210,
    n2401,
    n2379,
    n2489
  );


  xor
  g2642
  (
    n2647,
    n2535,
    n2370,
    n2406,
    n2390
  );


  xor
  g2643
  (
    n2657,
    n2506,
    n2393,
    n2508,
    n2517
  );


  and
  g2644
  (
    n2667,
    n2384,
    n2365,
    n2376,
    n2393
  );


  xor
  g2645
  (
    n2595,
    n2406,
    n2378,
    n2371,
    n2479
  );


  xnor
  g2646
  (
    n2641,
    n2372,
    n2392,
    n2381,
    n2498
  );


  or
  g2647
  (
    n2669,
    n1428,
    n2552,
    n2547,
    n2405
  );


  nand
  g2648
  (
    n2620,
    n2077,
    n2467,
    n2541,
    n2497
  );


  xnor
  g2649
  (
    n2676,
    n2399,
    n2548,
    n2084,
    n2378
  );


  xor
  g2650
  (
    n2623,
    n2387,
    n2395,
    n2487,
    n2385
  );


  xor
  g2651
  (
    n2637,
    n2382,
    n2539,
    n2488,
    n2555
  );


  or
  g2652
  (
    n2626,
    n2383,
    n2556,
    n2387,
    n2391
  );


  and
  g2653
  (
    n2615,
    n2408,
    n2490,
    n504,
    n2401
  );


  nor
  g2654
  (
    n2688,
    n2611,
    n2587,
    n2595,
    n2613
  );


  xnor
  g2655
  (
    n2684,
    n2619,
    n2615,
    n2594,
    n2564
  );


  xor
  g2656
  (
    n2679,
    n2589,
    n2599,
    n2577,
    n2605
  );


  nor
  g2657
  (
    n2687,
    n2576,
    n2588,
    n2583,
    n2612
  );


  or
  g2658
  (
    n2686,
    n2572,
    n2582,
    n2603,
    n2568
  );


  or
  g2659
  (
    n2693,
    n2575,
    n2563,
    n2578,
    n2601
  );


  nor
  g2660
  (
    n2689,
    n2597,
    n2621,
    n2608,
    n2567
  );


  xor
  g2661
  (
    n2691,
    n2562,
    n2584,
    n2581,
    n2609
  );


  and
  g2662
  (
    n2683,
    n2593,
    n2618,
    n2565,
    n2566
  );


  nand
  g2663
  (
    n2690,
    n2586,
    n2602,
    n2600,
    n2590
  );


  xor
  g2664
  (
    n2692,
    n2598,
    n2610,
    n2617,
    n2616
  );


  or
  g2665
  (
    n2685,
    n2620,
    n2579,
    n2607,
    n2580
  );


  nor
  g2666
  (
    n2680,
    n2585,
    n2614,
    n2596,
    n2592
  );


  xor
  g2667
  (
    n2682,
    n2606,
    n2569,
    n2574,
    n2570
  );


  or
  g2668
  (
    n2681,
    n2604,
    n2571,
    n2591,
    n2573
  );


  or
  g2669
  (
    n2698,
    n2623,
    n2644,
    n2629,
    n2654
  );


  nand
  g2670
  (
    n2694,
    n2649,
    n2645,
    n2636,
    n2643
  );


  nor
  g2671
  (
    n2702,
    n2630,
    n2641,
    n2691,
    n2642
  );


  nor
  g2672
  (
    n2696,
    n2683,
    n2686,
    n2682,
    n2632
  );


  xnor
  g2673
  (
    n2703,
    n2684,
    n2626,
    n2652,
    n2655
  );


  or
  g2674
  (
    n2705,
    n2693,
    n2648,
    n2631,
    n2633
  );


  nand
  g2675
  (
    n2697,
    n2086,
    n2689,
    n2692,
    n2634
  );


  or
  g2676
  (
    n2704,
    n2639,
    n2624,
    n2647,
    n2640
  );


  nor
  g2677
  (
    n2699,
    n2650,
    n2622,
    n2688,
    n2637
  );


  xnor
  g2678
  (
    n2695,
    n2625,
    n2635,
    n2638,
    n2685
  );


  xnor
  g2679
  (
    n2701,
    n2690,
    n2651,
    n2628,
    n2656
  );


  nand
  g2680
  (
    n2700,
    n2646,
    n2627,
    n2653,
    n2687
  );


  nor
  g2681
  (
    n2706,
    n1429,
    n2694
  );


  buf
  g2682
  (
    n2708,
    n2706
  );


  buf
  g2683
  (
    n2707,
    n2706
  );


  and
  g2684
  (
    n2715,
    n2663,
    n2659,
    n2673,
    n2658
  );


  nand
  g2685
  (
    n2709,
    n2670,
    n2707,
    n2662,
    n2674
  );


  xor
  g2686
  (
    n2716,
    n2677,
    n2708,
    n2664,
    n2669
  );


  xor
  g2687
  (
    n2711,
    n2668,
    n2672,
    n2708,
    n2088
  );


  xor
  g2688
  (
    n2714,
    n2676,
    n2708,
    n2657,
    n2707
  );


  xor
  g2689
  (
    n2710,
    n2087,
    n2707,
    n2665,
    n2666
  );


  and
  g2690
  (
    n2713,
    n2661,
    n2667,
    n2707,
    n2671
  );


  or
  g2691
  (
    n2712,
    n2675,
    n2678,
    n2660,
    n2708
  );


  and
  g2692
  (
    n2729,
    n1483,
    n2705,
    n1488,
    n2711
  );


  xnor
  g2693
  (
    n2735,
    n1467,
    n2704,
    n2714,
    n1462
  );


  and
  g2694
  (
    n2737,
    n1472,
    n1449,
    n2715,
    n1447
  );


  nand
  g2695
  (
    n2743,
    n1456,
    n2703,
    n1498,
    n1499
  );


  xnor
  g2696
  (
    n2724,
    n1476,
    n1508,
    n1439,
    n1474
  );


  nor
  g2697
  (
    n2745,
    n2713,
    n1459,
    n2711,
    n1481
  );


  or
  g2698
  (
    n2733,
    n1471,
    n1454,
    n1448,
    n1468
  );


  and
  g2699
  (
    n2738,
    n1431,
    n2699,
    n2702,
    n1446
  );


  or
  g2700
  (
    n2742,
    n2711,
    n1460,
    n1443,
    n2709
  );


  xnor
  g2701
  (
    n2727,
    n2715,
    n1441,
    n1485,
    n1502
  );


  nor
  g2702
  (
    n2722,
    n1469,
    n1496,
    n1444,
    n1432
  );


  xor
  g2703
  (
    n2725,
    n2710,
    n1477,
    n1466,
    n2709
  );


  or
  g2704
  (
    n2734,
    n1455,
    n2716,
    n2695
  );


  or
  g2705
  (
    n2741,
    n2712,
    n1504,
    n1509,
    n1507
  );


  nor
  g2706
  (
    n2740,
    n1436,
    n2716,
    n2229,
    n2701
  );


  nor
  g2707
  (
    n2747,
    n1464,
    n1486,
    n2698,
    n2715
  );


  or
  g2708
  (
    n2731,
    n2697,
    n1495,
    n2229,
    n1463
  );


  nand
  g2709
  (
    n2721,
    n2715,
    n1473,
    n1430,
    n1457
  );


  xor
  g2710
  (
    n2730,
    n1452,
    n1470,
    n2710,
    n2712
  );


  nor
  g2711
  (
    n2720,
    n1484,
    n2716,
    n1479,
    n2714
  );


  nand
  g2712
  (
    n2732,
    n2709,
    n1510,
    n1465,
    n1494
  );


  nor
  g2713
  (
    n2748,
    n1482,
    n1438,
    n1442,
    n1453
  );


  and
  g2714
  (
    n2717,
    n2710,
    n2713,
    n1503,
    n2712
  );


  or
  g2715
  (
    n2719,
    n1458,
    n1492,
    n1433,
    n2713
  );


  and
  g2716
  (
    n2746,
    n2710,
    n1480,
    n1461,
    n2711
  );


  and
  g2717
  (
    n2723,
    n1478,
    n1491,
    n2714,
    n1500
  );


  nor
  g2718
  (
    n2736,
    n1487,
    n1437,
    n1435,
    n1434
  );


  xnor
  g2719
  (
    n2744,
    n1501,
    n2714,
    n1489,
    n1440
  );


  xor
  g2720
  (
    n2728,
    n1493,
    n1450,
    n1445,
    n1451
  );


  or
  g2721
  (
    n2726,
    n1490,
    n2712,
    n1475,
    n2700
  );


  and
  g2722
  (
    n2718,
    n1497,
    n2229,
    n2709,
    n1506
  );


  xor
  g2723
  (
    n2739,
    n2713,
    n2229,
    n2696,
    n1505
  );


  and
  g2724
  (
    n2772,
    n2180,
    n2165,
    n2119,
    n2184
  );


  nand
  g2725
  (
    n2752,
    n2743,
    n2144,
    n2186,
    n2738
  );


  xor
  g2726
  (
    n2770,
    n2102,
    n2176,
    n2117,
    n2161
  );


  xor
  g2727
  (
    n2765,
    n2089,
    n2133,
    n2100,
    n2147
  );


  xor
  g2728
  (
    n2767,
    n2171,
    n2143,
    n2128,
    n2155
  );


  nand
  g2729
  (
    n2750,
    n2718,
    n2735,
    n2725,
    n2748
  );


  and
  g2730
  (
    n2757,
    n2135,
    n2098,
    n2152,
    n2094
  );


  xnor
  g2731
  (
    n2777,
    n2104,
    n2134,
    n2173,
    n2131
  );


  xor
  g2732
  (
    n2759,
    n2717,
    n2737,
    n2163,
    n2121
  );


  xnor
  g2733
  (
    n2776,
    n2136,
    n2187,
    n2744,
    n2113
  );


  xor
  g2734
  (
    n2773,
    n2174,
    n2733,
    n2154,
    n2742
  );


  nor
  g2735
  (
    n2769,
    n2092,
    n2731,
    n2123,
    n2170
  );


  xnor
  g2736
  (
    n2768,
    n2149,
    n2146,
    n2167,
    n2746
  );


  xor
  g2737
  (
    n2755,
    n2109,
    n2101,
    n2721,
    n2115
  );


  nor
  g2738
  (
    n2763,
    n2748,
    n2175,
    n2126,
    n2090
  );


  nand
  g2739
  (
    n2758,
    n2734,
    n2726,
    n2720,
    n2157
  );


  nand
  g2740
  (
    n2778,
    n2732,
    n2747,
    n2160,
    n2145
  );


  and
  g2741
  (
    n2753,
    n2096,
    n2169,
    n2105,
    n2730
  );


  and
  g2742
  (
    n2761,
    n2741,
    n2166,
    n2736,
    n2097
  );


  or
  g2743
  (
    n2779,
    n2138,
    n2150,
    n2132,
    n2185
  );


  and
  g2744
  (
    n2762,
    n2116,
    n2183,
    n2172,
    n2122
  );


  xnor
  g2745
  (
    n2766,
    n2107,
    n2148,
    n2719,
    n2093
  );


  and
  g2746
  (
    n2780,
    n2178,
    n2179,
    n2103,
    n2153
  );


  nand
  g2747
  (
    n2760,
    n2162,
    n2111,
    n2164,
    n2095
  );


  xnor
  g2748
  (
    n2781,
    n2141,
    n2118,
    n2112,
    n2740
  );


  or
  g2749
  (
    n2764,
    n2108,
    n2177,
    n2156,
    n2114
  );


  and
  g2750
  (
    n2774,
    n2729,
    n2139,
    n2127,
    n2106
  );


  xnor
  g2751
  (
    n2754,
    n2140,
    n2129,
    n2739,
    n2110
  );


  xnor
  g2752
  (
    n2749,
    n2137,
    n2723,
    n2125,
    n2728
  );


  xnor
  g2753
  (
    n2756,
    n2091,
    n2158,
    n2182,
    n2724
  );


  nand
  g2754
  (
    n2771,
    n2151,
    n2727,
    n2181,
    n2745
  );


  xnor
  g2755
  (
    n2751,
    n2159,
    n2120,
    n2130,
    n2142
  );


  nand
  g2756
  (
    n2775,
    n2168,
    n2124,
    n2722,
    n2099
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1552,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n2261,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n2329,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n2459,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1153,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n753,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n710,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n2034,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n240,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n2326,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n943,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n544,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n469,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n2635,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n905,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n447,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


