

module Stat_100_48
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n125,
  n122,
  n115,
  n131,
  n116,
  n111,
  n106,
  n130,
  n105,
  n119,
  n128,
  n102,
  n123,
  n120,
  n129,
  n107,
  n124,
  n127,
  n117,
  n104,
  n114,
  n101,
  n113,
  n110,
  n112,
  n103,
  n121,
  n132,
  n109,
  n126,
  n108,
  n118
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n125;output n122;output n115;output n131;output n116;output n111;output n106;output n130;output n105;output n119;output n128;output n102;output n123;output n120;output n129;output n107;output n124;output n127;output n117;output n104;output n114;output n101;output n113;output n110;output n112;output n103;output n121;output n132;output n109;output n126;output n108;output n118;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    KeyWire_0_18,
    n4
  );


  buf
  g1
  (
    KeyWire_0_26,
    n2
  );


  not
  g2
  (
    KeyWire_0_5,
    n4
  );


  not
  g3
  (
    n39,
    n3
  );


  not
  g4
  (
    n33,
    n1
  );


  not
  g5
  (
    KeyWire_0_58,
    n3
  );


  not
  g6
  (
    n37,
    n1
  );


  not
  g7
  (
    KeyWire_0_38,
    n2
  );


  buf
  g8
  (
    KeyWire_0_12,
    n1
  );


  xnor
  g9
  (
    KeyWire_0_16,
    n2,
    n3
  );


  buf
  g10
  (
    KeyWire_0_15,
    n37
  );


  buf
  g11
  (
    KeyWire_0_63,
    n40
  );


  buf
  g12
  (
    KeyWire_0_28,
    n34
  );


  buf
  g13
  (
    n45,
    n37
  );


  buf
  g14
  (
    KeyWire_0_21,
    n34
  );


  not
  g15
  (
    n55,
    n40
  );


  not
  g16
  (
    KeyWire_0_54,
    n37
  );


  buf
  g17
  (
    KeyWire_0_6,
    n36
  );


  not
  g18
  (
    n58,
    n38
  );


  or
  g19
  (
    KeyWire_0_57,
    n40,
    n42,
    n36,
    n33
  );


  xor
  g20
  (
    n44,
    n38,
    n38,
    n33,
    n42
  );


  nand
  g21
  (
    KeyWire_0_11,
    n36,
    n39,
    n35
  );


  nand
  g22
  (
    n52,
    n40,
    n39,
    n37,
    n38
  );


  and
  g23
  (
    n49,
    n34,
    n42,
    n36,
    n41
  );


  or
  g24
  (
    KeyWire_0_10,
    n41,
    n33,
    n35,
    n39
  );


  nand
  g25
  (
    KeyWire_0_45,
    n39,
    n42,
    n41
  );


  nor
  g26
  (
    n62,
    n15,
    n13,
    n45
  );


  nor
  g27
  (
    KeyWire_0_13,
    n10,
    n49,
    n7
  );


  or
  g28
  (
    KeyWire_0_27,
    n5,
    n24,
    n22
  );


  xor
  g29
  (
    KeyWire_0_40,
    n53,
    n49,
    n28
  );


  xnor
  g30
  (
    KeyWire_0_4,
    n12,
    n45,
    n10
  );


  or
  g31
  (
    n60,
    n54,
    n25,
    n45
  );


  and
  g32
  (
    n73,
    n30,
    n21,
    n12
  );


  xnor
  g33
  (
    KeyWire_0_46,
    n14,
    n58,
    n26
  );


  nor
  g34
  (
    KeyWire_0_34,
    n31,
    n22,
    n13
  );


  nand
  g35
  (
    KeyWire_0_61,
    n26,
    n47
  );


  and
  g36
  (
    n67,
    n15,
    n43,
    n46
  );


  and
  g37
  (
    KeyWire_0_47,
    n21,
    n9,
    n48
  );


  or
  g38
  (
    n84,
    n58,
    n28,
    n43
  );


  xnor
  g39
  (
    KeyWire_0_44,
    n23,
    n19,
    n57
  );


  or
  g40
  (
    KeyWire_0_30,
    n8,
    n27,
    n9
  );


  nand
  g41
  (
    n61,
    n52,
    n17,
    n53
  );


  and
  g42
  (
    KeyWire_0_56,
    n11,
    n16
  );


  nand
  g43
  (
    n66,
    n48,
    n18,
    n51
  );


  xnor
  g44
  (
    KeyWire_0_2,
    n26,
    n31,
    n22
  );


  nor
  g45
  (
    n81,
    n31,
    n27,
    n44
  );


  or
  g46
  (
    n63,
    n46,
    n25,
    n7
  );


  or
  g47
  (
    KeyWire_0_53,
    n30,
    n25,
    n58
  );


  xnor
  g48
  (
    n87,
    n52,
    n6,
    n55
  );


  or
  g49
  (
    KeyWire_0_20,
    n29,
    n23,
    n20,
    n56
  );


  and
  g50
  (
    KeyWire_0_39,
    n11,
    n56,
    n57,
    n23
  );


  or
  g51
  (
    KeyWire_0_37,
    n18,
    n56,
    n11,
    n16
  );


  xnor
  g52
  (
    KeyWire_0_31,
    n20,
    n27,
    n14,
    n22
  );


  nand
  g53
  (
    KeyWire_0_41,
    n50,
    n14,
    n6,
    n52
  );


  nand
  g54
  (
    KeyWire_0_32,
    n23,
    n58,
    n18,
    n43
  );


  nand
  g55
  (
    n99,
    n26,
    n47,
    n20,
    n51
  );


  xor
  g56
  (
    n64,
    n8,
    n21,
    n5,
    n55
  );


  xor
  g57
  (
    n100,
    n17,
    n30,
    n13,
    n25
  );


  and
  g58
  (
    KeyWire_0_49,
    n15,
    n44,
    n32,
    n50
  );


  xnor
  g59
  (
    n72,
    n28,
    n32,
    n10,
    n50
  );


  xnor
  g60
  (
    KeyWire_0_29,
    n29,
    n17,
    n57,
    n30
  );


  nor
  g61
  (
    KeyWire_0_48,
    n31,
    n55,
    n46,
    n6
  );


  or
  g62
  (
    n75,
    n24,
    n48,
    n7,
    n8
  );


  nor
  g63
  (
    n91,
    n49,
    n19,
    n54,
    n9
  );


  nor
  g64
  (
    n90,
    n29,
    n4,
    n20,
    n24
  );


  xnor
  g65
  (
    n76,
    n51,
    n44,
    n12,
    n54
  );


  or
  g66
  (
    KeyWire_0_25,
    n24,
    n27,
    n19,
    n29
  );


  xnor
  g67
  (
    n86,
    n28,
    n21,
    n53,
    n5
  );


  nor
  g68
  (
    KeyWire_0_8,
    n81,
    n69,
    n91
  );


  xnor
  g69
  (
    KeyWire_0_52,
    n88,
    n66,
    n67,
    n71
  );


  nor
  g70
  (
    KeyWire_0_50,
    n62,
    n84,
    n86,
    n74
  );


  xor
  g71
  (
    n126,
    n100,
    n93,
    n83,
    n97
  );


  xnor
  g72
  (
    KeyWire_0_36,
    n70,
    n70,
    n90,
    n92
  );


  or
  g73
  (
    KeyWire_0_1,
    n92,
    n97,
    n59,
    n77
  );


  xnor
  g74
  (
    KeyWire_0_7,
    n73,
    n81,
    n68,
    n79
  );


  or
  g75
  (
    KeyWire_0_43,
    n98,
    n65,
    n76,
    n80
  );


  nor
  g76
  (
    KeyWire_0_9,
    n72,
    n85,
    n64,
    n95
  );


  xnor
  g77
  (
    KeyWire_0_14,
    n91,
    n82,
    n90,
    n61
  );


  nor
  g78
  (
    KeyWire_0_19,
    n62,
    n94,
    n86,
    n71
  );


  or
  g79
  (
    KeyWire_0_0,
    n84,
    n99,
    n94,
    n63
  );


  nor
  g80
  (
    KeyWire_0_17,
    n79,
    n74,
    n75,
    n78
  );


  xor
  g81
  (
    KeyWire_0_24,
    n85,
    n93,
    n78,
    n61
  );


  nor
  g82
  (
    n106,
    n69,
    n82,
    n70,
    n65
  );


  nand
  g83
  (
    KeyWire_0_59,
    n60,
    n83,
    n32,
    n87
  );


  xor
  g84
  (
    n130,
    n67,
    n81,
    n99,
    n89
  );


  nor
  g85
  (
    n123,
    n95,
    n92,
    n88,
    n100
  );


  xnor
  g86
  (
    KeyWire_0_33,
    n96,
    n94,
    n60,
    n83
  );


  xnor
  g87
  (
    KeyWire_0_35,
    n68,
    n80,
    n64
  );


  xor
  g88
  (
    n128,
    n93,
    n66,
    n61,
    n100
  );


  nor
  g89
  (
    n129,
    n99,
    n63,
    n59
  );


  xnor
  g90
  (
    KeyWire_0_3,
    n84,
    n90,
    n62,
    n69
  );


  xor
  g91
  (
    KeyWire_0_55,
    n77,
    n75,
    n73,
    n96
  );


  xnor
  g92
  (
    KeyWire_0_62,
    n98,
    n71,
    n87,
    n64
  );


  xnor
  g93
  (
    KeyWire_0_22,
    n87,
    n72,
    n78,
    n75
  );


  xnor
  g94
  (
    KeyWire_0_60,
    n85,
    n74,
    n76,
    n79
  );


  nor
  g95
  (
    KeyWire_0_23,
    n68,
    n96,
    n76,
    n97
  );


  xor
  g96
  (
    n120,
    n66,
    n88,
    n89,
    n65
  );


  nand
  g97
  (
    KeyWire_0_51,
    n60,
    n73,
    n86,
    n98
  );


  or
  g98
  (
    KeyWire_0_42,
    n32,
    n72,
    n67,
    n89
  );


  and
  g99
  (
    n127,
    n59,
    n77,
    n82,
    n95
  );


  xor
  KeyGate_0_0
  (
    n125,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n118,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n77,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n114,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n79,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n41,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n51,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n119,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n109,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n101,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n57,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n43,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n35,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n89,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n122,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n50,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n38,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n102,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n34,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n111,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n59,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n47,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n108,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n116,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n107,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n65,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n40,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n85,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n46,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n68,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n80,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n97,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n98,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n105,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n88,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n104,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n112,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n74,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n42,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n96,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n94,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n78,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n110,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n113,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n69,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n54,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n71,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n70,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n92,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n95,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n131,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n103,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n115,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n82,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n48,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n121,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n83,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n56,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n36,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n132,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n117,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n93,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n124,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n53,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


