

module Stat_2149_33_13
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n2004,
  n2003,
  n2011,
  n2015,
  n2013,
  n2014,
  n2012,
  n2010,
  n2009,
  n2001,
  n2002,
  n2008,
  n2005,
  n2007,
  n2027,
  n2176,
  n2177,
  n2175,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n2004;
  output n2003;
  output n2011;
  output n2015;
  output n2013;
  output n2014;
  output n2012;
  output n2010;
  output n2009;
  output n2001;
  output n2002;
  output n2008;
  output n2005;
  output n2007;
  output n2027;
  output n2176;
  output n2177;
  output n2175;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2006;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n80,
    n2
  );


  buf
  g1
  (
    n131,
    n11
  );


  not
  g2
  (
    n110,
    n13
  );


  buf
  g3
  (
    n38,
    n26
  );


  buf
  g4
  (
    n30,
    n3
  );


  not
  g5
  (
    n106,
    n15
  );


  not
  g6
  (
    n57,
    n20
  );


  not
  g7
  (
    n52,
    n8
  );


  buf
  g8
  (
    n112,
    n7
  );


  buf
  g9
  (
    n60,
    n10
  );


  not
  g10
  (
    n70,
    n16
  );


  buf
  g11
  (
    n41,
    n27
  );


  buf
  g12
  (
    n39,
    n6
  );


  not
  g13
  (
    n76,
    n18
  );


  buf
  g14
  (
    n75,
    n21
  );


  buf
  g15
  (
    n91,
    n7
  );


  buf
  g16
  (
    n93,
    n19
  );


  buf
  g17
  (
    n111,
    n9
  );


  buf
  g18
  (
    n94,
    n27
  );


  not
  g19
  (
    n95,
    n19
  );


  buf
  g20
  (
    n56,
    n3
  );


  not
  g21
  (
    n130,
    n1
  );


  not
  g22
  (
    n31,
    n17
  );


  buf
  g23
  (
    n44,
    n17
  );


  not
  g24
  (
    n107,
    n17
  );


  not
  g25
  (
    n115,
    n15
  );


  buf
  g26
  (
    n33,
    n26
  );


  not
  g27
  (
    n46,
    n20
  );


  buf
  g28
  (
    n68,
    n20
  );


  not
  g29
  (
    n87,
    n11
  );


  not
  g30
  (
    n118,
    n24
  );


  not
  g31
  (
    n71,
    n1
  );


  buf
  g32
  (
    n133,
    n21
  );


  buf
  g33
  (
    n138,
    n15
  );


  not
  g34
  (
    n73,
    n7
  );


  not
  g35
  (
    n102,
    n9
  );


  buf
  g36
  (
    n126,
    n9
  );


  not
  g37
  (
    n127,
    n8
  );


  buf
  g38
  (
    n96,
    n2
  );


  not
  g39
  (
    n48,
    n7
  );


  buf
  g40
  (
    n47,
    n5
  );


  buf
  g41
  (
    n104,
    n17
  );


  buf
  g42
  (
    n40,
    n1
  );


  buf
  g43
  (
    n114,
    n22
  );


  not
  g44
  (
    n51,
    n5
  );


  not
  g45
  (
    n43,
    n13
  );


  not
  g46
  (
    n83,
    n1
  );


  buf
  g47
  (
    n66,
    n13
  );


  buf
  g48
  (
    n113,
    n24
  );


  not
  g49
  (
    n45,
    n4
  );


  not
  g50
  (
    n64,
    n25
  );


  not
  g51
  (
    n109,
    n24
  );


  buf
  g52
  (
    n122,
    n24
  );


  not
  g53
  (
    n54,
    n3
  );


  buf
  g54
  (
    n129,
    n6
  );


  not
  g55
  (
    n136,
    n18
  );


  buf
  g56
  (
    n32,
    n23
  );


  not
  g57
  (
    n61,
    n10
  );


  not
  g58
  (
    n77,
    n14
  );


  not
  g59
  (
    n90,
    n8
  );


  not
  g60
  (
    n42,
    n18
  );


  not
  g61
  (
    n74,
    n22
  );


  not
  g62
  (
    KeyWire_0_6,
    n28
  );


  not
  g63
  (
    n117,
    n12
  );


  buf
  g64
  (
    n81,
    n16
  );


  not
  g65
  (
    n86,
    n10
  );


  not
  g66
  (
    n78,
    n19
  );


  not
  g67
  (
    n55,
    n5
  );


  not
  g68
  (
    n50,
    n23
  );


  not
  g69
  (
    n36,
    n23
  );


  not
  g70
  (
    n89,
    n4
  );


  not
  g71
  (
    n34,
    n4
  );


  buf
  g72
  (
    n72,
    n26
  );


  buf
  g73
  (
    n53,
    n10
  );


  buf
  g74
  (
    n105,
    n6
  );


  buf
  g75
  (
    n65,
    n5
  );


  not
  g76
  (
    n35,
    n21
  );


  buf
  g77
  (
    n69,
    n25
  );


  buf
  g78
  (
    n123,
    n12
  );


  not
  g79
  (
    n88,
    n13
  );


  not
  g80
  (
    n124,
    n12
  );


  not
  g81
  (
    n82,
    n18
  );


  not
  g82
  (
    n137,
    n26
  );


  buf
  g83
  (
    n92,
    n6
  );


  not
  g84
  (
    n101,
    n21
  );


  buf
  g85
  (
    n100,
    n23
  );


  buf
  g86
  (
    n67,
    n15
  );


  not
  g87
  (
    n49,
    n27
  );


  not
  g88
  (
    n128,
    n22
  );


  buf
  g89
  (
    n99,
    n8
  );


  buf
  g90
  (
    n37,
    n27
  );


  buf
  g91
  (
    n132,
    n14
  );


  buf
  g92
  (
    n134,
    n2
  );


  buf
  g93
  (
    n58,
    n12
  );


  not
  g94
  (
    n59,
    n9
  );


  not
  g95
  (
    n63,
    n11
  );


  buf
  g96
  (
    n108,
    n25
  );


  not
  g97
  (
    n97,
    n14
  );


  buf
  g98
  (
    n29,
    n14
  );


  buf
  g99
  (
    n116,
    n4
  );


  not
  g100
  (
    n62,
    n28
  );


  buf
  g101
  (
    n98,
    n2
  );


  not
  g102
  (
    n121,
    n3
  );


  not
  g103
  (
    KeyWire_0_4,
    n16
  );


  not
  g104
  (
    n119,
    n20
  );


  buf
  g105
  (
    n85,
    n16
  );


  not
  g106
  (
    n84,
    n22
  );


  buf
  g107
  (
    n103,
    n25
  );


  not
  g108
  (
    n125,
    n11
  );


  buf
  g109
  (
    n135,
    n19
  );


  not
  g110
  (
    KeyWire_0_22,
    n55
  );


  not
  g111
  (
    n571,
    n120
  );


  buf
  g112
  (
    n325,
    n63
  );


  buf
  g113
  (
    n361,
    n59
  );


  not
  g114
  (
    n332,
    n56
  );


  buf
  g115
  (
    KeyWire_0_7,
    n115
  );


  not
  g116
  (
    n484,
    n129
  );


  buf
  g117
  (
    n462,
    n75
  );


  not
  g118
  (
    n167,
    n102
  );


  not
  g119
  (
    n384,
    n29
  );


  buf
  g120
  (
    n330,
    n32
  );


  buf
  g121
  (
    n492,
    n76
  );


  buf
  g122
  (
    n510,
    n107
  );


  not
  g123
  (
    n188,
    n60
  );


  buf
  g124
  (
    n248,
    n60
  );


  buf
  g125
  (
    n441,
    n46
  );


  not
  g126
  (
    n172,
    n99
  );


  buf
  g127
  (
    n414,
    n83
  );


  not
  g128
  (
    n430,
    n45
  );


  not
  g129
  (
    n435,
    n114
  );


  buf
  g130
  (
    n190,
    n119
  );


  not
  g131
  (
    n569,
    n39
  );


  buf
  g132
  (
    n146,
    n137
  );


  buf
  g133
  (
    n181,
    n109
  );


  buf
  g134
  (
    n380,
    n70
  );


  not
  g135
  (
    n401,
    n130
  );


  not
  g136
  (
    n357,
    n81
  );


  buf
  g137
  (
    n388,
    n120
  );


  not
  g138
  (
    n195,
    n112
  );


  not
  g139
  (
    n452,
    n49
  );


  not
  g140
  (
    n300,
    n102
  );


  not
  g141
  (
    n262,
    n133
  );


  not
  g142
  (
    n561,
    n82
  );


  buf
  g143
  (
    n198,
    n136
  );


  not
  g144
  (
    n545,
    n122
  );


  buf
  g145
  (
    n511,
    n51
  );


  not
  g146
  (
    n533,
    n58
  );


  not
  g147
  (
    n392,
    n44
  );


  buf
  g148
  (
    n540,
    n94
  );


  buf
  g149
  (
    n327,
    n134
  );


  not
  g150
  (
    n417,
    n88
  );


  not
  g151
  (
    n199,
    n136
  );


  not
  g152
  (
    n428,
    n137
  );


  buf
  g153
  (
    n372,
    n116
  );


  buf
  g154
  (
    n398,
    n103
  );


  not
  g155
  (
    n301,
    n103
  );


  buf
  g156
  (
    n211,
    n118
  );


  not
  g157
  (
    n311,
    n93
  );


  not
  g158
  (
    n310,
    n44
  );


  buf
  g159
  (
    n535,
    n113
  );


  not
  g160
  (
    n293,
    n77
  );


  not
  g161
  (
    n425,
    n123
  );


  buf
  g162
  (
    n315,
    n124
  );


  not
  g163
  (
    n214,
    n47
  );


  buf
  g164
  (
    n189,
    n90
  );


  buf
  g165
  (
    n180,
    n118
  );


  not
  g166
  (
    n221,
    n53
  );


  buf
  g167
  (
    n256,
    n123
  );


  not
  g168
  (
    n220,
    n88
  );


  buf
  g169
  (
    n234,
    n70
  );


  not
  g170
  (
    n449,
    n47
  );


  buf
  g171
  (
    n192,
    n59
  );


  not
  g172
  (
    n455,
    n36
  );


  buf
  g173
  (
    n153,
    n111
  );


  not
  g174
  (
    n481,
    n51
  );


  buf
  g175
  (
    n404,
    n78
  );


  buf
  g176
  (
    n314,
    n48
  );


  buf
  g177
  (
    n150,
    n122
  );


  buf
  g178
  (
    n247,
    n126
  );


  buf
  g179
  (
    n562,
    n29
  );


  buf
  g180
  (
    n513,
    n34
  );


  not
  g181
  (
    n451,
    n68
  );


  buf
  g182
  (
    n148,
    n119
  );


  buf
  g183
  (
    n419,
    n80
  );


  buf
  g184
  (
    n526,
    n76
  );


  buf
  g185
  (
    n208,
    n39
  );


  not
  g186
  (
    n304,
    n57
  );


  buf
  g187
  (
    n573,
    n51
  );


  buf
  g188
  (
    n166,
    n69
  );


  buf
  g189
  (
    n207,
    n66
  );


  not
  g190
  (
    n478,
    n42
  );


  not
  g191
  (
    n399,
    n134
  );


  buf
  g192
  (
    n469,
    n114
  );


  buf
  g193
  (
    n439,
    n35
  );


  buf
  g194
  (
    n556,
    n65
  );


  not
  g195
  (
    n555,
    n73
  );


  buf
  g196
  (
    n296,
    n107
  );


  not
  g197
  (
    n292,
    n116
  );


  not
  g198
  (
    n193,
    n123
  );


  not
  g199
  (
    n215,
    n104
  );


  not
  g200
  (
    n285,
    n109
  );


  buf
  g201
  (
    n164,
    n112
  );


  buf
  g202
  (
    n197,
    n89
  );


  buf
  g203
  (
    n313,
    n92
  );


  not
  g204
  (
    n253,
    n95
  );


  not
  g205
  (
    n260,
    n87
  );


  buf
  g206
  (
    n483,
    n30
  );


  buf
  g207
  (
    n173,
    n105
  );


  buf
  g208
  (
    n159,
    n64
  );


  buf
  g209
  (
    n379,
    n118
  );


  not
  g210
  (
    n223,
    n79
  );


  not
  g211
  (
    n385,
    n63
  );


  buf
  g212
  (
    n218,
    n69
  );


  buf
  g213
  (
    n222,
    n100
  );


  buf
  g214
  (
    n567,
    n110
  );


  not
  g215
  (
    n203,
    n87
  );


  not
  g216
  (
    n386,
    n98
  );


  not
  g217
  (
    n496,
    n73
  );


  not
  g218
  (
    n261,
    n54
  );


  not
  g219
  (
    n502,
    n33
  );


  not
  g220
  (
    n495,
    n88
  );


  not
  g221
  (
    n468,
    n82
  );


  not
  g222
  (
    n318,
    n70
  );


  buf
  g223
  (
    n394,
    n48
  );


  not
  g224
  (
    n324,
    n97
  );


  not
  g225
  (
    n499,
    n47
  );


  not
  g226
  (
    n497,
    n35
  );


  not
  g227
  (
    n171,
    n72
  );


  not
  g228
  (
    n346,
    n46
  );


  buf
  g229
  (
    n420,
    n51
  );


  not
  g230
  (
    n354,
    n111
  );


  not
  g231
  (
    n219,
    n98
  );


  not
  g232
  (
    n368,
    n47
  );


  buf
  g233
  (
    n393,
    n76
  );


  not
  g234
  (
    n160,
    n77
  );


  not
  g235
  (
    KeyWire_0_14,
    n115
  );


  not
  g236
  (
    n305,
    n65
  );


  not
  g237
  (
    n551,
    n125
  );


  not
  g238
  (
    n338,
    n106
  );


  not
  g239
  (
    n470,
    n78
  );


  buf
  g240
  (
    n429,
    n137
  );


  buf
  g241
  (
    n212,
    n43
  );


  buf
  g242
  (
    n410,
    n38
  );


  buf
  g243
  (
    KeyWire_0_2,
    n93
  );


  not
  g244
  (
    n174,
    n44
  );


  buf
  g245
  (
    n453,
    n116
  );


  buf
  g246
  (
    n515,
    n71
  );


  not
  g247
  (
    n466,
    n52
  );


  buf
  g248
  (
    n523,
    n66
  );


  not
  g249
  (
    n202,
    n68
  );


  not
  g250
  (
    n213,
    n55
  );


  buf
  g251
  (
    KeyWire_0_30,
    n80
  );


  buf
  g252
  (
    n447,
    n99
  );


  buf
  g253
  (
    n572,
    n131
  );


  not
  g254
  (
    n443,
    n38
  );


  not
  g255
  (
    n426,
    n61
  );


  buf
  g256
  (
    n438,
    n114
  );


  buf
  g257
  (
    n383,
    n45
  );


  buf
  g258
  (
    n520,
    n128
  );


  not
  g259
  (
    n151,
    n89
  );


  not
  g260
  (
    n161,
    n82
  );


  buf
  g261
  (
    n149,
    n56
  );


  buf
  g262
  (
    n272,
    n136
  );


  not
  g263
  (
    n390,
    n52
  );


  not
  g264
  (
    n140,
    n59
  );


  buf
  g265
  (
    n507,
    n130
  );


  not
  g266
  (
    n459,
    n33
  );


  not
  g267
  (
    n415,
    n37
  );


  buf
  g268
  (
    n235,
    n117
  );


  buf
  g269
  (
    n446,
    n118
  );


  not
  g270
  (
    n498,
    n106
  );


  not
  g271
  (
    n352,
    n85
  );


  buf
  g272
  (
    n351,
    n125
  );


  not
  g273
  (
    n370,
    n91
  );


  not
  g274
  (
    n475,
    n91
  );


  not
  g275
  (
    n157,
    n34
  );


  not
  g276
  (
    n431,
    n49
  );


  not
  g277
  (
    n505,
    n122
  );


  buf
  g278
  (
    n243,
    n89
  );


  buf
  g279
  (
    n490,
    n101
  );


  not
  g280
  (
    n387,
    n84
  );


  buf
  g281
  (
    n432,
    n74
  );


  not
  g282
  (
    n152,
    n58
  );


  not
  g283
  (
    n139,
    n67
  );


  not
  g284
  (
    n504,
    n128
  );


  not
  g285
  (
    n263,
    n61
  );


  not
  g286
  (
    n266,
    n48
  );


  buf
  g287
  (
    n440,
    n63
  );


  buf
  g288
  (
    n344,
    n108
  );


  buf
  g289
  (
    n559,
    n111
  );


  buf
  g290
  (
    n395,
    n104
  );


  not
  g291
  (
    n491,
    n85
  );


  buf
  g292
  (
    n308,
    n67
  );


  buf
  g293
  (
    n550,
    n126
  );


  not
  g294
  (
    n391,
    n106
  );


  buf
  g295
  (
    n282,
    n50
  );


  not
  g296
  (
    n375,
    n29
  );


  buf
  g297
  (
    n227,
    n129
  );


  not
  g298
  (
    n382,
    n107
  );


  buf
  g299
  (
    n554,
    n95
  );


  not
  g300
  (
    n489,
    n95
  );


  buf
  g301
  (
    n237,
    n75
  );


  buf
  g302
  (
    n542,
    n108
  );


  not
  g303
  (
    n158,
    n105
  );


  not
  g304
  (
    n179,
    n40
  );


  not
  g305
  (
    n348,
    n78
  );


  buf
  g306
  (
    n480,
    n135
  );


  not
  g307
  (
    n450,
    n29
  );


  buf
  g308
  (
    n230,
    n43
  );


  buf
  g309
  (
    n184,
    n34
  );


  buf
  g310
  (
    n465,
    n86
  );


  buf
  g311
  (
    n170,
    n96
  );


  not
  g312
  (
    KeyWire_0_12,
    n83
  );


  not
  g313
  (
    n290,
    n90
  );


  not
  g314
  (
    n275,
    n65
  );


  buf
  g315
  (
    n331,
    n117
  );


  buf
  g316
  (
    n416,
    n135
  );


  not
  g317
  (
    n412,
    n46
  );


  not
  g318
  (
    n279,
    n69
  );


  not
  g319
  (
    n362,
    n133
  );


  buf
  g320
  (
    n177,
    n117
  );


  buf
  g321
  (
    n365,
    n37
  );


  not
  g322
  (
    KeyWire_0_29,
    n81
  );


  not
  g323
  (
    n397,
    n131
  );


  buf
  g324
  (
    n283,
    n113
  );


  buf
  g325
  (
    n303,
    n60
  );


  buf
  g326
  (
    n200,
    n93
  );


  not
  g327
  (
    n503,
    n48
  );


  buf
  g328
  (
    n321,
    n53
  );


  buf
  g329
  (
    n236,
    n104
  );


  not
  g330
  (
    n270,
    n84
  );


  not
  g331
  (
    n512,
    n135
  );


  buf
  g332
  (
    n360,
    n86
  );


  buf
  g333
  (
    n413,
    n107
  );


  buf
  g334
  (
    n216,
    n82
  );


  buf
  g335
  (
    n196,
    n36
  );


  not
  g336
  (
    n474,
    n101
  );


  not
  g337
  (
    n349,
    n96
  );


  not
  g338
  (
    n543,
    n113
  );


  not
  g339
  (
    n210,
    n106
  );


  buf
  g340
  (
    n165,
    n69
  );


  not
  g341
  (
    n359,
    n58
  );


  buf
  g342
  (
    n527,
    n60
  );


  buf
  g343
  (
    n224,
    n112
  );


  not
  g344
  (
    n232,
    n73
  );


  buf
  g345
  (
    n464,
    n88
  );


  buf
  g346
  (
    n405,
    n79
  );


  buf
  g347
  (
    n467,
    n32
  );


  not
  g348
  (
    n544,
    n71
  );


  buf
  g349
  (
    n422,
    n95
  );


  buf
  g350
  (
    n541,
    n37
  );


  not
  g351
  (
    n553,
    n44
  );


  not
  g352
  (
    n141,
    n132
  );


  not
  g353
  (
    n145,
    n94
  );


  not
  g354
  (
    n493,
    n108
  );


  buf
  g355
  (
    n355,
    n31
  );


  not
  g356
  (
    n205,
    n120
  );


  buf
  g357
  (
    n326,
    n138
  );


  buf
  g358
  (
    n546,
    n94
  );


  buf
  g359
  (
    n244,
    n56
  );


  buf
  g360
  (
    n538,
    n105
  );


  buf
  g361
  (
    n280,
    n66
  );


  not
  g362
  (
    n336,
    n122
  );


  not
  g363
  (
    n231,
    n49
  );


  not
  g364
  (
    n154,
    n103
  );


  buf
  g365
  (
    n487,
    n119
  );


  buf
  g366
  (
    n233,
    n61
  );


  not
  g367
  (
    n460,
    n100
  );


  not
  g368
  (
    n565,
    n126
  );


  not
  g369
  (
    n284,
    n30
  );


  buf
  g370
  (
    n444,
    n49
  );


  not
  g371
  (
    n517,
    n102
  );


  not
  g372
  (
    n518,
    n45
  );


  buf
  g373
  (
    n350,
    n124
  );


  buf
  g374
  (
    n353,
    n41
  );


  not
  g375
  (
    n521,
    n99
  );


  buf
  g376
  (
    n183,
    n84
  );


  not
  g377
  (
    n306,
    n132
  );


  not
  g378
  (
    n374,
    n127
  );


  buf
  g379
  (
    n276,
    n30
  );


  not
  g380
  (
    n536,
    n109
  );


  not
  g381
  (
    n500,
    n98
  );


  not
  g382
  (
    n519,
    n133
  );


  not
  g383
  (
    n277,
    n124
  );


  not
  g384
  (
    n400,
    n113
  );


  buf
  g385
  (
    n516,
    n110
  );


  buf
  g386
  (
    n156,
    n73
  );


  buf
  g387
  (
    n264,
    n68
  );


  not
  g388
  (
    n378,
    n40
  );


  buf
  g389
  (
    n524,
    n111
  );


  not
  g390
  (
    n281,
    n131
  );


  buf
  g391
  (
    n340,
    n132
  );


  buf
  g392
  (
    n525,
    n136
  );


  not
  g393
  (
    n265,
    n36
  );


  not
  g394
  (
    n229,
    n100
  );


  not
  g395
  (
    n278,
    n84
  );


  not
  g396
  (
    n328,
    n54
  );


  not
  g397
  (
    n454,
    n101
  );


  buf
  g398
  (
    n477,
    n55
  );


  not
  g399
  (
    n514,
    n121
  );


  not
  g400
  (
    n427,
    n74
  );


  buf
  g401
  (
    n522,
    n68
  );


  buf
  g402
  (
    n341,
    n91
  );


  not
  g403
  (
    n269,
    n64
  );


  buf
  g404
  (
    n287,
    n31
  );


  buf
  g405
  (
    n201,
    n70
  );


  buf
  g406
  (
    n457,
    n31
  );


  not
  g407
  (
    n403,
    n121
  );


  not
  g408
  (
    KeyWire_0_18,
    n125
  );


  buf
  g409
  (
    n539,
    n128
  );


  not
  g410
  (
    n286,
    n104
  );


  not
  g411
  (
    n437,
    n43
  );


  buf
  g412
  (
    n408,
    n55
  );


  not
  g413
  (
    n409,
    n97
  );


  buf
  g414
  (
    n337,
    n92
  );


  buf
  g415
  (
    n143,
    n57
  );


  not
  g416
  (
    n482,
    n63
  );


  buf
  g417
  (
    n257,
    n41
  );


  buf
  g418
  (
    n288,
    n115
  );


  buf
  g419
  (
    n163,
    n54
  );


  buf
  g420
  (
    n373,
    n101
  );


  not
  g421
  (
    n471,
    n93
  );


  not
  g422
  (
    n381,
    n85
  );


  not
  g423
  (
    n320,
    n105
  );


  not
  g424
  (
    n547,
    n81
  );


  not
  g425
  (
    n294,
    n32
  );


  not
  g426
  (
    n267,
    n42
  );


  not
  g427
  (
    n309,
    n90
  );


  not
  g428
  (
    n376,
    n94
  );


  not
  g429
  (
    n434,
    n35
  );


  buf
  g430
  (
    n246,
    n109
  );


  not
  g431
  (
    n508,
    n53
  );


  not
  g432
  (
    n176,
    n80
  );


  not
  g433
  (
    n366,
    n127
  );


  buf
  g434
  (
    n144,
    n129
  );


  buf
  g435
  (
    n162,
    n131
  );


  buf
  g436
  (
    n485,
    n127
  );


  not
  g437
  (
    n274,
    n89
  );


  buf
  g438
  (
    n363,
    n112
  );


  buf
  g439
  (
    n473,
    n120
  );


  not
  g440
  (
    n549,
    n127
  );


  not
  g441
  (
    n552,
    n52
  );


  not
  g442
  (
    n185,
    n50
  );


  buf
  g443
  (
    n529,
    n100
  );


  buf
  g444
  (
    n259,
    n46
  );


  buf
  g445
  (
    n532,
    n62
  );


  buf
  g446
  (
    n240,
    n77
  );


  buf
  g447
  (
    n436,
    n92
  );


  not
  g448
  (
    n407,
    n42
  );


  buf
  g449
  (
    n548,
    n85
  );


  buf
  g450
  (
    n442,
    n71
  );


  not
  g451
  (
    n570,
    n86
  );


  not
  g452
  (
    n178,
    n52
  );


  not
  g453
  (
    n323,
    n99
  );


  not
  g454
  (
    n418,
    n110
  );


  buf
  g455
  (
    n206,
    n53
  );


  not
  g456
  (
    n317,
    n74
  );


  not
  g457
  (
    n563,
    n96
  );


  buf
  g458
  (
    n463,
    n38
  );


  buf
  g459
  (
    n312,
    n134
  );


  not
  g460
  (
    n297,
    n75
  );


  not
  g461
  (
    n343,
    n98
  );


  not
  g462
  (
    n225,
    n121
  );


  not
  g463
  (
    n377,
    n137
  );


  buf
  g464
  (
    n339,
    n81
  );


  not
  g465
  (
    n345,
    n67
  );


  buf
  g466
  (
    n252,
    n66
  );


  buf
  g467
  (
    n322,
    n38
  );


  buf
  g468
  (
    n448,
    n41
  );


  not
  g469
  (
    n242,
    n57
  );


  not
  g470
  (
    n501,
    n97
  );


  buf
  g471
  (
    n568,
    n35
  );


  buf
  g472
  (
    n209,
    n123
  );


  buf
  g473
  (
    n421,
    n79
  );


  not
  g474
  (
    n187,
    n74
  );


  not
  g475
  (
    n424,
    n130
  );


  not
  g476
  (
    n250,
    n64
  );


  buf
  g477
  (
    n364,
    n97
  );


  buf
  g478
  (
    n191,
    n116
  );


  buf
  g479
  (
    n271,
    n128
  );


  not
  g480
  (
    n194,
    n45
  );


  buf
  g481
  (
    n268,
    n50
  );


  not
  g482
  (
    n334,
    n124
  );


  not
  g483
  (
    n147,
    n83
  );


  not
  g484
  (
    n254,
    n39
  );


  not
  g485
  (
    n168,
    n56
  );


  buf
  g486
  (
    n186,
    n50
  );


  not
  g487
  (
    n371,
    n40
  );


  not
  g488
  (
    n169,
    n77
  );


  not
  g489
  (
    n530,
    n119
  );


  buf
  g490
  (
    n367,
    n62
  );


  buf
  g491
  (
    n369,
    n133
  );


  buf
  g492
  (
    n445,
    n65
  );


  not
  g493
  (
    n509,
    n129
  );


  buf
  g494
  (
    n486,
    n132
  );


  not
  g495
  (
    n389,
    n33
  );


  not
  g496
  (
    n142,
    n62
  );


  not
  g497
  (
    n358,
    n30
  );


  buf
  g498
  (
    n329,
    n58
  );


  buf
  g499
  (
    n531,
    n54
  );


  buf
  g500
  (
    n488,
    n61
  );


  not
  g501
  (
    n217,
    n33
  );


  buf
  g502
  (
    n411,
    n87
  );


  not
  g503
  (
    n564,
    n64
  );


  not
  g504
  (
    n302,
    n79
  );


  not
  g505
  (
    n433,
    n108
  );


  buf
  g506
  (
    n494,
    n72
  );


  not
  g507
  (
    n566,
    n40
  );


  not
  g508
  (
    n241,
    n78
  );


  not
  g509
  (
    n406,
    n37
  );


  not
  g510
  (
    n333,
    n130
  );


  not
  g511
  (
    n534,
    n41
  );


  not
  g512
  (
    KeyWire_0_5,
    n31
  );


  buf
  g513
  (
    n175,
    n43
  );


  not
  g514
  (
    n402,
    n72
  );


  not
  g515
  (
    n558,
    n103
  );


  not
  g516
  (
    n182,
    n87
  );


  not
  g517
  (
    n347,
    n75
  );


  buf
  g518
  (
    n273,
    n36
  );


  not
  g519
  (
    n461,
    n96
  );


  buf
  g520
  (
    n249,
    n121
  );


  not
  g521
  (
    n291,
    n90
  );


  buf
  g522
  (
    n251,
    n32
  );


  not
  g523
  (
    n479,
    n57
  );


  not
  g524
  (
    n458,
    n134
  );


  buf
  g525
  (
    n476,
    n67
  );


  not
  g526
  (
    n537,
    n138
  );


  buf
  g527
  (
    n245,
    n71
  );


  buf
  g528
  (
    n506,
    n39
  );


  not
  g529
  (
    n255,
    n83
  );


  not
  g530
  (
    n204,
    n115
  );


  not
  g531
  (
    n295,
    n102
  );


  buf
  g532
  (
    n289,
    n126
  );


  buf
  g533
  (
    n319,
    n72
  );


  buf
  g534
  (
    n396,
    n80
  );


  buf
  g535
  (
    n239,
    n86
  );


  not
  g536
  (
    n528,
    n92
  );


  buf
  g537
  (
    n238,
    n62
  );


  not
  g538
  (
    n226,
    n42
  );


  not
  g539
  (
    n557,
    n76
  );


  not
  g540
  (
    n456,
    n135
  );


  not
  g541
  (
    n155,
    n117
  );


  buf
  g542
  (
    n335,
    n125
  );


  buf
  g543
  (
    n560,
    n91
  );


  xor
  g544
  (
    n299,
    n34,
    n59,
    n110,
    n114
  );


  buf
  g545
  (
    n638,
    n477
  );


  not
  g546
  (
    n772,
    n299
  );


  buf
  g547
  (
    n1135,
    n411
  );


  buf
  g548
  (
    n1287,
    n491
  );


  not
  g549
  (
    n1270,
    n263
  );


  not
  g550
  (
    n1003,
    n359
  );


  not
  g551
  (
    n752,
    n307
  );


  not
  g552
  (
    n997,
    n310
  );


  buf
  g553
  (
    n1259,
    n438
  );


  buf
  g554
  (
    n1188,
    n317
  );


  not
  g555
  (
    n1179,
    n162
  );


  not
  g556
  (
    n951,
    n468
  );


  buf
  g557
  (
    n642,
    n254
  );


  buf
  g558
  (
    n1426,
    n384
  );


  not
  g559
  (
    n1187,
    n308
  );


  buf
  g560
  (
    KeyWire_0_23,
    n425
  );


  not
  g561
  (
    n633,
    n492
  );


  buf
  g562
  (
    n687,
    n166
  );


  buf
  g563
  (
    n643,
    n234
  );


  buf
  g564
  (
    n878,
    n397
  );


  buf
  g565
  (
    n973,
    n176
  );


  not
  g566
  (
    n627,
    n428
  );


  not
  g567
  (
    n1493,
    n418
  );


  buf
  g568
  (
    n707,
    n418
  );


  not
  g569
  (
    n1377,
    n469
  );


  buf
  g570
  (
    n1269,
    n451
  );


  not
  g571
  (
    n1407,
    n259
  );


  buf
  g572
  (
    n1038,
    n253
  );


  buf
  g573
  (
    n749,
    n191
  );


  buf
  g574
  (
    n1467,
    n146
  );


  not
  g575
  (
    n1554,
    n282
  );


  buf
  g576
  (
    n1221,
    n370
  );


  not
  g577
  (
    n1042,
    n347
  );


  buf
  g578
  (
    n794,
    n270
  );


  not
  g579
  (
    n832,
    n366
  );


  not
  g580
  (
    n1171,
    n298
  );


  not
  g581
  (
    n802,
    n156
  );


  not
  g582
  (
    n1499,
    n277
  );


  buf
  g583
  (
    n765,
    n384
  );


  buf
  g584
  (
    n1119,
    n315
  );


  not
  g585
  (
    n854,
    n303
  );


  buf
  g586
  (
    n888,
    n458
  );


  buf
  g587
  (
    n587,
    n485
  );


  not
  g588
  (
    n1545,
    n459
  );


  not
  g589
  (
    n1002,
    n395
  );


  buf
  g590
  (
    n1223,
    n278
  );


  buf
  g591
  (
    n726,
    n503
  );


  buf
  g592
  (
    n1552,
    n385
  );


  buf
  g593
  (
    n708,
    n360
  );


  buf
  g594
  (
    n1611,
    n361
  );


  not
  g595
  (
    n1061,
    n446
  );


  buf
  g596
  (
    n579,
    n334
  );


  not
  g597
  (
    n801,
    n432
  );


  not
  g598
  (
    n676,
    n283
  );


  not
  g599
  (
    n1263,
    n220
  );


  not
  g600
  (
    n1564,
    n272
  );


  not
  g601
  (
    n1340,
    n220
  );


  not
  g602
  (
    n1433,
    n390
  );


  not
  g603
  (
    n1265,
    n398
  );


  buf
  g604
  (
    n913,
    n492
  );


  buf
  g605
  (
    n817,
    n256
  );


  not
  g606
  (
    n1448,
    n434
  );


  buf
  g607
  (
    n679,
    n311
  );


  not
  g608
  (
    n1629,
    n375
  );


  buf
  g609
  (
    n1509,
    n285
  );


  buf
  g610
  (
    n791,
    n303
  );


  buf
  g611
  (
    n601,
    n174
  );


  buf
  g612
  (
    n1484,
    n155
  );


  not
  g613
  (
    n1160,
    n351
  );


  buf
  g614
  (
    n1122,
    n298
  );


  not
  g615
  (
    n905,
    n294
  );


  buf
  g616
  (
    n1214,
    n168
  );


  buf
  g617
  (
    n688,
    n272
  );


  buf
  g618
  (
    n1144,
    n338
  );


  not
  g619
  (
    n1030,
    n505
  );


  buf
  g620
  (
    n655,
    n274
  );


  buf
  g621
  (
    n1024,
    n402
  );


  buf
  g622
  (
    n1610,
    n342
  );


  not
  g623
  (
    n1051,
    n421
  );


  not
  g624
  (
    n1117,
    n369
  );


  buf
  g625
  (
    n1514,
    n304
  );


  not
  g626
  (
    KeyWire_0_10,
    n383
  );


  buf
  g627
  (
    n1346,
    n429
  );


  buf
  g628
  (
    n892,
    n351
  );


  buf
  g629
  (
    n703,
    n296
  );


  buf
  g630
  (
    n816,
    n276
  );


  buf
  g631
  (
    n871,
    n278
  );


  not
  g632
  (
    n1374,
    n252
  );


  not
  g633
  (
    n1558,
    n328
  );


  not
  g634
  (
    n833,
    n359
  );


  buf
  g635
  (
    n1078,
    n353
  );


  buf
  g636
  (
    KeyWire_0_1,
    n284
  );


  not
  g637
  (
    n1034,
    n339
  );


  not
  g638
  (
    n1085,
    n334
  );


  not
  g639
  (
    n721,
    n489
  );


  not
  g640
  (
    n744,
    n293
  );


  not
  g641
  (
    n1388,
    n327
  );


  buf
  g642
  (
    n593,
    n359
  );


  buf
  g643
  (
    n1320,
    n506
  );


  buf
  g644
  (
    n729,
    n499
  );


  not
  g645
  (
    n733,
    n253
  );


  buf
  g646
  (
    n1113,
    n474
  );


  buf
  g647
  (
    n1148,
    n179
  );


  not
  g648
  (
    n1413,
    n170
  );


  not
  g649
  (
    n1627,
    n422
  );


  not
  g650
  (
    n1485,
    n353
  );


  not
  g651
  (
    n1440,
    n258
  );


  not
  g652
  (
    n1566,
    n324
  );


  not
  g653
  (
    n1460,
    n316
  );


  not
  g654
  (
    n1011,
    n252
  );


  buf
  g655
  (
    n796,
    n181
  );


  not
  g656
  (
    n1649,
    n316
  );


  buf
  g657
  (
    n1563,
    n229
  );


  buf
  g658
  (
    n1432,
    n329
  );


  not
  g659
  (
    n1017,
    n322
  );


  not
  g660
  (
    n1075,
    n422
  );


  buf
  g661
  (
    n947,
    n346
  );


  buf
  g662
  (
    n1419,
    n493
  );


  buf
  g663
  (
    n640,
    n370
  );


  not
  g664
  (
    n1181,
    n499
  );


  buf
  g665
  (
    n1057,
    n306
  );


  not
  g666
  (
    n699,
    n256
  );


  not
  g667
  (
    n992,
    n442
  );


  buf
  g668
  (
    n641,
    n290
  );


  not
  g669
  (
    n1022,
    n470
  );


  buf
  g670
  (
    n1095,
    n417
  );


  buf
  g671
  (
    n647,
    n152
  );


  buf
  g672
  (
    n1020,
    n317
  );


  not
  g673
  (
    n1193,
    n319
  );


  buf
  g674
  (
    n1530,
    n301
  );


  buf
  g675
  (
    n1533,
    n245
  );


  not
  g676
  (
    n1012,
    n347
  );


  not
  g677
  (
    n1495,
    n207
  );


  buf
  g678
  (
    n800,
    n491
  );


  buf
  g679
  (
    n1196,
    n337
  );


  buf
  g680
  (
    n1162,
    n351
  );


  buf
  g681
  (
    n1508,
    n260
  );


  buf
  g682
  (
    n1539,
    n296
  );


  buf
  g683
  (
    n1121,
    n348
  );


  buf
  g684
  (
    n1202,
    n469
  );


  buf
  g685
  (
    n1476,
    n269
  );


  not
  g686
  (
    n1099,
    n355
  );


  buf
  g687
  (
    n1624,
    n227
  );


  buf
  g688
  (
    n953,
    n334
  );


  not
  g689
  (
    n847,
    n225
  );


  not
  g690
  (
    n691,
    n251
  );


  buf
  g691
  (
    n846,
    n331
  );


  not
  g692
  (
    n827,
    n264
  );


  not
  g693
  (
    n842,
    n452
  );


  not
  g694
  (
    n1520,
    n430
  );


  buf
  g695
  (
    n1050,
    n407
  );


  buf
  g696
  (
    n1466,
    n314
  );


  buf
  g697
  (
    n909,
    n411
  );


  not
  g698
  (
    n1216,
    n385
  );


  buf
  g699
  (
    n669,
    n255
  );


  buf
  g700
  (
    n1067,
    n414
  );


  buf
  g701
  (
    n969,
    n431
  );


  not
  g702
  (
    n1654,
    n413
  );


  not
  g703
  (
    n1178,
    n260
  );


  not
  g704
  (
    n1542,
    n338
  );


  not
  g705
  (
    n1456,
    n383
  );


  not
  g706
  (
    n684,
    n344
  );


  buf
  g707
  (
    n1507,
    n399
  );


  not
  g708
  (
    n773,
    n183
  );


  not
  g709
  (
    n843,
    n324
  );


  not
  g710
  (
    n1199,
    n397
  );


  not
  g711
  (
    n1069,
    n450
  );


  not
  g712
  (
    n853,
    n348
  );


  buf
  g713
  (
    n799,
    n158
  );


  not
  g714
  (
    n1065,
    n346
  );


  not
  g715
  (
    n797,
    n436
  );


  buf
  g716
  (
    n1190,
    n230
  );


  not
  g717
  (
    n884,
    n402
  );


  not
  g718
  (
    n1275,
    n492
  );


  buf
  g719
  (
    n789,
    n273
  );


  not
  g720
  (
    n852,
    n284
  );


  not
  g721
  (
    n1428,
    n413
  );


  buf
  g722
  (
    n883,
    n417
  );


  buf
  g723
  (
    n1568,
    n449
  );


  not
  g724
  (
    n872,
    n446
  );


  buf
  g725
  (
    n666,
    n331
  );


  buf
  g726
  (
    n1583,
    n496
  );


  not
  g727
  (
    n1389,
    n333
  );


  buf
  g728
  (
    n1302,
    n261
  );


  buf
  g729
  (
    n889,
    n476
  );


  buf
  g730
  (
    n683,
    n481
  );


  buf
  g731
  (
    n1289,
    n469
  );


  not
  g732
  (
    n861,
    n487
  );


  buf
  g733
  (
    n682,
    n275
  );


  not
  g734
  (
    n1540,
    n433
  );


  buf
  g735
  (
    n960,
    n173
  );


  buf
  g736
  (
    n1204,
    n314
  );


  buf
  g737
  (
    n989,
    n293
  );


  buf
  g738
  (
    n1070,
    n347
  );


  not
  g739
  (
    n1436,
    n483
  );


  not
  g740
  (
    n1560,
    n339
  );


  not
  g741
  (
    n1532,
    n193
  );


  buf
  g742
  (
    n977,
    n372
  );


  not
  g743
  (
    n646,
    n267
  );


  not
  g744
  (
    n742,
    n244
  );


  not
  g745
  (
    n837,
    n196
  );


  not
  g746
  (
    n1201,
    n502
  );


  not
  g747
  (
    n1597,
    n205
  );


  not
  g748
  (
    n959,
    n248
  );


  buf
  g749
  (
    n1446,
    n378
  );


  buf
  g750
  (
    n1043,
    n330
  );


  buf
  g751
  (
    n1208,
    n314
  );


  not
  g752
  (
    n1515,
    n279
  );


  not
  g753
  (
    n1305,
    n341
  );


  buf
  g754
  (
    n720,
    n291
  );


  not
  g755
  (
    n1161,
    n437
  );


  buf
  g756
  (
    n1329,
    n467
  );


  buf
  g757
  (
    n1536,
    n391
  );


  buf
  g758
  (
    n1096,
    n458
  );


  not
  g759
  (
    n1553,
    n313
  );


  not
  g760
  (
    n1608,
    n306
  );


  not
  g761
  (
    n1115,
    n498
  );


  not
  g762
  (
    n748,
    n366
  );


  not
  g763
  (
    n1548,
    n338
  );


  not
  g764
  (
    n984,
    n373
  );


  not
  g765
  (
    n1079,
    n280
  );


  not
  g766
  (
    n776,
    n455
  );


  buf
  g767
  (
    n1276,
    n398
  );


  buf
  g768
  (
    n1157,
    n463
  );


  buf
  g769
  (
    n1429,
    n345
  );


  not
  g770
  (
    n1307,
    n472
  );


  not
  g771
  (
    n1124,
    n255
  );


  not
  g772
  (
    n1247,
    n424
  );


  buf
  g773
  (
    n656,
    n500
  );


  buf
  g774
  (
    n1209,
    n344
  );


  not
  g775
  (
    n808,
    n476
  );


  not
  g776
  (
    n1631,
    n379
  );


  buf
  g777
  (
    n829,
    n432
  );


  buf
  g778
  (
    n840,
    n247
  );


  buf
  g779
  (
    n1296,
    n283
  );


  not
  g780
  (
    n758,
    n295
  );


  not
  g781
  (
    n732,
    n506
  );


  not
  g782
  (
    n746,
    n411
  );


  buf
  g783
  (
    n1524,
    n268
  );


  buf
  g784
  (
    n1120,
    n392
  );


  not
  g785
  (
    n1225,
    n494
  );


  not
  g786
  (
    n899,
    n458
  );


  not
  g787
  (
    n624,
    n423
  );


  not
  g788
  (
    n974,
    n180
  );


  buf
  g789
  (
    n1251,
    n380
  );


  not
  g790
  (
    n1384,
    n495
  );


  buf
  g791
  (
    n1471,
    n249
  );


  buf
  g792
  (
    n1543,
    n419
  );


  not
  g793
  (
    n615,
    n147
  );


  not
  g794
  (
    n722,
    n292
  );


  not
  g795
  (
    n1430,
    n380
  );


  not
  g796
  (
    n1322,
    n262
  );


  buf
  g797
  (
    n1310,
    n340
  );


  buf
  g798
  (
    n753,
    n326
  );


  buf
  g799
  (
    n589,
    n194
  );


  buf
  g800
  (
    n730,
    n497
  );


  buf
  g801
  (
    KeyWire_0_28,
    n471
  );


  buf
  g802
  (
    n1315,
    n254
  );


  buf
  g803
  (
    n694,
    n280
  );


  not
  g804
  (
    n626,
    n439
  );


  not
  g805
  (
    n1210,
    n141
  );


  not
  g806
  (
    n1084,
    n204
  );


  buf
  g807
  (
    n657,
    n412
  );


  buf
  g808
  (
    n1222,
    n335
  );


  buf
  g809
  (
    n1379,
    n292
  );


  not
  g810
  (
    n771,
    n364
  );


  buf
  g811
  (
    n914,
    n379
  );


  not
  g812
  (
    n1267,
    n368
  );


  buf
  g813
  (
    n900,
    n506
  );


  buf
  g814
  (
    n1596,
    n182
  );


  buf
  g815
  (
    n686,
    n394
  );


  not
  g816
  (
    n716,
    n264
  );


  not
  g817
  (
    n918,
    n489
  );


  not
  g818
  (
    n954,
    n476
  );


  buf
  g819
  (
    n1437,
    n430
  );


  not
  g820
  (
    n1584,
    n251
  );


  not
  g821
  (
    n1279,
    n398
  );


  not
  g822
  (
    n1298,
    n388
  );


  not
  g823
  (
    n1237,
    n250
  );


  buf
  g824
  (
    n671,
    n456
  );


  buf
  g825
  (
    n1444,
    n192
  );


  buf
  g826
  (
    n825,
    n318
  );


  not
  g827
  (
    n1072,
    n310
  );


  not
  g828
  (
    n1080,
    n486
  );


  not
  g829
  (
    n1383,
    n462
  );


  buf
  g830
  (
    n1090,
    n392
  );


  buf
  g831
  (
    n632,
    n410
  );


  not
  g832
  (
    n958,
    n384
  );


  not
  g833
  (
    n792,
    n304
  );


  not
  g834
  (
    n950,
    n257
  );


  buf
  g835
  (
    n1130,
    n453
  );


  not
  g836
  (
    n782,
    n441
  );


  buf
  g837
  (
    n790,
    n419
  );


  buf
  g838
  (
    n1571,
    n376
  );


  not
  g839
  (
    n980,
    n505
  );


  buf
  g840
  (
    n830,
    n497
  );


  not
  g841
  (
    n713,
    n338
  );


  not
  g842
  (
    n1349,
    n256
  );


  buf
  g843
  (
    n1104,
    n502
  );


  buf
  g844
  (
    n844,
    n339
  );


  not
  g845
  (
    n1640,
    n181
  );


  not
  g846
  (
    n1290,
    n260
  );


  not
  g847
  (
    n979,
    n237
  );


  buf
  g848
  (
    n1342,
    n400
  );


  buf
  g849
  (
    n1401,
    n328
  );


  buf
  g850
  (
    n929,
    n450
  );


  buf
  g851
  (
    n762,
    n345
  );


  buf
  g852
  (
    n976,
    n262
  );


  buf
  g853
  (
    n981,
    n504
  );


  buf
  g854
  (
    n1449,
    n355
  );


  buf
  g855
  (
    n709,
    n302
  );


  buf
  g856
  (
    n1353,
    n418
  );


  buf
  g857
  (
    n1273,
    n444
  );


  not
  g858
  (
    n1128,
    n250
  );


  buf
  g859
  (
    n941,
    n330
  );


  not
  g860
  (
    n1612,
    n381
  );


  not
  g861
  (
    n780,
    n279
  );


  not
  g862
  (
    n940,
    n189
  );


  buf
  g863
  (
    n920,
    n457
  );


  buf
  g864
  (
    n1537,
    n445
  );


  buf
  g865
  (
    n818,
    n470
  );


  not
  g866
  (
    n723,
    n393
  );


  buf
  g867
  (
    n674,
    n227
  );


  buf
  g868
  (
    n1395,
    n173
  );


  buf
  g869
  (
    n1111,
    n401
  );


  not
  g870
  (
    n1350,
    n319
  );


  buf
  g871
  (
    n1232,
    n396
  );


  buf
  g872
  (
    n1093,
    n386
  );


  not
  g873
  (
    n1513,
    n309
  );


  not
  g874
  (
    n1100,
    n289
  );


  buf
  g875
  (
    n1459,
    n336
  );


  buf
  g876
  (
    n1458,
    n484
  );


  not
  g877
  (
    n1029,
    n351
  );


  not
  g878
  (
    n779,
    n386
  );


  not
  g879
  (
    n1112,
    n393
  );


  not
  g880
  (
    n1546,
    n280
  );


  not
  g881
  (
    n1323,
    n396
  );


  not
  g882
  (
    n754,
    n199
  );


  buf
  g883
  (
    n1137,
    n302
  );


  not
  g884
  (
    n1600,
    n473
  );


  not
  g885
  (
    n991,
    n433
  );


  not
  g886
  (
    n665,
    n165
  );


  not
  g887
  (
    n1139,
    n442
  );


  not
  g888
  (
    n583,
    n307
  );


  not
  g889
  (
    n1258,
    n444
  );


  not
  g890
  (
    n944,
    n447
  );


  buf
  g891
  (
    n806,
    n406
  );


  buf
  g892
  (
    n724,
    n426
  );


  buf
  g893
  (
    n577,
    n360
  );


  not
  g894
  (
    n933,
    n235
  );


  buf
  g895
  (
    n604,
    n434
  );


  buf
  g896
  (
    n591,
    n426
  );


  not
  g897
  (
    n1044,
    n259
  );


  not
  g898
  (
    n1174,
    n406
  );


  buf
  g899
  (
    n935,
    n503
  );


  not
  g900
  (
    n798,
    n435
  );


  buf
  g901
  (
    n1573,
    n364
  );


  not
  g902
  (
    n1400,
    n413
  );


  buf
  g903
  (
    n1625,
    n410
  );


  buf
  g904
  (
    n1601,
    n342
  );


  not
  g905
  (
    n1632,
    n482
  );


  buf
  g906
  (
    n783,
    n241
  );


  buf
  g907
  (
    n1589,
    n188
  );


  not
  g908
  (
    n644,
    n420
  );


  not
  g909
  (
    n1132,
    n473
  );


  not
  g910
  (
    n1277,
    n142
  );


  buf
  g911
  (
    n1522,
    n274
  );


  not
  g912
  (
    n606,
    n363
  );


  buf
  g913
  (
    n1131,
    n353
  );


  not
  g914
  (
    n1559,
    n461
  );


  not
  g915
  (
    n751,
    n165
  );


  not
  g916
  (
    n660,
    n494
  );


  buf
  g917
  (
    n1510,
    n379
  );


  not
  g918
  (
    n1009,
    n447
  );


  not
  g919
  (
    n693,
    n202
  );


  buf
  g920
  (
    n1382,
    n297
  );


  buf
  g921
  (
    n916,
    n400
  );


  buf
  g922
  (
    n1058,
    n458
  );


  buf
  g923
  (
    n1045,
    n400
  );


  buf
  g924
  (
    n704,
    n352
  );


  buf
  g925
  (
    n1580,
    n170
  );


  buf
  g926
  (
    n826,
    n464
  );


  buf
  g927
  (
    n1217,
    n453
  );


  not
  g928
  (
    n1261,
    n319
  );


  buf
  g929
  (
    n585,
    n455
  );


  buf
  g930
  (
    n1393,
    n374
  );


  buf
  g931
  (
    n896,
    n484
  );


  not
  g932
  (
    n1227,
    n468
  );


  not
  g933
  (
    n845,
    n326
  );


  buf
  g934
  (
    n1005,
    n388
  );


  buf
  g935
  (
    n1420,
    n477
  );


  not
  g936
  (
    n1073,
    n379
  );


  not
  g937
  (
    n1047,
    n190
  );


  not
  g938
  (
    n982,
    n502
  );


  buf
  g939
  (
    n1488,
    n260
  );


  buf
  g940
  (
    n651,
    n467
  );


  buf
  g941
  (
    n811,
    n304
  );


  buf
  g942
  (
    n1218,
    n360
  );


  not
  g943
  (
    n1013,
    n452
  );


  not
  g944
  (
    n957,
    n504
  );


  not
  g945
  (
    n1588,
    n414
  );


  not
  g946
  (
    n1150,
    n343
  );


  not
  g947
  (
    n1511,
    n404
  );


  buf
  g948
  (
    n955,
    n198
  );


  buf
  g949
  (
    n1363,
    n394
  );


  buf
  g950
  (
    n1411,
    n434
  );


  not
  g951
  (
    n1197,
    n479
  );


  buf
  g952
  (
    n922,
    n175
  );


  not
  g953
  (
    n1033,
    n423
  );


  not
  g954
  (
    n1620,
    n313
  );


  buf
  g955
  (
    n1087,
    n504
  );


  not
  g956
  (
    n804,
    n399
  );


  buf
  g957
  (
    n1416,
    n451
  );


  buf
  g958
  (
    n1587,
    n453
  );


  buf
  g959
  (
    n639,
    n331
  );


  buf
  g960
  (
    n868,
    n454
  );


  not
  g961
  (
    n743,
    n299
  );


  not
  g962
  (
    n661,
    n409
  );


  buf
  g963
  (
    n1308,
    n478
  );


  not
  g964
  (
    n670,
    n285
  );


  not
  g965
  (
    n1091,
    n363
  );


  not
  g966
  (
    n1306,
    n236
  );


  not
  g967
  (
    n1191,
    n201
  );


  buf
  g968
  (
    n1235,
    n470
  );


  not
  g969
  (
    n620,
    n383
  );


  buf
  g970
  (
    n1239,
    n224
  );


  buf
  g971
  (
    n927,
    n427
  );


  buf
  g972
  (
    n815,
    n246
  );


  not
  g973
  (
    n1504,
    n247
  );


  not
  g974
  (
    n1301,
    n334
  );


  not
  g975
  (
    n1385,
    n307
  );


  buf
  g976
  (
    n1619,
    n448
  );


  buf
  g977
  (
    n1167,
    n285
  );


  buf
  g978
  (
    n986,
    n339
  );


  buf
  g979
  (
    n1652,
    n370
  );


  not
  g980
  (
    n1538,
    n213
  );


  not
  g981
  (
    n1442,
    n435
  );


  not
  g982
  (
    n1408,
    n261
  );


  buf
  g983
  (
    n893,
    n327
  );


  not
  g984
  (
    n968,
    n364
  );


  buf
  g985
  (
    n1646,
    n482
  );


  not
  g986
  (
    n697,
    n159
  );


  buf
  g987
  (
    n1102,
    n488
  );


  not
  g988
  (
    n696,
    n332
  );


  not
  g989
  (
    n1361,
    n415
  );


  buf
  g990
  (
    n1271,
    n327
  );


  not
  g991
  (
    n1284,
    n183
  );


  not
  g992
  (
    n1396,
    n261
  );


  not
  g993
  (
    n1234,
    n473
  );


  not
  g994
  (
    n1572,
    n479
  );


  not
  g995
  (
    n1316,
    n387
  );


  buf
  g996
  (
    n614,
    n323
  );


  not
  g997
  (
    n698,
    n193
  );


  not
  g998
  (
    n1439,
    n349
  );


  buf
  g999
  (
    n1489,
    n382
  );


  buf
  g1000
  (
    n1282,
    n352
  );


  not
  g1001
  (
    n1101,
    n457
  );


  not
  g1002
  (
    n586,
    n457
  );


  buf
  g1003
  (
    n1074,
    n268
  );


  buf
  g1004
  (
    n770,
    n280
  );


  buf
  g1005
  (
    n1375,
    n402
  );


  not
  g1006
  (
    n983,
    n397
  );


  not
  g1007
  (
    n1286,
    n166
  );


  buf
  g1008
  (
    n737,
    n459
  );


  buf
  g1009
  (
    n705,
    n375
  );


  not
  g1010
  (
    n1339,
    n374
  );


  not
  g1011
  (
    n1630,
    n285
  );


  not
  g1012
  (
    n1355,
    n484
  );


  not
  g1013
  (
    n600,
    n239
  );


  not
  g1014
  (
    n1336,
    n348
  );


  not
  g1015
  (
    n1642,
    n230
  );


  not
  g1016
  (
    n831,
    n286
  );


  buf
  g1017
  (
    n1211,
    n274
  );


  buf
  g1018
  (
    n1206,
    n257
  );


  buf
  g1019
  (
    n1412,
    n244
  );


  not
  g1020
  (
    n895,
    n275
  );


  not
  g1021
  (
    n1392,
    n463
  );


  buf
  g1022
  (
    n851,
    n156
  );


  not
  g1023
  (
    n1081,
    n276
  );


  buf
  g1024
  (
    KeyWire_0_9,
    n333
  );


  buf
  g1025
  (
    n1366,
    n347
  );


  not
  g1026
  (
    n747,
    n488
  );


  not
  g1027
  (
    n760,
    n313
  );


  not
  g1028
  (
    n685,
    n365
  );


  not
  g1029
  (
    n1506,
    n289
  );


  buf
  g1030
  (
    n1519,
    n218
  );


  not
  g1031
  (
    n1365,
    n413
  );


  buf
  g1032
  (
    n1195,
    n441
  );


  not
  g1033
  (
    n803,
    n343
  );


  not
  g1034
  (
    n1189,
    n256
  );


  buf
  g1035
  (
    n1634,
    n422
  );


  buf
  g1036
  (
    n1274,
    n195
  );


  not
  g1037
  (
    n1592,
    n424
  );


  buf
  g1038
  (
    n1593,
    n311
  );


  buf
  g1039
  (
    n1125,
    n365
  );


  buf
  g1040
  (
    n936,
    n416
  );


  not
  g1041
  (
    n867,
    n259
  );


  not
  g1042
  (
    n1257,
    n424
  );


  not
  g1043
  (
    n1557,
    n289
  );


  buf
  g1044
  (
    n648,
    n225
  );


  not
  g1045
  (
    n1337,
    n372
  );


  not
  g1046
  (
    n1586,
    n358
  );


  not
  g1047
  (
    n814,
    n447
  );


  buf
  g1048
  (
    n1372,
    n315
  );


  buf
  g1049
  (
    n971,
    n303
  );


  not
  g1050
  (
    n1487,
    n206
  );


  not
  g1051
  (
    n634,
    n375
  );


  not
  g1052
  (
    n1605,
    n462
  );


  buf
  g1053
  (
    n1606,
    n162
  );


  buf
  g1054
  (
    n1097,
    n349
  );


  not
  g1055
  (
    n668,
    n271
  );


  not
  g1056
  (
    n1590,
    n485
  );


  not
  g1057
  (
    n1578,
    n286
  );


  not
  g1058
  (
    n672,
    n245
  );


  not
  g1059
  (
    n1041,
    n251
  );


  not
  g1060
  (
    n1421,
    n226
  );


  not
  g1061
  (
    n1242,
    n429
  );


  not
  g1062
  (
    n1371,
    n291
  );


  buf
  g1063
  (
    n1481,
    n445
  );


  not
  g1064
  (
    n681,
    n369
  );


  buf
  g1065
  (
    n1457,
    n149
  );


  not
  g1066
  (
    n1126,
    n371
  );


  buf
  g1067
  (
    n1198,
    n178
  );


  buf
  g1068
  (
    n1299,
    n232
  );


  buf
  g1069
  (
    n1358,
    n352
  );


  not
  g1070
  (
    n1082,
    n344
  );


  not
  g1071
  (
    n821,
    n390
  );


  buf
  g1072
  (
    n1123,
    n373
  );


  buf
  g1073
  (
    n735,
    n477
  );


  buf
  g1074
  (
    n1410,
    n395
  );


  buf
  g1075
  (
    n630,
    n286
  );


  not
  g1076
  (
    n882,
    n376
  );


  buf
  g1077
  (
    n1230,
    n239
  );


  buf
  g1078
  (
    n873,
    n463
  );


  buf
  g1079
  (
    n1129,
    n438
  );


  buf
  g1080
  (
    n1356,
    n358
  );


  not
  g1081
  (
    n1262,
    n371
  );


  not
  g1082
  (
    n1406,
    n486
  );


  not
  g1083
  (
    n1528,
    n483
  );


  buf
  g1084
  (
    n1184,
    n409
  );


  not
  g1085
  (
    n999,
    n342
  );


  buf
  g1086
  (
    n1445,
    n455
  );


  buf
  g1087
  (
    KeyWire_0_8,
    n311
  );


  buf
  g1088
  (
    n1417,
    n382
  );


  not
  g1089
  (
    n1638,
    n396
  );


  not
  g1090
  (
    n795,
    n348
  );


  not
  g1091
  (
    n1381,
    n336
  );


  buf
  g1092
  (
    n1330,
    n335
  );


  not
  g1093
  (
    n1354,
    n449
  );


  buf
  g1094
  (
    n1402,
    n473
  );


  buf
  g1095
  (
    n924,
    n451
  );


  buf
  g1096
  (
    n1294,
    n198
  );


  buf
  g1097
  (
    n625,
    n253
  );


  buf
  g1098
  (
    n807,
    n184
  );


  buf
  g1099
  (
    n985,
    n421
  );


  not
  g1100
  (
    n1231,
    n233
  );


  not
  g1101
  (
    n1462,
    n315
  );


  buf
  g1102
  (
    n897,
    n332
  );


  not
  g1103
  (
    n1153,
    n322
  );


  buf
  g1104
  (
    n1016,
    n248
  );


  buf
  g1105
  (
    n949,
    n270
  );


  buf
  g1106
  (
    n1378,
    n250
  );


  buf
  g1107
  (
    n654,
    n291
  );


  buf
  g1108
  (
    n1454,
    n481
  );


  buf
  g1109
  (
    n1317,
    n273
  );


  buf
  g1110
  (
    n1149,
    n441
  );


  not
  g1111
  (
    n987,
    n420
  );


  buf
  g1112
  (
    n715,
    n475
  );


  not
  g1113
  (
    n1328,
    n264
  );


  buf
  g1114
  (
    n1386,
    n290
  );


  not
  g1115
  (
    n894,
    n479
  );


  buf
  g1116
  (
    n1496,
    n357
  );


  not
  g1117
  (
    n967,
    n385
  );


  not
  g1118
  (
    n1529,
    n148
  );


  buf
  g1119
  (
    n1465,
    n454
  );


  not
  g1120
  (
    n1617,
    n261
  );


  buf
  g1121
  (
    n1200,
    n277
  );


  not
  g1122
  (
    n1391,
    n381
  );


  not
  g1123
  (
    n628,
    n405
  );


  buf
  g1124
  (
    n1486,
    n179
  );


  buf
  g1125
  (
    n738,
    n464
  );


  buf
  g1126
  (
    n1173,
    n502
  );


  not
  g1127
  (
    n1059,
    n200
  );


  buf
  g1128
  (
    n1639,
    n363
  );


  not
  g1129
  (
    n1526,
    n501
  );


  not
  g1130
  (
    n653,
    n304
  );


  buf
  g1131
  (
    n942,
    n501
  );


  not
  g1132
  (
    n1203,
    n358
  );


  buf
  g1133
  (
    n823,
    n203
  );


  not
  g1134
  (
    n906,
    n207
  );


  buf
  g1135
  (
    n590,
    n474
  );


  not
  g1136
  (
    n1224,
    n319
  );


  not
  g1137
  (
    n1023,
    n404
  );


  buf
  g1138
  (
    n1168,
    n232
  );


  not
  g1139
  (
    n1362,
    n406
  );


  not
  g1140
  (
    n759,
    n328
  );


  buf
  g1141
  (
    n637,
    n309
  );


  not
  g1142
  (
    n890,
    n494
  );


  buf
  g1143
  (
    n1414,
    n377
  );


  buf
  g1144
  (
    n712,
    n445
  );


  buf
  g1145
  (
    n1046,
    n288
  );


  not
  g1146
  (
    n1064,
    n366
  );


  buf
  g1147
  (
    n1505,
    n274
  );


  not
  g1148
  (
    n1534,
    n434
  );


  not
  g1149
  (
    n1453,
    n320
  );


  buf
  g1150
  (
    n635,
    n276
  );


  not
  g1151
  (
    n1422,
    n138
  );


  not
  g1152
  (
    n1469,
    n275
  );


  not
  g1153
  (
    n1105,
    n167
  );


  not
  g1154
  (
    n1404,
    n376
  );


  not
  g1155
  (
    n848,
    n432
  );


  buf
  g1156
  (
    n1158,
    n491
  );


  not
  g1157
  (
    n1136,
    n174
  );


  not
  g1158
  (
    n1574,
    n356
  );


  not
  g1159
  (
    n750,
    n282
  );


  buf
  g1160
  (
    n1598,
    n308
  );


  buf
  g1161
  (
    n1106,
    n341
  );


  buf
  g1162
  (
    n849,
    n345
  );


  buf
  g1163
  (
    KeyWire_0_17,
    n167
  );


  buf
  g1164
  (
    n652,
    n245
  );


  buf
  g1165
  (
    n881,
    n329
  );


  buf
  g1166
  (
    n777,
    n449
  );


  buf
  g1167
  (
    n1194,
    n271
  );


  buf
  g1168
  (
    n910,
    n427
  );


  buf
  g1169
  (
    n1618,
    n180
  );


  not
  g1170
  (
    n1341,
    n437
  );


  not
  g1171
  (
    n1474,
    n283
  );


  buf
  g1172
  (
    n931,
    n192
  );


  not
  g1173
  (
    n1180,
    n496
  );


  buf
  g1174
  (
    n856,
    n178
  );


  not
  g1175
  (
    n1645,
    n474
  );


  buf
  g1176
  (
    n1450,
    n415
  );


  buf
  g1177
  (
    n1278,
    n287
  );


  buf
  g1178
  (
    n1228,
    n291
  );


  not
  g1179
  (
    n1561,
    n420
  );


  not
  g1180
  (
    n1364,
    n350
  );


  buf
  g1181
  (
    n988,
    n278
  );


  buf
  g1182
  (
    n1060,
    n296
  );


  buf
  g1183
  (
    n1164,
    n312
  );


  not
  g1184
  (
    n875,
    n397
  );


  buf
  g1185
  (
    n1256,
    n305
  );


  not
  g1186
  (
    n1145,
    n446
  );


  buf
  g1187
  (
    n869,
    n427
  );


  not
  g1188
  (
    n1272,
    n153
  );


  not
  g1189
  (
    n1415,
    n425
  );


  not
  g1190
  (
    n1480,
    n321
  );


  buf
  g1191
  (
    KeyWire_0_21,
    n255
  );


  not
  g1192
  (
    n740,
    n373
  );


  buf
  g1193
  (
    n1134,
    n294
  );


  buf
  g1194
  (
    n1418,
    n257
  );


  not
  g1195
  (
    n1525,
    n310
  );


  not
  g1196
  (
    n595,
    n352
  );


  buf
  g1197
  (
    n1004,
    n354
  );


  not
  g1198
  (
    n1018,
    n463
  );


  buf
  g1199
  (
    n1321,
    n315
  );


  buf
  g1200
  (
    n1443,
    n391
  );


  not
  g1201
  (
    n1243,
    n389
  );


  buf
  g1202
  (
    n937,
    n160
  );


  not
  g1203
  (
    n886,
    n403
  );


  buf
  g1204
  (
    n1233,
    n252
  );


  buf
  g1205
  (
    n1019,
    n454
  );


  buf
  g1206
  (
    n915,
    n197
  );


  not
  g1207
  (
    n996,
    n341
  );


  not
  g1208
  (
    n1565,
    n262
  );


  not
  g1209
  (
    n1053,
    n224
  );


  not
  g1210
  (
    n1207,
    n416
  );


  buf
  g1211
  (
    KeyWire_0_27,
    n258
  );


  buf
  g1212
  (
    n1240,
    n249
  );


  buf
  g1213
  (
    n582,
    n487
  );


  not
  g1214
  (
    n1477,
    n505
  );


  buf
  g1215
  (
    n1483,
    n417
  );


  not
  g1216
  (
    n575,
    n233
  );


  buf
  g1217
  (
    n1603,
    n377
  );


  not
  g1218
  (
    n592,
    n212
  );


  not
  g1219
  (
    n1527,
    n388
  );


  not
  g1220
  (
    n828,
    n440
  );


  not
  g1221
  (
    n788,
    n250
  );


  buf
  g1222
  (
    n1501,
    n465
  );


  not
  g1223
  (
    n912,
    n317
  );


  not
  g1224
  (
    n1512,
    n495
  );


  not
  g1225
  (
    n1360,
    n440
  );


  buf
  g1226
  (
    n1517,
    n196
  );


  not
  g1227
  (
    n1156,
    n392
  );


  buf
  g1228
  (
    n725,
    n417
  );


  not
  g1229
  (
    n1521,
    n495
  );


  buf
  g1230
  (
    n902,
    n350
  );


  not
  g1231
  (
    n1604,
    n431
  );


  not
  g1232
  (
    n1063,
    n480
  );


  buf
  g1233
  (
    n1482,
    n464
  );


  buf
  g1234
  (
    n1461,
    n503
  );


  buf
  g1235
  (
    n1464,
    n169
  );


  not
  g1236
  (
    n1028,
    n460
  );


  not
  g1237
  (
    n649,
    n273
  );


  not
  g1238
  (
    n1254,
    n288
  );


  buf
  g1239
  (
    n1498,
    n294
  );


  not
  g1240
  (
    n1479,
    n454
  );


  buf
  g1241
  (
    n766,
    n209
  );


  buf
  g1242
  (
    n1040,
    n263
  );


  buf
  g1243
  (
    n1118,
    n236
  );


  not
  g1244
  (
    n1427,
    n481
  );


  buf
  g1245
  (
    n1491,
    n300
  );


  buf
  g1246
  (
    n964,
    n242
  );


  not
  g1247
  (
    n1248,
    n403
  );


  buf
  g1248
  (
    n1213,
    n259
  );


  buf
  g1249
  (
    n1219,
    n195
  );


  buf
  g1250
  (
    n1140,
    n157
  );


  buf
  g1251
  (
    n692,
    n387
  );


  buf
  g1252
  (
    n629,
    n292
  );


  not
  g1253
  (
    KeyWire_0_16,
    n465
  );


  not
  g1254
  (
    n616,
    n435
  );


  not
  g1255
  (
    n677,
    n364
  );


  buf
  g1256
  (
    n1068,
    n489
  );


  buf
  g1257
  (
    n1089,
    n292
  );


  buf
  g1258
  (
    n581,
    n218
  );


  not
  g1259
  (
    n1653,
    n332
  );


  not
  g1260
  (
    n1052,
    n267
  );


  not
  g1261
  (
    n907,
    n429
  );


  not
  g1262
  (
    n1647,
    n177
  );


  buf
  g1263
  (
    n727,
    n164
  );


  not
  g1264
  (
    n998,
    n143
  );


  not
  g1265
  (
    n1026,
    n204
  );


  buf
  g1266
  (
    n739,
    n184
  );


  buf
  g1267
  (
    n1303,
    n414
  );


  buf
  g1268
  (
    n903,
    n282
  );


  buf
  g1269
  (
    n734,
    n281
  );


  not
  g1270
  (
    n812,
    n362
  );


  not
  g1271
  (
    n1348,
    n219
  );


  buf
  g1272
  (
    n1006,
    n197
  );


  buf
  g1273
  (
    n1576,
    n217
  );


  not
  g1274
  (
    n923,
    n320
  );


  buf
  g1275
  (
    n841,
    n490
  );


  buf
  g1276
  (
    n1351,
    n501
  );


  not
  g1277
  (
    n1447,
    n415
  );


  buf
  g1278
  (
    n1579,
    n341
  );


  buf
  g1279
  (
    n1622,
    n445
  );


  not
  g1280
  (
    n1335,
    n493
  );


  buf
  g1281
  (
    n1648,
    n423
  );


  not
  g1282
  (
    n1643,
    n294
  );


  buf
  g1283
  (
    n925,
    n194
  );


  buf
  g1284
  (
    n578,
    n325
  );


  not
  g1285
  (
    n835,
    n161
  );


  buf
  g1286
  (
    n1037,
    n324
  );


  not
  g1287
  (
    n850,
    n157
  );


  buf
  g1288
  (
    n755,
    n377
  );


  not
  g1289
  (
    n645,
    n219
  );


  not
  g1290
  (
    n1155,
    n295
  );


  not
  g1291
  (
    n1127,
    n238
  );


  buf
  g1292
  (
    n1031,
    n423
  );


  not
  g1293
  (
    n1326,
    n330
  );


  not
  g1294
  (
    n736,
    n249
  );


  not
  g1295
  (
    n1325,
    n336
  );


  not
  g1296
  (
    n1594,
    n392
  );


  buf
  g1297
  (
    n1549,
    n381
  );


  not
  g1298
  (
    n1409,
    n353
  );


  not
  g1299
  (
    n1394,
    n305
  );


  not
  g1300
  (
    n1021,
    n506
  );


  buf
  g1301
  (
    n963,
    n297
  );


  not
  g1302
  (
    n891,
    n401
  );


  buf
  g1303
  (
    n901,
    n322
  );


  buf
  g1304
  (
    n1226,
    n265
  );


  buf
  g1305
  (
    n1249,
    n264
  );


  not
  g1306
  (
    n1015,
    n386
  );


  not
  g1307
  (
    n728,
    n414
  );


  not
  g1308
  (
    n621,
    n299
  );


  not
  g1309
  (
    n1555,
    n287
  );


  not
  g1310
  (
    n658,
    n433
  );


  buf
  g1311
  (
    n1293,
    n329
  );


  not
  g1312
  (
    n675,
    n268
  );


  not
  g1313
  (
    n908,
    n431
  );


  buf
  g1314
  (
    n594,
    n475
  );


  not
  g1315
  (
    n1599,
    n235
  );


  not
  g1316
  (
    n1516,
    n185
  );


  buf
  g1317
  (
    n859,
    n429
  );


  not
  g1318
  (
    n785,
    n240
  );


  not
  g1319
  (
    n1352,
    n468
  );


  buf
  g1320
  (
    n1268,
    n272
  );


  not
  g1321
  (
    n1472,
    n478
  );


  buf
  g1322
  (
    n623,
    n305
  );


  not
  g1323
  (
    n1098,
    n350
  );


  buf
  g1324
  (
    n898,
    n439
  );


  not
  g1325
  (
    n1027,
    n323
  );


  buf
  g1326
  (
    n612,
    n408
  );


  not
  g1327
  (
    n879,
    n211
  );


  buf
  g1328
  (
    n1369,
    n378
  );


  buf
  g1329
  (
    n1380,
    n186
  );


  not
  g1330
  (
    n1569,
    n342
  );


  not
  g1331
  (
    n978,
    n442
  );


  buf
  g1332
  (
    n1327,
    n221
  );


  buf
  g1333
  (
    n943,
    n302
  );


  not
  g1334
  (
    n819,
    n210
  );


  buf
  g1335
  (
    n1455,
    n443
  );


  buf
  g1336
  (
    n745,
    n245
  );


  buf
  g1337
  (
    n576,
    n480
  );


  not
  g1338
  (
    n1334,
    n370
  );


  buf
  g1339
  (
    n1628,
    n298
  );


  buf
  g1340
  (
    n1116,
    n321
  );


  buf
  g1341
  (
    n887,
    n273
  );


  buf
  g1342
  (
    n874,
    n343
  );


  not
  g1343
  (
    n607,
    n498
  );


  buf
  g1344
  (
    n741,
    n255
  );


  not
  g1345
  (
    n919,
    n265
  );


  buf
  g1346
  (
    n917,
    n453
  );


  buf
  g1347
  (
    n580,
    n320
  );


  buf
  g1348
  (
    n602,
    n477
  );


  not
  g1349
  (
    n613,
    n484
  );


  not
  g1350
  (
    n1295,
    n487
  );


  not
  g1351
  (
    n1387,
    n503
  );


  buf
  g1352
  (
    n1212,
    n410
  );


  not
  g1353
  (
    n855,
    n493
  );


  buf
  g1354
  (
    n1138,
    n160
  );


  not
  g1355
  (
    n1220,
    n321
  );


  buf
  g1356
  (
    n1497,
    n185
  );


  not
  g1357
  (
    n764,
    n428
  );


  buf
  g1358
  (
    n618,
    n316
  );


  not
  g1359
  (
    n1502,
    n296
  );


  not
  g1360
  (
    n948,
    n461
  );


  not
  g1361
  (
    n1370,
    n270
  );


  not
  g1362
  (
    n1032,
    n358
  );


  not
  g1363
  (
    n1347,
    n335
  );


  not
  g1364
  (
    n1470,
    n466
  );


  buf
  g1365
  (
    n1585,
    n306
  );


  buf
  g1366
  (
    n1280,
    n365
  );


  buf
  g1367
  (
    n793,
    n216
  );


  not
  g1368
  (
    n1088,
    n469
  );


  buf
  g1369
  (
    n1405,
    n313
  );


  buf
  g1370
  (
    n1390,
    n462
  );


  not
  g1371
  (
    n1007,
    n487
  );


  buf
  g1372
  (
    n838,
    n266
  );


  buf
  g1373
  (
    n1159,
    n281
  );


  buf
  g1374
  (
    n1451,
    n490
  );


  buf
  g1375
  (
    n809,
    n276
  );


  buf
  g1376
  (
    n667,
    n286
  );


  not
  g1377
  (
    n1172,
    n301
  );


  not
  g1378
  (
    n1338,
    n460
  );


  buf
  g1379
  (
    n1367,
    n217
  );


  buf
  g1380
  (
    n617,
    n333
  );


  buf
  g1381
  (
    n778,
    n440
  );


  not
  g1382
  (
    n1651,
    n145
  );


  buf
  g1383
  (
    n1241,
    n401
  );


  not
  g1384
  (
    n605,
    n139
  );


  buf
  g1385
  (
    n1518,
    n212
  );


  not
  g1386
  (
    n597,
    n425
  );


  not
  g1387
  (
    n636,
    n214
  );


  not
  g1388
  (
    n1636,
    n376
  );


  buf
  g1389
  (
    n1616,
    n345
  );


  buf
  g1390
  (
    n1637,
    n340
  );


  not
  g1391
  (
    n757,
    n471
  );


  buf
  g1392
  (
    n1010,
    n442
  );


  buf
  g1393
  (
    n588,
    n400
  );


  buf
  g1394
  (
    n1633,
    n391
  );


  not
  g1395
  (
    n1368,
    n327
  );


  buf
  g1396
  (
    n990,
    n248
  );


  not
  g1397
  (
    n1283,
    n449
  );


  not
  g1398
  (
    n1077,
    n324
  );


  not
  g1399
  (
    n1062,
    n329
  );


  not
  g1400
  (
    n695,
    n408
  );


  not
  g1401
  (
    n598,
    n277
  );


  buf
  g1402
  (
    n1094,
    n412
  );


  buf
  g1403
  (
    n1500,
    n288
  );


  buf
  g1404
  (
    n939,
    n478
  );


  buf
  g1405
  (
    n1141,
    n267
  );


  not
  g1406
  (
    n1582,
    n271
  );


  not
  g1407
  (
    n1478,
    n377
  );


  buf
  g1408
  (
    n1281,
    n288
  );


  not
  g1409
  (
    n1001,
    n470
  );


  buf
  g1410
  (
    n932,
    n432
  );


  buf
  g1411
  (
    n1054,
    n246
  );


  not
  g1412
  (
    n1551,
    n266
  );


  buf
  g1413
  (
    n1595,
    n357
  );


  not
  g1414
  (
    n1035,
    n430
  );


  buf
  g1415
  (
    n860,
    n381
  );


  not
  g1416
  (
    n689,
    n246
  );


  not
  g1417
  (
    n1152,
    n443
  );


  not
  g1418
  (
    n1253,
    n208
  );


  not
  g1419
  (
    n784,
    n326
  );


  buf
  g1420
  (
    n994,
    n246
  );


  buf
  g1421
  (
    n956,
    n215
  );


  buf
  g1422
  (
    n877,
    n450
  );


  buf
  g1423
  (
    n1399,
    n279
  );


  not
  g1424
  (
    n664,
    n140
  );


  buf
  g1425
  (
    n1244,
    n481
  );


  buf
  g1426
  (
    n921,
    n263
  );


  buf
  g1427
  (
    n1403,
    n471
  );


  buf
  g1428
  (
    n863,
    n419
  );


  buf
  g1429
  (
    n719,
    n362
  );


  not
  g1430
  (
    n1556,
    n399
  );


  buf
  g1431
  (
    n1170,
    n169
  );


  buf
  g1432
  (
    n1163,
    n480
  );


  not
  g1433
  (
    n1577,
    n262
  );


  buf
  g1434
  (
    n1169,
    n383
  );


  buf
  g1435
  (
    n1291,
    n408
  );


  not
  g1436
  (
    n926,
    n452
  );


  buf
  g1437
  (
    n1108,
    n507
  );


  buf
  g1438
  (
    n622,
    n299
  );


  buf
  g1439
  (
    n574,
    n231
  );


  not
  g1440
  (
    n1083,
    n418
  );


  not
  g1441
  (
    n1602,
    n460
  );


  buf
  g1442
  (
    n1550,
    n385
  );


  buf
  g1443
  (
    n767,
    n465
  );


  buf
  g1444
  (
    n584,
    n206
  );


  buf
  g1445
  (
    n1183,
    n238
  );


  buf
  g1446
  (
    n663,
    n284
  );


  not
  g1447
  (
    n1621,
    n407
  );


  buf
  g1448
  (
    n1048,
    n287
  );


  buf
  g1449
  (
    n1110,
    n466
  );


  buf
  g1450
  (
    n934,
    n208
  );


  buf
  g1451
  (
    n1641,
    n361
  );


  not
  g1452
  (
    n701,
    n202
  );


  not
  g1453
  (
    n1373,
    n427
  );


  not
  g1454
  (
    n1297,
    n223
  );


  not
  g1455
  (
    n1151,
    n374
  );


  buf
  g1456
  (
    n1175,
    n355
  );


  not
  g1457
  (
    n608,
    n390
  );


  buf
  g1458
  (
    n1055,
    n226
  );


  not
  g1459
  (
    n1103,
    n461
  );


  not
  g1460
  (
    n1541,
    n237
  );


  not
  g1461
  (
    n952,
    n357
  );


  not
  g1462
  (
    n1314,
    n490
  );


  not
  g1463
  (
    n1609,
    n244
  );


  not
  g1464
  (
    n1357,
    n460
  );


  buf
  g1465
  (
    n1650,
    n398
  );


  not
  g1466
  (
    n1182,
    n247
  );


  not
  g1467
  (
    n928,
    n426
  );


  not
  g1468
  (
    n710,
    n332
  );


  not
  g1469
  (
    n839,
    n501
  );


  not
  g1470
  (
    n774,
    n436
  );


  buf
  g1471
  (
    n631,
    n354
  );


  not
  g1472
  (
    n1288,
    n222
  );


  not
  g1473
  (
    n659,
    n306
  );


  buf
  g1474
  (
    n1441,
    n253
  );


  buf
  g1475
  (
    n961,
    n321
  );


  buf
  g1476
  (
    n619,
    n412
  );


  not
  g1477
  (
    n1434,
    n497
  );


  buf
  g1478
  (
    n1318,
    n439
  );


  not
  g1479
  (
    n805,
    n420
  );


  not
  g1480
  (
    n1397,
    n269
  );


  buf
  g1481
  (
    n717,
    n361
  );


  not
  g1482
  (
    n690,
    n393
  );


  buf
  g1483
  (
    n768,
    n281
  );


  buf
  g1484
  (
    n1146,
    n307
  );


  buf
  g1485
  (
    n1425,
    n394
  );


  not
  g1486
  (
    n1613,
    n378
  );


  buf
  g1487
  (
    n1229,
    n486
  );


  buf
  g1488
  (
    n834,
    n176
  );


  buf
  g1489
  (
    n1575,
    n314
  );


  buf
  g1490
  (
    n1614,
    n172
  );


  not
  g1491
  (
    n1490,
    n171
  );


  buf
  g1492
  (
    n810,
    n283
  );


  not
  g1493
  (
    n870,
    n440
  );


  buf
  g1494
  (
    n1236,
    n498
  );


  buf
  g1495
  (
    n1025,
    n369
  );


  not
  g1496
  (
    n1246,
    n491
  );


  buf
  g1497
  (
    n995,
    n474
  );


  not
  g1498
  (
    n1036,
    n325
  );


  buf
  g1499
  (
    n966,
    n325
  );


  buf
  g1500
  (
    n1398,
    n366
  );


  buf
  g1501
  (
    n673,
    n354
  );


  buf
  g1502
  (
    n650,
    n265
  );


  buf
  g1503
  (
    n1176,
    n325
  );


  not
  g1504
  (
    n706,
    n249
  );


  not
  g1505
  (
    n1071,
    n410
  );


  not
  g1506
  (
    n1423,
    n367
  );


  not
  g1507
  (
    n972,
    n466
  );


  not
  g1508
  (
    n596,
    n316
  );


  not
  g1509
  (
    n1547,
    n479
  );


  buf
  g1510
  (
    n678,
    n263
  );


  not
  g1511
  (
    n1473,
    n436
  );


  not
  g1512
  (
    n1635,
    n189
  );


  not
  g1513
  (
    n904,
    n344
  );


  buf
  g1514
  (
    n1142,
    n426
  );


  not
  g1515
  (
    n1463,
    n387
  );


  buf
  g1516
  (
    n1311,
    n190
  );


  buf
  g1517
  (
    n1304,
    n231
  );


  not
  g1518
  (
    n1324,
    n311
  );


  not
  g1519
  (
    n858,
    n467
  );


  not
  g1520
  (
    n1313,
    n248
  );


  buf
  g1521
  (
    n945,
    n308
  );


  not
  g1522
  (
    n1014,
    n478
  );


  not
  g1523
  (
    n756,
    n318
  );


  buf
  g1524
  (
    n1250,
    n375
  );


  buf
  g1525
  (
    n1345,
    n415
  );


  not
  g1526
  (
    n1438,
    n450
  );


  buf
  g1527
  (
    n1492,
    n168
  );


  not
  g1528
  (
    n731,
    n271
  );


  buf
  g1529
  (
    n1039,
    n483
  );


  not
  g1530
  (
    n1264,
    n380
  );


  buf
  g1531
  (
    n1544,
    n284
  );


  not
  g1532
  (
    n880,
    n363
  );


  not
  g1533
  (
    n965,
    n356
  );


  not
  g1534
  (
    n611,
    n456
  );


  not
  g1535
  (
    n1331,
    n482
  );


  not
  g1536
  (
    n1166,
    n365
  );


  buf
  g1537
  (
    n1531,
    n437
  );


  not
  g1538
  (
    n1644,
    n320
  );


  not
  g1539
  (
    n865,
    n215
  );


  buf
  g1540
  (
    n970,
    n300
  );


  buf
  g1541
  (
    n1591,
    n448
  );


  not
  g1542
  (
    n946,
    n300
  );


  buf
  g1543
  (
    n1008,
    n318
  );


  buf
  g1544
  (
    n1133,
    n251
  );


  not
  g1545
  (
    n1107,
    n268
  );


  not
  g1546
  (
    n711,
    n485
  );


  not
  g1547
  (
    n1468,
    n504
  );


  not
  g1548
  (
    n603,
    n340
  );


  buf
  g1549
  (
    n1503,
    n405
  );


  buf
  g1550
  (
    n1066,
    n451
  );


  buf
  g1551
  (
    n609,
    n333
  );


  buf
  g1552
  (
    n787,
    n372
  );


  buf
  g1553
  (
    n822,
    n447
  );


  buf
  g1554
  (
    n763,
    n350
  );


  not
  g1555
  (
    n1626,
    n221
  );


  not
  g1556
  (
    n1086,
    n356
  );


  not
  g1557
  (
    n1435,
    n428
  );


  not
  g1558
  (
    n786,
    n467
  );


  not
  g1559
  (
    n1615,
    n389
  );


  not
  g1560
  (
    n599,
    n278
  );


  buf
  g1561
  (
    n1300,
    n403
  );


  buf
  g1562
  (
    n1238,
    n290
  );


  buf
  g1563
  (
    n1000,
    n448
  );


  buf
  g1564
  (
    n1319,
    n496
  );


  buf
  g1565
  (
    n864,
    n444
  );


  not
  g1566
  (
    n680,
    n371
  );


  buf
  g1567
  (
    n761,
    n404
  );


  buf
  g1568
  (
    n1570,
    n438
  );


  buf
  g1569
  (
    n1245,
    n317
  );


  not
  g1570
  (
    n1177,
    n495
  );


  and
  g1571
  (
    n1655,
    n161,
    n211,
    n356,
    n438
  );


  xnor
  g1572
  (
    n1494,
    n497,
    n382,
    n496,
    n367
  );


  nand
  g1573
  (
    n862,
    n407,
    n430,
    n369,
    n298
  );


  nor
  g1574
  (
    n1215,
    n200,
    n309,
    n403,
    n163
  );


  nor
  g1575
  (
    n1109,
    n367,
    n265,
    n301,
    n455
  );


  nor
  g1576
  (
    n1376,
    n362,
    n175,
    n401,
    n210
  );


  or
  g1577
  (
    n1114,
    n483,
    n312,
    n328,
    n269
  );


  xnor
  g1578
  (
    n1431,
    n158,
    n480,
    n330,
    n269
  );


  nor
  g1579
  (
    n1452,
    n267,
    n505,
    n229,
    n374
  );


  nor
  g1580
  (
    n1523,
    n373,
    n500,
    n421,
    n359
  );


  xnor
  g1581
  (
    n975,
    n404,
    n187,
    n312,
    n372
  );


  nor
  g1582
  (
    n824,
    n318,
    n472,
    n411,
    n475
  );


  or
  g1583
  (
    n714,
    n216,
    n368,
    n490,
    n389
  );


  nor
  g1584
  (
    n876,
    n441,
    n382,
    n337,
    n393
  );


  nor
  g1585
  (
    n1252,
    n472,
    n443,
    n346,
    n154
  );


  nand
  g1586
  (
    n1186,
    n254,
    n425,
    n448,
    n357
  );


  xor
  g1587
  (
    n1292,
    n159,
    n424,
    n367,
    n391
  );


  nand
  g1588
  (
    n1424,
    n243,
    n433,
    n475,
    n456
  );


  xor
  g1589
  (
    n1147,
    n222,
    n310,
    n151,
    n466
  );


  or
  g1590
  (
    n1344,
    n464,
    n465,
    n290,
    n355
  );


  or
  g1591
  (
    n702,
    n199,
    n254,
    n337,
    n297
  );


  xnor
  g1592
  (
    n1535,
    n498,
    n459,
    n247,
    n293
  );


  xor
  g1593
  (
    n1143,
    n277,
    n407,
    n163,
    n349
  );


  xor
  g1594
  (
    n1332,
    n323,
    n396,
    n472,
    n295
  );


  nor
  g1595
  (
    n1192,
    n395,
    n387,
    n389,
    n272
  );


  xnor
  g1596
  (
    n1343,
    n214,
    n155,
    n409,
    n459
  );


  nand
  g1597
  (
    n1285,
    n164,
    n258,
    n228,
    n408
  );


  or
  g1598
  (
    n1567,
    n326,
    n144,
    n172,
    n293
  );


  or
  g1599
  (
    n775,
    n435,
    n203,
    n266,
    n499
  );


  xor
  g1600
  (
    n1260,
    n252,
    n302,
    n213,
    n488
  );


  xnor
  g1601
  (
    n700,
    n187,
    n266,
    n171,
    n489
  );


  xnor
  g1602
  (
    n1581,
    n371,
    n346,
    n471,
    n488
  );


  xor
  g1603
  (
    n930,
    n308,
    n309,
    n354,
    n279
  );


  or
  g1604
  (
    n1092,
    n419,
    n452,
    n412,
    n499
  );


  or
  g1605
  (
    n1056,
    n191,
    n305,
    n456,
    n500
  );


  xor
  g1606
  (
    n1266,
    n303,
    n209,
    n336,
    n297
  );


  nand
  g1607
  (
    n857,
    n405,
    n138,
    n422,
    n340
  );


  xnor
  g1608
  (
    n820,
    n462,
    n301,
    n349,
    n380
  );


  or
  g1609
  (
    n1255,
    n228,
    n312,
    n493,
    n335
  );


  xnor
  g1610
  (
    n885,
    n386,
    n282,
    n150,
    n322
  );


  nand
  g1611
  (
    n993,
    n436,
    n399,
    n507,
    n368
  );


  xor
  g1612
  (
    n813,
    n406,
    n258,
    n431,
    n485
  );


  xnor
  g1613
  (
    n1623,
    n384,
    n457,
    n343,
    n241
  );


  or
  g1614
  (
    n1475,
    n409,
    n421,
    n289,
    n378
  );


  and
  g1615
  (
    n866,
    n182,
    n188,
    n494,
    n444
  );


  xnor
  g1616
  (
    n1165,
    n486,
    n281,
    n395,
    n476
  );


  nand
  g1617
  (
    n718,
    n388,
    n295,
    n201,
    n360
  );


  nand
  g1618
  (
    KeyWire_0_31,
    n402,
    n492,
    n482,
    n416
  );


  and
  g1619
  (
    n911,
    n243,
    n468,
    n205,
    n287
  );


  nand
  g1620
  (
    n1359,
    n443,
    n394,
    n428,
    n331
  );


  xor
  g1621
  (
    n769,
    n500,
    n405,
    n439,
    n368
  );


  or
  g1622
  (
    n1049,
    n361,
    n437,
    n177,
    n362
  );


  and
  g1623
  (
    n781,
    n461,
    n242,
    n240,
    n300
  );


  xnor
  g1624
  (
    n1309,
    n390,
    n234,
    n337,
    n270
  );


  nand
  g1625
  (
    n1185,
    n257,
    n223,
    n416,
    n446
  );


  xnor
  g1626
  (
    n1154,
    n323,
    n244,
    n186,
    n275
  );


  xnor
  g1627
  (
    n1893,
    n1407,
    n614,
    n1409,
    n1206
  );


  or
  g1628
  (
    n1925,
    n1071,
    n615,
    n1280,
    n708
  );


  xor
  g1629
  (
    n1728,
    n1607,
    n1438,
    n1403,
    n1308
  );


  xor
  g1630
  (
    n1908,
    n545,
    n1055,
    n1531,
    n1429
  );


  xor
  g1631
  (
    n1809,
    n1588,
    n569,
    n1237,
    n541
  );


  and
  g1632
  (
    n1891,
    n757,
    n748,
    n1067,
    n691
  );


  nor
  g1633
  (
    n1716,
    n963,
    n1184,
    n1470,
    n838
  );


  xnor
  g1634
  (
    n1942,
    n802,
    n700,
    n860,
    n903
  );


  xnor
  g1635
  (
    n1778,
    n752,
    n889,
    n559,
    n1436
  );


  or
  g1636
  (
    n1856,
    n951,
    n1513,
    n1105,
    n1213
  );


  or
  g1637
  (
    n1820,
    n1354,
    n1381,
    n1503,
    n1271
  );


  and
  g1638
  (
    n1664,
    n559,
    n1239,
    n893,
    n1589
  );


  nand
  g1639
  (
    n1873,
    n900,
    n531,
    n1561,
    n547
  );


  nand
  g1640
  (
    n1827,
    n602,
    n1463,
    n1427,
    n552
  );


  or
  g1641
  (
    n1876,
    n880,
    n948,
    n1343,
    n529
  );


  nor
  g1642
  (
    n1730,
    n715,
    n1501,
    n534,
    n1113
  );


  xor
  g1643
  (
    n1732,
    n1433,
    n1051,
    n1246,
    n910
  );


  and
  g1644
  (
    n1890,
    n556,
    n756,
    n551,
    n1388
  );


  nand
  g1645
  (
    n1813,
    n1574,
    n682,
    n688,
    n527
  );


  or
  g1646
  (
    n1864,
    n508,
    n1360,
    n586,
    n544
  );


  nand
  g1647
  (
    n1862,
    n1248,
    n1182,
    n1192,
    n535
  );


  nand
  g1648
  (
    n1945,
    n1514,
    n565,
    n1525,
    n558
  );


  or
  g1649
  (
    n1738,
    n517,
    n913,
    n994,
    n858
  );


  and
  g1650
  (
    KeyWire_0_15,
    n1181,
    n1201,
    n735,
    n1143
  );


  nand
  g1651
  (
    n1914,
    n1139,
    n803,
    n550,
    n531
  );


  xnor
  g1652
  (
    n1806,
    n1147,
    n1145,
    n1315,
    n1205
  );


  and
  g1653
  (
    n1805,
    n1008,
    n837,
    n697,
    n1459
  );


  nand
  g1654
  (
    n1741,
    n1200,
    n1536,
    n1088,
    n797
  );


  nor
  g1655
  (
    n1757,
    n746,
    n1332,
    n1521,
    n1411
  );


  xnor
  g1656
  (
    n1760,
    n513,
    n689,
    n1496,
    n1049
  );


  xnor
  g1657
  (
    n1794,
    n1202,
    n1598,
    n1207,
    n706
  );


  nand
  g1658
  (
    n1743,
    n1254,
    n543,
    n1408,
    n549
  );


  xor
  g1659
  (
    n1929,
    n1163,
    n890,
    n507,
    n1177
  );


  xor
  g1660
  (
    n1769,
    n778,
    n1001,
    n510,
    n1507
  );


  nand
  g1661
  (
    n1814,
    n1210,
    n1204,
    n695,
    n1465
  );


  and
  g1662
  (
    n1754,
    n1357,
    n1477,
    n1069,
    n606
  );


  nor
  g1663
  (
    n1679,
    n551,
    n1242,
    n1196,
    n1223
  );


  xor
  g1664
  (
    n1709,
    n1327,
    n1535,
    n564,
    n978
  );


  nand
  g1665
  (
    n1676,
    n1080,
    n1258,
    n1518,
    n1461
  );


  and
  g1666
  (
    n1681,
    n514,
    n865,
    n1211,
    n1547
  );


  nor
  g1667
  (
    n1735,
    n1156,
    n1290,
    n887,
    n1570
  );


  nand
  g1668
  (
    n1901,
    n810,
    n592,
    n546,
    n1291
  );


  nor
  g1669
  (
    n1686,
    n664,
    n817,
    n1270,
    n1064
  );


  xor
  g1670
  (
    n1711,
    n539,
    n526,
    n535,
    n1033
  );


  nor
  g1671
  (
    n1838,
    n829,
    n852,
    n699,
    n971
  );


  nand
  g1672
  (
    n1699,
    n513,
    n1014,
    n1367,
    n539
  );


  and
  g1673
  (
    n1882,
    n598,
    n909,
    n894,
    n1344
  );


  nor
  g1674
  (
    n1960,
    n1041,
    n535,
    n565,
    n509
  );


  xor
  g1675
  (
    n1782,
    n966,
    n672,
    n1331,
    n995
  );


  nor
  g1676
  (
    n1958,
    n1121,
    n635,
    n623,
    n1379
  );


  xor
  g1677
  (
    n1956,
    n515,
    n764,
    n1347,
    n1095
  );


  xnor
  g1678
  (
    n1853,
    n647,
    n848,
    n828,
    n1288
  );


  or
  g1679
  (
    n1957,
    n806,
    n1552,
    n1262,
    n1126
  );


  and
  g1680
  (
    n1829,
    n1148,
    n891,
    n749,
    n1544
  );


  and
  g1681
  (
    n1911,
    n509,
    n1212,
    n805,
    n768
  );


  or
  g1682
  (
    n1719,
    n1530,
    n518,
    n1311,
    n1078
  );


  and
  g1683
  (
    n1823,
    n524,
    n1479,
    n1369,
    n545
  );


  xnor
  g1684
  (
    n1858,
    n1593,
    n997,
    n625,
    n1310
  );


  xnor
  g1685
  (
    n1811,
    n1091,
    n621,
    n785,
    n552
  );


  or
  g1686
  (
    n1896,
    n530,
    n1128,
    n1303,
    n1557
  );


  and
  g1687
  (
    n1780,
    n551,
    n545,
    n876,
    n1592
  );


  xor
  g1688
  (
    n1788,
    n605,
    n1222,
    n915,
    n1572
  );


  and
  g1689
  (
    n1791,
    n1397,
    n638,
    n526,
    n1543
  );


  xnor
  g1690
  (
    n1768,
    n1251,
    n1434,
    n892,
    n1172
  );


  xor
  g1691
  (
    n1726,
    n546,
    n518,
    n1233,
    n954
  );


  and
  g1692
  (
    n1656,
    n1522,
    n1187,
    n525,
    n1125
  );


  xor
  g1693
  (
    n1944,
    n540,
    n704,
    n1000,
    n554
  );


  nor
  g1694
  (
    n1867,
    n899,
    n710,
    n1102,
    n944
  );


  xnor
  g1695
  (
    n1954,
    n1556,
    n517,
    n631,
    n888
  );


  nor
  g1696
  (
    n1690,
    n1371,
    n1460,
    n917,
    n637
  );


  or
  g1697
  (
    n1961,
    n762,
    n886,
    n885,
    n1442
  );


  or
  g1698
  (
    n1963,
    n1273,
    n1165,
    n1019,
    n1319
  );


  and
  g1699
  (
    n1669,
    n1261,
    n1099,
    n1101,
    n680
  );


  nor
  g1700
  (
    n1887,
    n1219,
    n533,
    n1214,
    n759
  );


  nor
  g1701
  (
    n1841,
    n1416,
    n1450,
    n1399,
    n1027
  );


  nor
  g1702
  (
    n1915,
    n717,
    n1474,
    n1068,
    n564
  );


  nor
  g1703
  (
    n1804,
    n552,
    n550,
    n1505,
    n607
  );


  and
  g1704
  (
    KeyWire_0_19,
    n984,
    n713,
    n517,
    n1578
  );


  nand
  g1705
  (
    n1787,
    n564,
    n1188,
    n1284,
    n675
  );


  and
  g1706
  (
    n1712,
    n541,
    n942,
    n1337,
    n1137
  );


  and
  g1707
  (
    n1830,
    n1401,
    n1155,
    n510,
    n1045
  );


  or
  g1708
  (
    n1935,
    n1282,
    n1036,
    n1523,
    n780
  );


  xor
  g1709
  (
    n1912,
    n1092,
    n1455,
    n1151,
    n619
  );


  and
  g1710
  (
    n1872,
    n1435,
    n1065,
    n1604,
    n839
  );


  nand
  g1711
  (
    n1949,
    n569,
    n617,
    n1256,
    n1278
  );


  nand
  g1712
  (
    n1817,
    n1353,
    n929,
    n1185,
    n977
  );


  and
  g1713
  (
    n1668,
    n630,
    n914,
    n1255,
    n763
  );


  xnor
  g1714
  (
    n1696,
    n832,
    n1502,
    n822,
    n1035
  );


  nand
  g1715
  (
    n1678,
    n1026,
    n576,
    n769,
    n653
  );


  nand
  g1716
  (
    n1865,
    n976,
    n1224,
    n546,
    n1410
  );


  nor
  g1717
  (
    n1724,
    n520,
    n703,
    n898,
    n729
  );


  xor
  g1718
  (
    n1680,
    n527,
    n1456,
    n539,
    n1558
  );


  nor
  g1719
  (
    n1874,
    n1473,
    n671,
    n935,
    n1186
  );


  and
  g1720
  (
    n1907,
    n1596,
    n1272,
    n730,
    n801
  );


  and
  g1721
  (
    n1878,
    n1425,
    n1393,
    n1484,
    n941
  );


  or
  g1722
  (
    n1799,
    n582,
    n1142,
    n720,
    n1516
  );


  nor
  g1723
  (
    n1884,
    n813,
    n1216,
    n799,
    n820
  );


  and
  g1724
  (
    n1842,
    n724,
    n590,
    n959,
    n1312
  );


  nor
  g1725
  (
    n1847,
    n520,
    n1325,
    n524,
    n1573
  );


  and
  g1726
  (
    n1670,
    n1002,
    n1046,
    n1526,
    n1231
  );


  xor
  g1727
  (
    n1926,
    n1372,
    n528,
    n783,
    n513
  );


  xnor
  g1728
  (
    n1752,
    n609,
    n1333,
    n549,
    n1532
  );


  nand
  g1729
  (
    n1753,
    n1517,
    n516,
    n1448,
    n754
  );


  and
  g1730
  (
    n1698,
    n1220,
    n597,
    n767,
    n1096
  );


  and
  g1731
  (
    n1746,
    n1383,
    n1153,
    n869,
    n1447
  );


  or
  g1732
  (
    n1930,
    n1400,
    n1039,
    n1395,
    n574
  );


  or
  g1733
  (
    n1871,
    n1351,
    n874,
    n622,
    n1412
  );


  or
  g1734
  (
    n1703,
    n516,
    n1136,
    n815,
    n776
  );


  and
  g1735
  (
    n1950,
    n896,
    n1396,
    n1235,
    n1488
  );


  xnor
  g1736
  (
    n1665,
    n1377,
    n1490,
    n1585,
    n1605
  );


  and
  g1737
  (
    n1705,
    n511,
    n524,
    n1267,
    n1286
  );


  and
  g1738
  (
    n1729,
    n544,
    n539,
    n575,
    n928
  );


  nand
  g1739
  (
    n1750,
    n1082,
    n770,
    n1402,
    n1074
  );


  or
  g1740
  (
    n1916,
    n519,
    n1225,
    n1253,
    n543
  );


  and
  g1741
  (
    n1919,
    n846,
    n745,
    n808,
    n1493
  );


  xor
  g1742
  (
    n1938,
    n1160,
    n845,
    n1560,
    n562
  );


  xnor
  g1743
  (
    KeyWire_0_3,
    n1349,
    n857,
    n538,
    n508
  );


  xnor
  g1744
  (
    n1706,
    n1443,
    n873,
    n775,
    n855
  );


  xnor
  g1745
  (
    n1927,
    n694,
    n1227,
    n1313,
    n676
  );


  xnor
  g1746
  (
    n1821,
    n553,
    n809,
    n1150,
    n1240
  );


  nor
  g1747
  (
    n1940,
    n1582,
    n534,
    n732,
    n1324
  );


  or
  g1748
  (
    n1685,
    n1510,
    n1375,
    n1464,
    n612
  );


  nand
  g1749
  (
    n1815,
    n992,
    n546,
    n532,
    n1419
  );


  or
  g1750
  (
    n1766,
    n519,
    n921,
    n1478,
    n737
  );


  nor
  g1751
  (
    n1900,
    n811,
    n1335,
    n561,
    n1118
  );


  xnor
  g1752
  (
    n1855,
    n1116,
    n1029,
    n723,
    n932
  );


  and
  g1753
  (
    n1727,
    n667,
    n834,
    n1208,
    n626
  );


  and
  g1754
  (
    n1803,
    n1169,
    n879,
    n1594,
    n847
  );


  or
  g1755
  (
    n1868,
    n818,
    n1385,
    n636,
    n1167
  );


  nor
  g1756
  (
    n1660,
    n559,
    n542,
    n1555,
    n541
  );


  xnor
  g1757
  (
    n1843,
    n1066,
    n1159,
    n772,
    n739
  );


  nand
  g1758
  (
    n1967,
    n1489,
    n1376,
    n1345,
    n1601
  );


  and
  g1759
  (
    n1765,
    n1032,
    n982,
    n854,
    n1083
  );


  xor
  g1760
  (
    n1913,
    n955,
    n511,
    n1162,
    n1392
  );


  xnor
  g1761
  (
    n1895,
    n633,
    n1564,
    n827,
    n1287
  );


  or
  g1762
  (
    n1824,
    n515,
    n938,
    n532,
    n1330
  );


  xor
  g1763
  (
    n1968,
    n998,
    n1323,
    n1334,
    n525
  );


  xor
  g1764
  (
    n1795,
    n736,
    n1174,
    n980,
    n744
  );


  or
  g1765
  (
    n1683,
    n793,
    n601,
    n1052,
    n1296
  );


  xnor
  g1766
  (
    n1953,
    n702,
    n1072,
    n537,
    n849
  );


  nand
  g1767
  (
    n1722,
    n514,
    n1164,
    n934,
    n1017
  );


  and
  g1768
  (
    n1835,
    n556,
    n547,
    n532,
    n1384
  );


  and
  g1769
  (
    n1673,
    n973,
    n510,
    n1130,
    n1355
  );


  nor
  g1770
  (
    n1937,
    n777,
    n1413,
    n1079,
    n1540
  );


  xor
  g1771
  (
    n1845,
    n1554,
    n591,
    n877,
    n1281
  );


  xor
  g1772
  (
    n1941,
    n1506,
    n765,
    n1314,
    n872
  );


  nor
  g1773
  (
    n1920,
    n537,
    n620,
    n1548,
    n1166
  );


  xnor
  g1774
  (
    n1905,
    n513,
    n1018,
    n520,
    n530
  );


  xor
  g1775
  (
    n1854,
    n1299,
    n1199,
    n518,
    n1541
  );


  and
  g1776
  (
    n1691,
    n958,
    n553,
    n1428,
    n1269
  );


  xnor
  g1777
  (
    n1798,
    n918,
    n833,
    n923,
    n1306
  );


  nor
  g1778
  (
    n1807,
    n1404,
    n509,
    n686,
    n669
  );


  nor
  g1779
  (
    n1875,
    n1587,
    n1243,
    n1329,
    n867
  );


  and
  g1780
  (
    n1774,
    n866,
    n1595,
    n594,
    n1171
  );


  xor
  g1781
  (
    n1658,
    n709,
    n1062,
    n1189,
    n1048
  );


  and
  g1782
  (
    n1870,
    n1061,
    n796,
    n791,
    n1317
  );


  nand
  g1783
  (
    n1800,
    n679,
    n842,
    n1031,
    n1120
  );


  nor
  g1784
  (
    n1965,
    n1512,
    n523,
    n1034,
    n707
  );


  xor
  g1785
  (
    n1888,
    n925,
    n1576,
    n1117,
    n670
  );


  and
  g1786
  (
    n1904,
    n742,
    n904,
    n698,
    n611
  );


  and
  g1787
  (
    n1692,
    n1366,
    n1476,
    n557,
    n1426
  );


  or
  g1788
  (
    n1737,
    n527,
    n1382,
    n541,
    n655
  );


  and
  g1789
  (
    n1955,
    n919,
    n643,
    n512,
    n905
  );


  nand
  g1790
  (
    n1851,
    n510,
    n1567,
    n999,
    n1259
  );


  nor
  g1791
  (
    n1695,
    n1338,
    n1124,
    n537,
    n1050
  );


  or
  g1792
  (
    n1971,
    n719,
    n881,
    n650,
    n1274
  );


  and
  g1793
  (
    n1966,
    n1057,
    n712,
    n1328,
    n555
  );


  nand
  g1794
  (
    n1863,
    n711,
    n1106,
    n738,
    n1075
  );


  xor
  g1795
  (
    n1898,
    n1519,
    n1346,
    n1063,
    n654
  );


  or
  g1796
  (
    KeyWire_0_25,
    n949,
    n1292,
    n961,
    n581
  );


  nor
  g1797
  (
    n1918,
    n521,
    n538,
    n577,
    n560
  );


  xor
  g1798
  (
    n1663,
    n1378,
    n1252,
    n786,
    n1504
  );


  xor
  g1799
  (
    n1834,
    n726,
    n1011,
    n908,
    n1581
  );


  xor
  g1800
  (
    n1700,
    n1430,
    n1316,
    n844,
    n1406
  );


  or
  g1801
  (
    n1702,
    n1134,
    n1264,
    n530,
    n1417
  );


  and
  g1802
  (
    n1707,
    n823,
    n662,
    n787,
    n1363
  );


  xor
  g1803
  (
    n1849,
    n1146,
    n536,
    n544,
    n985
  );


  or
  g1804
  (
    n1952,
    n1021,
    n657,
    n646,
    n1135
  );


  xor
  g1805
  (
    n1826,
    n911,
    n1215,
    n1423,
    n530
  );


  and
  g1806
  (
    n1713,
    n1364,
    n734,
    n1571,
    n1307
  );


  nand
  g1807
  (
    n1785,
    n969,
    n1230,
    n972,
    n1114
  );


  xor
  g1808
  (
    n1751,
    n945,
    n523,
    n589,
    n1144
  );


  nand
  g1809
  (
    n1902,
    n540,
    n596,
    n826,
    n836
  );


  xor
  g1810
  (
    n1792,
    n1498,
    n1586,
    n526,
    n1158
  );


  nand
  g1811
  (
    n1959,
    n1275,
    n1391,
    n558,
    n1268
  );


  or
  g1812
  (
    n1825,
    n1431,
    n525,
    n1265,
    n1468
  );


  nand
  g1813
  (
    n1749,
    n1449,
    n595,
    n1133,
    n1276
  );


  or
  g1814
  (
    n1693,
    n569,
    n1515,
    n562,
    n1260
  );


  and
  g1815
  (
    n1866,
    n1497,
    n798,
    n549,
    n1195
  );


  nand
  g1816
  (
    n1770,
    n986,
    n1483,
    n564,
    n1437
  );


  nor
  g1817
  (
    n1922,
    n1446,
    n790,
    n1533,
    n673
  );


  xor
  g1818
  (
    n1923,
    n584,
    n1418,
    n957,
    n940
  );


  xnor
  g1819
  (
    n1869,
    n931,
    n751,
    n566,
    n1054
  );


  nand
  g1820
  (
    n1933,
    n553,
    n579,
    n960,
    n556
  );


  nand
  g1821
  (
    n1802,
    n550,
    n947,
    n1453,
    n1538
  );


  or
  g1822
  (
    n1948,
    n548,
    n1495,
    n610,
    n1482
  );


  nor
  g1823
  (
    n1934,
    n1221,
    n1520,
    n524,
    n1348
  );


  xnor
  g1824
  (
    n1859,
    n608,
    n831,
    n1568,
    n521
  );


  xnor
  g1825
  (
    n1861,
    n523,
    n795,
    n521,
    n1109
  );


  xor
  g1826
  (
    n1725,
    n1342,
    n1583,
    n533,
    n1194
  );


  nand
  g1827
  (
    n1943,
    n1414,
    n629,
    n561,
    n1534
  );


  xor
  g1828
  (
    n1877,
    n536,
    n1294,
    n906,
    n512
  );


  xor
  g1829
  (
    n1761,
    n1457,
    n1122,
    n516,
    n560
  );


  xor
  g1830
  (
    n1767,
    n821,
    n548,
    n1094,
    n1180
  );


  xnor
  g1831
  (
    n1808,
    n1365,
    n1129,
    n755,
    n1042
  );


  or
  g1832
  (
    n1659,
    n1451,
    n563,
    n656,
    n683
  );


  nand
  g1833
  (
    n1818,
    n1236,
    n604,
    n651,
    n685
  );


  xor
  g1834
  (
    n1715,
    n1003,
    n1087,
    n788,
    n1362
  );


  xnor
  g1835
  (
    n1836,
    n554,
    n568,
    n536,
    n1546
  );


  xnor
  g1836
  (
    n1832,
    n645,
    n1140,
    n937,
    n1245
  );


  xor
  g1837
  (
    n1970,
    n693,
    n563,
    n658,
    n519
  );


  nor
  g1838
  (
    n1975,
    n1100,
    n761,
    n819,
    n538
  );


  nand
  g1839
  (
    n1928,
    n996,
    n1141,
    n1295,
    n1326
  );


  or
  g1840
  (
    n1848,
    n946,
    n642,
    n533,
    n1013
  );


  nor
  g1841
  (
    n1733,
    n1104,
    n853,
    n554,
    n648
  );


  nand
  g1842
  (
    n1931,
    n830,
    n987,
    n850,
    n1386
  );


  and
  g1843
  (
    n1764,
    n640,
    n603,
    n1038,
    n1320
  );


  and
  g1844
  (
    n1852,
    n1352,
    n1597,
    n1492,
    n1298
  );


  and
  g1845
  (
    n1921,
    n1152,
    n557,
    n1175,
    n1108
  );


  xor
  g1846
  (
    n1762,
    n824,
    n1509,
    n1350,
    n627
  );


  or
  g1847
  (
    n1759,
    n953,
    n871,
    n1545,
    n1373
  );


  or
  g1848
  (
    n1773,
    n660,
    n560,
    n568,
    n727
  );


  nor
  g1849
  (
    n1910,
    n740,
    n1070,
    n812,
    n1539
  );


  xor
  g1850
  (
    n1903,
    n784,
    n1304,
    n907,
    n916
  );


  xor
  g1851
  (
    n1917,
    n553,
    n1138,
    n1123,
    n1015
  );


  nand
  g1852
  (
    n1721,
    n1606,
    n1110,
    n728,
    n1336
  );


  xnor
  g1853
  (
    n1973,
    n902,
    n684,
    n1132,
    n547
  );


  nor
  g1854
  (
    n1748,
    n1575,
    n1250,
    n549,
    n1305
  );


  or
  g1855
  (
    n1694,
    n1161,
    n725,
    n548,
    n884
  );


  and
  g1856
  (
    n1897,
    n1603,
    n1309,
    n1602,
    n1405
  );


  xnor
  g1857
  (
    n1710,
    n979,
    n1389,
    n639,
    n599
  );


  nor
  g1858
  (
    n1939,
    n1579,
    n1368,
    n766,
    n1183
  );


  xnor
  g1859
  (
    n1899,
    n862,
    n659,
    n1283,
    n1257
  );


  and
  g1860
  (
    n1964,
    n859,
    n1422,
    n1524,
    n1058
  );


  xor
  g1861
  (
    n1771,
    n528,
    n1550,
    n841,
    n518
  );


  and
  g1862
  (
    n1894,
    n936,
    n522,
    n632,
    n1010
  );


  and
  g1863
  (
    n1846,
    n663,
    n1228,
    n1559,
    n1209
  );


  and
  g1864
  (
    n1677,
    n1190,
    n975,
    n1193,
    n964
  );


  nand
  g1865
  (
    n1744,
    n1244,
    n779,
    n509,
    n1485
  );


  nor
  g1866
  (
    n1739,
    n558,
    n950,
    n760,
    n517
  );


  nor
  g1867
  (
    n1687,
    n567,
    n895,
    n652,
    n528
  );


  nor
  g1868
  (
    n1889,
    n644,
    n1370,
    n529,
    n864
  );


  nor
  g1869
  (
    n1936,
    n578,
    n721,
    n814,
    n1444
  );


  nand
  g1870
  (
    n1883,
    n613,
    n983,
    n514,
    n974
  );


  nand
  g1871
  (
    n1701,
    n1356,
    n993,
    n1563,
    n1030
  );


  and
  g1872
  (
    n1671,
    n970,
    n580,
    n1247,
    n515
  );


  and
  g1873
  (
    n1734,
    n600,
    n1127,
    n568,
    n661
  );


  xor
  g1874
  (
    n1736,
    n952,
    n566,
    n1458,
    n924
  );


  xor
  g1875
  (
    n1688,
    n1600,
    n1481,
    n1380,
    n1056
  );


  nor
  g1876
  (
    n1708,
    n807,
    n668,
    n641,
    n1020
  );


  nand
  g1877
  (
    n1886,
    n542,
    n1115,
    n789,
    n851
  );


  xor
  g1878
  (
    n1781,
    n634,
    n556,
    n1077,
    n1300
  );


  nor
  g1879
  (
    n1951,
    n1060,
    n1119,
    n1387,
    n1420
  );


  nand
  g1880
  (
    n1755,
    n956,
    n1486,
    n535,
    n563
  );


  xnor
  g1881
  (
    n1969,
    n1599,
    n1421,
    n1084,
    n840
  );


  xor
  g1882
  (
    n1674,
    n1005,
    n649,
    n1318,
    n794
  );


  nor
  g1883
  (
    n1790,
    n1157,
    n1302,
    n1341,
    n511
  );


  and
  g1884
  (
    n1718,
    n561,
    n1608,
    n558,
    n1487
  );


  and
  g1885
  (
    n1812,
    n1475,
    n1040,
    n665,
    n1390
  );


  or
  g1886
  (
    n1657,
    n516,
    n1263,
    n551,
    n550
  );


  nor
  g1887
  (
    n1881,
    n690,
    n696,
    n1452,
    n1086
  );


  xor
  g1888
  (
    n1775,
    n1241,
    n1107,
    n967,
    n965
  );


  nand
  g1889
  (
    n1731,
    n1500,
    n562,
    n1203,
    n1179
  );


  xnor
  g1890
  (
    n1880,
    n531,
    n981,
    n701,
    n1112
  );


  nor
  g1891
  (
    n1840,
    n943,
    n512,
    n533,
    n1218
  );


  xnor
  g1892
  (
    n1789,
    n1569,
    n1081,
    n792,
    n1226
  );


  xnor
  g1893
  (
    n1844,
    n1432,
    n1234,
    n542,
    n705
  );


  xnor
  g1894
  (
    n1892,
    n687,
    n1176,
    n1022,
    n555
  );


  nor
  g1895
  (
    n1779,
    n692,
    n1089,
    n747,
    n1168
  );


  xnor
  g1896
  (
    n1672,
    n512,
    n540,
    n1577,
    n543
  );


  xor
  g1897
  (
    n1946,
    n681,
    n1424,
    n927,
    n1103
  );


  or
  g1898
  (
    n1822,
    n548,
    n1007,
    n1277,
    n743
  );


  or
  g1899
  (
    n1747,
    n1037,
    n677,
    n835,
    n552
  );


  nor
  g1900
  (
    n1763,
    n1197,
    n1198,
    n554,
    n1361
  );


  xnor
  g1901
  (
    n1974,
    n989,
    n1415,
    n962,
    n1454
  );


  nor
  g1902
  (
    n1772,
    n1111,
    n991,
    n1238,
    n522
  );


  and
  g1903
  (
    n1689,
    n1047,
    n563,
    n1466,
    n534
  );


  nand
  g1904
  (
    n1833,
    n1359,
    n1076,
    n1494,
    n1321
  );


  or
  g1905
  (
    n1837,
    n618,
    n733,
    n1016,
    n875
  );


  or
  g1906
  (
    n1786,
    n678,
    n1178,
    n1131,
    n557
  );


  nand
  g1907
  (
    n1756,
    n1580,
    n628,
    n1471,
    n1028
  );


  xnor
  g1908
  (
    n1976,
    n714,
    n718,
    n753,
    n861
  );


  xnor
  g1909
  (
    n1666,
    n532,
    n1012,
    n1149,
    n560
  );


  xor
  g1910
  (
    n1797,
    n566,
    n1491,
    n1289,
    n567
  );


  nand
  g1911
  (
    n1860,
    n1154,
    n1009,
    n1025,
    n1024
  );


  nand
  g1912
  (
    n1742,
    n1279,
    n511,
    n1394,
    n716
  );


  xnor
  g1913
  (
    n1801,
    n566,
    n870,
    n536,
    n1004
  );


  nand
  g1914
  (
    n1745,
    n731,
    n816,
    n1462,
    n1301
  );


  xnor
  g1915
  (
    n1684,
    n562,
    n567,
    n583,
    n559
  );


  xnor
  g1916
  (
    n1661,
    n528,
    n774,
    n1374,
    n1085
  );


  nor
  g1917
  (
    n1831,
    n920,
    n525,
    n1499,
    n520
  );


  xor
  g1918
  (
    n1839,
    n758,
    n555,
    n1528,
    n804
  );


  or
  g1919
  (
    n1932,
    n557,
    n529,
    n912,
    n531
  );


  xnor
  g1920
  (
    n1675,
    n856,
    n1059,
    n1358,
    n588
  );


  xor
  g1921
  (
    n1662,
    n1469,
    n1266,
    n519,
    n968
  );


  xor
  g1922
  (
    n1906,
    n1090,
    n781,
    n1508,
    n933
  );


  and
  g1923
  (
    n1828,
    n565,
    n741,
    n616,
    n555
  );


  xnor
  g1924
  (
    n1947,
    n1191,
    n1467,
    n1097,
    n514
  );


  nand
  g1925
  (
    n1697,
    n1565,
    n930,
    n565,
    n522
  );


  and
  g1926
  (
    n1714,
    n1073,
    n1173,
    n926,
    n1445
  );


  or
  g1927
  (
    n1810,
    n507,
    n863,
    n1472,
    n534
  );


  nor
  g1928
  (
    n1793,
    n990,
    n1285,
    n1340,
    n567
  );


  and
  g1929
  (
    n1885,
    n1566,
    n545,
    n1590,
    n825
  );


  xor
  g1930
  (
    n1962,
    n1023,
    n939,
    n1297,
    n1480
  );


  xnor
  g1931
  (
    n1796,
    n1398,
    n1044,
    n587,
    n585
  );


  nand
  g1932
  (
    n1717,
    n901,
    n1043,
    n547,
    n521
  );


  xor
  g1933
  (
    n1784,
    n868,
    n988,
    n1249,
    n508
  );


  xor
  g1934
  (
    n1850,
    n1549,
    n1562,
    n674,
    n1542
  );


  and
  g1935
  (
    n1776,
    n568,
    n782,
    n540,
    n1527
  );


  or
  g1936
  (
    n1819,
    n1553,
    n882,
    n544,
    n800
  );


  xnor
  g1937
  (
    KeyWire_0_13,
    n1053,
    n1217,
    n561,
    n1339
  );


  xor
  g1938
  (
    n1682,
    n922,
    n1232,
    n1511,
    n750
  );


  nand
  g1939
  (
    n1857,
    n508,
    n1322,
    n883,
    n624
  );


  xor
  g1940
  (
    n1972,
    n1098,
    n722,
    n538,
    n878
  );


  nor
  g1941
  (
    n1909,
    n1093,
    n1439,
    n1529,
    n843
  );


  or
  g1942
  (
    n1758,
    n1293,
    n771,
    n1441,
    n593
  );


  xnor
  g1943
  (
    n1924,
    n1537,
    n1229,
    n543,
    n523
  );


  xnor
  g1944
  (
    n1720,
    n1591,
    n527,
    n1170,
    n1440
  );


  xnor
  g1945
  (
    n1740,
    n522,
    n1551,
    n897,
    n773
  );


  nand
  g1946
  (
    n1667,
    n526,
    n1006,
    n529,
    n542
  );


  xor
  g1947
  (
    n1704,
    n537,
    n666,
    n515,
    n1584
  );


  buf
  g1948
  (
    n1978,
    n1656
  );


  not
  g1949
  (
    n1977,
    n1657
  );


  xor
  g1950
  (
    n1985,
    n1678,
    n1669,
    n1977,
    n1677
  );


  xor
  g1951
  (
    n1979,
    n1670,
    n1977,
    n1661,
    n1672
  );


  and
  g1952
  (
    n1984,
    n1665,
    n1662,
    n1977,
    n1978
  );


  and
  g1953
  (
    n1983,
    n1681,
    n1674,
    n1671,
    n1660
  );


  and
  g1954
  (
    n1986,
    n1666,
    n1978,
    n1667
  );


  and
  g1955
  (
    n1980,
    n1663,
    n1675,
    n1668,
    n1664
  );


  nand
  g1956
  (
    n1981,
    n1659,
    n1978,
    n1977,
    n1679
  );


  nand
  g1957
  (
    n1982,
    n1673,
    n1658,
    n1676,
    n1680
  );


  and
  g1958
  (
    n1988,
    n1694,
    n1983,
    n1692
  );


  nand
  g1959
  (
    n1989,
    n1693,
    n1684,
    n1683,
    n1682
  );


  xor
  g1960
  (
    n1991,
    n1979,
    n1981,
    n1691,
    n1688
  );


  nand
  g1961
  (
    n1987,
    n1686,
    n1687,
    n1689,
    n1695
  );


  nor
  g1962
  (
    n1990,
    n1982,
    n1685,
    n1980,
    n1690
  );


  buf
  g1963
  (
    n1992,
    n1697
  );


  not
  g1964
  (
    n1993,
    n1696
  );


  xor
  g1965
  (
    n1994,
    n1698,
    n1989,
    n1990,
    n1701
  );


  nand
  g1966
  (
    n1995,
    n1700,
    n1988,
    n1987,
    n1699
  );


  buf
  g1967
  (
    n1999,
    n1993
  );


  not
  g1968
  (
    KeyWire_0_24,
    n1995
  );


  buf
  g1969
  (
    n1996,
    n1994
  );


  buf
  g1970
  (
    n1998,
    n1992
  );


  nor
  g1971
  (
    n2007,
    n1731,
    n1707,
    n1730,
    n1727
  );


  or
  g1972
  (
    n2010,
    n1705,
    n1702,
    n1714,
    n1996
  );


  xor
  g1973
  (
    n2012,
    n1996,
    n1708,
    n1721,
    n1717
  );


  xor
  g1974
  (
    n2000,
    n1719,
    n1996,
    n1724,
    n1720
  );


  and
  g1975
  (
    n2002,
    n1709,
    n1736,
    n1997,
    n1745
  );


  or
  g1976
  (
    n2008,
    n1741,
    n1999,
    n1746,
    n1742
  );


  xor
  g1977
  (
    KeyWire_0_20,
    n1747,
    n1999,
    n1715,
    n1998
  );


  nand
  g1978
  (
    n2014,
    n1998,
    n1997,
    n1748
  );


  nand
  g1979
  (
    n2004,
    n1998,
    n1728,
    n1713,
    n1723
  );


  nand
  g1980
  (
    n2009,
    n1743,
    n1733,
    n1740,
    n1744
  );


  xor
  g1981
  (
    n2005,
    n1998,
    n1999,
    n1703,
    n1738
  );


  xnor
  g1982
  (
    n2001,
    n1725,
    n1711,
    n1996,
    n1704
  );


  xor
  g1983
  (
    n2011,
    n1732,
    n1718,
    n1749,
    n1710
  );


  or
  g1984
  (
    n2003,
    n1999,
    n1726,
    n1712,
    n1716
  );


  or
  g1985
  (
    n2013,
    n1722,
    n1997,
    n1729,
    n1706
  );


  xnor
  g1986
  (
    n2015,
    n1734,
    n1735,
    n1737,
    n1739
  );


  xnor
  g1987
  (
    n2016,
    n569,
    n570,
    n2014
  );


  nand
  g1988
  (
    n2018,
    n1754,
    n2016,
    n1752,
    n1753
  );


  nor
  g1989
  (
    n2017,
    n2016,
    n1755,
    n1750,
    n1751
  );


  xor
  g1990
  (
    n2019,
    n1759,
    n2017,
    n1760
  );


  xnor
  g1991
  (
    n2020,
    n1757,
    n1756,
    n1758,
    n2017
  );


  nor
  g1992
  (
    n2021,
    n1761,
    n2019,
    n1762
  );


  and
  g1993
  (
    n2023,
    n1991,
    n1986,
    n2021,
    n1984
  );


  nand
  g1994
  (
    n2022,
    n1991,
    n1991,
    n1985,
    n2021
  );


  buf
  g1995
  (
    n2024,
    n1764
  );


  buf
  g1996
  (
    n2025,
    n1765
  );


  xor
  g1997
  (
    n2026,
    n2022,
    n1763,
    n2023
  );


  not
  g1998
  (
    n2027,
    n2024
  );


  buf
  g1999
  (
    n2028,
    n2025
  );


  and
  g2000
  (
    n2029,
    n2028,
    n570,
    n2015
  );


  nor
  g2001
  (
    n2033,
    n1771,
    n1774,
    n1767,
    n1773
  );


  and
  g2002
  (
    n2031,
    n1772,
    n1776,
    n1775,
    n1768
  );


  xor
  g2003
  (
    KeyWire_0_11,
    n1770,
    n2029
  );


  xor
  g2004
  (
    n2032,
    n1777,
    n2029,
    n1766,
    n1769
  );


  not
  g2005
  (
    n2035,
    n1779
  );


  xor
  g2006
  (
    n2034,
    n2031,
    n1778,
    n2030
  );


  not
  g2007
  (
    n2036,
    n2034
  );


  not
  g2008
  (
    n2037,
    n2034
  );


  xor
  g2009
  (
    n2045,
    n2034,
    n2019,
    n2036,
    n2025
  );


  nand
  g2010
  (
    n2044,
    n2035,
    n2035,
    n2037,
    n2034
  );


  and
  g2011
  (
    n2038,
    n2035,
    n2018,
    n2020,
    n2037
  );


  xnor
  g2012
  (
    n2043,
    n2018,
    n2037,
    n2020
  );


  nand
  g2013
  (
    n2040,
    n571,
    n2020,
    n2036
  );


  or
  g2014
  (
    n2041,
    n2018,
    n571,
    n2035,
    n2017
  );


  xor
  g2015
  (
    n2042,
    n572,
    n571,
    n2037
  );


  xnor
  g2016
  (
    n2039,
    n1780,
    n2018,
    n2036,
    n2017
  );


  and
  g2017
  (
    n2051,
    n1615,
    n2041,
    n2038,
    n1648
  );


  xnor
  g2018
  (
    n2047,
    n1635,
    n1790,
    n1805,
    n1789
  );


  xor
  g2019
  (
    n2048,
    n1636,
    n1785,
    n1614,
    n1618
  );


  xnor
  g2020
  (
    n2053,
    n2044,
    n1621,
    n2039,
    n1620
  );


  nand
  g2021
  (
    n2065,
    n1619,
    n1783,
    n1787,
    n573
  );


  xor
  g2022
  (
    n2077,
    n1613,
    n2032,
    n1627,
    n2038
  );


  nor
  g2023
  (
    n2057,
    n2042,
    n2025,
    n1807,
    n1788
  );


  or
  g2024
  (
    n2059,
    n1804,
    n1991,
    n2040,
    n2044
  );


  or
  g2025
  (
    n2074,
    n1611,
    n1610,
    n2040,
    n2033
  );


  xnor
  g2026
  (
    n2072,
    n2044,
    n2038,
    n2043,
    n1646
  );


  nor
  g2027
  (
    n2071,
    n1653,
    n2039,
    n2033,
    n2041
  );


  xor
  g2028
  (
    n2062,
    n1617,
    n1643,
    n1630,
    n28
  );


  and
  g2029
  (
    n2070,
    n2043,
    n1622,
    n572,
    n1639
  );


  xnor
  g2030
  (
    n2054,
    n1647,
    n1651,
    n1800,
    n2039
  );


  nand
  g2031
  (
    n2068,
    n1786,
    n2026,
    n1644,
    n1791
  );


  xor
  g2032
  (
    n2061,
    n2045,
    n1801,
    n2039,
    n1637
  );


  nand
  g2033
  (
    n2058,
    n1625,
    n2042,
    n1642,
    n1624
  );


  nor
  g2034
  (
    n2075,
    n1628,
    n1797,
    n1649,
    n2045
  );


  xnor
  g2035
  (
    n2060,
    n1812,
    n1794,
    n2041,
    n28
  );


  and
  g2036
  (
    n2076,
    n573,
    n1798,
    n1811,
    n1631
  );


  nand
  g2037
  (
    n2069,
    n1640,
    n1633,
    n1655,
    n573
  );


  nor
  g2038
  (
    n2064,
    n1799,
    n1616,
    n2044,
    n1782
  );


  nand
  g2039
  (
    n2050,
    n2026,
    n1650,
    n573,
    n1641
  );


  xor
  g2040
  (
    n2055,
    n2038,
    n1792,
    n1796,
    n2045
  );


  xnor
  g2041
  (
    n2056,
    n2043,
    n1612,
    n1793,
    n2041
  );


  nor
  g2042
  (
    n2052,
    n1634,
    n2045,
    n1654,
    n1806
  );


  nand
  g2043
  (
    n2049,
    n572,
    n2040,
    n2042,
    n1795
  );


  xnor
  g2044
  (
    KeyWire_0_0,
    n1784,
    n1781,
    n1632,
    n2042
  );


  xor
  g2045
  (
    n2067,
    n1629,
    n1652,
    n1802,
    n1609
  );


  nand
  g2046
  (
    n2063,
    n2040,
    n1626,
    n1803,
    n572
  );


  nand
  g2047
  (
    n2046,
    n1623,
    n2043,
    n1808,
    n2025
  );


  or
  g2048
  (
    n2066,
    n1810,
    n1645,
    n1809,
    n1638
  );


  or
  g2049
  (
    n2127,
    n1820,
    n1953,
    n1822,
    n2061
  );


  xor
  g2050
  (
    n2108,
    n2071,
    n1962,
    n1951,
    n1824
  );


  or
  g2051
  (
    n2114,
    n1894,
    n1845,
    n1835,
    n2075
  );


  xnor
  g2052
  (
    n2117,
    n1898,
    n1908,
    n1913,
    n1909
  );


  and
  g2053
  (
    n2110,
    n1860,
    n1968,
    n2064,
    n2076
  );


  xor
  g2054
  (
    n2132,
    n1872,
    n1931,
    n1922,
    n2071
  );


  or
  g2055
  (
    n2095,
    n2058,
    n2073,
    n1846,
    n2077
  );


  or
  g2056
  (
    n2083,
    n1959,
    n1926,
    n1937,
    n2068
  );


  xor
  g2057
  (
    n2100,
    n1904,
    n1892,
    n1832,
    n1955
  );


  or
  g2058
  (
    n2093,
    n2066,
    n2072,
    n1932,
    n1842
  );


  xnor
  g2059
  (
    n2097,
    n2026,
    n1879,
    n1945,
    n1973
  );


  nand
  g2060
  (
    n2099,
    n1827,
    n2074,
    n1944,
    n1890
  );


  nor
  g2061
  (
    n2106,
    n1972,
    n1867,
    n2077,
    n1865
  );


  xnor
  g2062
  (
    n2078,
    n1928,
    n2074,
    n1923,
    n1837
  );


  nor
  g2063
  (
    n2125,
    n1881,
    n2062,
    n1821,
    n2072
  );


  xor
  g2064
  (
    n2090,
    n1957,
    n2048,
    n1875,
    n1963
  );


  nor
  g2065
  (
    n2092,
    n1940,
    n1933,
    n1954,
    n1814
  );


  xnor
  g2066
  (
    n2124,
    n1813,
    n2071,
    n2077,
    n1900
  );


  nor
  g2067
  (
    n2098,
    n1838,
    n2053,
    n1884,
    n1943
  );


  nor
  g2068
  (
    n2123,
    n1917,
    n1836,
    n1895,
    n1960
  );


  xor
  g2069
  (
    n2088,
    n2077,
    n2056,
    n1966,
    n2072
  );


  xnor
  g2070
  (
    n2111,
    n1942,
    n1901,
    n1914,
    n1903
  );


  xnor
  g2071
  (
    n2126,
    n1885,
    n2046,
    n1877,
    n2075
  );


  xnor
  g2072
  (
    n2107,
    n1907,
    n2070,
    n1887
  );


  and
  g2073
  (
    n2121,
    n2069,
    n1878,
    n1965,
    n1852
  );


  nand
  g2074
  (
    n2131,
    n1869,
    n1870,
    n2065,
    n1839
  );


  nor
  g2075
  (
    n2079,
    n1906,
    n1947,
    n2069,
    n1847
  );


  nand
  g2076
  (
    n2091,
    n1833,
    n1850,
    n1936,
    n1823
  );


  or
  g2077
  (
    n2089,
    n2072,
    n1844,
    n2073,
    n2074
  );


  and
  g2078
  (
    n2128,
    n1974,
    n1934,
    n1848,
    n1863
  );


  xnor
  g2079
  (
    n2096,
    n1916,
    n1902,
    n1918,
    n1915
  );


  or
  g2080
  (
    n2120,
    n2063,
    n1817,
    n1896,
    n1964
  );


  and
  g2081
  (
    n2101,
    n1899,
    n1828,
    n1882,
    n1946
  );


  xor
  g2082
  (
    n2119,
    n1950,
    n2073,
    n1876,
    n1920
  );


  xnor
  g2083
  (
    n2105,
    n1970,
    n1949,
    n2059,
    n1929
  );


  nor
  g2084
  (
    n2080,
    n2075,
    n1841,
    n1834,
    n2060
  );


  and
  g2085
  (
    n2129,
    n1921,
    n1969,
    n1905,
    n2049
  );


  nand
  g2086
  (
    n2081,
    n1961,
    n1831,
    n1911,
    n1866
  );


  or
  g2087
  (
    n2084,
    n2067,
    n2054,
    n2026,
    n2050
  );


  xnor
  g2088
  (
    n2112,
    n1897,
    n2073,
    n1854,
    n1888
  );


  nor
  g2089
  (
    n2103,
    n1829,
    n1971,
    n1840,
    n1889
  );


  xnor
  g2090
  (
    n2113,
    n1912,
    n1868,
    n1830,
    n1880
  );


  or
  g2091
  (
    n2118,
    n1891,
    n1956,
    n2047,
    n1855
  );


  nand
  g2092
  (
    n2086,
    n1818,
    n1843,
    n1938,
    n1952
  );


  and
  g2093
  (
    n2082,
    n2057,
    n1859,
    n1927,
    n1819
  );


  xor
  g2094
  (
    n2085,
    n1886,
    n1883,
    n1871,
    n1967
  );


  or
  g2095
  (
    n2122,
    n2055,
    n1919,
    n1910,
    n2076
  );


  or
  g2096
  (
    n2104,
    n1815,
    n1826,
    n1941,
    n1935
  );


  and
  g2097
  (
    n2130,
    n1825,
    n1861,
    n1856,
    n1930
  );


  and
  g2098
  (
    n2094,
    n1853,
    n2075,
    n1851,
    n2052
  );


  and
  g2099
  (
    n2116,
    n1858,
    n1939,
    n2076,
    n2051
  );


  nand
  g2100
  (
    n2102,
    n1873,
    n1975,
    n1864,
    n1893
  );


  nand
  g2101
  (
    n2109,
    n1849,
    n2076,
    n1924,
    n1958
  );


  or
  g2102
  (
    n2087,
    n2071,
    n1925,
    n1948,
    n2074
  );


  nor
  g2103
  (
    n2115,
    n1857,
    n1816,
    n1862,
    n1874
  );


  buf
  g2104
  (
    n2134,
    n2078
  );


  not
  g2105
  (
    n2133,
    n2079
  );


  nor
  g2106
  (
    n2138,
    n2082,
    n2093,
    n2133,
    n2091
  );


  xor
  g2107
  (
    n2142,
    n2094,
    n2083,
    n2081,
    n2103
  );


  nand
  g2108
  (
    n2140,
    n2133,
    n2134,
    n2097,
    n2080
  );


  nor
  g2109
  (
    n2135,
    n2134,
    n2089,
    n2098,
    n2086
  );


  and
  g2110
  (
    n2137,
    n2133,
    n2101,
    n2085,
    n2088
  );


  and
  g2111
  (
    n2141,
    n2133,
    n2084,
    n2096,
    n2134
  );


  xor
  g2112
  (
    n2136,
    n2092,
    n2095,
    n2102,
    n2090
  );


  xor
  g2113
  (
    n2139,
    n2087,
    n2100,
    n2134,
    n2099
  );


  nor
  g2114
  (
    n2147,
    n2135,
    n2105,
    n2110,
    n2140
  );


  and
  g2115
  (
    n2146,
    n2138,
    n2108,
    n2142
  );


  and
  g2116
  (
    n2145,
    n2142,
    n2139,
    n2111,
    n2136
  );


  and
  g2117
  (
    n2143,
    n2142,
    n2107,
    n2137,
    n2109
  );


  xor
  g2118
  (
    n2144,
    n2112,
    n2106,
    n2104,
    n2141
  );


  buf
  g2119
  (
    n2148,
    n2143
  );


  not
  g2120
  (
    n2149,
    n2143
  );


  and
  g2121
  (
    n2154,
    n2115,
    n2126,
    n2120,
    n2148
  );


  or
  g2122
  (
    n2156,
    n2116,
    n2118,
    n2145,
    n2123
  );


  nand
  g2123
  (
    n2153,
    n2121,
    n2148,
    n2122,
    n2149
  );


  nand
  g2124
  (
    n2151,
    n2148,
    n2144,
    n2125,
    n2149
  );


  nor
  g2125
  (
    n2157,
    n2148,
    n2114,
    n2149,
    n2145
  );


  xnor
  g2126
  (
    n2150,
    n2113,
    n2144
  );


  nor
  g2127
  (
    n2155,
    n2124,
    n2117,
    n2127,
    n2149
  );


  nand
  g2128
  (
    n2152,
    n2128,
    n2119,
    n2145
  );


  not
  g2129
  (
    n2158,
    n2150
  );


  nor
  g2130
  (
    n2159,
    n2152,
    n2151,
    n1976,
    n2158
  );


  nand
  g2131
  (
    n2162,
    n2151,
    n2158,
    n2152
  );


  and
  g2132
  (
    n2161,
    n2158,
    n2150,
    n2151,
    n2152
  );


  nor
  g2133
  (
    n2160,
    n2150,
    n2150,
    n2151,
    n2152
  );


  xnor
  g2134
  (
    n2174,
    n2157,
    n2146,
    n2154
  );


  xor
  g2135
  (
    n2163,
    n2160,
    n2132,
    n2155
  );


  xnor
  g2136
  (
    n2170,
    n2161,
    n2154,
    n2129,
    n2147
  );


  nand
  g2137
  (
    n2169,
    n2160,
    n2157,
    n2162,
    n2153
  );


  and
  g2138
  (
    KeyWire_0_26,
    n2160,
    n2159,
    n2153,
    n2147
  );


  nor
  g2139
  (
    n2172,
    n2154,
    n2147,
    n2160,
    n2162
  );


  nor
  g2140
  (
    n2164,
    n2146,
    n2153,
    n2162,
    n2156
  );


  xnor
  g2141
  (
    n2173,
    n2161,
    n2153,
    n2159,
    n2155
  );


  nand
  g2142
  (
    n2171,
    n2146,
    n2155,
    n2156,
    n2159
  );


  nor
  g2143
  (
    n2166,
    n2131,
    n2159,
    n2157,
    n2130
  );


  or
  g2144
  (
    n2167,
    n2157,
    n2156,
    n2161
  );


  or
  g2145
  (
    n2168,
    n2161,
    n2162,
    n2147,
    n2146
  );


  xor
  g2146
  (
    n2176,
    n2167,
    n2168,
    n2171,
    n2170
  );


  and
  g2147
  (
    n2175,
    n2166,
    n2169,
    n2165,
    n2173
  );


  xor
  g2148
  (
    n2177,
    n2163,
    n2174,
    n2164,
    n2172
  );


  xnor
  KeyGate_0_0
  (
    n2073,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1076,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n298,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1816,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n120,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n356,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n79,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n258,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n662,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1205,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n962,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n2030,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n307,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1777,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n342,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1723,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1312,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n938,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n316,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1783,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n2006,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n836,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n472,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1607,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1997,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1879,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n2165,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1333,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1562,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n228,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n423,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n610,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

