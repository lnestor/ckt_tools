

module Stat_100_65
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n90,
  n122,
  n125,
  n128,
  n131,
  n108,
  n102,
  n120,
  n105,
  n130,
  n115,
  n112,
  n121,
  n107,
  n117,
  n114,
  n113,
  n126,
  n119,
  n124,
  n111,
  n106,
  n123,
  n127,
  n104,
  n118,
  n129,
  n132,
  n109,
  n110,
  n116,
  n103,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n90;
  output n122;
  output n125;
  output n128;
  output n131;
  output n108;
  output n102;
  output n120;
  output n105;
  output n130;
  output n115;
  output n112;
  output n121;
  output n107;
  output n117;
  output n114;
  output n113;
  output n126;
  output n119;
  output n124;
  output n111;
  output n106;
  output n123;
  output n127;
  output n104;
  output n118;
  output n129;
  output n132;
  output n109;
  output n110;
  output n116;
  output n103;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n40,
    n25
  );


  not
  g1
  (
    n34,
    n23
  );


  buf
  g2
  (
    n41,
    n1
  );


  buf
  g3
  (
    KeyWire_0_56,
    n6
  );


  buf
  g4
  (
    n38,
    n19
  );


  buf
  g5
  (
    KeyWire_0_28,
    n13
  );


  buf
  g6
  (
    KeyWire_0_32,
    n31
  );


  buf
  g7
  (
    n37,
    n30
  );


  not
  g8
  (
    KeyWire_0_29,
    n21
  );


  buf
  g9
  (
    n33,
    n8
  );


  not
  g10
  (
    KeyWire_0_44,
    n9
  );


  not
  g11
  (
    n45,
    n4
  );


  not
  g12
  (
    KeyWire_0_4,
    n20
  );


  buf
  g13
  (
    KeyWire_0_47,
    n7
  );


  and
  g14
  (
    KeyWire_0_50,
    n26,
    n22
  );


  nor
  g15
  (
    KeyWire_0_63,
    n18,
    n32,
    n3,
    n24
  );


  and
  g16
  (
    n49,
    n11,
    n16,
    n29,
    n10
  );


  nand
  g17
  (
    KeyWire_0_6,
    n28,
    n27,
    n15,
    n17
  );


  xnor
  g18
  (
    n47,
    n14,
    n2,
    n12,
    n5
  );


  not
  g19
  (
    n58,
    n34
  );


  not
  g20
  (
    n81,
    n44
  );


  buf
  g21
  (
    KeyWire_0_37,
    n42
  );


  buf
  g22
  (
    KeyWire_0_3,
    n41
  );


  not
  g23
  (
    KeyWire_0_22,
    n39
  );


  not
  g24
  (
    n76,
    n42
  );


  not
  g25
  (
    KeyWire_0_13,
    n46
  );


  buf
  g26
  (
    KeyWire_0_35,
    n48
  );


  not
  g27
  (
    KeyWire_0_25,
    n44
  );


  buf
  g28
  (
    n66,
    n44
  );


  not
  g29
  (
    KeyWire_0_51,
    n45
  );


  buf
  g30
  (
    KeyWire_0_55,
    n36
  );


  not
  g31
  (
    KeyWire_0_36,
    n33
  );


  not
  g32
  (
    KeyWire_0_59,
    n36
  );


  buf
  g33
  (
    n71,
    n39
  );


  not
  g34
  (
    KeyWire_0_33,
    n40
  );


  buf
  g35
  (
    KeyWire_0_62,
    n46
  );


  buf
  g36
  (
    KeyWire_0_26,
    n47
  );


  not
  g37
  (
    n63,
    n40
  );


  buf
  g38
  (
    n78,
    n36
  );


  buf
  g39
  (
    KeyWire_0_18,
    n34
  );


  buf
  g40
  (
    n55,
    n37
  );


  not
  g41
  (
    KeyWire_0_10,
    n37
  );


  not
  g42
  (
    KeyWire_0_40,
    n47
  );


  not
  g43
  (
    n77,
    n35
  );


  buf
  g44
  (
    KeyWire_0_0,
    n38
  );


  not
  g45
  (
    KeyWire_0_20,
    n43
  );


  not
  g46
  (
    KeyWire_0_11,
    n38
  );


  buf
  g47
  (
    KeyWire_0_7,
    n42
  );


  buf
  g48
  (
    n82,
    n45
  );


  buf
  g49
  (
    KeyWire_0_45,
    n33
  );


  not
  g50
  (
    KeyWire_0_1,
    n34
  );


  not
  g51
  (
    n59,
    n38
  );


  not
  g52
  (
    n60,
    n33
  );


  nand
  g53
  (
    KeyWire_0_53,
    n45,
    n47,
    n41
  );


  xor
  g54
  (
    KeyWire_0_60,
    n40,
    n35,
    n37,
    n39
  );


  and
  g55
  (
    KeyWire_0_31,
    n35,
    n46,
    n43
  );


  not
  g56
  (
    KeyWire_0_57,
    n54
  );


  buf
  g57
  (
    n90,
    n53
  );


  nand
  g58
  (
    KeyWire_0_38,
    n52,
    n53
  );


  buf
  g59
  (
    KeyWire_0_48,
    n91
  );


  not
  g60
  (
    n93,
    n90
  );


  or
  g61
  (
    n98,
    n57,
    n54
  );


  and
  g62
  (
    KeyWire_0_49,
    n51,
    n93,
    n55,
    n48
  );


  xnor
  g63
  (
    KeyWire_0_41,
    n92,
    n57,
    n55,
    n54
  );


  and
  g64
  (
    n97,
    n49,
    n56,
    n50,
    n57
  );


  nor
  g65
  (
    KeyWire_0_16,
    n92,
    n51,
    n50,
    n55
  );


  xor
  g66
  (
    n95,
    n49,
    n49,
    n51,
    n50
  );


  xor
  g67
  (
    KeyWire_0_61,
    n93,
    n92,
    n56
  );


  xor
  g68
  (
    KeyWire_0_54,
    n56,
    n93,
    n48
  );


  nand
  g69
  (
    KeyWire_0_19,
    n87,
    n71,
    n97,
    n72
  );


  or
  g70
  (
    KeyWire_0_12,
    n100,
    n83,
    n68,
    n96
  );


  xnor
  g71
  (
    n123,
    n58,
    n100,
    n67,
    n86
  );


  nor
  g72
  (
    KeyWire_0_46,
    n95,
    n100,
    n66
  );


  nand
  g73
  (
    KeyWire_0_9,
    n88,
    n84,
    n85,
    n74
  );


  and
  g74
  (
    KeyWire_0_43,
    n98,
    n63,
    n101,
    n69
  );


  or
  g75
  (
    KeyWire_0_24,
    n77,
    n71,
    n64,
    n62
  );


  and
  g76
  (
    KeyWire_0_42,
    n83,
    n65,
    n99,
    n95
  );


  xor
  g77
  (
    KeyWire_0_5,
    n72,
    n96,
    n95,
    n73
  );


  nor
  g78
  (
    n131,
    n80,
    n97,
    n70,
    n87
  );


  xor
  g79
  (
    KeyWire_0_23,
    n101,
    n82,
    n86,
    n68
  );


  nor
  g80
  (
    n116,
    n77,
    n67,
    n78,
    n85
  );


  nor
  g81
  (
    n104,
    n98,
    n97,
    n74,
    n76
  );


  xnor
  g82
  (
    KeyWire_0_58,
    n86,
    n99,
    n59,
    n79
  );


  or
  g83
  (
    KeyWire_0_27,
    n58,
    n58,
    n59,
    n88
  );


  or
  g84
  (
    KeyWire_0_52,
    n59,
    n74,
    n72,
    n65
  );


  nand
  g85
  (
    KeyWire_0_17,
    n61,
    n94,
    n80,
    n75
  );


  and
  g86
  (
    KeyWire_0_14,
    n71,
    n69,
    n65,
    n79
  );


  nor
  g87
  (
    n105,
    n94,
    n95,
    n82,
    n84
  );


  and
  g88
  (
    KeyWire_0_2,
    n96,
    n94,
    n63,
    n87
  );


  xor
  g89
  (
    n119,
    n99,
    n61,
    n62,
    n81
  );


  xor
  g90
  (
    KeyWire_0_21,
    n83,
    n78,
    n98,
    n77
  );


  xnor
  g91
  (
    n127,
    n73,
    n78,
    n64,
    n70
  );


  xor
  g92
  (
    KeyWire_0_8,
    n99,
    n76,
    n96,
    n88
  );


  nor
  g93
  (
    KeyWire_0_30,
    n84,
    n70,
    n101,
    n80
  );


  or
  g94
  (
    n118,
    n60,
    n68,
    n81
  );


  xnor
  g95
  (
    KeyWire_0_39,
    n62,
    n75,
    n97,
    n82
  );


  xor
  g96
  (
    KeyWire_0_15,
    n75,
    n67,
    n63,
    n79
  );


  or
  g97
  (
    KeyWire_0_34,
    n73,
    n66,
    n76,
    n64
  );


  xnor
  g98
  (
    n124,
    n85,
    n61,
    n101,
    n69
  );


  xor
  g99
  (
    n120,
    n100,
    n60,
    n98
  );


  xor
  KeyGate_0_0
  (
    n69,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n61,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n106,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n52,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n35,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n117,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n43,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n54,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n114,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n121,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n73,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n70,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n132,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n62,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n103,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n110,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n99,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n112,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n88,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n109,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n75,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n102,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n87,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n125,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n107,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n56,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n67,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n111,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n46,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n51,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n108,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n65,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n50,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n84,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n129,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n64,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n57,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n85,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n91,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n122,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n53,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n100,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n130,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n128,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n42,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n80,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n115,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n44,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n92,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n94,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n39,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n68,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n126,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n72,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n96,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n83,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n36,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n89,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n113,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n86,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n79,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n101,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n74,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n48,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

