

module Stat_100_44
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n113,
  n114,
  n123,
  n105,
  n101,
  n122,
  n111,
  n115,
  n119,
  n110,
  n131,
  n103,
  n107,
  n109,
  n129,
  n116,
  n106,
  n128,
  n132,
  n130,
  n125,
  n120,
  n117,
  n118,
  n126,
  n127,
  n104,
  n121,
  n108,
  n102,
  n124
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n112;output n113;output n114;output n123;output n105;output n101;output n122;output n111;output n115;output n119;output n110;output n131;output n103;output n107;output n109;output n129;output n116;output n106;output n128;output n132;output n130;output n125;output n120;output n117;output n118;output n126;output n127;output n104;output n121;output n108;output n102;output n124;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    KeyWire_0_58,
    n19
  );


  buf
  g1
  (
    n88,
    n21
  );


  not
  g2
  (
    KeyWire_0_18,
    n22
  );


  not
  g3
  (
    KeyWire_0_62,
    n18
  );


  buf
  g4
  (
    KeyWire_0_3,
    n31
  );


  buf
  g5
  (
    KeyWire_0_48,
    n6
  );


  not
  g6
  (
    KeyWire_0_23,
    n1
  );


  not
  g7
  (
    n72,
    n25
  );


  not
  g8
  (
    KeyWire_0_56,
    n8
  );


  buf
  g9
  (
    n70,
    n28
  );


  buf
  g10
  (
    KeyWire_0_12,
    n26
  );


  not
  g11
  (
    KeyWire_0_1,
    n32
  );


  buf
  g12
  (
    n37,
    n20
  );


  not
  g13
  (
    KeyWire_0_13,
    n27
  );


  buf
  g14
  (
    n84,
    n23
  );


  not
  g15
  (
    KeyWire_0_27,
    n15
  );


  not
  g16
  (
    n50,
    n13
  );


  not
  g17
  (
    n49,
    n27
  );


  buf
  g18
  (
    KeyWire_0_6,
    n3
  );


  not
  g19
  (
    KeyWire_0_32,
    n29
  );


  buf
  g20
  (
    KeyWire_0_28,
    n11
  );


  not
  g21
  (
    n34,
    n29
  );


  buf
  g22
  (
    KeyWire_0_30,
    n14
  );


  not
  g23
  (
    n52,
    n4
  );


  not
  g24
  (
    n38,
    n27
  );


  buf
  g25
  (
    n68,
    n23
  );


  not
  g26
  (
    n85,
    n30
  );


  not
  g27
  (
    n73,
    n25
  );


  buf
  g28
  (
    KeyWire_0_55,
    n24
  );


  not
  g29
  (
    n55,
    n5
  );


  buf
  g30
  (
    KeyWire_0_8,
    n16
  );


  not
  g31
  (
    KeyWire_0_21,
    n28
  );


  not
  g32
  (
    KeyWire_0_9,
    n21
  );


  buf
  g33
  (
    n66,
    n9
  );


  buf
  g34
  (
    n76,
    n17
  );


  not
  g35
  (
    n56,
    n29
  );


  buf
  g36
  (
    KeyWire_0_16,
    n21
  );


  buf
  g37
  (
    KeyWire_0_54,
    n32
  );


  not
  g38
  (
    KeyWire_0_49,
    n31
  );


  buf
  g39
  (
    KeyWire_0_34,
    n26
  );


  buf
  g40
  (
    n58,
    n7
  );


  not
  g41
  (
    n57,
    n24
  );


  not
  g42
  (
    KeyWire_0_14,
    n10
  );


  buf
  g43
  (
    KeyWire_0_39,
    n30
  );


  buf
  g44
  (
    KeyWire_0_26,
    n26
  );


  buf
  g45
  (
    n54,
    n31
  );


  buf
  g46
  (
    KeyWire_0_2,
    n12
  );


  buf
  g47
  (
    n64,
    n23
  );


  buf
  g48
  (
    KeyWire_0_41,
    n30
  );


  buf
  g49
  (
    KeyWire_0_51,
    n25
  );


  buf
  g50
  (
    KeyWire_0_53,
    n22
  );


  buf
  g51
  (
    KeyWire_0_22,
    n24
  );


  buf
  g52
  (
    KeyWire_0_25,
    n22
  );


  buf
  g53
  (
    KeyWire_0_20,
    n28
  );


  buf
  g54
  (
    KeyWire_0_7,
    n32
  );


  buf
  g55
  (
    KeyWire_0_40,
    n2
  );


  buf
  g56
  (
    KeyWire_0_43,
    n38
  );


  not
  g57
  (
    KeyWire_0_10,
    n36
  );


  buf
  g58
  (
    n89,
    n34
  );


  and
  g59
  (
    KeyWire_0_47,
    n33,
    n35,
    n37
  );


  not
  g60
  (
    n95,
    n91
  );


  buf
  g61
  (
    KeyWire_0_63,
    n90
  );


  buf
  g62
  (
    KeyWire_0_17,
    n92
  );


  buf
  g63
  (
    KeyWire_0_0,
    n92
  );


  not
  g64
  (
    n97,
    n92
  );


  not
  g65
  (
    KeyWire_0_45,
    n91
  );


  not
  g66
  (
    n94,
    n91
  );


  buf
  g67
  (
    KeyWire_0_15,
    n89
  );


  xnor
  g68
  (
    n127,
    n98,
    n75,
    n97,
    n54
  );


  xor
  g69
  (
    KeyWire_0_11,
    n69,
    n56,
    n62,
    n85
  );


  or
  g70
  (
    n126,
    n88,
    n76,
    n63,
    n68
  );


  and
  g71
  (
    KeyWire_0_33,
    n100,
    n96,
    n45,
    n93
  );


  xnor
  g72
  (
    KeyWire_0_24,
    n74,
    n51,
    n52,
    n76
  );


  and
  g73
  (
    KeyWire_0_42,
    n84,
    n99,
    n66
  );


  xnor
  g74
  (
    KeyWire_0_60,
    n82,
    n44,
    n86,
    n88
  );


  and
  g75
  (
    n114,
    n96,
    n98,
    n75,
    n70
  );


  xor
  g76
  (
    KeyWire_0_50,
    n81,
    n53,
    n66,
    n97
  );


  nand
  g77
  (
    KeyWire_0_36,
    n71,
    n73,
    n79
  );


  and
  g78
  (
    n123,
    n79,
    n72,
    n88
  );


  nand
  g79
  (
    n124,
    n43,
    n71,
    n95,
    n85
  );


  xnor
  g80
  (
    KeyWire_0_59,
    n100,
    n81,
    n60,
    n94
  );


  and
  g81
  (
    KeyWire_0_19,
    n87,
    n66,
    n42,
    n86
  );


  nand
  g82
  (
    KeyWire_0_35,
    n93,
    n69,
    n94,
    n77
  );


  xnor
  g83
  (
    n111,
    n76,
    n67,
    n70,
    n80
  );


  xnor
  g84
  (
    KeyWire_0_31,
    n83,
    n82,
    n95,
    n77
  );


  xnor
  g85
  (
    KeyWire_0_4,
    n99,
    n94,
    n82,
    n65
  );


  or
  g86
  (
    KeyWire_0_61,
    n98,
    n79,
    n49,
    n68
  );


  xnor
  g87
  (
    KeyWire_0_52,
    n80,
    n50,
    n93,
    n68
  );


  nand
  g88
  (
    KeyWire_0_5,
    n78,
    n99,
    n95,
    n41
  );


  or
  g89
  (
    KeyWire_0_46,
    n98,
    n78,
    n61,
    n100
  );


  nand
  g90
  (
    KeyWire_0_37,
    n80,
    n40,
    n94,
    n78
  );


  or
  g91
  (
    KeyWire_0_44,
    n59,
    n48,
    n97,
    n58
  );


  nand
  g92
  (
    n105,
    n86,
    n46,
    n84,
    n81
  );


  xnor
  g93
  (
    KeyWire_0_29,
    n97,
    n67,
    n39,
    n64
  );


  xor
  g94
  (
    KeyWire_0_57,
    n95,
    n75,
    n47,
    n70
  );


  and
  g95
  (
    n120,
    n57,
    n87,
    n73,
    n96
  );


  or
  g96
  (
    n130,
    n55,
    n69,
    n87,
    n100
  );


  nand
  g97
  (
    KeyWire_0_38,
    n74,
    n85,
    n84,
    n96
  );


  nand
  g98
  (
    n106,
    n93,
    n67,
    n77,
    n74
  );


  or
  g99
  (
    n102,
    n71,
    n83,
    n72
  );


  xor
  KeyGate_0_0
  (
    n100,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n78,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n47,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n77,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n109,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n101,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n48,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n59,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n43,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n86,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n92,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n103,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n82,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n46,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n41,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n99,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n61,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n98,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n39,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n104,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n42,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n80,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n87,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n71,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n113,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n53,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n69,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n63,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n33,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n122,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n51,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n107,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n60,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n128,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n83,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n132,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n117,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n131,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n116,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n40,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n67,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n62,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n129,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n91,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n112,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n96,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n110,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n90,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n65,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n79,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n125,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n81,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n121,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n44,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n35,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n36,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n75,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n108,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n45,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n119,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n118,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n115,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n74,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n93,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


