// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_43 written by SynthGen on 2021/04/05 11:08:37
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_43 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n108, n118, n127, n131, n124, n115, n125, n116,
 n101, n126, n129, n111, n112, n110, n120, n123,
 n104, n130, n113, n132, n128, n102, n114, n119,
 n109, n121, n122, n105, n106, n107, n117, n103);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n108, n118, n127, n131, n124, n115, n125, n116,
 n101, n126, n129, n111, n112, n110, n120, n123,
 n104, n130, n113, n132, n128, n102, n114, n119,
 n109, n121, n122, n105, n106, n107, n117, n103;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

not  g0 (n43, n3);
not  g1 (n46, n4);
not  g2 (n33, n2);
buf  g3 (n39, n2);
not  g4 (n44, n2);
not  g5 (n47, n1);
not  g6 (n38, n1);
not  g7 (n35, n3);
not  g8 (n36, n3);
not  g9 (n37, n3);
not  g10 (n40, n4);
not  g11 (n45, n1);
buf  g12 (n34, n4);
not  g13 (n41, n1);
buf  g14 (n42, n2);
buf  g15 (n55, n7);
not  g16 (n76, n44);
not  g17 (n49, n24);
not  g18 (n57, n27);
not  g19 (n63, n38);
buf  g20 (n73, n35);
or   g21 (n79, n12, n9, n13);
xnor g22 (n89, n34, n24, n8, n7);
nand g23 (n88, n38, n5, n22, n21);
xor  g24 (n78, n29, n11, n31, n39);
xor  g25 (n51, n37, n30, n20, n43);
and  g26 (n92, n23, n20, n14, n44);
xnor g27 (n48, n27, n10, n34, n15);
nand g28 (n71, n39, n19, n17, n37);
nand g29 (n72, n34, n15, n29, n31);
xnor g30 (n64, n41, n37, n6, n26);
nor  g31 (n75, n22, n22, n30, n35);
nand g32 (n77, n29, n44, n18, n17);
nand g33 (n56, n33, n29, n10, n17);
xor  g34 (n53, n43, n28, n41, n14);
or   g35 (n81, n32, n21, n42, n26);
or   g36 (n91, n17, n12, n30, n26);
nand g37 (n61, n16, n9, n26, n43);
xor  g38 (n52, n31, n42, n20, n30);
xnor g39 (n82, n21, n19, n6, n5);
and  g40 (n84, n45, n16, n9, n23);
xor  g41 (n86, n18, n18, n24, n36);
xor  g42 (n80, n44, n11, n5, n25);
nor  g43 (n67, n45, n40, n19, n42);
and  g44 (n62, n25, n12, n38, n22);
xor  g45 (n87, n32, n42, n8, n35);
nor  g46 (n83, n40, n14, n15, n7);
and  g47 (n66, n23, n15, n37, n32);
and  g48 (n90, n28, n5, n25, n41);
nand g49 (n68, n16, n23, n31, n34);
and  g50 (n50, n16, n45, n6, n10);
or   g51 (n59, n39, n9, n25, n7);
nor  g52 (n60, n36, n40, n35, n38);
xor  g53 (n54, n14, n28, n36);
nor  g54 (n58, n21, n40, n27, n43);
nand g55 (n69, n41, n8, n28);
nand g56 (n70, n18, n27, n11);
xnor g57 (n65, n12, n13, n24);
nand g58 (n85, n39, n4, n10, n6);
and  g59 (n74, n20, n45, n19, n32);
buf  g60 (n97, n51);
not  g61 (n100, n47);
not  g62 (n95, n48);
not  g63 (n99, n50);
xor  g64 (n96, n47, n58, n46);
nand g65 (n93, n47, n49, n57, n53);
xnor g66 (n94, n56, n46, n52);
nor  g67 (n98, n47, n59, n54, n55);
or   g68 (n102, n90, n75, n87, n83);
xor  g69 (n104, n96, n90, n79, n89);
xnor g70 (n106, n67, n72, n60, n90);
nand g71 (n130, n81, n61, n84, n93);
nor  g72 (n113, n85, n73, n77, n93);
xnor g73 (n122, n97, n80, n83, n89);
xor  g74 (n109, n85, n95, n99, n90);
xor  g75 (n118, n99, n89, n77, n68);
or   g76 (n117, n75, n74, n78, n92);
xnor g77 (n125, n81, n76, n72, n85);
nor  g78 (n123, n85, n77, n82, n92);
nor  g79 (n114, n89, n76, n70, n64);
nand g80 (n128, n100, n74, n96, n95);
xnor g81 (n129, n83, n75, n93, n73);
xnor g82 (n107, n96, n88, n95, n79);
xnor g83 (n127, n80, n65, n81, n73);
xor  g84 (n112, n86, n87, n91, n97);
or   g85 (n111, n100, n82, n66, n72);
nor  g86 (n126, n100, n96, n93, n92);
xnor g87 (n116, n94, n95, n62, n86);
or   g88 (n131, n79, n78, n98, n81);
nand g89 (n101, n84, n94, n72, n88);
xor  g90 (n105, n91, n77, n97, n71);
xnor g91 (n110, n98, n86, n99, n97);
xor  g92 (n124, n91, n82, n74, n76);
or   g93 (n132, n94, n94, n87, n76);
xnor g94 (n115, n86, n88, n78, n82);
nand g95 (n108, n63, n73, n99, n80);
and  g96 (n103, n74, n79, n84, n91);
nand g97 (n119, n92, n88, n80, n98);
and  g98 (n121, n87, n75, n100, n69);
or   g99 (n120, n83, n84, n98, n78);
endmodule
