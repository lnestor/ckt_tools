

module Stat_1684_57_8
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n1145,
  n1171,
  n1162,
  n1154,
  n1164,
  n1174,
  n1177,
  n1153,
  n1235,
  n1234,
  n1557,
  n1552,
  n1558,
  n1553,
  n1559,
  n1554,
  n1701,
  n1703,
  n1702,
  n1705,
  n1713
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1145;output n1171;output n1162;output n1154;output n1164;output n1174;output n1177;output n1153;output n1235;output n1234;output n1557;output n1552;output n1558;output n1553;output n1559;output n1554;output n1701;output n1703;output n1702;output n1705;output n1713;
  wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1163;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1172;wire n1173;wire n1175;wire n1176;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1555;wire n1556;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1704;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n47,
    n21
  );


  buf
  g1
  (
    n96,
    n20
  );


  buf
  g2
  (
    n66,
    n29
  );


  not
  g3
  (
    n92,
    n19
  );


  buf
  g4
  (
    n137,
    n18
  );


  not
  g5
  (
    n144,
    n6
  );


  buf
  g6
  (
    n123,
    n6
  );


  buf
  g7
  (
    n43,
    n17
  );


  not
  g8
  (
    n114,
    n21
  );


  buf
  g9
  (
    n91,
    n17
  );


  buf
  g10
  (
    n94,
    n19
  );


  not
  g11
  (
    n112,
    n7
  );


  buf
  g12
  (
    n64,
    n23
  );


  not
  g13
  (
    n132,
    n1
  );


  buf
  g14
  (
    n126,
    n14
  );


  not
  g15
  (
    n46,
    n10
  );


  buf
  g16
  (
    n48,
    n14
  );


  buf
  g17
  (
    n74,
    n19
  );


  buf
  g18
  (
    n31,
    n25
  );


  buf
  g19
  (
    n51,
    n10
  );


  buf
  g20
  (
    n134,
    n7
  );


  buf
  g21
  (
    n53,
    n2
  );


  buf
  g22
  (
    n117,
    n6
  );


  not
  g23
  (
    n65,
    n26
  );


  buf
  g24
  (
    n34,
    n7
  );


  buf
  g25
  (
    n40,
    n26
  );


  not
  g26
  (
    n76,
    n26
  );


  buf
  g27
  (
    n105,
    n8
  );


  buf
  g28
  (
    n32,
    n5
  );


  buf
  g29
  (
    n56,
    n18
  );


  not
  g30
  (
    n107,
    n29
  );


  buf
  g31
  (
    n82,
    n16
  );


  buf
  g32
  (
    n59,
    n4
  );


  not
  g33
  (
    n75,
    n3
  );


  not
  g34
  (
    n90,
    n16
  );


  not
  g35
  (
    n83,
    n11
  );


  not
  g36
  (
    n111,
    n1
  );


  not
  g37
  (
    n88,
    n3
  );


  buf
  g38
  (
    n143,
    n8
  );


  buf
  g39
  (
    n100,
    n16
  );


  not
  g40
  (
    n129,
    n24
  );


  not
  g41
  (
    n49,
    n18
  );


  buf
  g42
  (
    n99,
    n4
  );


  buf
  g43
  (
    n145,
    n27
  );


  not
  g44
  (
    n86,
    n10
  );


  buf
  g45
  (
    n125,
    n2
  );


  not
  g46
  (
    n55,
    n11
  );


  not
  g47
  (
    n85,
    n1
  );


  not
  g48
  (
    n61,
    n19
  );


  not
  g49
  (
    n72,
    n17
  );


  not
  g50
  (
    n109,
    n9
  );


  not
  g51
  (
    n140,
    n15
  );


  not
  g52
  (
    n122,
    n18
  );


  not
  g53
  (
    n57,
    n15
  );


  not
  g54
  (
    n38,
    n4
  );


  not
  g55
  (
    n128,
    n25
  );


  not
  g56
  (
    n133,
    n5
  );


  buf
  g57
  (
    n33,
    n16
  );


  not
  g58
  (
    n95,
    n14
  );


  not
  g59
  (
    n79,
    n20
  );


  not
  g60
  (
    n124,
    n13
  );


  not
  g61
  (
    n142,
    n29
  );


  not
  g62
  (
    n69,
    n21
  );


  buf
  g63
  (
    n50,
    n9
  );


  not
  g64
  (
    n68,
    n22
  );


  buf
  g65
  (
    n135,
    n12
  );


  not
  g66
  (
    n71,
    n22
  );


  not
  g67
  (
    n116,
    n23
  );


  buf
  g68
  (
    n54,
    n23
  );


  not
  g69
  (
    n101,
    n8
  );


  not
  g70
  (
    n36,
    n12
  );


  buf
  g71
  (
    n60,
    n13
  );


  not
  g72
  (
    n119,
    n3
  );


  buf
  g73
  (
    KeyWire_0_12,
    n28
  );


  not
  g74
  (
    n118,
    n28
  );


  not
  g75
  (
    n41,
    n26
  );


  not
  g76
  (
    n67,
    n23
  );


  buf
  g77
  (
    n108,
    n15
  );


  buf
  g78
  (
    n127,
    n13
  );


  buf
  g79
  (
    n45,
    n25
  );


  not
  g80
  (
    n81,
    n24
  );


  not
  g81
  (
    n84,
    n5
  );


  not
  g82
  (
    n120,
    n15
  );


  not
  g83
  (
    n63,
    n24
  );


  buf
  g84
  (
    n141,
    n22
  );


  buf
  g85
  (
    n78,
    n24
  );


  not
  g86
  (
    n73,
    n13
  );


  not
  g87
  (
    n110,
    n11
  );


  not
  g88
  (
    n103,
    n29
  );


  not
  g89
  (
    n93,
    n17
  );


  buf
  g90
  (
    n113,
    n3
  );


  not
  g91
  (
    n62,
    n28
  );


  not
  g92
  (
    n52,
    n10
  );


  buf
  g93
  (
    n70,
    n20
  );


  buf
  g94
  (
    KeyWire_0_17,
    n2
  );


  not
  g95
  (
    n121,
    n28
  );


  buf
  g96
  (
    n87,
    n27
  );


  buf
  g97
  (
    n98,
    n22
  );


  not
  g98
  (
    n77,
    n4
  );


  buf
  g99
  (
    n80,
    n27
  );


  not
  g100
  (
    n42,
    n25
  );


  not
  g101
  (
    n115,
    n9
  );


  not
  g102
  (
    n139,
    n21
  );


  not
  g103
  (
    n35,
    n1
  );


  not
  g104
  (
    n30,
    n27
  );


  buf
  g105
  (
    KeyWire_0_14,
    n7
  );


  buf
  g106
  (
    n106,
    n2
  );


  buf
  g107
  (
    n104,
    n12
  );


  not
  g108
  (
    n44,
    n6
  );


  buf
  g109
  (
    n130,
    n5
  );


  not
  g110
  (
    n97,
    n14
  );


  buf
  g111
  (
    n131,
    n8
  );


  not
  g112
  (
    n102,
    n12
  );


  not
  g113
  (
    n89,
    n9
  );


  not
  g114
  (
    n136,
    n11
  );


  buf
  g115
  (
    n138,
    n20
  );


  buf
  g116
  (
    n367,
    n57
  );


  buf
  g117
  (
    n525,
    n84
  );


  buf
  g118
  (
    n241,
    n74
  );


  not
  g119
  (
    n154,
    n110
  );


  not
  g120
  (
    n260,
    n82
  );


  not
  g121
  (
    n225,
    n132
  );


  not
  g122
  (
    n333,
    n32
  );


  buf
  g123
  (
    n362,
    n125
  );


  not
  g124
  (
    n325,
    n142
  );


  not
  g125
  (
    n353,
    n72
  );


  not
  g126
  (
    n340,
    n126
  );


  not
  g127
  (
    n151,
    n89
  );


  not
  g128
  (
    n237,
    n132
  );


  not
  g129
  (
    n196,
    n125
  );


  buf
  g130
  (
    n398,
    n108
  );


  not
  g131
  (
    n257,
    n64
  );


  not
  g132
  (
    n560,
    n56
  );


  not
  g133
  (
    n312,
    n97
  );


  buf
  g134
  (
    n542,
    n107
  );


  buf
  g135
  (
    n566,
    n103
  );


  not
  g136
  (
    n556,
    n100
  );


  buf
  g137
  (
    n267,
    n125
  );


  not
  g138
  (
    n538,
    n127
  );


  buf
  g139
  (
    n388,
    n53
  );


  not
  g140
  (
    n450,
    n72
  );


  not
  g141
  (
    n193,
    n141
  );


  not
  g142
  (
    n483,
    n67
  );


  not
  g143
  (
    n549,
    n34
  );


  not
  g144
  (
    n471,
    n95
  );


  not
  g145
  (
    n210,
    n140
  );


  buf
  g146
  (
    n463,
    n37
  );


  buf
  g147
  (
    n183,
    n133
  );


  buf
  g148
  (
    n270,
    n77
  );


  not
  g149
  (
    n247,
    n94
  );


  not
  g150
  (
    n360,
    n57
  );


  buf
  g151
  (
    n551,
    n69
  );


  buf
  g152
  (
    n261,
    n102
  );


  not
  g153
  (
    n147,
    n140
  );


  not
  g154
  (
    n293,
    n35
  );


  buf
  g155
  (
    n171,
    n142
  );


  buf
  g156
  (
    n350,
    n61
  );


  buf
  g157
  (
    n508,
    n79
  );


  buf
  g158
  (
    n440,
    n75
  );


  not
  g159
  (
    n331,
    n117
  );


  not
  g160
  (
    n491,
    n60
  );


  buf
  g161
  (
    n443,
    n107
  );


  buf
  g162
  (
    n243,
    n68
  );


  not
  g163
  (
    n596,
    n33
  );


  buf
  g164
  (
    n164,
    n102
  );


  not
  g165
  (
    n368,
    n131
  );


  buf
  g166
  (
    n249,
    n112
  );


  not
  g167
  (
    n413,
    n99
  );


  not
  g168
  (
    n266,
    n35
  );


  buf
  g169
  (
    n271,
    n97
  );


  buf
  g170
  (
    n386,
    n85
  );


  not
  g171
  (
    n304,
    n132
  );


  not
  g172
  (
    n289,
    n88
  );


  buf
  g173
  (
    n191,
    n41
  );


  buf
  g174
  (
    n373,
    n139
  );


  buf
  g175
  (
    n390,
    n131
  );


  not
  g176
  (
    n263,
    n45
  );


  buf
  g177
  (
    n153,
    n128
  );


  buf
  g178
  (
    n274,
    n67
  );


  buf
  g179
  (
    n295,
    n129
  );


  not
  g180
  (
    n215,
    n79
  );


  not
  g181
  (
    n516,
    n48
  );


  not
  g182
  (
    n518,
    n83
  );


  not
  g183
  (
    n514,
    n91
  );


  buf
  g184
  (
    n434,
    n144
  );


  not
  g185
  (
    n348,
    n81
  );


  buf
  g186
  (
    n207,
    n113
  );


  not
  g187
  (
    n364,
    n41
  );


  buf
  g188
  (
    n506,
    n61
  );


  buf
  g189
  (
    n519,
    n94
  );


  buf
  g190
  (
    n476,
    n96
  );


  not
  g191
  (
    n269,
    n115
  );


  not
  g192
  (
    n321,
    n97
  );


  buf
  g193
  (
    n453,
    n64
  );


  buf
  g194
  (
    n588,
    n118
  );


  not
  g195
  (
    n157,
    n46
  );


  not
  g196
  (
    n320,
    n37
  );


  not
  g197
  (
    n166,
    n33
  );


  not
  g198
  (
    n279,
    n35
  );


  buf
  g199
  (
    n580,
    n120
  );


  not
  g200
  (
    n258,
    n116
  );


  buf
  g201
  (
    n490,
    n124
  );


  not
  g202
  (
    n250,
    n88
  );


  buf
  g203
  (
    n593,
    n59
  );


  not
  g204
  (
    n280,
    n43
  );


  not
  g205
  (
    n239,
    n67
  );


  not
  g206
  (
    n167,
    n103
  );


  not
  g207
  (
    n475,
    n97
  );


  not
  g208
  (
    n392,
    n47
  );


  buf
  g209
  (
    n235,
    n39
  );


  not
  g210
  (
    n494,
    n89
  );


  not
  g211
  (
    n452,
    n123
  );


  buf
  g212
  (
    n406,
    n136
  );


  not
  g213
  (
    n176,
    n71
  );


  not
  g214
  (
    n276,
    n78
  );


  not
  g215
  (
    n488,
    n74
  );


  not
  g216
  (
    n517,
    n105
  );


  buf
  g217
  (
    n173,
    n133
  );


  not
  g218
  (
    n217,
    n139
  );


  buf
  g219
  (
    n165,
    n53
  );


  buf
  g220
  (
    n532,
    n45
  );


  not
  g221
  (
    n430,
    n73
  );


  buf
  g222
  (
    n464,
    n96
  );


  not
  g223
  (
    n534,
    n36
  );


  not
  g224
  (
    KeyWire_0_0,
    n128
  );


  buf
  g225
  (
    n179,
    n31
  );


  not
  g226
  (
    n457,
    n100
  );


  not
  g227
  (
    n446,
    n105
  );


  not
  g228
  (
    n567,
    n98
  );


  not
  g229
  (
    n211,
    n58
  );


  not
  g230
  (
    n273,
    n145
  );


  buf
  g231
  (
    n444,
    n122
  );


  not
  g232
  (
    n427,
    n82
  );


  not
  g233
  (
    n423,
    n114
  );


  not
  g234
  (
    n418,
    n54
  );


  not
  g235
  (
    n482,
    n119
  );


  buf
  g236
  (
    n294,
    n95
  );


  not
  g237
  (
    n318,
    n75
  );


  buf
  g238
  (
    n161,
    n50
  );


  buf
  g239
  (
    n579,
    n39
  );


  buf
  g240
  (
    n282,
    n59
  );


  buf
  g241
  (
    n485,
    n55
  );


  buf
  g242
  (
    n302,
    n118
  );


  not
  g243
  (
    n449,
    n106
  );


  not
  g244
  (
    n428,
    n45
  );


  buf
  g245
  (
    n592,
    n31
  );


  not
  g246
  (
    n172,
    n39
  );


  not
  g247
  (
    n507,
    n85
  );


  buf
  g248
  (
    n358,
    n111
  );


  buf
  g249
  (
    n572,
    n32
  );


  not
  g250
  (
    n334,
    n107
  );


  not
  g251
  (
    n550,
    n145
  );


  not
  g252
  (
    n512,
    n131
  );


  buf
  g253
  (
    n437,
    n38
  );


  not
  g254
  (
    n431,
    n104
  );


  buf
  g255
  (
    n349,
    n35
  );


  buf
  g256
  (
    n425,
    n60
  );


  buf
  g257
  (
    n410,
    n135
  );


  buf
  g258
  (
    n474,
    n68
  );


  not
  g259
  (
    n332,
    n40
  );


  not
  g260
  (
    n600,
    n130
  );


  not
  g261
  (
    n382,
    n72
  );


  not
  g262
  (
    n578,
    n36
  );


  buf
  g263
  (
    n223,
    n58
  );


  not
  g264
  (
    n315,
    n99
  );


  buf
  g265
  (
    n565,
    n56
  );


  not
  g266
  (
    n497,
    n110
  );


  buf
  g267
  (
    n585,
    n44
  );


  buf
  g268
  (
    n231,
    n77
  );


  not
  g269
  (
    n194,
    n76
  );


  buf
  g270
  (
    n394,
    n37
  );


  not
  g271
  (
    n272,
    n138
  );


  buf
  g272
  (
    n277,
    n34
  );


  not
  g273
  (
    n355,
    n85
  );


  buf
  g274
  (
    n376,
    n64
  );


  buf
  g275
  (
    n533,
    n105
  );


  not
  g276
  (
    n470,
    n116
  );


  buf
  g277
  (
    n416,
    n48
  );


  not
  g278
  (
    n404,
    n102
  );


  not
  g279
  (
    n393,
    n44
  );


  buf
  g280
  (
    n552,
    n88
  );


  buf
  g281
  (
    n501,
    n128
  );


  not
  g282
  (
    n541,
    n124
  );


  buf
  g283
  (
    n149,
    n99
  );


  not
  g284
  (
    n341,
    n66
  );


  buf
  g285
  (
    n181,
    n38
  );


  buf
  g286
  (
    n445,
    n120
  );


  buf
  g287
  (
    n503,
    n50
  );


  buf
  g288
  (
    n384,
    n63
  );


  not
  g289
  (
    n454,
    n119
  );


  buf
  g290
  (
    n292,
    n67
  );


  buf
  g291
  (
    n442,
    n71
  );


  buf
  g292
  (
    n213,
    n105
  );


  not
  g293
  (
    n264,
    n78
  );


  not
  g294
  (
    n229,
    n56
  );


  buf
  g295
  (
    n298,
    n117
  );


  not
  g296
  (
    n553,
    n69
  );


  buf
  g297
  (
    n544,
    n86
  );


  buf
  g298
  (
    n493,
    n75
  );


  not
  g299
  (
    n421,
    n92
  );


  buf
  g300
  (
    n182,
    n102
  );


  not
  g301
  (
    n219,
    n145
  );


  not
  g302
  (
    n528,
    n143
  );


  not
  g303
  (
    n426,
    n138
  );


  buf
  g304
  (
    n226,
    n93
  );


  not
  g305
  (
    n300,
    n54
  );


  buf
  g306
  (
    n597,
    n104
  );


  not
  g307
  (
    n162,
    n81
  );


  not
  g308
  (
    n220,
    n39
  );


  buf
  g309
  (
    n422,
    n86
  );


  not
  g310
  (
    n547,
    n64
  );


  buf
  g311
  (
    n594,
    n56
  );


  not
  g312
  (
    n366,
    n78
  );


  buf
  g313
  (
    n439,
    n93
  );


  buf
  g314
  (
    n352,
    n134
  );


  buf
  g315
  (
    n356,
    n120
  );


  buf
  g316
  (
    n511,
    n60
  );


  not
  g317
  (
    n351,
    n100
  );


  buf
  g318
  (
    n316,
    n55
  );


  not
  g319
  (
    n570,
    n137
  );


  not
  g320
  (
    n526,
    n51
  );


  not
  g321
  (
    n248,
    n114
  );


  not
  g322
  (
    n308,
    n62
  );


  buf
  g323
  (
    n401,
    n50
  );


  buf
  g324
  (
    n199,
    n84
  );


  buf
  g325
  (
    n458,
    n91
  );


  not
  g326
  (
    n344,
    n134
  );


  buf
  g327
  (
    n178,
    n33
  );


  not
  g328
  (
    n381,
    n110
  );


  buf
  g329
  (
    n288,
    n101
  );


  not
  g330
  (
    n346,
    n93
  );


  buf
  g331
  (
    n584,
    n98
  );


  buf
  g332
  (
    n252,
    n57
  );


  buf
  g333
  (
    n451,
    n77
  );


  buf
  g334
  (
    n152,
    n77
  );


  not
  g335
  (
    n411,
    n75
  );


  not
  g336
  (
    n177,
    n30
  );


  not
  g337
  (
    n537,
    n41
  );


  not
  g338
  (
    n540,
    n117
  );


  buf
  g339
  (
    n407,
    n121
  );


  buf
  g340
  (
    n343,
    n40
  );


  buf
  g341
  (
    n399,
    n100
  );


  buf
  g342
  (
    n405,
    n60
  );


  buf
  g343
  (
    n548,
    n81
  );


  buf
  g344
  (
    n265,
    n108
  );


  buf
  g345
  (
    n326,
    n115
  );


  not
  g346
  (
    n203,
    n135
  );


  buf
  g347
  (
    n189,
    n30
  );


  not
  g348
  (
    n230,
    n122
  );


  buf
  g349
  (
    n371,
    n94
  );


  not
  g350
  (
    n502,
    n66
  );


  not
  g351
  (
    n383,
    n112
  );


  buf
  g352
  (
    n509,
    n126
  );


  not
  g353
  (
    n268,
    n90
  );


  not
  g354
  (
    n562,
    n59
  );


  not
  g355
  (
    n286,
    n130
  );


  not
  g356
  (
    n221,
    n61
  );


  buf
  g357
  (
    n198,
    n93
  );


  not
  g358
  (
    n290,
    n127
  );


  buf
  g359
  (
    n543,
    n98
  );


  buf
  g360
  (
    n159,
    n101
  );


  buf
  g361
  (
    n424,
    n92
  );


  buf
  g362
  (
    n233,
    n141
  );


  not
  g363
  (
    n253,
    n51
  );


  not
  g364
  (
    n484,
    n43
  );


  not
  g365
  (
    KeyWire_0_29,
    n143
  );


  buf
  g366
  (
    n190,
    n49
  );


  not
  g367
  (
    n586,
    n126
  );


  not
  g368
  (
    n150,
    n44
  );


  buf
  g369
  (
    n574,
    n37
  );


  not
  g370
  (
    n313,
    n47
  );


  buf
  g371
  (
    n520,
    n123
  );


  buf
  g372
  (
    n587,
    n125
  );


  not
  g373
  (
    n531,
    n52
  );


  not
  g374
  (
    n380,
    n42
  );


  not
  g375
  (
    n322,
    n41
  );


  not
  g376
  (
    n414,
    n54
  );


  not
  g377
  (
    n323,
    n70
  );


  not
  g378
  (
    n459,
    n114
  );


  not
  g379
  (
    n499,
    n115
  );


  buf
  g380
  (
    n468,
    n95
  );


  buf
  g381
  (
    n432,
    n111
  );


  buf
  g382
  (
    n208,
    n122
  );


  buf
  g383
  (
    n573,
    n71
  );


  buf
  g384
  (
    n400,
    n65
  );


  not
  g385
  (
    n224,
    n80
  );


  buf
  g386
  (
    n415,
    n48
  );


  not
  g387
  (
    n598,
    n83
  );


  not
  g388
  (
    n436,
    n63
  );


  not
  g389
  (
    n546,
    n126
  );


  not
  g390
  (
    n319,
    n90
  );


  buf
  g391
  (
    n296,
    n130
  );


  not
  g392
  (
    n500,
    n109
  );


  not
  g393
  (
    n256,
    n111
  );


  not
  g394
  (
    n200,
    n53
  );


  buf
  g395
  (
    n187,
    n50
  );


  not
  g396
  (
    n456,
    n129
  );


  not
  g397
  (
    n192,
    n133
  );


  buf
  g398
  (
    n559,
    n121
  );


  not
  g399
  (
    n389,
    n66
  );


  buf
  g400
  (
    KeyWire_0_23,
    n103
  );


  not
  g401
  (
    n378,
    n46
  );


  buf
  g402
  (
    n513,
    n92
  );


  not
  g403
  (
    n186,
    n51
  );


  buf
  g404
  (
    n466,
    n55
  );


  not
  g405
  (
    n524,
    n99
  );


  buf
  g406
  (
    n336,
    n68
  );


  buf
  g407
  (
    n487,
    n96
  );


  buf
  g408
  (
    n591,
    n137
  );


  not
  g409
  (
    n420,
    n31
  );


  buf
  g410
  (
    n455,
    n145
  );


  not
  g411
  (
    n412,
    n36
  );


  buf
  g412
  (
    n480,
    n73
  );


  not
  g413
  (
    n309,
    n104
  );


  not
  g414
  (
    n216,
    n122
  );


  buf
  g415
  (
    n195,
    n128
  );


  buf
  g416
  (
    n460,
    n107
  );


  not
  g417
  (
    n184,
    n62
  );


  buf
  g418
  (
    n174,
    n121
  );


  not
  g419
  (
    n515,
    n70
  );


  not
  g420
  (
    n409,
    n140
  );


  buf
  g421
  (
    n467,
    n58
  );


  not
  g422
  (
    n338,
    n112
  );


  buf
  g423
  (
    n254,
    n136
  );


  not
  g424
  (
    n510,
    n33
  );


  buf
  g425
  (
    n281,
    n136
  );


  not
  g426
  (
    n201,
    n123
  );


  not
  g427
  (
    n595,
    n139
  );


  not
  g428
  (
    n403,
    n57
  );


  not
  g429
  (
    n461,
    n47
  );


  buf
  g430
  (
    n175,
    n40
  );


  buf
  g431
  (
    n576,
    n118
  );


  buf
  g432
  (
    n568,
    n52
  );


  buf
  g433
  (
    n204,
    n34
  );


  buf
  g434
  (
    n299,
    n136
  );


  not
  g435
  (
    n481,
    n71
  );


  not
  g436
  (
    n330,
    n124
  );


  not
  g437
  (
    n354,
    n96
  );


  buf
  g438
  (
    n365,
    n123
  );


  not
  g439
  (
    n244,
    n98
  );


  buf
  g440
  (
    n402,
    n89
  );


  buf
  g441
  (
    n307,
    n111
  );


  not
  g442
  (
    n155,
    n30
  );


  not
  g443
  (
    n554,
    n79
  );


  not
  g444
  (
    n245,
    n143
  );


  buf
  g445
  (
    n387,
    n80
  );


  buf
  g446
  (
    n435,
    n141
  );


  not
  g447
  (
    n287,
    n58
  );


  buf
  g448
  (
    n535,
    n72
  );


  buf
  g449
  (
    n438,
    n74
  );


  buf
  g450
  (
    n169,
    n109
  );


  buf
  g451
  (
    n545,
    n43
  );


  not
  g452
  (
    n297,
    n30
  );


  buf
  g453
  (
    n504,
    n40
  );


  not
  g454
  (
    n582,
    n101
  );


  buf
  g455
  (
    n495,
    n138
  );


  buf
  g456
  (
    n205,
    n137
  );


  not
  g457
  (
    n188,
    n127
  );


  not
  g458
  (
    n234,
    n129
  );


  buf
  g459
  (
    n522,
    n38
  );


  not
  g460
  (
    n214,
    n65
  );


  not
  g461
  (
    n462,
    n138
  );


  not
  g462
  (
    n251,
    n95
  );


  not
  g463
  (
    n328,
    n135
  );


  buf
  g464
  (
    n539,
    n142
  );


  buf
  g465
  (
    n206,
    n118
  );


  buf
  g466
  (
    n291,
    n134
  );


  buf
  g467
  (
    n284,
    n108
  );


  buf
  g468
  (
    n324,
    n78
  );


  buf
  g469
  (
    n303,
    n79
  );


  buf
  g470
  (
    n255,
    n61
  );


  not
  g471
  (
    n521,
    n124
  );


  not
  g472
  (
    n347,
    n83
  );


  buf
  g473
  (
    n575,
    n104
  );


  buf
  g474
  (
    n590,
    n106
  );


  buf
  g475
  (
    n228,
    n70
  );


  buf
  g476
  (
    n377,
    n45
  );


  not
  g477
  (
    n465,
    n32
  );


  not
  g478
  (
    n283,
    n62
  );


  buf
  g479
  (
    n339,
    n49
  );


  not
  g480
  (
    n564,
    n53
  );


  not
  g481
  (
    n555,
    n144
  );


  buf
  g482
  (
    n275,
    n90
  );


  not
  g483
  (
    n492,
    n117
  );


  buf
  g484
  (
    n361,
    n119
  );


  buf
  g485
  (
    n477,
    n76
  );


  not
  g486
  (
    n429,
    n73
  );


  buf
  g487
  (
    n306,
    n92
  );


  buf
  g488
  (
    n561,
    n112
  );


  not
  g489
  (
    n227,
    n91
  );


  buf
  g490
  (
    n530,
    n51
  );


  not
  g491
  (
    n498,
    n82
  );


  not
  g492
  (
    n314,
    n142
  );


  not
  g493
  (
    n337,
    n129
  );


  not
  g494
  (
    n238,
    n66
  );


  buf
  g495
  (
    n391,
    n140
  );


  not
  g496
  (
    n305,
    n141
  );


  buf
  g497
  (
    n345,
    n62
  );


  not
  g498
  (
    KeyWire_0_13,
    n76
  );


  buf
  g499
  (
    n148,
    n86
  );


  not
  g500
  (
    n240,
    n94
  );


  not
  g501
  (
    n583,
    n42
  );


  not
  g502
  (
    n329,
    n59
  );


  not
  g503
  (
    n357,
    n106
  );


  not
  g504
  (
    n218,
    n34
  );


  buf
  g505
  (
    n523,
    n91
  );


  not
  g506
  (
    n417,
    n87
  );


  buf
  g507
  (
    n571,
    n109
  );


  not
  g508
  (
    n478,
    n43
  );


  buf
  g509
  (
    n527,
    n109
  );


  not
  g510
  (
    n335,
    n103
  );


  not
  g511
  (
    n486,
    n87
  );


  buf
  g512
  (
    n359,
    n121
  );


  not
  g513
  (
    n311,
    n63
  );


  not
  g514
  (
    n469,
    n130
  );


  buf
  g515
  (
    n301,
    n113
  );


  buf
  g516
  (
    n379,
    n69
  );


  buf
  g517
  (
    n599,
    n80
  );


  buf
  g518
  (
    n395,
    n85
  );


  buf
  g519
  (
    n577,
    n135
  );


  buf
  g520
  (
    n236,
    n76
  );


  not
  g521
  (
    n558,
    n108
  );


  not
  g522
  (
    n278,
    n38
  );


  buf
  g523
  (
    n385,
    n55
  );


  not
  g524
  (
    n374,
    n90
  );


  buf
  g525
  (
    n479,
    n48
  );


  not
  g526
  (
    n472,
    n68
  );


  not
  g527
  (
    n496,
    n113
  );


  not
  g528
  (
    n327,
    n115
  );


  not
  g529
  (
    n163,
    n84
  );


  buf
  g530
  (
    n342,
    n143
  );


  buf
  g531
  (
    n569,
    n70
  );


  not
  g532
  (
    n317,
    n49
  );


  buf
  g533
  (
    n581,
    n82
  );


  buf
  g534
  (
    n536,
    n137
  );


  buf
  g535
  (
    n160,
    n133
  );


  not
  g536
  (
    n158,
    n83
  );


  buf
  g537
  (
    n372,
    n87
  );


  not
  g538
  (
    n369,
    n87
  );


  buf
  g539
  (
    n448,
    n47
  );


  not
  g540
  (
    n433,
    n52
  );


  buf
  g541
  (
    n209,
    n65
  );


  not
  g542
  (
    n242,
    n73
  );


  not
  g543
  (
    n232,
    n119
  );


  not
  g544
  (
    n505,
    n42
  );


  buf
  g545
  (
    n156,
    n69
  );


  not
  g546
  (
    n180,
    n139
  );


  buf
  g547
  (
    n419,
    n89
  );


  buf
  g548
  (
    n202,
    n144
  );


  buf
  g549
  (
    n370,
    n110
  );


  not
  g550
  (
    n168,
    n106
  );


  not
  g551
  (
    n146,
    n127
  );


  buf
  g552
  (
    n489,
    n63
  );


  not
  g553
  (
    n259,
    n116
  );


  not
  g554
  (
    n473,
    n101
  );


  not
  g555
  (
    n557,
    n81
  );


  buf
  g556
  (
    n529,
    n46
  );


  not
  g557
  (
    n285,
    n80
  );


  not
  g558
  (
    n408,
    n114
  );


  buf
  g559
  (
    n447,
    n88
  );


  not
  g560
  (
    n363,
    n49
  );


  not
  g561
  (
    n375,
    n132
  );


  buf
  g562
  (
    KeyWire_0_27,
    n42
  );


  not
  g563
  (
    n197,
    n36
  );


  not
  g564
  (
    n397,
    n65
  );


  not
  g565
  (
    n262,
    n74
  );


  buf
  g566
  (
    n310,
    n31
  );


  not
  g567
  (
    n170,
    n116
  );


  nor
  g568
  (
    n396,
    n46,
    n54,
    n120,
    n86
  );


  nand
  g569
  (
    n563,
    n134,
    n44,
    n144,
    n32
  );


  xnor
  g570
  (
    n212,
    n52,
    n113,
    n131,
    n84
  );


  xor
  g571
  (
    n607,
    n147,
    n154,
    n168,
    n196
  );


  and
  g572
  (
    n621,
    n214,
    n170,
    n156,
    n233
  );


  or
  g573
  (
    n628,
    n218,
    n188,
    n260,
    n161
  );


  or
  g574
  (
    n612,
    n146,
    n157,
    n255,
    n251
  );


  nand
  g575
  (
    n611,
    n257,
    n160,
    n252,
    n231
  );


  xnor
  g576
  (
    n619,
    n229,
    n205,
    n237,
    n265
  );


  nor
  g577
  (
    n629,
    n199,
    n208,
    n195,
    n179
  );


  xor
  g578
  (
    n626,
    n159,
    n212,
    n200,
    n151
  );


  nor
  g579
  (
    n613,
    n150,
    n165,
    n230,
    n193
  );


  xor
  g580
  (
    n616,
    n213,
    n153,
    n235,
    n167
  );


  nor
  g581
  (
    n623,
    n176,
    n222,
    n262,
    n244
  );


  nand
  g582
  (
    n605,
    n250,
    n259,
    n152,
    n210
  );


  xor
  g583
  (
    n601,
    n184,
    n240,
    n264,
    n225
  );


  and
  g584
  (
    n615,
    n245,
    n253,
    n207,
    n261
  );


  and
  g585
  (
    n630,
    n221,
    n185,
    n227,
    n166
  );


  and
  g586
  (
    n618,
    n173,
    n186,
    n246,
    n194
  );


  nand
  g587
  (
    n631,
    n238,
    n239,
    n216,
    n175
  );


  nand
  g588
  (
    n609,
    n169,
    n198,
    n183,
    n249
  );


  and
  g589
  (
    n606,
    n211,
    n174,
    n148,
    n254
  );


  xnor
  g590
  (
    n617,
    n190,
    n220,
    n228,
    n224
  );


  and
  g591
  (
    n627,
    n162,
    n206,
    n226,
    n217
  );


  xnor
  g592
  (
    n614,
    n234,
    n202,
    n149,
    n248
  );


  nor
  g593
  (
    n603,
    n164,
    n242,
    n219,
    n189
  );


  or
  g594
  (
    n608,
    n191,
    n241,
    n155,
    n197
  );


  xnor
  g595
  (
    n624,
    n268,
    n236,
    n232,
    n177
  );


  xor
  g596
  (
    n622,
    n203,
    n178,
    n204,
    n209
  );


  and
  g597
  (
    n625,
    n192,
    n172,
    n263,
    n171
  );


  nand
  g598
  (
    n610,
    n258,
    n267,
    n266,
    n223
  );


  or
  g599
  (
    n620,
    n180,
    n182,
    n158,
    n201
  );


  nor
  g600
  (
    n602,
    n163,
    n215,
    n247,
    n181
  );


  and
  g601
  (
    n604,
    n269,
    n187,
    n243,
    n256
  );


  xnor
  g602
  (
    n636,
    n286,
    n607,
    n277,
    n275
  );


  xor
  g603
  (
    n633,
    n605,
    n276,
    n274,
    n287
  );


  xnor
  g604
  (
    n634,
    n288,
    n284,
    n282,
    n270
  );


  xor
  g605
  (
    n637,
    n281,
    n272,
    n280,
    n606
  );


  nand
  g606
  (
    n638,
    n278,
    n289,
    n602,
    n603
  );


  xor
  g607
  (
    n635,
    n604,
    n273,
    n283,
    n290
  );


  nor
  g608
  (
    n632,
    n285,
    n279,
    n601,
    n271
  );


  buf
  g609
  (
    n640,
    n635
  );


  not
  g610
  (
    n653,
    n636
  );


  buf
  g611
  (
    n644,
    n634
  );


  buf
  g612
  (
    n646,
    n634
  );


  buf
  g613
  (
    n650,
    n634
  );


  buf
  g614
  (
    n651,
    n634
  );


  buf
  g615
  (
    n649,
    n637
  );


  buf
  g616
  (
    n652,
    n636
  );


  not
  g617
  (
    n639,
    n632
  );


  not
  g618
  (
    n643,
    n635
  );


  buf
  g619
  (
    n645,
    n635
  );


  buf
  g620
  (
    n648,
    n633
  );


  buf
  g621
  (
    n642,
    n636
  );


  buf
  g622
  (
    n641,
    n636
  );


  not
  g623
  (
    n647,
    n635
  );


  nor
  g624
  (
    n660,
    n614,
    n612,
    n646,
    n639
  );


  and
  g625
  (
    n655,
    n618,
    n626,
    n628,
    n627
  );


  nand
  g626
  (
    n659,
    n630,
    n625,
    n615,
    n645
  );


  and
  g627
  (
    n657,
    n619,
    n644,
    n640,
    n608
  );


  xnor
  g628
  (
    n656,
    n616,
    n610,
    n631,
    n623
  );


  nand
  g629
  (
    n661,
    n621,
    n620,
    n611,
    n609
  );


  or
  g630
  (
    n658,
    n641,
    n642,
    n622,
    n613
  );


  xnor
  g631
  (
    n654,
    n643,
    n617,
    n624,
    n629
  );


  not
  g632
  (
    n662,
    n638
  );


  not
  g633
  (
    n669,
    n656
  );


  buf
  g634
  (
    n668,
    n637
  );


  buf
  g635
  (
    n667,
    n637
  );


  buf
  g636
  (
    n666,
    n655
  );


  not
  g637
  (
    n665,
    n661
  );


  nand
  g638
  (
    n663,
    n657,
    n654,
    n637,
    n658
  );


  or
  g639
  (
    n664,
    n659,
    n660,
    n638
  );


  nor
  g640
  (
    n690,
    n668,
    n349,
    n304,
    n320
  );


  nand
  g641
  (
    n688,
    n665,
    n662,
    n299,
    n305
  );


  xor
  g642
  (
    n693,
    n326,
    n303,
    n664,
    n369
  );


  or
  g643
  (
    n686,
    n308,
    n333,
    n358,
    n331
  );


  nor
  g644
  (
    n684,
    n327,
    n321,
    n316,
    n346
  );


  or
  g645
  (
    n694,
    n296,
    n325,
    n371,
    n667
  );


  and
  g646
  (
    n682,
    n662,
    n345,
    n314,
    n364
  );


  nand
  g647
  (
    n675,
    n376,
    n378,
    n302,
    n668
  );


  xnor
  g648
  (
    n674,
    n307,
    n347,
    n356,
    n666
  );


  nand
  g649
  (
    n696,
    n362,
    n310,
    n663,
    n669
  );


  and
  g650
  (
    n681,
    n666,
    n324,
    n348,
    n315
  );


  xnor
  g651
  (
    n689,
    n312,
    n354,
    n664,
    n311
  );


  xor
  g652
  (
    n672,
    n361,
    n669,
    n664,
    n335
  );


  or
  g653
  (
    n680,
    n366,
    n336,
    n351,
    n343
  );


  nor
  g654
  (
    n676,
    n295,
    n360,
    n365,
    n292
  );


  nand
  g655
  (
    n677,
    n667,
    n309,
    n301,
    n662
  );


  xor
  g656
  (
    n670,
    n297,
    n352,
    n344,
    n375
  );


  nor
  g657
  (
    n692,
    n668,
    n330,
    n665,
    n328
  );


  and
  g658
  (
    n698,
    n337,
    n374,
    n353,
    n379
  );


  xnor
  g659
  (
    n695,
    n664,
    n294,
    n350,
    n668
  );


  or
  g660
  (
    n683,
    n368,
    n367,
    n667,
    n359
  );


  nand
  g661
  (
    n691,
    n313,
    n372,
    n665,
    n306
  );


  or
  g662
  (
    n671,
    n319,
    n300,
    n298,
    n322
  );


  nand
  g663
  (
    n679,
    n355,
    n293,
    n332,
    n329
  );


  or
  g664
  (
    n687,
    n662,
    n373,
    n666,
    n342
  );


  nand
  g665
  (
    n699,
    n363,
    n323,
    n377,
    n341
  );


  xnor
  g666
  (
    n673,
    n340,
    n380,
    n663,
    n317
  );


  nor
  g667
  (
    n678,
    n370,
    n663,
    n339,
    n291
  );


  and
  g668
  (
    KeyWire_0_26,
    n667,
    n357,
    n666,
    n665
  );


  xnor
  g669
  (
    n685,
    n663,
    n334,
    n338,
    n318
  );


  not
  g670
  (
    n702,
    n671
  );


  buf
  g671
  (
    n713,
    n670
  );


  buf
  g672
  (
    n714,
    n670
  );


  buf
  g673
  (
    n712,
    n673
  );


  buf
  g674
  (
    n706,
    n670
  );


  buf
  g675
  (
    n709,
    n672
  );


  not
  g676
  (
    n704,
    n673
  );


  buf
  g677
  (
    n710,
    n672
  );


  buf
  g678
  (
    n705,
    n672
  );


  buf
  g679
  (
    n703,
    n671
  );


  buf
  g680
  (
    n700,
    n671
  );


  buf
  g681
  (
    n711,
    n673
  );


  not
  g682
  (
    n707,
    n672
  );


  not
  g683
  (
    n701,
    n670
  );


  buf
  g684
  (
    n708,
    n671
  );


  buf
  g685
  (
    KeyWire_0_15,
    n679
  );


  not
  g686
  (
    n765,
    n678
  );


  not
  g687
  (
    n722,
    n681
  );


  not
  g688
  (
    n734,
    n685
  );


  not
  g689
  (
    n757,
    n684
  );


  buf
  g690
  (
    n752,
    n707
  );


  not
  g691
  (
    n749,
    n700
  );


  buf
  g692
  (
    KeyWire_0_31,
    n706
  );


  buf
  g693
  (
    n720,
    n678
  );


  buf
  g694
  (
    n741,
    n673
  );


  not
  g695
  (
    n756,
    n703
  );


  not
  g696
  (
    n750,
    n702
  );


  not
  g697
  (
    n732,
    n669
  );


  not
  g698
  (
    n743,
    n682
  );


  buf
  g699
  (
    n747,
    n701
  );


  buf
  g700
  (
    n715,
    n679
  );


  not
  g701
  (
    n726,
    n682
  );


  not
  g702
  (
    n740,
    n708
  );


  buf
  g703
  (
    n762,
    n675
  );


  buf
  g704
  (
    n718,
    n677
  );


  buf
  g705
  (
    n735,
    n683
  );


  buf
  g706
  (
    n745,
    n707
  );


  buf
  g707
  (
    n733,
    n705
  );


  buf
  g708
  (
    n738,
    n676
  );


  not
  g709
  (
    n730,
    n708
  );


  buf
  g710
  (
    n731,
    n638
  );


  not
  g711
  (
    n753,
    n709
  );


  buf
  g712
  (
    n728,
    n704
  );


  not
  g713
  (
    n754,
    n703
  );


  not
  g714
  (
    n727,
    n707
  );


  not
  g715
  (
    n764,
    n702
  );


  not
  g716
  (
    n760,
    n684
  );


  not
  g717
  (
    n759,
    n712
  );


  not
  g718
  (
    n737,
    n674
  );


  and
  g719
  (
    n746,
    n678,
    n705,
    n680,
    n700
  );


  or
  g720
  (
    n742,
    n711,
    n707,
    n681,
    n680
  );


  and
  g721
  (
    n723,
    n681,
    n684,
    n701,
    n711
  );


  and
  g722
  (
    n744,
    n712,
    n685,
    n704,
    n700
  );


  nand
  g723
  (
    n721,
    n685,
    n676,
    n704,
    n675
  );


  and
  g724
  (
    n758,
    n706,
    n678,
    n704,
    n712
  );


  or
  g725
  (
    n719,
    n680,
    n710,
    n709,
    n677
  );


  and
  g726
  (
    n748,
    n682,
    n675,
    n701
  );


  nand
  g727
  (
    n755,
    n703,
    n683,
    n702,
    n684
  );


  or
  g728
  (
    n729,
    n679,
    n703,
    n674,
    n677
  );


  xor
  g729
  (
    n725,
    n706,
    n710,
    n702,
    n669
  );


  nand
  g730
  (
    n763,
    n706,
    n705,
    n700,
    n711
  );


  xor
  g731
  (
    n751,
    n709,
    n701,
    n711,
    n676
  );


  xnor
  g732
  (
    n739,
    n710,
    n676,
    n682,
    n681
  );


  xnor
  g733
  (
    n761,
    n683,
    n709,
    n708,
    n705
  );


  xor
  g734
  (
    n716,
    n708,
    n710,
    n683,
    n677
  );


  xnor
  g735
  (
    n717,
    n674,
    n674,
    n680,
    n679
  );


  xor
  g736
  (
    n790,
    n531,
    n503,
    n719,
    n744
  );


  and
  g737
  (
    n797,
    n408,
    n737,
    n443,
    n763
  );


  or
  g738
  (
    n898,
    n404,
    n529,
    n423,
    n688
  );


  and
  g739
  (
    n804,
    n400,
    n689,
    n447,
    n698
  );


  nand
  g740
  (
    n769,
    n523,
    n697,
    n467,
    n429
  );


  or
  g741
  (
    n772,
    n726,
    n443,
    n452,
    n470
  );


  nor
  g742
  (
    n795,
    n471,
    n440,
    n746,
    n542
  );


  xnor
  g743
  (
    n782,
    n482,
    n721,
    n761,
    n429
  );


  xor
  g744
  (
    n836,
    n475,
    n419,
    n500,
    n758
  );


  or
  g745
  (
    n911,
    n750,
    n427,
    n471,
    n761
  );


  nand
  g746
  (
    n874,
    n484,
    n501,
    n493,
    n756
  );


  or
  g747
  (
    n794,
    n500,
    n477,
    n453,
    n429
  );


  xnor
  g748
  (
    n817,
    n747,
    n481,
    n417,
    n735
  );


  xor
  g749
  (
    n877,
    n695,
    n718,
    n508,
    n534
  );


  nor
  g750
  (
    n767,
    n439,
    n436,
    n416,
    n719
  );


  and
  g751
  (
    n905,
    n459,
    n734,
    n762,
    n497
  );


  xnor
  g752
  (
    n876,
    n450,
    n725,
    n448,
    n715
  );


  nor
  g753
  (
    n946,
    n390,
    n431,
    n733,
    n745
  );


  nor
  g754
  (
    n776,
    n716,
    n519,
    n531,
    n479
  );


  or
  g755
  (
    n909,
    n761,
    n426,
    n690,
    n729
  );


  xnor
  g756
  (
    n948,
    n764,
    n729,
    n517,
    n418
  );


  xnor
  g757
  (
    n904,
    n690,
    n463,
    n453,
    n441
  );


  or
  g758
  (
    n964,
    n524,
    n694,
    n422,
    n540
  );


  nor
  g759
  (
    n880,
    n397,
    n686,
    n727,
    n695
  );


  or
  g760
  (
    n936,
    n539,
    n498,
    n504,
    n730
  );


  xnor
  g761
  (
    n785,
    n466,
    n507,
    n526,
    n425
  );


  xor
  g762
  (
    n824,
    n457,
    n751,
    n530,
    n734
  );


  nor
  g763
  (
    n916,
    n494,
    n538,
    n754,
    n720
  );


  xnor
  g764
  (
    n897,
    n510,
    n438,
    n441,
    n734
  );


  nand
  g765
  (
    n969,
    n745,
    n500,
    n431,
    n462
  );


  nor
  g766
  (
    n933,
    n486,
    n435,
    n698,
    n756
  );


  and
  g767
  (
    n925,
    n737,
    n472,
    n517,
    n503
  );


  xnor
  g768
  (
    n770,
    n487,
    n439,
    n498,
    n717
  );


  nand
  g769
  (
    n914,
    n716,
    n724,
    n528,
    n722
  );


  nand
  g770
  (
    n830,
    n449,
    n517,
    n471,
    n442
  );


  nor
  g771
  (
    n822,
    n472,
    n723,
    n509,
    n457
  );


  xor
  g772
  (
    n837,
    n437,
    n430,
    n387,
    n736
  );


  xnor
  g773
  (
    n787,
    n424,
    n757,
    n505,
    n464
  );


  or
  g774
  (
    n811,
    n469,
    n458,
    n528,
    n483
  );


  and
  g775
  (
    n807,
    n413,
    n508,
    n490,
    n693
  );


  and
  g776
  (
    n951,
    n459,
    n519,
    n391,
    n415
  );


  xnor
  g777
  (
    n955,
    n418,
    n755,
    n721,
    n693
  );


  nand
  g778
  (
    n917,
    n739,
    n497,
    n754,
    n396
  );


  or
  g779
  (
    n882,
    n748,
    n492,
    n528,
    n753
  );


  and
  g780
  (
    n862,
    n742,
    n516,
    n447,
    n542
  );


  xor
  g781
  (
    n820,
    n487,
    n520,
    n468,
    n493
  );


  nor
  g782
  (
    n959,
    n523,
    n523,
    n699,
    n475
  );


  or
  g783
  (
    n789,
    n499,
    n538,
    n733,
    n399
  );


  nor
  g784
  (
    n921,
    n473,
    n462,
    n533
  );


  or
  g785
  (
    n828,
    n422,
    n528,
    n728,
    n493
  );


  xor
  g786
  (
    n900,
    n514,
    n418,
    n727,
    n737
  );


  nand
  g787
  (
    n930,
    n409,
    n485,
    n736,
    n487
  );


  or
  g788
  (
    n857,
    n759,
    n747,
    n537,
    n512
  );


  nand
  g789
  (
    n886,
    n537,
    n765,
    n760,
    n726
  );


  or
  g790
  (
    n810,
    n415,
    n454,
    n448,
    n762
  );


  nand
  g791
  (
    n869,
    n489,
    n738,
    n429,
    n473
  );


  and
  g792
  (
    n884,
    n540,
    n451,
    n718,
    n495
  );


  nand
  g793
  (
    n952,
    n693,
    n424,
    n418,
    n478
  );


  nor
  g794
  (
    n966,
    n541,
    n508,
    n753,
    n698
  );


  or
  g795
  (
    n913,
    n513,
    n417,
    n536,
    n730
  );


  or
  g796
  (
    n929,
    n686,
    n691,
    n478,
    n545
  );


  and
  g797
  (
    n931,
    n461,
    n729,
    n497,
    n442
  );


  and
  g798
  (
    n935,
    n685,
    n525,
    n491,
    n444
  );


  xnor
  g799
  (
    n902,
    n518,
    n481,
    n498,
    n466
  );


  xor
  g800
  (
    n812,
    n410,
    n421,
    n512,
    n686
  );


  or
  g801
  (
    n901,
    n476,
    n519,
    n499,
    n464
  );


  and
  g802
  (
    n864,
    n466,
    n537,
    n485,
    n381
  );


  nor
  g803
  (
    n829,
    n759,
    n515,
    n430,
    n725
  );


  nor
  g804
  (
    n919,
    n697,
    n393,
    n479,
    n414
  );


  xnor
  g805
  (
    n808,
    n717,
    n490,
    n454,
    n735
  );


  nor
  g806
  (
    n890,
    n527,
    n422,
    n416,
    n759
  );


  nand
  g807
  (
    n887,
    n449,
    n743,
    n498,
    n474
  );


  xor
  g808
  (
    n831,
    n435,
    n432,
    n526,
    n484
  );


  nand
  g809
  (
    n907,
    n763,
    n461,
    n478,
    n750
  );


  nor
  g810
  (
    n796,
    n733,
    n740,
    n511,
    n460
  );


  nor
  g811
  (
    n849,
    n764,
    n750,
    n448,
    n412
  );


  or
  g812
  (
    n803,
    n759,
    n743,
    n694,
    n729
  );


  nand
  g813
  (
    n863,
    n505,
    n734,
    n445,
    n738
  );


  xnor
  g814
  (
    n844,
    n465,
    n692,
    n697
  );


  xor
  g815
  (
    n814,
    n469,
    n433,
    n740,
    n464
  );


  xnor
  g816
  (
    n816,
    n489,
    n688,
    n432,
    n544
  );


  nor
  g817
  (
    n798,
    n736,
    n444,
    n525,
    n463
  );


  xor
  g818
  (
    n793,
    n522,
    n492,
    n431,
    n742
  );


  nor
  g819
  (
    n865,
    n440,
    n488,
    n446,
    n727
  );


  xor
  g820
  (
    n842,
    n435,
    n533,
    n722,
    n747
  );


  nand
  g821
  (
    n920,
    n543,
    n752,
    n455,
    n720
  );


  nor
  g822
  (
    n826,
    n757,
    n472,
    n758,
    n691
  );


  or
  g823
  (
    n792,
    n382,
    n741,
    n537,
    n521
  );


  xnor
  g824
  (
    n894,
    n433,
    n488,
    n451,
    n437
  );


  nand
  g825
  (
    n768,
    n746,
    n763,
    n524,
    n420
  );


  xor
  g826
  (
    n815,
    n444,
    n717,
    n459,
    n751
  );


  xor
  g827
  (
    n852,
    n715,
    n694,
    n692,
    n454
  );


  or
  g828
  (
    n859,
    n510,
    n541,
    n533,
    n690
  );


  nor
  g829
  (
    n840,
    n751,
    n765,
    n748,
    n507
  );


  xnor
  g830
  (
    n823,
    n521,
    n490,
    n476,
    n403
  );


  nand
  g831
  (
    KeyWire_0_16,
    n473,
    n502,
    n415,
    n715
  );


  and
  g832
  (
    n893,
    n736,
    n427,
    n440,
    n742
  );


  nor
  g833
  (
    n777,
    n507,
    n755,
    n691,
    n495
  );


  nor
  g834
  (
    n924,
    n748,
    n541,
    n757,
    n535
  );


  nand
  g835
  (
    n888,
    n508,
    n695,
    n719,
    n463
  );


  or
  g836
  (
    n806,
    n471,
    n483,
    n436,
    n501
  );


  or
  g837
  (
    n791,
    n505,
    n754,
    n476,
    n423
  );


  nor
  g838
  (
    n775,
    n510,
    n694,
    n506,
    n491
  );


  nand
  g839
  (
    n821,
    n522,
    n446,
    n402,
    n509
  );


  xnor
  g840
  (
    n885,
    n526,
    n486,
    n538,
    n492
  );


  and
  g841
  (
    n847,
    n395,
    n718,
    n406,
    n536
  );


  xor
  g842
  (
    n932,
    n424,
    n439,
    n764,
    n454
  );


  nand
  g843
  (
    n866,
    n689,
    n452,
    n465,
    n470
  );


  nand
  g844
  (
    KeyWire_0_4,
    n451,
    n422,
    n728,
    n763
  );


  nand
  g845
  (
    n871,
    n445,
    n520,
    n536,
    n730
  );


  and
  g846
  (
    n818,
    n728,
    n456,
    n752,
    n423
  );


  or
  g847
  (
    n968,
    n748,
    n758,
    n746,
    n449
  );


  nand
  g848
  (
    n835,
    n467,
    n527,
    n513,
    n442
  );


  or
  g849
  (
    n962,
    n481,
    n497,
    n521,
    n480
  );


  xnor
  g850
  (
    n873,
    n725,
    n474,
    n506,
    n496
  );


  and
  g851
  (
    n944,
    n544,
    n415,
    n726,
    n425
  );


  nor
  g852
  (
    n827,
    n696,
    n419,
    n532,
    n544
  );


  nor
  g853
  (
    n870,
    n443,
    n532,
    n749,
    n488
  );


  or
  g854
  (
    n954,
    n495,
    n520,
    n464,
    n461
  );


  xor
  g855
  (
    n912,
    n721,
    n741,
    n401,
    n383
  );


  xor
  g856
  (
    n773,
    n731,
    n470,
    n485,
    n434
  );


  or
  g857
  (
    n934,
    n527,
    n449,
    n452,
    n389
  );


  or
  g858
  (
    n875,
    n468,
    n425,
    n716,
    n388
  );


  nand
  g859
  (
    n788,
    n437,
    n419,
    n455,
    n752
  );


  xor
  g860
  (
    n802,
    n426,
    n738,
    n750,
    n474
  );


  or
  g861
  (
    n834,
    n501,
    n428,
    n765,
    n747
  );


  xor
  g862
  (
    n843,
    n515,
    n534,
    n755,
    n439
  );


  xnor
  g863
  (
    n774,
    n512,
    n692,
    n420,
    n511
  );


  xnor
  g864
  (
    n949,
    n411,
    n458,
    n722,
    n540
  );


  and
  g865
  (
    n861,
    n478,
    n495,
    n717,
    n740
  );


  xor
  g866
  (
    n963,
    n687,
    n486,
    n732,
    n435
  );


  xor
  g867
  (
    n891,
    n474,
    n430,
    n526,
    n724
  );


  or
  g868
  (
    n805,
    n699,
    n518,
    n500,
    n487
  );


  or
  g869
  (
    n956,
    n758,
    n457,
    n428,
    n441
  );


  nand
  g870
  (
    n853,
    n420,
    n470,
    n448,
    n516
  );


  or
  g871
  (
    n848,
    n539,
    n492,
    n732,
    n543
  );


  or
  g872
  (
    n927,
    n494,
    n434,
    n723,
    n535
  );


  and
  g873
  (
    n915,
    n739,
    n753,
    n384,
    n529
  );


  or
  g874
  (
    n953,
    n504,
    n507,
    n693,
    n720
  );


  and
  g875
  (
    n957,
    n732,
    n456,
    n483,
    n686
  );


  and
  g876
  (
    n781,
    n427,
    n436,
    n484,
    n517
  );


  xnor
  g877
  (
    n928,
    n516,
    n536,
    n741,
    n479
  );


  or
  g878
  (
    n896,
    n461,
    n489,
    n455,
    n735
  );


  xnor
  g879
  (
    n771,
    n503,
    n751,
    n691,
    n433
  );


  nand
  g880
  (
    n960,
    n446,
    n442,
    n731,
    n696
  );


  xnor
  g881
  (
    n868,
    n525,
    n460,
    n516,
    n687
  );


  nand
  g882
  (
    KeyWire_0_6,
    n720,
    n419,
    n446,
    n757
  );


  xor
  g883
  (
    n841,
    n447,
    n491,
    n468,
    n760
  );


  and
  g884
  (
    n854,
    n688,
    n425,
    n743,
    n522
  );


  or
  g885
  (
    n778,
    n484,
    n719,
    n756,
    n398
  );


  and
  g886
  (
    n918,
    n437,
    n513,
    n692,
    n764
  );


  xnor
  g887
  (
    n860,
    n438,
    n509,
    n426,
    n453
  );


  or
  g888
  (
    n923,
    n530,
    n499,
    n480,
    n523
  );


  nor
  g889
  (
    n867,
    n493,
    n417,
    n465,
    n475
  );


  xor
  g890
  (
    n856,
    n434,
    n489,
    n531,
    n530
  );


  xor
  g891
  (
    n833,
    n499,
    n723,
    n741,
    n530
  );


  and
  g892
  (
    n872,
    n761,
    n731,
    n494,
    n762
  );


  and
  g893
  (
    n892,
    n440,
    n472,
    n538,
    n476
  );


  xor
  g894
  (
    n942,
    n744,
    n732,
    n496,
    n718
  );


  xor
  g895
  (
    n958,
    n534,
    n690,
    n749,
    n689
  );


  or
  g896
  (
    n922,
    n721,
    n737,
    n466,
    n695
  );


  xnor
  g897
  (
    n938,
    n436,
    n749,
    n431,
    n469
  );


  or
  g898
  (
    n784,
    n467,
    n432,
    n749,
    n482
  );


  nand
  g899
  (
    n878,
    n451,
    n515,
    n727,
    n509
  );


  or
  g900
  (
    n943,
    n724,
    n386,
    n426,
    n428
  );


  or
  g901
  (
    n813,
    n532,
    n503,
    n756,
    n743
  );


  and
  g902
  (
    n940,
    n696,
    n724,
    n445,
    n752
  );


  xnor
  g903
  (
    KeyWire_0_30,
    n458,
    n739,
    n428,
    n699
  );


  xnor
  g904
  (
    n809,
    n427,
    n453,
    n452,
    n543
  );


  and
  g905
  (
    n910,
    n522,
    n525,
    n545,
    n527
  );


  and
  g906
  (
    n801,
    n491,
    n514,
    n455,
    n465
  );


  xnor
  g907
  (
    n926,
    n441,
    n519,
    n543,
    n520
  );


  xnor
  g908
  (
    n825,
    n424,
    n511,
    n535,
    n531
  );


  or
  g909
  (
    n895,
    n725,
    n434,
    n521,
    n462
  );


  and
  g910
  (
    n832,
    n481,
    n745,
    n423,
    n458
  );


  or
  g911
  (
    n903,
    n430,
    n753,
    n765,
    n696
  );


  xnor
  g912
  (
    n783,
    n755,
    n460,
    n754,
    n480
  );


  nand
  g913
  (
    n850,
    n733,
    n467,
    n421,
    n518
  );


  nor
  g914
  (
    n961,
    n502,
    n506,
    n416,
    n438
  );


  and
  g915
  (
    n858,
    n715,
    n477,
    n735,
    n728
  );


  or
  g916
  (
    n908,
    n502,
    n542,
    n529,
    n450
  );


  nand
  g917
  (
    n800,
    n514,
    n539,
    n501,
    n468
  );


  xor
  g918
  (
    n937,
    n722,
    n417,
    n744,
    n513
  );


  or
  g919
  (
    n879,
    n490,
    n511,
    n504,
    n479
  );


  and
  g920
  (
    n965,
    n745,
    n698,
    n532,
    n740
  );


  and
  g921
  (
    n945,
    n407,
    n535,
    n687,
    n416
  );


  nor
  g922
  (
    n779,
    n438,
    n502,
    n529,
    n485
  );


  xor
  g923
  (
    n799,
    n510,
    n746,
    n524,
    n486
  );


  or
  g924
  (
    n851,
    n488,
    n477,
    n394,
    n716
  );


  nor
  g925
  (
    n950,
    n482,
    n742,
    n539,
    n456
  );


  xnor
  g926
  (
    n819,
    n512,
    n542,
    n421,
    n723
  );


  or
  g927
  (
    n766,
    n726,
    n506,
    n444,
    n392
  );


  and
  g928
  (
    n906,
    n496,
    n504,
    n760,
    n450
  );


  nand
  g929
  (
    n883,
    n760,
    n541,
    n432,
    n762
  );


  nor
  g930
  (
    n947,
    n445,
    n744,
    n420,
    n463
  );


  and
  g931
  (
    n839,
    n540,
    n475,
    n385,
    n689
  );


  xnor
  g932
  (
    n967,
    n496,
    n447,
    n524,
    n480
  );


  or
  g933
  (
    n881,
    n494,
    n433,
    n469,
    n456
  );


  nand
  g934
  (
    n941,
    n457,
    n477,
    n460,
    n739
  );


  or
  g935
  (
    n845,
    n405,
    n459,
    n505,
    n687
  );


  xor
  g936
  (
    n899,
    n514,
    n482,
    n483,
    n515
  );


  xor
  g937
  (
    n889,
    n730,
    n731,
    n688,
    n534
  );


  xnor
  g938
  (
    n939,
    n473,
    n518,
    n533,
    n443
  );


  or
  g939
  (
    n786,
    n738,
    n544,
    n421,
    n450
  );


  buf
  g940
  (
    n1020,
    n810
  );


  not
  g941
  (
    n1001,
    n847
  );


  buf
  g942
  (
    n1018,
    n817
  );


  buf
  g943
  (
    n975,
    n650
  );


  not
  g944
  (
    n992,
    n652
  );


  not
  g945
  (
    n993,
    n831
  );


  buf
  g946
  (
    n1004,
    n792
  );


  buf
  g947
  (
    n984,
    n834
  );


  buf
  g948
  (
    n982,
    n787
  );


  not
  g949
  (
    n1014,
    n778
  );


  not
  g950
  (
    n1022,
    n799
  );


  not
  g951
  (
    n1010,
    n781
  );


  not
  g952
  (
    n1000,
    n712
  );


  buf
  g953
  (
    n986,
    n829
  );


  not
  g954
  (
    n985,
    n819
  );


  buf
  g955
  (
    n995,
    n820
  );


  not
  g956
  (
    n1007,
    n816
  );


  not
  g957
  (
    n1021,
    n804
  );


  buf
  g958
  (
    n976,
    n774
  );


  not
  g959
  (
    n1016,
    n714
  );


  buf
  g960
  (
    n1011,
    n815
  );


  not
  g961
  (
    n1012,
    n822
  );


  not
  g962
  (
    n1015,
    n806
  );


  not
  g963
  (
    n991,
    n845
  );


  buf
  g964
  (
    n981,
    n839
  );


  not
  g965
  (
    n1003,
    n803
  );


  not
  g966
  (
    n1019,
    n843
  );


  buf
  g967
  (
    n1009,
    n824
  );


  not
  g968
  (
    n983,
    n828
  );


  not
  g969
  (
    n1005,
    n794
  );


  buf
  g970
  (
    n997,
    n840
  );


  buf
  g971
  (
    n979,
    n713
  );


  not
  g972
  (
    n978,
    n842
  );


  buf
  g973
  (
    n971,
    n851
  );


  not
  g974
  (
    n1006,
    n832
  );


  nor
  g975
  (
    n1008,
    n653,
    n651,
    n714
  );


  xor
  g976
  (
    n990,
    n800,
    n661,
    n775,
    n835
  );


  or
  g977
  (
    n970,
    n713,
    n661,
    n827,
    n782
  );


  nand
  g978
  (
    n994,
    n808,
    n790,
    n714,
    n809
  );


  or
  g979
  (
    n988,
    n767,
    n811,
    n791,
    n784
  );


  xnor
  g980
  (
    n972,
    n786,
    n849,
    n837,
    n850
  );


  xnor
  g981
  (
    n998,
    n793,
    n648,
    n714,
    n846
  );


  nand
  g982
  (
    n989,
    n788,
    n795,
    n661,
    n796
  );


  or
  g983
  (
    n980,
    n777,
    n769,
    n807,
    n826
  );


  xor
  g984
  (
    n977,
    n797,
    n841,
    n768,
    n779
  );


  nor
  g985
  (
    n996,
    n770,
    n821,
    n814,
    n785
  );


  xnor
  g986
  (
    n974,
    n805,
    n844,
    n647,
    n852
  );


  xor
  g987
  (
    n987,
    n766,
    n801,
    n771,
    n833
  );


  and
  g988
  (
    n1013,
    n783,
    n836,
    n798,
    n773
  );


  and
  g989
  (
    n1017,
    n812,
    n802,
    n813,
    n838
  );


  nor
  g990
  (
    n999,
    n776,
    n772,
    n713,
    n830
  );


  and
  g991
  (
    n1002,
    n649,
    n713,
    n789,
    n848
  );


  nand
  g992
  (
    n973,
    n818,
    n825,
    n780,
    n823
  );


  and
  g993
  (
    n1059,
    n964,
    n1013,
    n940,
    n914
  );


  and
  g994
  (
    n1093,
    n935,
    n935,
    n1019,
    n883
  );


  or
  g995
  (
    n1085,
    n901,
    n1003,
    n908,
    n929
  );


  nand
  g996
  (
    n1098,
    n949,
    n933,
    n938,
    n956
  );


  nor
  g997
  (
    n1032,
    n858,
    n910,
    n1021,
    n905
  );


  xnor
  g998
  (
    n1039,
    n1011,
    n877,
    n935,
    n928
  );


  nor
  g999
  (
    n1074,
    n943,
    n937,
    n957,
    n869
  );


  or
  g1000
  (
    n1025,
    n939,
    n907,
    n979,
    n970
  );


  xor
  g1001
  (
    n1071,
    n936,
    n950,
    n874,
    n885
  );


  xnor
  g1002
  (
    n1096,
    n854,
    n949,
    n943,
    n981
  );


  xnor
  g1003
  (
    n1072,
    n932,
    n960,
    n958,
    n954
  );


  nand
  g1004
  (
    n1035,
    n952,
    n950,
    n955,
    n992
  );


  xor
  g1005
  (
    n1031,
    n1015,
    n1017,
    n954,
    n942
  );


  xnor
  g1006
  (
    n1078,
    n965,
    n940,
    n945,
    n863
  );


  nand
  g1007
  (
    n1047,
    n956,
    n951,
    n1014,
    n987
  );


  or
  g1008
  (
    n1044,
    n1005,
    n958,
    n961,
    n952
  );


  nor
  g1009
  (
    n1037,
    n909,
    n934,
    n973,
    n1022
  );


  xor
  g1010
  (
    n1057,
    n934,
    n947,
    n994,
    n1017
  );


  xor
  g1011
  (
    n1063,
    n1006,
    n978,
    n856,
    n1002
  );


  xor
  g1012
  (
    n1083,
    n952,
    n894,
    n926,
    n985
  );


  or
  g1013
  (
    n1055,
    n1008,
    n957,
    n949,
    n865
  );


  xnor
  g1014
  (
    n1076,
    n963,
    n900,
    n853,
    n975
  );


  nand
  g1015
  (
    n1043,
    n933,
    n911,
    n855,
    n990
  );


  xnor
  g1016
  (
    n1053,
    n878,
    n958,
    n963,
    n956
  );


  nor
  g1017
  (
    n1065,
    n959,
    n918,
    n932,
    n965
  );


  or
  g1018
  (
    n1079,
    n984,
    n921,
    n946,
    n929
  );


  and
  g1019
  (
    n1024,
    n947,
    n895,
    n938,
    n1022
  );


  and
  g1020
  (
    n1049,
    n998,
    n943,
    n965,
    n879
  );


  and
  g1021
  (
    n1056,
    n951,
    n906,
    n948,
    n943
  );


  nand
  g1022
  (
    n1084,
    n986,
    n951,
    n958,
    n941
  );


  nand
  g1023
  (
    n1051,
    n923,
    n962,
    n964,
    n960
  );


  and
  g1024
  (
    n1095,
    n959,
    n966,
    n971,
    n988
  );


  nand
  g1025
  (
    KeyWire_0_8,
    n922,
    n966,
    n931,
    n889
  );


  nand
  g1026
  (
    n1058,
    n962,
    n941,
    n967,
    n937
  );


  nor
  g1027
  (
    n1023,
    n940,
    n942,
    n944,
    n897
  );


  xor
  g1028
  (
    n1068,
    n938,
    n966,
    n931,
    n1019
  );


  nor
  g1029
  (
    n1075,
    n1016,
    n1017,
    n948,
    n1020
  );


  xor
  g1030
  (
    n1034,
    n953,
    n927,
    n929,
    n946
  );


  nand
  g1031
  (
    n1041,
    n932,
    n939,
    n941,
    n997
  );


  nor
  g1032
  (
    n1052,
    n962,
    n944,
    n896,
    n1022
  );


  and
  g1033
  (
    n1082,
    n887,
    n962,
    n866,
    n951
  );


  xor
  g1034
  (
    n1040,
    n1016,
    n936,
    n995,
    n1021
  );


  and
  g1035
  (
    n1048,
    n972,
    n933,
    n948,
    n859
  );


  or
  g1036
  (
    n1054,
    n944,
    n955,
    n956,
    n946
  );


  xnor
  g1037
  (
    n1027,
    n999,
    n1007,
    n991,
    n1020
  );


  nor
  g1038
  (
    n1062,
    n1016,
    n938,
    n857,
    n1019
  );


  nand
  g1039
  (
    n1046,
    n1000,
    n955,
    n1018,
    n948
  );


  xor
  g1040
  (
    n1080,
    n891,
    n902,
    n989,
    n960
  );


  nand
  g1041
  (
    n1097,
    n965,
    n1017,
    n953,
    n959
  );


  nand
  g1042
  (
    n1060,
    n886,
    n941,
    n957,
    n1018
  );


  or
  g1043
  (
    n1069,
    n860,
    n933,
    n974,
    n917
  );


  nand
  g1044
  (
    n1091,
    n903,
    n892,
    n916,
    n955
  );


  nor
  g1045
  (
    n1028,
    n949,
    n940,
    n1015,
    n960
  );


  xor
  g1046
  (
    n1067,
    n929,
    n950,
    n1020
  );


  xor
  g1047
  (
    n1092,
    n945,
    n937,
    n934,
    n931
  );


  nand
  g1048
  (
    n1064,
    n925,
    n996,
    n982,
    n893
  );


  and
  g1049
  (
    n1073,
    n884,
    n1009,
    n947,
    n946
  );


  xor
  g1050
  (
    n1026,
    n930,
    n904,
    n953,
    n937
  );


  and
  g1051
  (
    n1081,
    n957,
    n924,
    n961,
    n1021
  );


  xnor
  g1052
  (
    n1033,
    n867,
    n875,
    n959,
    n942
  );


  nor
  g1053
  (
    n1099,
    n961,
    n977,
    n1020,
    n1021
  );


  nand
  g1054
  (
    n1036,
    n930,
    n935,
    n1010,
    n963
  );


  or
  g1055
  (
    n1061,
    n1016,
    n936,
    n872,
    n890
  );


  nor
  g1056
  (
    n1094,
    n961,
    n1022,
    n976,
    n964
  );


  and
  g1057
  (
    n1029,
    n939,
    n880,
    n881,
    n932
  );


  nand
  g1058
  (
    n1089,
    n964,
    n939,
    n898,
    n952
  );


  nor
  g1059
  (
    n1090,
    n954,
    n864,
    n861,
    n888
  );


  nand
  g1060
  (
    n1077,
    n1012,
    n882,
    n963,
    n966
  );


  nand
  g1061
  (
    n1030,
    n913,
    n993,
    n919,
    n1019
  );


  xnor
  g1062
  (
    n1070,
    n873,
    n947,
    n899,
    n1001
  );


  xor
  g1063
  (
    n1087,
    n983,
    n967,
    n953,
    n868
  );


  xnor
  g1064
  (
    n1088,
    n945,
    n967,
    n870,
    n931
  );


  nand
  g1065
  (
    n1038,
    n1018,
    n912,
    n934,
    n936
  );


  xor
  g1066
  (
    n1042,
    n930,
    n945,
    n876,
    n980
  );


  nor
  g1067
  (
    n1066,
    n944,
    n930,
    n1018,
    n915
  );


  nor
  g1068
  (
    n1050,
    n954,
    n871,
    n1004,
    n862
  );


  xnor
  g1069
  (
    n1086,
    n942,
    n920,
    n1015
  );


  not
  g1070
  (
    n1104,
    n1031
  );


  not
  g1071
  (
    n1106,
    n969
  );


  not
  g1072
  (
    n1109,
    n1028
  );


  buf
  g1073
  (
    n1101,
    n1029
  );


  nand
  g1074
  (
    n1111,
    n967,
    n1027
  );


  and
  g1075
  (
    n1110,
    n1025,
    n1023
  );


  and
  g1076
  (
    n1102,
    n1030,
    n968
  );


  nand
  g1077
  (
    n1108,
    n968,
    n1032
  );


  xor
  g1078
  (
    n1107,
    n968,
    n969
  );


  nor
  g1079
  (
    n1103,
    n969,
    n1026
  );


  or
  g1080
  (
    n1100,
    n1033,
    n968
  );


  xor
  g1081
  (
    n1105,
    n1024,
    n1034
  );


  or
  g1082
  (
    n1147,
    n1109,
    n1111,
    n1078,
    n1104
  );


  or
  g1083
  (
    n1120,
    n1064,
    n1104,
    n1050,
    n1076
  );


  nand
  g1084
  (
    n1125,
    n1056,
    n1040,
    n1064,
    n1052
  );


  xor
  g1085
  (
    n1123,
    n1108,
    n1103,
    n1071,
    n1038
  );


  xor
  g1086
  (
    n1114,
    n1075,
    n1074,
    n1077,
    n1111
  );


  nand
  g1087
  (
    n1136,
    n1110,
    n1070,
    n1043,
    n1039
  );


  nor
  g1088
  (
    n1117,
    n1060,
    n1070,
    n1069,
    n1048
  );


  or
  g1089
  (
    n1128,
    n1067,
    n1067,
    n1062,
    n1065
  );


  nor
  g1090
  (
    n1116,
    n1065,
    n1108,
    n1111,
    n1071
  );


  and
  g1091
  (
    n1144,
    n1110,
    n1078,
    n1056,
    n1111
  );


  or
  g1092
  (
    n1122,
    n1107,
    n1073,
    n1109,
    n1058
  );


  nand
  g1093
  (
    n1145,
    n1066,
    n1057,
    n1044,
    n1104
  );


  nand
  g1094
  (
    n1138,
    n1069,
    n1101,
    n1067,
    n1073
  );


  and
  g1095
  (
    n1140,
    n1105,
    n1058,
    n1064,
    n1062
  );


  xor
  g1096
  (
    n1129,
    n1076,
    n1108,
    n1073,
    n1049
  );


  xnor
  g1097
  (
    n1150,
    n1109,
    n1061,
    n1103,
    n1059
  );


  xor
  g1098
  (
    n1133,
    n1060,
    n1076,
    n1056
  );


  and
  g1099
  (
    n1131,
    n1074,
    n1079,
    n1072,
    n1061
  );


  xor
  g1100
  (
    n1142,
    n1109,
    n1107,
    n1108
  );


  xor
  g1101
  (
    n1119,
    n1075,
    n1057,
    n1051,
    n1106
  );


  nor
  g1102
  (
    n1135,
    n1060,
    n1070,
    n1072,
    n1047
  );


  nor
  g1103
  (
    n1127,
    n1053,
    n1072,
    n1057,
    n1037
  );


  xnor
  g1104
  (
    n1141,
    n1063,
    n1102,
    n1105,
    n1062
  );


  xor
  g1105
  (
    n1137,
    n1106,
    n1075,
    n1110,
    n1042
  );


  nor
  g1106
  (
    n1121,
    n1107,
    n1071,
    n1069,
    n1078
  );


  xnor
  g1107
  (
    n1148,
    n1104,
    n1103,
    n1106
  );


  xnor
  g1108
  (
    n1118,
    n1079,
    n1059,
    n1045,
    n1065
  );


  nor
  g1109
  (
    n1130,
    n1056,
    n1100,
    n1110,
    n1057
  );


  xor
  g1110
  (
    n1149,
    n1058,
    n1072,
    n1055,
    n1064
  );


  xnor
  g1111
  (
    n1146,
    n1071,
    n1059,
    n1041,
    n1068
  );


  or
  g1112
  (
    n1115,
    n1073,
    n1036,
    n1070,
    n1069
  );


  nor
  g1113
  (
    n1134,
    n1075,
    n1066,
    n1065,
    n1074
  );


  or
  g1114
  (
    n1124,
    n1062,
    n1106,
    n1068
  );


  or
  g1115
  (
    n1112,
    n1061,
    n1077,
    n1063,
    n1105
  );


  xnor
  g1116
  (
    n1126,
    n1079,
    n1061,
    n1066,
    n1054
  );


  or
  g1117
  (
    n1143,
    n1063,
    n1063,
    n1058,
    n1035
  );


  nor
  g1118
  (
    n1132,
    n1060,
    n699,
    n1105,
    n1078
  );


  or
  g1119
  (
    n1139,
    n1046,
    n1066,
    n1077
  );


  xor
  g1120
  (
    n1113,
    n1068,
    n1074,
    n1067,
    n1059
  );


  xnor
  g1121
  (
    n1153,
    n1113,
    n1118,
    n1092,
    n1095
  );


  nand
  g1122
  (
    n1151,
    n1087,
    n1083,
    n1094,
    n1123
  );


  xor
  g1123
  (
    n1160,
    n1116,
    n1112,
    n1115,
    n1121
  );


  and
  g1124
  (
    n1154,
    n1080,
    n1082,
    n1096,
    n1122
  );


  or
  g1125
  (
    n1165,
    n1086,
    n1084,
    n1117
  );


  nand
  g1126
  (
    n1157,
    n1120,
    n1083,
    n1088,
    n1091
  );


  and
  g1127
  (
    n1161,
    n1090,
    n1116,
    n1093,
    n1123
  );


  xor
  g1128
  (
    n1152,
    n1117,
    n1114,
    n1094,
    n1115
  );


  xor
  g1129
  (
    n1167,
    n1086,
    n1090,
    n1093,
    n1081
  );


  xor
  g1130
  (
    KeyWire_0_19,
    n1121,
    n1091,
    n1114,
    n1115
  );


  xor
  g1131
  (
    n1162,
    n1086,
    n1082,
    n1084,
    n1114
  );


  and
  g1132
  (
    n1163,
    n1117,
    n1119,
    n1121,
    n1088
  );


  xor
  g1133
  (
    n1175,
    n1120,
    n1085,
    n1087,
    n1114
  );


  and
  g1134
  (
    n1169,
    n1082,
    n1119,
    n1121,
    n1096
  );


  xnor
  g1135
  (
    n1156,
    n1085,
    n1120,
    n1081
  );


  or
  g1136
  (
    KeyWire_0_9,
    n1080,
    n1085,
    n1096,
    n1118
  );


  xnor
  g1137
  (
    n1155,
    n1122,
    n1085,
    n1090,
    n1092
  );


  xnor
  g1138
  (
    n1168,
    n1088,
    n1087,
    n1089
  );


  nor
  g1139
  (
    n1170,
    n1092,
    n1116,
    n1122,
    n1093
  );


  or
  g1140
  (
    n1177,
    n1093,
    n1086,
    n1079,
    n1091
  );


  xor
  g1141
  (
    n1171,
    n1116,
    n1094,
    n1080
  );


  nor
  g1142
  (
    n1158,
    n1122,
    n1088,
    n1089,
    n1090
  );


  xnor
  g1143
  (
    n1159,
    n1080,
    n1119,
    n1087,
    n1095
  );


  and
  g1144
  (
    n1174,
    n1095,
    n1092,
    n1120,
    n1089
  );


  nand
  g1145
  (
    n1172,
    n1118,
    n1091,
    n1082,
    n1095
  );


  nor
  g1146
  (
    n1176,
    n1083,
    n1083,
    n1081,
    n1084
  );


  xor
  g1147
  (
    n1164,
    n1115,
    n1118,
    n1084,
    n1119
  );


  not
  g1148
  (
    n1185,
    n1128
  );


  buf
  g1149
  (
    n1184,
    n1127
  );


  not
  g1150
  (
    n1179,
    n1124
  );


  nand
  g1151
  (
    n1192,
    n1162,
    n1171
  );


  or
  g1152
  (
    n1178,
    n1130,
    n1129,
    n1158,
    n1128
  );


  and
  g1153
  (
    n1190,
    n1123,
    n1126,
    n1127,
    n1129
  );


  and
  g1154
  (
    n1186,
    n1172,
    n1125,
    n1131
  );


  xnor
  g1155
  (
    n1193,
    n1125,
    n1129,
    n1127
  );


  nor
  g1156
  (
    n1183,
    n1124,
    n1124,
    n1165,
    n1132
  );


  or
  g1157
  (
    n1191,
    n1130,
    n1126,
    n1131,
    n1163
  );


  nand
  g1158
  (
    n1180,
    n1167,
    n1170,
    n1124,
    n1128
  );


  xor
  g1159
  (
    n1189,
    n1128,
    n1125,
    n1131,
    n1130
  );


  nor
  g1160
  (
    n1181,
    n1126,
    n1125,
    n1173,
    n1123
  );


  and
  g1161
  (
    n1182,
    n1126,
    n1168,
    n1130,
    n1161
  );


  xnor
  g1162
  (
    n1187,
    n1169,
    n1159,
    n1129,
    n1132
  );


  xnor
  g1163
  (
    n1188,
    n1132,
    n1166,
    n1160,
    n1164
  );


  not
  g1164
  (
    n1204,
    n1134
  );


  not
  g1165
  (
    n1205,
    n1132
  );


  buf
  g1166
  (
    n1196,
    n1190
  );


  not
  g1167
  (
    n1201,
    n1190
  );


  buf
  g1168
  (
    n1210,
    n1191
  );


  not
  g1169
  (
    n1202,
    n1133
  );


  buf
  g1170
  (
    n1211,
    n1184
  );


  buf
  g1171
  (
    n1194,
    n1182
  );


  buf
  g1172
  (
    n1197,
    n1191
  );


  buf
  g1173
  (
    n1199,
    n1133
  );


  buf
  g1174
  (
    n1203,
    n1134
  );


  not
  g1175
  (
    n1207,
    n1190
  );


  buf
  g1176
  (
    n1195,
    n1185
  );


  not
  g1177
  (
    n1212,
    n1178
  );


  not
  g1178
  (
    n1213,
    n1133
  );


  buf
  g1179
  (
    n1200,
    n1181
  );


  and
  g1180
  (
    n1198,
    n1191,
    n1183
  );


  nor
  g1181
  (
    n1208,
    n1133,
    n1189,
    n1179,
    n1188
  );


  and
  g1182
  (
    n1209,
    n1180,
    n1135,
    n1191,
    n1186
  );


  and
  g1183
  (
    n1206,
    n1187,
    n1190,
    n1134
  );


  not
  g1184
  (
    n1225,
    n1098
  );


  buf
  g1185
  (
    n1221,
    n1097
  );


  not
  g1186
  (
    n1223,
    n1195
  );


  not
  g1187
  (
    n1217,
    n1098
  );


  not
  g1188
  (
    n1224,
    n1197
  );


  not
  g1189
  (
    n1218,
    n1097
  );


  not
  g1190
  (
    n1215,
    n1096
  );


  buf
  g1191
  (
    n1216,
    n1098
  );


  and
  g1192
  (
    n1222,
    n1196,
    n1195
  );


  and
  g1193
  (
    n1226,
    n1196,
    n1196,
    n1194,
    n1097
  );


  xnor
  g1194
  (
    n1220,
    n1194,
    n1099,
    n1195
  );


  nand
  g1195
  (
    n1219,
    n1196,
    n1097,
    n1194,
    n1195
  );


  nor
  g1196
  (
    n1214,
    n1194,
    n1098,
    n1099
  );


  or
  g1197
  (
    n1237,
    n1198,
    n1215,
    n1216
  );


  nand
  g1198
  (
    n1231,
    n1205,
    n969,
    n1214,
    n1198
  );


  and
  g1199
  (
    n1236,
    n1216,
    n1204,
    n1201,
    n1214
  );


  nor
  g1200
  (
    n1228,
    n1197,
    n1203,
    n1205,
    n1214
  );


  nand
  g1201
  (
    n1233,
    n1204,
    n1203,
    n1202,
    n1205
  );


  xor
  g1202
  (
    n1229,
    n1202,
    n1199,
    n1201,
    n1214
  );


  or
  g1203
  (
    n1234,
    n1200,
    n1200,
    n1201,
    n1204
  );


  or
  g1204
  (
    n1227,
    n1204,
    n1199,
    n1203,
    n1205
  );


  nor
  g1205
  (
    n1232,
    n1201,
    n1215,
    n1216
  );


  nand
  g1206
  (
    n1238,
    n1197,
    n1200,
    n1215,
    n1198
  );


  or
  g1207
  (
    n1235,
    n1198,
    n1202,
    n1197
  );


  or
  g1208
  (
    n1230,
    n1199,
    n1199,
    n1200,
    n1203
  );


  and
  g1209
  (
    n1246,
    n1233,
    n1236,
    n1229,
    n1142
  );


  xor
  g1210
  (
    n1244,
    n1235,
    n1237,
    n1140
  );


  or
  g1211
  (
    n1245,
    n1238,
    n1139,
    n1231,
    n1138
  );


  xnor
  g1212
  (
    n1241,
    n1140,
    n1141,
    n1136,
    n1137
  );


  nor
  g1213
  (
    KeyWire_0_22,
    n1135,
    n1139,
    n1141,
    n1142
  );


  or
  g1214
  (
    n1239,
    n1141,
    n1139,
    n1137,
    n1136
  );


  nor
  g1215
  (
    n1242,
    n1137,
    n1136,
    n1138,
    n1135
  );


  or
  g1216
  (
    n1248,
    n1230,
    n1135,
    n1141,
    n1142
  );


  nand
  g1217
  (
    n1247,
    n1138,
    n1138,
    n1137,
    n1140
  );


  xnor
  g1218
  (
    n1243,
    n1139,
    n1234,
    n1232,
    n1136
  );


  buf
  g1219
  (
    n1254,
    n1147
  );


  not
  g1220
  (
    n1260,
    n1242
  );


  not
  g1221
  (
    n1258,
    n1143
  );


  nand
  g1222
  (
    n1255,
    n1143,
    n1245,
    n1149
  );


  or
  g1223
  (
    n1257,
    n1143,
    n1142,
    n1148
  );


  and
  g1224
  (
    n1249,
    n1245,
    n1145,
    n1147
  );


  or
  g1225
  (
    n1252,
    n1146,
    n1148,
    n1244,
    n1246
  );


  nor
  g1226
  (
    n1250,
    n1146,
    n1243,
    n1148,
    n1241
  );


  or
  g1227
  (
    n1256,
    n1245,
    n1143,
    n1145,
    n1144
  );


  xor
  g1228
  (
    n1253,
    n1144,
    n1144,
    n1146,
    n1147
  );


  nand
  g1229
  (
    n1259,
    n1240,
    n1239,
    n1146,
    n1245
  );


  xor
  g1230
  (
    n1251,
    n1246,
    n1145,
    n1144
  );


  and
  g1231
  (
    n1264,
    n1249,
    n1254,
    n1257
  );


  nor
  g1232
  (
    n1268,
    n1256,
    n1175,
    n1251,
    n1249
  );


  or
  g1233
  (
    n1267,
    n1174,
    n1254,
    n1255,
    n1251
  );


  nor
  g1234
  (
    KeyWire_0_18,
    n1251,
    n1253,
    n1257,
    n1177
  );


  nand
  g1235
  (
    n1263,
    n1254,
    n1176,
    n1252,
    n1249
  );


  xor
  g1236
  (
    n1269,
    n1250,
    n1252,
    n1255,
    n1253
  );


  nand
  g1237
  (
    n1262,
    n1255,
    n1255,
    n1256,
    n1252
  );


  xor
  g1238
  (
    n1261,
    n1253,
    n1256,
    n1252,
    n1250
  );


  xnor
  g1239
  (
    n1270,
    n1249,
    n1251,
    n1250,
    n1254
  );


  xnor
  g1240
  (
    n1266,
    n1256,
    n1250,
    n1253,
    n1257
  );


  and
  g1241
  (
    n1271,
    n1149,
    n1150
  );


  nor
  g1242
  (
    n1272,
    n1149,
    n1149,
    n1261,
    n1262
  );


  buf
  g1243
  (
    n1275,
    n1206
  );


  not
  g1244
  (
    n1276,
    n1206
  );


  buf
  g1245
  (
    n1273,
    n1271
  );


  buf
  g1246
  (
    n1277,
    n1272
  );


  xnor
  g1247
  (
    n1280,
    n1271,
    n1207
  );


  or
  g1248
  (
    n1279,
    n1272,
    n1271
  );


  or
  g1249
  (
    n1278,
    n1271,
    n1272
  );


  not
  g1250
  (
    n1274,
    n1206
  );


  buf
  g1251
  (
    n1301,
    n1222
  );


  buf
  g1252
  (
    n1288,
    n1221
  );


  buf
  g1253
  (
    n1285,
    n1217
  );


  not
  g1254
  (
    n1304,
    n1274
  );


  not
  g1255
  (
    n1312,
    n1224
  );


  not
  g1256
  (
    n1299,
    n1277
  );


  buf
  g1257
  (
    n1282,
    n1222
  );


  buf
  g1258
  (
    n1307,
    n1222
  );


  not
  g1259
  (
    n1298,
    n1273
  );


  buf
  g1260
  (
    n1284,
    n1192
  );


  not
  g1261
  (
    n1290,
    n1224
  );


  not
  g1262
  (
    n1291,
    n1221
  );


  buf
  g1263
  (
    n1293,
    n1192
  );


  buf
  g1264
  (
    n1311,
    n1275
  );


  buf
  g1265
  (
    n1286,
    n1226
  );


  buf
  g1266
  (
    n1283,
    n1225
  );


  xnor
  g1267
  (
    n1287,
    n1220,
    n1279,
    n1278,
    n1276
  );


  xnor
  g1268
  (
    n1294,
    n1217,
    n1222,
    n1219,
    n1221
  );


  nor
  g1269
  (
    n1292,
    n1278,
    n1273,
    n1276,
    n1223
  );


  xnor
  g1270
  (
    n1296,
    n1277,
    n1219,
    n1226,
    n1276
  );


  nand
  g1271
  (
    n1309,
    n1277,
    n1221,
    n1279,
    n1218
  );


  xor
  g1272
  (
    n1306,
    n1217,
    n1218,
    n1220,
    n1280
  );


  or
  g1273
  (
    n1300,
    n1275,
    n1192,
    n1226
  );


  or
  g1274
  (
    n1303,
    n1218,
    n1219,
    n1220,
    n1275
  );


  or
  g1275
  (
    n1281,
    n1278,
    n1224,
    n1280,
    n1276
  );


  nor
  g1276
  (
    n1295,
    n1274,
    n1280,
    n1223,
    n1193
  );


  and
  g1277
  (
    n1305,
    n1274,
    n1279,
    n1273
  );


  nand
  g1278
  (
    n1289,
    n1280,
    n1275,
    n1220,
    n1225
  );


  xor
  g1279
  (
    n1297,
    n1193,
    n1223
  );


  xor
  g1280
  (
    n1308,
    n1278,
    n1225,
    n1219
  );


  nor
  g1281
  (
    n1302,
    n1218,
    n1224,
    n1277,
    n1274
  );


  xnor
  g1282
  (
    KeyWire_0_20,
    n1217,
    n1193,
    n1226,
    n1279
  );


  and
  g1283
  (
    n1318,
    n1211,
    n1210,
    n1207
  );


  xnor
  g1284
  (
    n1316,
    n1281,
    n1210,
    n1208,
    n1213
  );


  nor
  g1285
  (
    n1320,
    n1209,
    n1213,
    n1282,
    n1208
  );


  xnor
  g1286
  (
    n1319,
    n1208,
    n1209,
    n1212,
    n1281
  );


  nor
  g1287
  (
    n1317,
    n1281,
    n1209,
    n1282
  );


  and
  g1288
  (
    n1313,
    n1212,
    n1212,
    n1211,
    n1282
  );


  nor
  g1289
  (
    n1315,
    n1208,
    n1281,
    n1212,
    n1282
  );


  nand
  g1290
  (
    n1321,
    n1210,
    n1211,
    n1207
  );


  xnor
  g1291
  (
    n1314,
    n1211,
    n1213,
    n1283
  );


  xor
  g1292
  (
    n1330,
    n1287,
    n1288,
    n1290
  );


  nand
  g1293
  (
    n1326,
    n1319,
    n1285,
    n1258
  );


  and
  g1294
  (
    n1334,
    n1318,
    n1321,
    n1288
  );


  or
  g1295
  (
    n1322,
    n1289,
    n1286,
    n1292
  );


  nor
  g1296
  (
    n1337,
    n1290,
    n1315,
    n1285
  );


  xnor
  g1297
  (
    n1333,
    n1285,
    n1318
  );


  nand
  g1298
  (
    n1342,
    n1284,
    n1321,
    n1318
  );


  or
  g1299
  (
    n1339,
    n1259,
    n1295,
    n1289
  );


  xnor
  g1300
  (
    n1338,
    n1291,
    n1289,
    n1317
  );


  xnor
  g1301
  (
    n1323,
    n1317,
    n1290,
    n1289
  );


  xor
  g1302
  (
    n1341,
    n1293,
    n1294,
    n1259
  );


  nand
  g1303
  (
    n1343,
    n1258,
    n1286,
    n1291
  );


  or
  g1304
  (
    n1340,
    n1317,
    n1293,
    n1316,
    n1319
  );


  or
  g1305
  (
    n1331,
    n1320,
    n1259,
    n1292,
    n1286
  );


  xor
  g1306
  (
    n1335,
    n1292,
    n1320,
    n1293,
    n1258
  );


  nand
  g1307
  (
    n1329,
    n1294,
    n1287,
    n1258,
    n1286
  );


  xor
  g1308
  (
    n1345,
    n1291,
    n1320,
    n1319
  );


  and
  g1309
  (
    n1336,
    n1295,
    n1288,
    n1287,
    n1313
  );


  nand
  g1310
  (
    n1328,
    n1321,
    n1319,
    n1287,
    n1292
  );


  nor
  g1311
  (
    n1325,
    n1283,
    n1284,
    n1291
  );


  nand
  g1312
  (
    n1324,
    n1294,
    n1283,
    n1295,
    n1257
  );


  or
  g1313
  (
    n1344,
    n1314,
    n1288,
    n1290,
    n1259
  );


  nor
  g1314
  (
    n1327,
    n1321,
    n1284,
    n1295,
    n1283
  );


  xnor
  g1315
  (
    n1332,
    n1285,
    n1317,
    n1293,
    n1294
  );


  buf
  g1316
  (
    n1350,
    n1299
  );


  buf
  g1317
  (
    n1365,
    n1298
  );


  not
  g1318
  (
    n1349,
    n1324
  );


  not
  g1319
  (
    n1364,
    n1300
  );


  buf
  g1320
  (
    n1352,
    n1296
  );


  buf
  g1321
  (
    n1346,
    n1323
  );


  buf
  g1322
  (
    n1354,
    n1299
  );


  not
  g1323
  (
    n1363,
    n1300
  );


  buf
  g1324
  (
    n1348,
    n1324
  );


  not
  g1325
  (
    n1347,
    n1298
  );


  not
  g1326
  (
    n1362,
    n1300
  );


  buf
  g1327
  (
    n1358,
    n1323
  );


  nor
  g1328
  (
    n1360,
    n1323,
    n1296,
    n1297
  );


  and
  g1329
  (
    n1356,
    n1298,
    n1322,
    n1301,
    n1325
  );


  or
  g1330
  (
    n1355,
    n1322,
    n1301,
    n1323,
    n1297
  );


  xnor
  g1331
  (
    n1361,
    n1325,
    n1324,
    n1298
  );


  and
  g1332
  (
    n1357,
    n1299,
    n1297,
    n1301
  );


  and
  g1333
  (
    n1353,
    n1325,
    n1296,
    n1326
  );


  and
  g1334
  (
    n1359,
    n1326,
    n1299,
    n1322
  );


  nand
  g1335
  (
    n1351,
    n1325,
    n1326,
    n1296,
    n1300
  );


  buf
  g1336
  (
    n1403,
    n1360
  );


  buf
  g1337
  (
    n1412,
    n1365
  );


  xor
  g1338
  (
    n1406,
    n1349,
    n1351,
    n1305,
    n1333
  );


  and
  g1339
  (
    n1398,
    n1360,
    n1361,
    n1352,
    n1345
  );


  xnor
  g1340
  (
    n1370,
    n1260,
    n1339,
    n1328,
    n1360
  );


  xnor
  g1341
  (
    n1407,
    n1343,
    n1341,
    n1260,
    n1338
  );


  nor
  g1342
  (
    n1372,
    n1355,
    n1344,
    n1358,
    n1331
  );


  nand
  g1343
  (
    n1404,
    n1311,
    n1339,
    n1345,
    n1338
  );


  xnor
  g1344
  (
    n1383,
    n1346,
    n1327,
    n1350,
    n1337
  );


  nand
  g1345
  (
    n1419,
    n1248,
    n1363,
    n1350
  );


  xnor
  g1346
  (
    n1413,
    n1332,
    n1334,
    n1359,
    n1340
  );


  xor
  g1347
  (
    n1369,
    n1337,
    n1303,
    n1309,
    n1356
  );


  and
  g1348
  (
    n1385,
    n1264,
    n1353,
    n1333,
    n1334
  );


  and
  g1349
  (
    n1401,
    n1336,
    n1355,
    n1352,
    n1306
  );


  xor
  g1350
  (
    n1405,
    n1308,
    n1304,
    n1344,
    n1361
  );


  nand
  g1351
  (
    n1381,
    n1335,
    n1311,
    n1302,
    n1308
  );


  nand
  g1352
  (
    n1402,
    n1312,
    n1338,
    n1305,
    n1362
  );


  xnor
  g1353
  (
    n1422,
    n1330,
    n1351,
    n1346,
    n1340
  );


  nand
  g1354
  (
    n1387,
    n1312,
    n1364,
    n1357,
    n1365
  );


  xor
  g1355
  (
    n1418,
    n1336,
    n1303,
    n1247,
    n1329
  );


  xor
  g1356
  (
    n1392,
    n1365,
    n1341,
    n1329,
    n1362
  );


  nor
  g1357
  (
    n1371,
    n1312,
    n1303,
    n1348,
    n1248
  );


  or
  g1358
  (
    n1420,
    n1307,
    n1269,
    n1331,
    n1356
  );


  xnor
  g1359
  (
    n1416,
    n1348,
    n1359,
    n1307,
    n1328
  );


  nor
  g1360
  (
    n1374,
    n1302,
    n1334,
    n1328,
    n1356
  );


  nand
  g1361
  (
    n1397,
    n1357,
    n1327,
    n1338,
    n1358
  );


  xor
  g1362
  (
    n1379,
    n1260,
    n1359,
    n1311,
    n1363
  );


  or
  g1363
  (
    n1414,
    n1352,
    n1348,
    n1330,
    n1354
  );


  xor
  g1364
  (
    n1373,
    n1352,
    n1346,
    n1265,
    n1343
  );


  xor
  g1365
  (
    n1417,
    n1337,
    n1304,
    n1309,
    n1248
  );


  xor
  g1366
  (
    n1399,
    n1339,
    n1246,
    n1341,
    n1356
  );


  xor
  g1367
  (
    n1368,
    n1342,
    n1345,
    n1330,
    n1340
  );


  or
  g1368
  (
    n1386,
    n1350,
    n1335,
    n1332,
    n1329
  );


  xnor
  g1369
  (
    n1394,
    n1305,
    n1332,
    n1247,
    n1364
  );


  nor
  g1370
  (
    n1393,
    n1334,
    n1342,
    n1362,
    n1330
  );


  or
  g1371
  (
    n1367,
    n1364,
    n1361,
    n1349,
    n1351
  );


  xnor
  g1372
  (
    KeyWire_0_3,
    n1347,
    n1328,
    n1353,
    n1346
  );


  xnor
  g1373
  (
    n1400,
    n1357,
    n1303,
    n1310,
    n1347
  );


  xnor
  g1374
  (
    n1410,
    n1355,
    n1306,
    n1263
  );


  or
  g1375
  (
    n1378,
    n1247,
    n1308,
    n1358,
    n1361
  );


  and
  g1376
  (
    n1376,
    n1339,
    n1266,
    n1363,
    n1359
  );


  nand
  g1377
  (
    n1421,
    n1312,
    n1336,
    n1332,
    n1335
  );


  or
  g1378
  (
    n1380,
    n1268,
    n1267,
    n1343,
    n1246
  );


  xnor
  g1379
  (
    n1377,
    n1353,
    n1354,
    n1349,
    n1345
  );


  nor
  g1380
  (
    n1388,
    n1343,
    n1341,
    n1308,
    n1342
  );


  xnor
  g1381
  (
    n1391,
    n1340,
    n1307,
    n1329,
    n1348
  );


  xor
  g1382
  (
    n1390,
    n1351,
    n1309,
    n1355,
    n1302
  );


  xnor
  g1383
  (
    n1375,
    n1304,
    n1310,
    n1247,
    n1347
  );


  xor
  g1384
  (
    n1366,
    n1336,
    n1358,
    n1353,
    n1365
  );


  or
  g1385
  (
    n1395,
    n1362,
    n1309,
    n1305,
    n1333
  );


  xnor
  g1386
  (
    n1389,
    n1270,
    n1342,
    n1360,
    n1347
  );


  and
  g1387
  (
    n1384,
    n1304,
    n1357,
    n1248,
    n1333
  );


  nand
  g1388
  (
    KeyWire_0_21,
    n1311,
    n1335,
    n1306,
    n1327
  );


  xnor
  g1389
  (
    n1415,
    n1349,
    n1364,
    n1354,
    n1363
  );


  or
  g1390
  (
    n1396,
    n1327,
    n1354,
    n1307,
    n1344
  );


  xor
  g1391
  (
    n1411,
    n1331,
    n1310,
    n1337
  );


  xnor
  g1392
  (
    n1382,
    n1331,
    n1302,
    n1260,
    n1344
  );


  or
  g1393
  (
    n1442,
    n1375,
    n1378,
    n1395,
    n1393
  );


  xor
  g1394
  (
    n1429,
    n1387,
    n1390,
    n1386,
    n1369
  );


  or
  g1395
  (
    n1426,
    n1382,
    n1389,
    n1386,
    n1366
  );


  and
  g1396
  (
    n1436,
    n1390,
    n1384,
    n1394
  );


  xor
  g1397
  (
    n1435,
    n1384,
    n1379,
    n1391
  );


  nand
  g1398
  (
    n1423,
    n1381,
    n1383,
    n1388,
    n1393
  );


  xnor
  g1399
  (
    n1428,
    n1386,
    n1382,
    n1380,
    n1383
  );


  and
  g1400
  (
    n1431,
    n1384,
    n1373,
    n1389
  );


  nand
  g1401
  (
    n1424,
    n1389,
    n1388,
    n1387,
    n1379
  );


  nor
  g1402
  (
    n1430,
    n1383,
    n1386,
    n1391,
    n1390
  );


  xnor
  g1403
  (
    KeyWire_0_2,
    n1367,
    n1372,
    n1381,
    n1377
  );


  xor
  g1404
  (
    n1427,
    n1385,
    n1390,
    n1376,
    n1395
  );


  xor
  g1405
  (
    n1440,
    n1387,
    n1393,
    n1379,
    n1382
  );


  or
  g1406
  (
    n1432,
    n1394,
    n1385,
    n1392,
    n1391
  );


  nor
  g1407
  (
    n1438,
    n1388,
    n1383,
    n1380,
    n1381
  );


  xnor
  g1408
  (
    n1437,
    n1394,
    n1380,
    n1381,
    n1391
  );


  or
  g1409
  (
    n1433,
    n1382,
    n1393,
    n1392,
    n1371
  );


  nand
  g1410
  (
    n1425,
    n1387,
    n1392,
    n1394
  );


  xnor
  g1411
  (
    n1434,
    n1380,
    n1370,
    n1368,
    n1388
  );


  and
  g1412
  (
    n1439,
    n1385,
    n1385,
    n1395,
    n1374
  );


  buf
  g1413
  (
    n1443,
    n1427
  );


  buf
  g1414
  (
    n1448,
    n1429
  );


  not
  g1415
  (
    n1445,
    n1428
  );


  not
  g1416
  (
    n1449,
    n1423
  );


  not
  g1417
  (
    n1446,
    n1425
  );


  not
  g1418
  (
    n1450,
    n1426
  );


  not
  g1419
  (
    n1447,
    n1430
  );


  buf
  g1420
  (
    n1444,
    n1424
  );


  or
  g1421
  (
    n1467,
    n1402,
    n1410,
    n1448,
    n1443
  );


  xnor
  g1422
  (
    n1461,
    n1399,
    n1408,
    n1402,
    n1406
  );


  xor
  g1423
  (
    n1475,
    n1417,
    n1405,
    n1446,
    n1412
  );


  xor
  g1424
  (
    n1454,
    n1447,
    n1399,
    n1417,
    n1402
  );


  xnor
  g1425
  (
    n1482,
    n1396,
    n1445,
    n1408,
    n1409
  );


  xor
  g1426
  (
    n1472,
    n1404,
    n1412,
    n1400,
    n1406
  );


  nand
  g1427
  (
    n1451,
    n1443,
    n1418,
    n1398,
    n1401
  );


  nor
  g1428
  (
    n1477,
    n1450,
    n1450,
    n1448,
    n1418
  );


  or
  g1429
  (
    n1473,
    n1413,
    n1414,
    n1410,
    n1403
  );


  and
  g1430
  (
    n1466,
    n1412,
    n1449,
    n1409,
    n1404
  );


  xnor
  g1431
  (
    n1460,
    n1404,
    n1398,
    n1414,
    n1445
  );


  or
  g1432
  (
    n1479,
    n1415,
    n1413,
    n1400,
    n1406
  );


  xnor
  g1433
  (
    n1458,
    n1447,
    n1405,
    n1411,
    n1396
  );


  nor
  g1434
  (
    n1455,
    n1407,
    n1417,
    n1410,
    n1448
  );


  nand
  g1435
  (
    n1452,
    n1398,
    n1416,
    n1415,
    n1413
  );


  nor
  g1436
  (
    n1470,
    n1400,
    n1444,
    n1409,
    n1449
  );


  and
  g1437
  (
    n1471,
    n1395,
    n1416,
    n1409
  );


  nor
  g1438
  (
    n1457,
    n1406,
    n1399,
    n1405,
    n1397
  );


  or
  g1439
  (
    n1456,
    n1408,
    n1446,
    n1444,
    n1396
  );


  nor
  g1440
  (
    n1459,
    n1419,
    n1400,
    n1402,
    n1446
  );


  nor
  g1441
  (
    n1462,
    n1417,
    n1419,
    n1407
  );


  and
  g1442
  (
    KeyWire_0_7,
    n1446,
    n1408,
    n1401,
    n1403
  );


  nor
  g1443
  (
    n1463,
    n1411,
    n1416,
    n1405,
    n1397
  );


  xor
  g1444
  (
    n1469,
    n1447,
    n1448,
    n1398,
    n1415
  );


  nand
  g1445
  (
    n1480,
    n1413,
    n1444,
    n1450,
    n1445
  );


  or
  g1446
  (
    n1465,
    n1415,
    n1450,
    n1443,
    n1411
  );


  nand
  g1447
  (
    n1481,
    n1447,
    n1401,
    n1410,
    n1449
  );


  xor
  g1448
  (
    n1453,
    n1397,
    n1407,
    n1449,
    n1443
  );


  nand
  g1449
  (
    n1468,
    n1396,
    n1403,
    n1414,
    n1401
  );


  nand
  g1450
  (
    n1478,
    n1418,
    n1399,
    n1444,
    n1412
  );


  nor
  g1451
  (
    n1464,
    n1403,
    n1414,
    n1411,
    n1407
  );


  or
  g1452
  (
    n1476,
    n1404,
    n1445,
    n1397,
    n1418
  );


  nand
  g1453
  (
    n1489,
    n1436,
    n1452,
    n1440,
    n1451
  );


  or
  g1454
  (
    n1483,
    n1433,
    n1451,
    n1438,
    n1441
  );


  nand
  g1455
  (
    n1484,
    n1437,
    n1439,
    n1442
  );


  and
  g1456
  (
    n1485,
    n1439,
    n1442,
    n1451,
    n1431
  );


  or
  g1457
  (
    n1490,
    n1441,
    n1440,
    n1432
  );


  nor
  g1458
  (
    n1488,
    n1435,
    n1442,
    n1439,
    n1452
  );


  nand
  g1459
  (
    n1487,
    n1452,
    n1441,
    n1440,
    n1442
  );


  and
  g1460
  (
    n1486,
    n1451,
    n1434,
    n1452,
    n1441
  );


  buf
  g1461
  (
    n1492,
    n1483
  );


  not
  g1462
  (
    n1498,
    n1453
  );


  buf
  g1463
  (
    n1494,
    n1453
  );


  not
  g1464
  (
    n1495,
    n1488
  );


  not
  g1465
  (
    n1496,
    n1453
  );


  xnor
  g1466
  (
    n1497,
    n1454,
    n1486,
    n1487
  );


  nor
  g1467
  (
    n1493,
    n1453,
    n1454,
    n1485
  );


  nand
  g1468
  (
    KeyWire_0_25,
    n1490,
    n1454,
    n1489,
    n1484
  );


  or
  g1469
  (
    n1499,
    n1464,
    n1461,
    n1465,
    n1468
  );


  xor
  g1470
  (
    n1510,
    n1469,
    n1457,
    n1475
  );


  xnor
  g1471
  (
    n1513,
    n1498,
    n1422,
    n1497,
    n1463
  );


  and
  g1472
  (
    KeyWire_0_1,
    n1474,
    n1473,
    n1496,
    n1493
  );


  nand
  g1473
  (
    n1512,
    n1422,
    n1456,
    n1419,
    n1462
  );


  nand
  g1474
  (
    n1523,
    n1455,
    n1457,
    n1492,
    n1464
  );


  and
  g1475
  (
    n1504,
    n1471,
    n1464,
    n1461,
    n1468
  );


  nand
  g1476
  (
    n1503,
    n1460,
    n1468,
    n1470,
    n1461
  );


  and
  g1477
  (
    n1501,
    n1460,
    n1473,
    n1469,
    n1466
  );


  nand
  g1478
  (
    n1506,
    n1496,
    n1467,
    n1471,
    n1462
  );


  xnor
  g1479
  (
    n1502,
    n1468,
    n1420,
    n1459,
    n1457
  );


  xor
  g1480
  (
    n1516,
    n1463,
    n1421,
    n1496,
    n1469
  );


  xor
  g1481
  (
    n1525,
    n1461,
    n1422,
    n1467,
    n1492
  );


  nor
  g1482
  (
    n1524,
    n1495,
    n1462,
    n1466,
    n1491
  );


  and
  g1483
  (
    n1511,
    n1460,
    n1494,
    n1422,
    n1469
  );


  nand
  g1484
  (
    n1518,
    n1470,
    n1462,
    n1472,
    n1456
  );


  or
  g1485
  (
    n1530,
    n1474,
    n1491,
    n1472,
    n1464
  );


  or
  g1486
  (
    n1520,
    n1467,
    n1494,
    n1498,
    n1456
  );


  nor
  g1487
  (
    n1505,
    n1495,
    n1421,
    n1498,
    n1459
  );


  or
  g1488
  (
    n1527,
    n1459,
    n1475,
    n1497,
    n1456
  );


  and
  g1489
  (
    n1509,
    n1475,
    n1491,
    n1420,
    n1458
  );


  or
  g1490
  (
    n1507,
    n1494,
    n1455,
    n1493,
    n1497
  );


  nor
  g1491
  (
    n1517,
    n1420,
    n1492,
    n1455
  );


  and
  g1492
  (
    n1508,
    n1496,
    n1498,
    n1491,
    n1420
  );


  xor
  g1493
  (
    n1515,
    n1495,
    n1455,
    n1473
  );


  nor
  g1494
  (
    n1528,
    n1458,
    n1495,
    n1474,
    n1493
  );


  xnor
  g1495
  (
    n1529,
    n1459,
    n1465,
    n1497
  );


  and
  g1496
  (
    n1519,
    n1470,
    n1472,
    n1474,
    n1458
  );


  nand
  g1497
  (
    n1514,
    n1421,
    n1421,
    n1466,
    n1463
  );


  xor
  g1498
  (
    n1500,
    n1466,
    n1471,
    n1467
  );


  and
  g1499
  (
    n1526,
    n1493,
    n1458,
    n1472,
    n1465
  );


  xor
  g1500
  (
    n1522,
    n1470,
    n1463,
    n1494,
    n1460
  );


  buf
  g1501
  (
    n1532,
    n1499
  );


  buf
  g1502
  (
    n1531,
    n1500
  );


  buf
  g1503
  (
    n1533,
    n1501
  );


  nand
  g1504
  (
    n1537,
    n1503,
    n1508,
    n1533,
    n1512
  );


  xnor
  g1505
  (
    n1542,
    n1533,
    n1532,
    n1507
  );


  and
  g1506
  (
    n1541,
    n1509,
    n1532,
    n1531,
    n1511
  );


  xor
  g1507
  (
    KeyWire_0_28,
    n1513,
    n1510,
    n1512
  );


  xnor
  g1508
  (
    n1536,
    n1510,
    n1506,
    n1513,
    n1504
  );


  xnor
  g1509
  (
    KeyWire_0_11,
    n1531,
    n1509,
    n1513,
    n1533
  );


  or
  g1510
  (
    n1539,
    n1509,
    n1511
  );


  nor
  g1511
  (
    n1535,
    n1502,
    n1512,
    n1533,
    n1513
  );


  or
  g1512
  (
    n1534,
    n1509,
    n1512,
    n1505,
    n1510
  );


  nor
  g1513
  (
    n1548,
    n1518,
    n1534,
    n1514,
    n1515
  );


  xnor
  g1514
  (
    n1547,
    n1517,
    n1516,
    n1515
  );


  xor
  g1515
  (
    n1544,
    n1514,
    n1538,
    n1535,
    n1519
  );


  xor
  g1516
  (
    n1549,
    n1537,
    n1514,
    n1517,
    n1518
  );


  xor
  g1517
  (
    n1546,
    n1515,
    n1516,
    n1518,
    n1517
  );


  xnor
  g1518
  (
    n1543,
    n1517,
    n1515,
    n1540,
    n1514
  );


  or
  g1519
  (
    n1545,
    n1518,
    n1536,
    n1516,
    n1539
  );


  and
  g1520
  (
    n1554,
    n1478,
    n1544,
    n1476,
    n1480
  );


  or
  g1521
  (
    n1550,
    n1477,
    n1475,
    n1476,
    n1481
  );


  xnor
  g1522
  (
    n1553,
    n1477,
    n1480,
    n1476
  );


  and
  g1523
  (
    n1559,
    n1481,
    n1482,
    n1545
  );


  xor
  g1524
  (
    n1551,
    n1543,
    n1482,
    n1477,
    n1545
  );


  nand
  g1525
  (
    n1557,
    n1543,
    n1480,
    n1477,
    n1481
  );


  or
  g1526
  (
    n1552,
    n1479,
    n1478,
    n1544
  );


  or
  g1527
  (
    n1556,
    n1544,
    n1543,
    n1478,
    n1479
  );


  xnor
  g1528
  (
    n1558,
    n1478,
    n1482,
    n1543,
    n1476
  );


  or
  g1529
  (
    n1555,
    n1479,
    n1479,
    n1481,
    n1545
  );


  nor
  g1530
  (
    n1563,
    n1519,
    n1547,
    n1558
  );


  and
  g1531
  (
    n1561,
    n1557,
    n1546,
    n1556,
    n1519
  );


  xnor
  g1532
  (
    n1562,
    n1547,
    n1520,
    n1546
  );


  nor
  g1533
  (
    n1560,
    n1559,
    n1546,
    n1519,
    n1545
  );


  or
  g1534
  (
    n1566,
    n1563,
    n1561,
    n1522
  );


  nor
  g1535
  (
    n1564,
    n1523,
    n1521,
    n1522
  );


  xor
  g1536
  (
    n1567,
    n1520,
    n1521,
    n1523,
    n1522
  );


  nor
  g1537
  (
    n1565,
    n1562,
    n1520,
    n1523
  );


  and
  g1538
  (
    n1568,
    n1523,
    n1563,
    n1521,
    n1560
  );


  buf
  g1539
  (
    n1569,
    n1564
  );


  and
  g1540
  (
    n1570,
    n1565,
    n1524
  );


  and
  g1541
  (
    n1573,
    n1525,
    n1567,
    n1542
  );


  or
  g1542
  (
    n1571,
    n1525,
    n1570,
    n1542
  );


  nand
  g1543
  (
    n1572,
    n1541,
    n1566,
    n1542,
    n1568
  );


  nor
  g1544
  (
    n1574,
    n1542,
    n1524,
    n1569,
    n1541
  );


  nor
  g1545
  (
    n1575,
    n1541,
    n1570
  );


  xor
  g1546
  (
    n1577,
    n1528,
    n1526
  );


  xnor
  g1547
  (
    n1579,
    n1528,
    n1571,
    n1527
  );


  or
  g1548
  (
    n1578,
    n1525,
    n1527,
    n1526
  );


  or
  g1549
  (
    n1576,
    n1571,
    n1571,
    n1525,
    n1527
  );


  xor
  g1550
  (
    n1582,
    n1579,
    n1578,
    n1528,
    n1530
  );


  nand
  g1551
  (
    n1583,
    n1577,
    n546,
    n1529
  );


  and
  g1552
  (
    n1580,
    n547,
    n1530,
    n1579,
    n546
  );


  nor
  g1553
  (
    n1584,
    n1579,
    n546,
    n1530,
    n545
  );


  xnor
  g1554
  (
    n1585,
    n545,
    n1530,
    n1579,
    n1529
  );


  xor
  g1555
  (
    n1581,
    n1528,
    n547,
    n1529,
    n546
  );


  xnor
  g1556
  (
    n1597,
    n1584,
    n1572,
    n549,
    n554
  );


  nor
  g1557
  (
    n1587,
    n1584,
    n555,
    n548,
    n552
  );


  xnor
  g1558
  (
    n1595,
    n550,
    n1575,
    n1572,
    n551
  );


  xnor
  g1559
  (
    n1606,
    n1573,
    n561,
    n556,
    n550
  );


  xor
  g1560
  (
    n1598,
    n556,
    n1573
  );


  nand
  g1561
  (
    n1590,
    n551,
    n1574,
    n553,
    n557
  );


  xor
  g1562
  (
    n1603,
    n550,
    n551,
    n555,
    n548
  );


  xor
  g1563
  (
    n1594,
    n1580,
    n1575,
    n559,
    n1581
  );


  xor
  g1564
  (
    n1596,
    n552,
    n559,
    n1584,
    n1583
  );


  xor
  g1565
  (
    n1605,
    n553,
    n549,
    n1580,
    n555
  );


  xnor
  g1566
  (
    n1604,
    n1575,
    n558,
    n1581,
    n1585
  );


  or
  g1567
  (
    n1609,
    n556,
    n549,
    n559
  );


  and
  g1568
  (
    n1586,
    n1580,
    n553,
    n547,
    n548
  );


  xor
  g1569
  (
    n1593,
    n560,
    n547,
    n1585,
    n553
  );


  or
  g1570
  (
    n1592,
    n552,
    n554,
    n1574,
    n1582
  );


  nand
  g1571
  (
    n1588,
    n1581,
    n1582,
    n554,
    n560
  );


  nand
  g1572
  (
    n1600,
    n1572,
    n554,
    n1584,
    n1582
  );


  xor
  g1573
  (
    n1602,
    n1575,
    n557,
    n558
  );


  xor
  g1574
  (
    n1608,
    n550,
    n1582,
    n1583,
    n556
  );


  nand
  g1575
  (
    n1599,
    n552,
    n1581,
    n560,
    n1583
  );


  nor
  g1576
  (
    n1589,
    n548,
    n1572,
    n1580,
    n557
  );


  nor
  g1577
  (
    n1601,
    n551,
    n1574,
    n1585,
    n1583
  );


  and
  g1578
  (
    n1607,
    n559,
    n555,
    n1585,
    n557
  );


  or
  g1579
  (
    n1591,
    n561,
    n560,
    n1574,
    n558
  );


  or
  g1580
  (
    n1615,
    n562,
    n1600,
    n580,
    n564
  );


  xnor
  g1581
  (
    n1614,
    n579,
    n1603,
    n577,
    n575
  );


  nor
  g1582
  (
    n1611,
    n562,
    n579,
    n1599,
    n1601
  );


  xnor
  g1583
  (
    n1618,
    n579,
    n1548,
    n1601
  );


  nor
  g1584
  (
    n1631,
    n568,
    n570,
    n561
  );


  xnor
  g1585
  (
    n1612,
    n567,
    n569,
    n574,
    n576
  );


  or
  g1586
  (
    n1636,
    n1549,
    n574,
    n576,
    n1602
  );


  and
  g1587
  (
    n1633,
    n573,
    n578,
    n565,
    n561
  );


  nor
  g1588
  (
    KeyWire_0_5,
    n562,
    n580,
    n570
  );


  nand
  g1589
  (
    n1624,
    n569,
    n1603,
    n1547
  );


  xnor
  g1590
  (
    n1635,
    n1598,
    n1594,
    n575,
    n564
  );


  xor
  g1591
  (
    n1634,
    n572,
    n1589,
    n1600,
    n1586
  );


  and
  g1592
  (
    n1616,
    n565,
    n567,
    n571,
    n566
  );


  xnor
  g1593
  (
    n1629,
    n571,
    n1600,
    n1601,
    n1593
  );


  nor
  g1594
  (
    n1630,
    n1602,
    n571,
    n568,
    n580
  );


  nor
  g1595
  (
    n1617,
    n577,
    n568,
    n565,
    n567
  );


  xnor
  g1596
  (
    n1622,
    n1587,
    n572,
    n1549,
    n563
  );


  and
  g1597
  (
    n1627,
    n1588,
    n573,
    n1597
  );


  nand
  g1598
  (
    n1620,
    n578,
    n1591,
    n1600,
    n570
  );


  and
  g1599
  (
    n1610,
    n1549,
    n576,
    n577,
    n565
  );


  or
  g1600
  (
    KeyWire_0_24,
    n566,
    n571,
    n569,
    n1548
  );


  xor
  g1601
  (
    n1628,
    n573,
    n574,
    n578,
    n572
  );


  nand
  g1602
  (
    n1619,
    n563,
    n575,
    n567,
    n1601
  );


  or
  g1603
  (
    n1613,
    n568,
    n574,
    n564,
    n1602
  );


  xnor
  g1604
  (
    n1623,
    n1595,
    n1602,
    n577,
    n1590
  );


  xnor
  g1605
  (
    n1621,
    n576,
    n563,
    n562,
    n566
  );


  and
  g1606
  (
    n1638,
    n1549,
    n575,
    n563,
    n1596
  );


  nor
  g1607
  (
    n1625,
    n564,
    n578,
    n569,
    n579
  );


  nand
  g1608
  (
    n1626,
    n1548,
    n572,
    n566,
    n1592
  );


  nor
  g1609
  (
    n1654,
    n586,
    n1620
  );


  and
  g1610
  (
    n1641,
    n591,
    n594,
    n588,
    n1633
  );


  and
  g1611
  (
    n1657,
    n582,
    n592,
    n581
  );


  xnor
  g1612
  (
    n1646,
    n591,
    n1625,
    n593,
    n598
  );


  and
  g1613
  (
    n1658,
    n591,
    n583,
    n587,
    n597
  );


  or
  g1614
  (
    n1648,
    n588,
    n595,
    n1632,
    n586
  );


  and
  g1615
  (
    n1645,
    n584,
    n1623,
    n585,
    n590
  );


  nor
  g1616
  (
    n1644,
    n595,
    n1610,
    n1617,
    n1614
  );


  and
  g1617
  (
    n1660,
    n1630,
    n582,
    n583,
    n1619
  );


  xnor
  g1618
  (
    n1649,
    n589,
    n596,
    n594,
    n1616
  );


  or
  g1619
  (
    n1639,
    n589,
    n592,
    n595,
    n597
  );


  nor
  g1620
  (
    n1642,
    n1611,
    n588,
    n596,
    n581
  );


  xnor
  g1621
  (
    n1651,
    n593,
    n583,
    n1626,
    n1631
  );


  nor
  g1622
  (
    n1643,
    n593,
    n583,
    n590,
    n589
  );


  and
  g1623
  (
    n1653,
    n585,
    n587,
    n1622,
    n584
  );


  or
  g1624
  (
    n1655,
    n1624,
    n595,
    n1612,
    n598
  );


  xnor
  g1625
  (
    n1640,
    n1627,
    n591,
    n587,
    n1621
  );


  xnor
  g1626
  (
    n1662,
    n590,
    n581,
    n594,
    n1628
  );


  or
  g1627
  (
    n1661,
    n594,
    n593,
    n597
  );


  xnor
  g1628
  (
    n1652,
    n581,
    n585,
    n586,
    n1629
  );


  xor
  g1629
  (
    n1650,
    n590,
    n585,
    n586,
    n592
  );


  or
  g1630
  (
    n1656,
    n584,
    n587,
    n596,
    n1613
  );


  or
  g1631
  (
    n1647,
    n582,
    n589,
    n588,
    n1618
  );


  nand
  g1632
  (
    n1659,
    n596,
    n1615,
    n584,
    n582
  );


  xnor
  g1633
  (
    n1695,
    n1608,
    n1660,
    n1645,
    n1609
  );


  or
  g1634
  (
    n1692,
    n1609,
    n1658,
    n1659,
    n1651
  );


  and
  g1635
  (
    n1669,
    n1605,
    n1649,
    n1603,
    n1652
  );


  nand
  g1636
  (
    n1680,
    n1606,
    n1609,
    n1654
  );


  xor
  g1637
  (
    n1690,
    n1660,
    n599,
    n1662
  );


  or
  g1638
  (
    n1685,
    n1641,
    n1640,
    n1655,
    n1661
  );


  xor
  g1639
  (
    n1674,
    n1604,
    n598,
    n1660,
    n1606
  );


  xnor
  g1640
  (
    n1694,
    n1648,
    n1607,
    n1606
  );


  or
  g1641
  (
    n1684,
    n1650,
    n1654,
    n1651,
    n1646
  );


  xnor
  g1642
  (
    n1682,
    n1607,
    n599,
    n1661,
    n1653
  );


  nand
  g1643
  (
    n1673,
    n1650,
    n1639,
    n1642,
    n1649
  );


  and
  g1644
  (
    n1693,
    n1637,
    n1658,
    n1659,
    n1648
  );


  nand
  g1645
  (
    n1688,
    n1653,
    n1635,
    n1655,
    n1647
  );


  nor
  g1646
  (
    n1696,
    n1644,
    n1651,
    n598,
    n1604
  );


  xnor
  g1647
  (
    n1683,
    n600,
    n1662,
    n1644,
    n1650
  );


  xnor
  g1648
  (
    n1665,
    n1657,
    n1654,
    n1655,
    n1605
  );


  xnor
  g1649
  (
    n1671,
    n1656,
    n600,
    n1647,
    n1661
  );


  or
  g1650
  (
    n1681,
    n1646,
    n1643,
    n1605
  );


  nand
  g1651
  (
    n1687,
    n1658,
    n1645,
    n1652,
    n1640
  );


  and
  g1652
  (
    n1678,
    n1639,
    n1649,
    n1648,
    n1662
  );


  nor
  g1653
  (
    n1686,
    n599,
    n1649,
    n1641,
    n1655
  );


  nor
  g1654
  (
    n1663,
    n1646,
    n1656,
    n1644,
    n1150
  );


  nand
  g1655
  (
    n1668,
    n1653,
    n1640,
    n1642,
    n1662
  );


  nor
  g1656
  (
    n1670,
    n1652,
    n1651,
    n1654,
    n1656
  );


  and
  g1657
  (
    n1664,
    n1607,
    n1648,
    n1642,
    n1656
  );


  nand
  g1658
  (
    n1677,
    n1604,
    n1641,
    n1643,
    n1608
  );


  xnor
  g1659
  (
    n1676,
    n1608,
    n1657,
    n1641,
    n1640
  );


  xor
  g1660
  (
    n1689,
    n1657,
    n1645,
    n1642
  );


  nor
  g1661
  (
    n1691,
    n1605,
    n1661,
    n1646,
    n1652
  );


  nor
  g1662
  (
    n1666,
    n1604,
    n1644,
    n1643,
    n600
  );


  nor
  g1663
  (
    n1675,
    n1657,
    n1659,
    n1634,
    n1639
  );


  or
  g1664
  (
    n1672,
    n1647,
    n1647,
    n1658,
    n600
  );


  nor
  g1665
  (
    KeyWire_0_10,
    n1608,
    n1607,
    n1660,
    n1659
  );


  nor
  g1666
  (
    n1679,
    n1653,
    n1636,
    n1650,
    n1639
  );


  buf
  g1667
  (
    n1697,
    n1665
  );


  nand
  g1668
  (
    n1698,
    n1667,
    n1664,
    n1666,
    n1663
  );


  buf
  g1669
  (
    n1699,
    n1697
  );


  buf
  g1670
  (
    n1700,
    n1698
  );


  or
  g1671
  (
    n1705,
    n1673,
    n1681,
    n1677,
    n1674
  );


  xor
  g1672
  (
    n1701,
    n1700,
    n1678,
    n1670,
    n1699
  );


  and
  g1673
  (
    n1703,
    n1700,
    n1669,
    n1682,
    n1680
  );


  or
  g1674
  (
    n1704,
    n1675,
    n1700,
    n1672
  );


  xor
  g1675
  (
    n1702,
    n1676,
    n1671,
    n1668,
    n1679
  );


  nor
  g1676
  (
    n1706,
    n1705,
    n1684,
    n1683,
    n1638
  );


  nand
  g1677
  (
    n1707,
    n1706,
    n1706,
    n1694,
    n1691
  );


  xnor
  g1678
  (
    n1708,
    n1687,
    n1706,
    n1696,
    n1690
  );


  nor
  g1679
  (
    n1710,
    n1706,
    n1686,
    n1689,
    n1685
  );


  and
  g1680
  (
    n1709,
    n1695,
    n1692,
    n1688,
    n1693
  );


  not
  g1681
  (
    n1711,
    n1708
  );


  buf
  g1682
  (
    n1712,
    n1707
  );


  or
  g1683
  (
    n1713,
    n1710,
    n1711,
    n1712,
    n1709
  );


  xor
  KeyGate_0_0
  (
    n589,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1521,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1441,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1409,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n846,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n1632,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n838,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1474,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1045,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1166,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1667,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1538,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n58,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n222,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n39,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n736,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n780,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n37,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1265,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1173,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1310,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1408,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1240,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n441,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1637,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1491,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n697,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n246,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1540,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n185,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n855,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n724,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


