

module Stat_803_2716
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n698,
  n701,
  n689,
  n693,
  n794,
  n830,
  n820,
  n828,
  n819,
  n821,
  n825,
  n824,
  n823,
  n829,
  n827,
  n822,
  n826
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n698;output n701;output n689;output n693;output n794;output n830;output n820;output n828;output n819;output n821;output n825;output n824;output n823;output n829;output n827;output n822;output n826;
  wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n690;wire n691;wire n692;wire n694;wire n695;wire n696;wire n697;wire n699;wire n700;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  not
  g0
  (
    n80,
    n8
  );


  buf
  g1
  (
    n119,
    n16
  );


  not
  g2
  (
    n123,
    n5
  );


  not
  g3
  (
    n74,
    n23
  );


  buf
  g4
  (
    n88,
    n8
  );


  not
  g5
  (
    n77,
    n9
  );


  not
  g6
  (
    n107,
    n12
  );


  not
  g7
  (
    n47,
    n5
  );


  buf
  g8
  (
    n70,
    n18
  );


  buf
  g9
  (
    n65,
    n4
  );


  not
  g10
  (
    n97,
    n3
  );


  not
  g11
  (
    n46,
    n12
  );


  buf
  g12
  (
    n98,
    n6
  );


  buf
  g13
  (
    n109,
    n24
  );


  buf
  g14
  (
    n55,
    n14
  );


  not
  g15
  (
    n35,
    n7
  );


  buf
  g16
  (
    n89,
    n10
  );


  buf
  g17
  (
    n58,
    n2
  );


  buf
  g18
  (
    n45,
    n6
  );


  not
  g19
  (
    KeyWire_0_17,
    n22
  );


  not
  g20
  (
    n39,
    n2
  );


  buf
  g21
  (
    n76,
    n21
  );


  buf
  g22
  (
    n108,
    n8
  );


  not
  g23
  (
    KeyWire_0_62,
    n6
  );


  not
  g24
  (
    n53,
    n14
  );


  not
  g25
  (
    n103,
    n15
  );


  buf
  g26
  (
    n106,
    n14
  );


  buf
  g27
  (
    n44,
    n2
  );


  not
  g28
  (
    n82,
    n6
  );


  not
  g29
  (
    n68,
    n10
  );


  buf
  g30
  (
    n41,
    n1
  );


  buf
  g31
  (
    n50,
    n11
  );


  not
  g32
  (
    n96,
    n13
  );


  not
  g33
  (
    n36,
    n7
  );


  not
  g34
  (
    n59,
    n10
  );


  not
  g35
  (
    n75,
    n13
  );


  not
  g36
  (
    n126,
    n22
  );


  not
  g37
  (
    n85,
    n25
  );


  not
  g38
  (
    n64,
    n16
  );


  buf
  g39
  (
    KeyWire_0_20,
    n17
  );


  not
  g40
  (
    n118,
    n9
  );


  buf
  g41
  (
    KeyWire_0_32,
    n15
  );


  not
  g42
  (
    n81,
    n23
  );


  buf
  g43
  (
    n51,
    n21
  );


  buf
  g44
  (
    n124,
    n12
  );


  not
  g45
  (
    n69,
    n18
  );


  not
  g46
  (
    n56,
    n24
  );


  buf
  g47
  (
    n60,
    n12
  );


  buf
  g48
  (
    n113,
    n2
  );


  not
  g49
  (
    n62,
    n23
  );


  buf
  g50
  (
    n94,
    n19
  );


  buf
  g51
  (
    n30,
    n1
  );


  not
  g52
  (
    KeyWire_0_22,
    n21
  );


  buf
  g53
  (
    n48,
    n20
  );


  not
  g54
  (
    n117,
    n4
  );


  buf
  g55
  (
    KeyWire_0_15,
    n10
  );


  buf
  g56
  (
    n105,
    n1
  );


  not
  g57
  (
    n66,
    n13
  );


  not
  g58
  (
    n52,
    n20
  );


  not
  g59
  (
    n57,
    n4
  );


  buf
  g60
  (
    n91,
    n17
  );


  buf
  g61
  (
    n61,
    n4
  );


  buf
  g62
  (
    n84,
    n19
  );


  buf
  g63
  (
    n54,
    n13
  );


  not
  g64
  (
    KeyWire_0_26,
    n16
  );


  buf
  g65
  (
    n125,
    n17
  );


  buf
  g66
  (
    n33,
    n7
  );


  buf
  g67
  (
    n42,
    n7
  );


  buf
  g68
  (
    n86,
    n9
  );


  not
  g69
  (
    n83,
    n18
  );


  not
  g70
  (
    n40,
    n3
  );


  not
  g71
  (
    n31,
    n5
  );


  buf
  g72
  (
    n73,
    n19
  );


  buf
  g73
  (
    n95,
    n3
  );


  buf
  g74
  (
    n90,
    n11
  );


  not
  g75
  (
    n122,
    n20
  );


  buf
  g76
  (
    KeyWire_0_16,
    n25
  );


  not
  g77
  (
    KeyWire_0_21,
    n15
  );


  buf
  g78
  (
    KeyWire_0_52,
    n19
  );


  not
  g79
  (
    n34,
    n17
  );


  not
  g80
  (
    n115,
    n8
  );


  not
  g81
  (
    n37,
    n21
  );


  buf
  g82
  (
    KeyWire_0_46,
    n20
  );


  buf
  g83
  (
    n67,
    n15
  );


  not
  g84
  (
    n43,
    n23
  );


  buf
  g85
  (
    n100,
    n11
  );


  buf
  g86
  (
    n72,
    n14
  );


  buf
  g87
  (
    n101,
    n24
  );


  buf
  g88
  (
    KeyWire_0_13,
    n16
  );


  not
  g89
  (
    n99,
    n1
  );


  not
  g90
  (
    KeyWire_0_6,
    n24
  );


  buf
  g91
  (
    n32,
    n9
  );


  not
  g92
  (
    n116,
    n11
  );


  buf
  g93
  (
    KeyWire_0_1,
    n3
  );


  not
  g94
  (
    KeyWire_0_38,
    n5
  );


  not
  g95
  (
    n28,
    n22
  );


  not
  g96
  (
    n79,
    n18
  );


  buf
  g97
  (
    n102,
    n25
  );


  buf
  g98
  (
    n38,
    n22
  );


  buf
  g99
  (
    n169,
    n29
  );


  buf
  g100
  (
    n394,
    n30
  );


  buf
  g101
  (
    n207,
    n43
  );


  buf
  g102
  (
    n349,
    n67
  );


  buf
  g103
  (
    n320,
    n54
  );


  buf
  g104
  (
    n202,
    n50
  );


  buf
  g105
  (
    n257,
    n40
  );


  not
  g106
  (
    n290,
    n55
  );


  not
  g107
  (
    n385,
    n84
  );


  buf
  g108
  (
    n301,
    n89
  );


  not
  g109
  (
    n263,
    n97
  );


  not
  g110
  (
    n162,
    n32
  );


  buf
  g111
  (
    n293,
    n42
  );


  not
  g112
  (
    n152,
    n97
  );


  buf
  g113
  (
    n265,
    n44
  );


  buf
  g114
  (
    n194,
    n40
  );


  not
  g115
  (
    n363,
    n60
  );


  not
  g116
  (
    n333,
    n79
  );


  buf
  g117
  (
    n184,
    n64
  );


  buf
  g118
  (
    n392,
    n96
  );


  not
  g119
  (
    n187,
    n36
  );


  not
  g120
  (
    n221,
    n93
  );


  buf
  g121
  (
    n168,
    n89
  );


  buf
  g122
  (
    n277,
    n38
  );


  not
  g123
  (
    n155,
    n71
  );


  buf
  g124
  (
    KeyWire_0_24,
    n93
  );


  not
  g125
  (
    n241,
    n88
  );


  buf
  g126
  (
    n356,
    n30
  );


  buf
  g127
  (
    n147,
    n82
  );


  buf
  g128
  (
    n315,
    n79
  );


  buf
  g129
  (
    n188,
    n67
  );


  buf
  g130
  (
    n171,
    n72
  );


  not
  g131
  (
    n195,
    n43
  );


  buf
  g132
  (
    n170,
    n59
  );


  buf
  g133
  (
    KeyWire_0_49,
    n38
  );


  buf
  g134
  (
    n179,
    n82
  );


  buf
  g135
  (
    n323,
    n34
  );


  not
  g136
  (
    n208,
    n73
  );


  buf
  g137
  (
    n218,
    n32
  );


  buf
  g138
  (
    n390,
    n68
  );


  not
  g139
  (
    n410,
    n44
  );


  not
  g140
  (
    n236,
    n48
  );


  not
  g141
  (
    n283,
    n56
  );


  not
  g142
  (
    n159,
    n76
  );


  not
  g143
  (
    n373,
    n37
  );


  buf
  g144
  (
    KeyWire_0_44,
    n29
  );


  buf
  g145
  (
    n205,
    n92
  );


  buf
  g146
  (
    n346,
    n31
  );


  buf
  g147
  (
    n369,
    n57
  );


  buf
  g148
  (
    n300,
    n79
  );


  not
  g149
  (
    n381,
    n99
  );


  buf
  g150
  (
    n371,
    n67
  );


  not
  g151
  (
    n364,
    n57
  );


  buf
  g152
  (
    n255,
    n75
  );


  buf
  g153
  (
    n359,
    n60
  );


  not
  g154
  (
    n312,
    n83
  );


  not
  g155
  (
    n294,
    n55
  );


  buf
  g156
  (
    n134,
    n74
  );


  not
  g157
  (
    n271,
    n31
  );


  not
  g158
  (
    n180,
    n42
  );


  buf
  g159
  (
    n299,
    n95
  );


  buf
  g160
  (
    n386,
    n78
  );


  not
  g161
  (
    n302,
    n40
  );


  buf
  g162
  (
    n193,
    n72
  );


  buf
  g163
  (
    n225,
    n80
  );


  not
  g164
  (
    n228,
    n87
  );


  buf
  g165
  (
    n328,
    n54
  );


  buf
  g166
  (
    n166,
    n37
  );


  buf
  g167
  (
    n370,
    n65
  );


  buf
  g168
  (
    n259,
    n57
  );


  not
  g169
  (
    n274,
    n45
  );


  not
  g170
  (
    n230,
    n92
  );


  buf
  g171
  (
    n137,
    n52
  );


  buf
  g172
  (
    n128,
    n99
  );


  not
  g173
  (
    n192,
    n58
  );


  not
  g174
  (
    n148,
    n88
  );


  buf
  g175
  (
    n295,
    n72
  );


  not
  g176
  (
    n181,
    n32
  );


  buf
  g177
  (
    n269,
    n61
  );


  buf
  g178
  (
    n209,
    n30
  );


  not
  g179
  (
    n270,
    n46
  );


  buf
  g180
  (
    n331,
    n40
  );


  buf
  g181
  (
    n150,
    n33
  );


  not
  g182
  (
    n136,
    n94
  );


  not
  g183
  (
    n264,
    n96
  );


  buf
  g184
  (
    n345,
    n69
  );


  not
  g185
  (
    n232,
    n53
  );


  buf
  g186
  (
    n223,
    n88
  );


  buf
  g187
  (
    n324,
    n58
  );


  buf
  g188
  (
    n282,
    n48
  );


  buf
  g189
  (
    n336,
    n62
  );


  buf
  g190
  (
    n178,
    n98
  );


  not
  g191
  (
    n298,
    n69
  );


  not
  g192
  (
    n142,
    n39
  );


  not
  g193
  (
    n332,
    n80
  );


  not
  g194
  (
    n379,
    n78
  );


  buf
  g195
  (
    n201,
    n28
  );


  not
  g196
  (
    n376,
    n73
  );


  not
  g197
  (
    n189,
    n63
  );


  buf
  g198
  (
    n206,
    n35
  );


  buf
  g199
  (
    KeyWire_0_4,
    n66
  );


  buf
  g200
  (
    n297,
    n87
  );


  buf
  g201
  (
    n317,
    n61
  );


  buf
  g202
  (
    n341,
    n87
  );


  buf
  g203
  (
    n243,
    n54
  );


  buf
  g204
  (
    n186,
    n33
  );


  buf
  g205
  (
    n174,
    n67
  );


  buf
  g206
  (
    n337,
    n35
  );


  not
  g207
  (
    n139,
    n49
  );


  not
  g208
  (
    n304,
    n97
  );


  buf
  g209
  (
    n289,
    n29
  );


  buf
  g210
  (
    KeyWire_0_7,
    n86
  );


  buf
  g211
  (
    n260,
    n65
  );


  buf
  g212
  (
    n343,
    n95
  );


  buf
  g213
  (
    n327,
    n77
  );


  not
  g214
  (
    n316,
    n83
  );


  not
  g215
  (
    n211,
    n37
  );


  not
  g216
  (
    n391,
    n32
  );


  buf
  g217
  (
    n130,
    n70
  );


  buf
  g218
  (
    n388,
    n46
  );


  not
  g219
  (
    n144,
    n82
  );


  buf
  g220
  (
    n314,
    n56
  );


  buf
  g221
  (
    n351,
    n91
  );


  buf
  g222
  (
    n262,
    n37
  );


  buf
  g223
  (
    n239,
    n63
  );


  buf
  g224
  (
    n254,
    n92
  );


  buf
  g225
  (
    n272,
    n55
  );


  buf
  g226
  (
    n131,
    n50
  );


  buf
  g227
  (
    KeyWire_0_33,
    n91
  );


  not
  g228
  (
    n368,
    n84
  );


  buf
  g229
  (
    n252,
    n47
  );


  buf
  g230
  (
    n402,
    n96
  );


  not
  g231
  (
    n354,
    n74
  );


  not
  g232
  (
    n309,
    n46
  );


  buf
  g233
  (
    n384,
    n33
  );


  buf
  g234
  (
    n286,
    n77
  );


  not
  g235
  (
    n242,
    n85
  );


  not
  g236
  (
    n375,
    n28
  );


  not
  g237
  (
    n244,
    n63
  );


  buf
  g238
  (
    n352,
    n91
  );


  not
  g239
  (
    n382,
    n47
  );


  buf
  g240
  (
    n220,
    n90
  );


  buf
  g241
  (
    n306,
    n80
  );


  buf
  g242
  (
    n378,
    n78
  );


  not
  g243
  (
    n361,
    n85
  );


  buf
  g244
  (
    KeyWire_0_14,
    n34
  );


  buf
  g245
  (
    n129,
    n49
  );


  not
  g246
  (
    n231,
    n98
  );


  buf
  g247
  (
    n200,
    n75
  );


  buf
  g248
  (
    n401,
    n99
  );


  not
  g249
  (
    n127,
    n45
  );


  not
  g250
  (
    n279,
    n86
  );


  not
  g251
  (
    n350,
    n41
  );


  buf
  g252
  (
    n355,
    n66
  );


  buf
  g253
  (
    n338,
    n45
  );


  buf
  g254
  (
    n342,
    n96
  );


  buf
  g255
  (
    n387,
    n34
  );


  buf
  g256
  (
    n374,
    n51
  );


  buf
  g257
  (
    n226,
    n63
  );


  buf
  g258
  (
    n339,
    n42
  );


  buf
  g259
  (
    n308,
    n60
  );


  not
  g260
  (
    n393,
    n36
  );


  not
  g261
  (
    n249,
    n45
  );


  not
  g262
  (
    n358,
    n82
  );


  buf
  g263
  (
    KeyWire_0_50,
    n60
  );


  buf
  g264
  (
    n197,
    n71
  );


  not
  g265
  (
    n222,
    n53
  );


  not
  g266
  (
    n367,
    n59
  );


  buf
  g267
  (
    n268,
    n38
  );


  buf
  g268
  (
    n141,
    n94
  );


  not
  g269
  (
    n247,
    n41
  );


  buf
  g270
  (
    n140,
    n34
  );


  buf
  g271
  (
    n348,
    n66
  );


  buf
  g272
  (
    n353,
    n39
  );


  buf
  g273
  (
    n253,
    n69
  );


  not
  g274
  (
    n227,
    n90
  );


  not
  g275
  (
    n303,
    n64
  );


  not
  g276
  (
    n413,
    n95
  );


  not
  g277
  (
    n248,
    n98
  );


  buf
  g278
  (
    n234,
    n68
  );


  buf
  g279
  (
    n411,
    n81
  );


  buf
  g280
  (
    n143,
    n52
  );


  not
  g281
  (
    n377,
    n92
  );


  buf
  g282
  (
    n278,
    n64
  );


  buf
  g283
  (
    n344,
    n79
  );


  buf
  g284
  (
    n198,
    n84
  );


  not
  g285
  (
    n204,
    n93
  );


  buf
  g286
  (
    n276,
    n81
  );


  not
  g287
  (
    n224,
    n85
  );


  not
  g288
  (
    n291,
    n56
  );


  buf
  g289
  (
    n135,
    n59
  );


  buf
  g290
  (
    n365,
    n66
  );


  not
  g291
  (
    n360,
    n71
  );


  not
  g292
  (
    n172,
    n33
  );


  buf
  g293
  (
    n305,
    n81
  );


  buf
  g294
  (
    n214,
    n53
  );


  not
  g295
  (
    n215,
    n70
  );


  not
  g296
  (
    n176,
    n65
  );


  buf
  g297
  (
    n330,
    n89
  );


  buf
  g298
  (
    n389,
    n51
  );


  not
  g299
  (
    n213,
    n77
  );


  not
  g300
  (
    n167,
    n86
  );


  not
  g301
  (
    n199,
    n52
  );


  buf
  g302
  (
    n149,
    n43
  );


  not
  g303
  (
    n267,
    n28
  );


  buf
  g304
  (
    n372,
    n38
  );


  buf
  g305
  (
    n325,
    n89
  );


  not
  g306
  (
    n395,
    n98
  );


  buf
  g307
  (
    n326,
    n83
  );


  not
  g308
  (
    n321,
    n83
  );


  not
  g309
  (
    n292,
    n46
  );


  buf
  g310
  (
    n400,
    n95
  );


  not
  g311
  (
    n318,
    n47
  );


  not
  g312
  (
    n246,
    n36
  );


  buf
  g313
  (
    n133,
    n30
  );


  buf
  g314
  (
    n396,
    n44
  );


  not
  g315
  (
    n157,
    n74
  );


  not
  g316
  (
    n217,
    n58
  );


  not
  g317
  (
    n319,
    n50
  );


  buf
  g318
  (
    n409,
    n76
  );


  buf
  g319
  (
    n240,
    n55
  );


  not
  g320
  (
    n380,
    n76
  );


  not
  g321
  (
    KeyWire_0_57,
    n29
  );


  not
  g322
  (
    n407,
    n31
  );


  buf
  g323
  (
    n256,
    n41
  );


  buf
  g324
  (
    n160,
    n64
  );


  buf
  g325
  (
    n273,
    n70
  );


  buf
  g326
  (
    n158,
    n77
  );


  buf
  g327
  (
    n237,
    n36
  );


  buf
  g328
  (
    n163,
    n80
  );


  buf
  g329
  (
    n313,
    n62
  );


  not
  g330
  (
    KeyWire_0_5,
    n58
  );


  buf
  g331
  (
    n164,
    n59
  );


  buf
  g332
  (
    n357,
    n97
  );


  not
  g333
  (
    n412,
    n73
  );


  buf
  g334
  (
    n183,
    n93
  );


  not
  g335
  (
    n347,
    n49
  );


  buf
  g336
  (
    n175,
    n81
  );


  not
  g337
  (
    n132,
    n68
  );


  not
  g338
  (
    n296,
    n88
  );


  not
  g339
  (
    n154,
    n90
  );


  buf
  g340
  (
    n173,
    n90
  );


  not
  g341
  (
    n287,
    n91
  );


  buf
  g342
  (
    n190,
    n28
  );


  not
  g343
  (
    n185,
    n68
  );


  not
  g344
  (
    n405,
    n73
  );


  buf
  g345
  (
    n281,
    n48
  );


  buf
  g346
  (
    n310,
    n51
  );


  buf
  g347
  (
    n146,
    n53
  );


  not
  g348
  (
    n235,
    n85
  );


  not
  g349
  (
    KeyWire_0_11,
    n44
  );


  not
  g350
  (
    KeyWire_0_41,
    n69
  );


  buf
  g351
  (
    KeyWire_0_60,
    n54
  );


  not
  g352
  (
    n329,
    n78
  );


  not
  g353
  (
    n275,
    n94
  );


  buf
  g354
  (
    n340,
    n31
  );


  not
  g355
  (
    n156,
    n75
  );


  buf
  g356
  (
    n399,
    n94
  );


  not
  g357
  (
    n145,
    n41
  );


  buf
  g358
  (
    n216,
    n61
  );


  not
  g359
  (
    n151,
    n86
  );


  not
  g360
  (
    n233,
    n65
  );


  not
  g361
  (
    n261,
    n43
  );


  buf
  g362
  (
    n219,
    n39
  );


  buf
  g363
  (
    n266,
    n35
  );


  buf
  g364
  (
    n408,
    n70
  );


  not
  g365
  (
    KeyWire_0_27,
    n47
  );


  buf
  g366
  (
    n229,
    n49
  );


  not
  g367
  (
    n210,
    n57
  );


  not
  g368
  (
    n203,
    n84
  );


  buf
  g369
  (
    n288,
    n74
  );


  buf
  g370
  (
    KeyWire_0_0,
    n52
  );


  not
  g371
  (
    n280,
    n50
  );


  not
  g372
  (
    n138,
    n56
  );


  buf
  g373
  (
    n322,
    n51
  );


  not
  g374
  (
    n284,
    n35
  );


  not
  g375
  (
    n406,
    n76
  );


  buf
  g376
  (
    n191,
    n75
  );


  buf
  g377
  (
    n165,
    n61
  );


  not
  g378
  (
    n212,
    n62
  );


  not
  g379
  (
    n362,
    n71
  );


  buf
  g380
  (
    n366,
    n62
  );


  buf
  g381
  (
    n398,
    n72
  );


  buf
  g382
  (
    KeyWire_0_29,
    n48
  );


  buf
  g383
  (
    n397,
    n87
  );


  not
  g384
  (
    KeyWire_0_35,
    n39
  );


  buf
  g385
  (
    n403,
    n42
  );


  not
  g386
  (
    n430,
    n146
  );


  not
  g387
  (
    n423,
    n135
  );


  not
  g388
  (
    n431,
    n147
  );


  buf
  g389
  (
    n429,
    n151
  );


  not
  g390
  (
    n433,
    n152
  );


  buf
  g391
  (
    n421,
    n150
  );


  buf
  g392
  (
    KeyWire_0_3,
    n145
  );


  buf
  g393
  (
    n426,
    n133
  );


  buf
  g394
  (
    n422,
    n130
  );


  buf
  g395
  (
    n424,
    n134
  );


  not
  g396
  (
    n436,
    n140
  );


  not
  g397
  (
    n419,
    n144
  );


  buf
  g398
  (
    n427,
    n138
  );


  buf
  g399
  (
    n414,
    n132
  );


  buf
  g400
  (
    n420,
    n129
  );


  not
  g401
  (
    n435,
    n128
  );


  buf
  g402
  (
    n428,
    n137
  );


  not
  g403
  (
    n432,
    n131
  );


  not
  g404
  (
    n416,
    n142
  );


  not
  g405
  (
    n417,
    n136
  );


  buf
  g406
  (
    KeyWire_0_30,
    n149
  );


  not
  g407
  (
    n425,
    n143
  );


  buf
  g408
  (
    n418,
    n141
  );


  buf
  g409
  (
    n437,
    n127
  );


  buf
  g410
  (
    n438,
    n148
  );


  buf
  g411
  (
    n415,
    n139
  );


  nand
  g412
  (
    n474,
    n260,
    n177,
    n174,
    n197
  );


  xnor
  g413
  (
    n452,
    n239,
    n195,
    n266,
    n262
  );


  xnor
  g414
  (
    n533,
    n416,
    n155,
    n275,
    n425
  );


  nand
  g415
  (
    n524,
    n194,
    n284,
    n298,
    n430
  );


  nor
  g416
  (
    n503,
    n314,
    n183,
    n180,
    n298
  );


  or
  g417
  (
    n527,
    n269,
    n208,
    n251,
    n415
  );


  xor
  g418
  (
    n455,
    n237,
    n244,
    n204,
    n270
  );


  nor
  g419
  (
    n448,
    n295,
    n242,
    n250,
    n189
  );


  xnor
  g420
  (
    n479,
    n314,
    n429,
    n425,
    n439
  );


  xor
  g421
  (
    n523,
    n253,
    n424,
    n265
  );


  nor
  g422
  (
    KeyWire_0_12,
    n302,
    n437,
    n428,
    n198
  );


  xor
  g423
  (
    n493,
    n286,
    n291,
    n236,
    n312
  );


  and
  g424
  (
    n463,
    n437,
    n249,
    n303,
    n438
  );


  xor
  g425
  (
    n505,
    n272,
    n190,
    n431,
    n280
  );


  nand
  g426
  (
    n506,
    n309,
    n426,
    n157,
    n219
  );


  xor
  g427
  (
    n520,
    n222,
    n434,
    n303,
    n240
  );


  xnor
  g428
  (
    n515,
    n256,
    n214,
    n185,
    n300
  );


  nor
  g429
  (
    n532,
    n229,
    n289,
    n206,
    n249
  );


  nand
  g430
  (
    n528,
    n436,
    n275,
    n420,
    n418
  );


  and
  g431
  (
    n489,
    n223,
    n247,
    n189,
    n284
  );


  xor
  g432
  (
    n540,
    n311,
    n156,
    n435,
    n287
  );


  or
  g433
  (
    n497,
    n420,
    n239,
    n294,
    n283
  );


  xor
  g434
  (
    n501,
    n228,
    n261,
    n205,
    n252
  );


  xor
  g435
  (
    n539,
    n216,
    n260,
    n419,
    n425
  );


  nor
  g436
  (
    n480,
    n267,
    n301,
    n203,
    n432
  );


  xor
  g437
  (
    n478,
    n273,
    n261,
    n299,
    n256
  );


  and
  g438
  (
    n471,
    n271,
    n282,
    n428,
    n186
  );


  nand
  g439
  (
    n459,
    n422,
    n164,
    n304,
    n424
  );


  and
  g440
  (
    n472,
    n431,
    n163,
    n423,
    n427
  );


  xor
  g441
  (
    n457,
    n418,
    n417,
    n192,
    n421
  );


  and
  g442
  (
    n498,
    n421,
    n251,
    n434,
    n230
  );


  and
  g443
  (
    n488,
    n192,
    n435,
    n224,
    n198
  );


  or
  g444
  (
    n473,
    n180,
    n272,
    n226,
    n199
  );


  nand
  g445
  (
    n494,
    n181,
    n268,
    n175,
    n211
  );


  or
  g446
  (
    n442,
    n209,
    n212,
    n219,
    n439
  );


  nor
  g447
  (
    n504,
    n221,
    n201,
    n278,
    n257
  );


  xor
  g448
  (
    n484,
    n305,
    n211,
    n214,
    n171
  );


  or
  g449
  (
    n451,
    n286,
    n264,
    n296,
    n419
  );


  nand
  g450
  (
    n537,
    n215,
    n193,
    n207,
    n288
  );


  xnor
  g451
  (
    n464,
    n308,
    n292,
    n429,
    n433
  );


  or
  g452
  (
    n477,
    n308,
    n416,
    n306,
    n297
  );


  nor
  g453
  (
    n519,
    n184,
    n154,
    n310,
    n199
  );


  xor
  g454
  (
    n440,
    n184,
    n257,
    n422,
    n235
  );


  xnor
  g455
  (
    n486,
    n414,
    n196,
    n438,
    n417
  );


  and
  g456
  (
    n460,
    n233,
    n267,
    n208,
    n244
  );


  xnor
  g457
  (
    n514,
    n283,
    n417,
    n234,
    n217
  );


  xor
  g458
  (
    n444,
    n315,
    n188,
    n187,
    n289
  );


  xor
  g459
  (
    n453,
    n414,
    n243,
    n161,
    n202
  );


  nand
  g460
  (
    n535,
    n241,
    n427,
    n309,
    n224
  );


  nand
  g461
  (
    n462,
    n271,
    n282,
    n218,
    n212
  );


  nand
  g462
  (
    n482,
    n246,
    n248,
    n238,
    n172
  );


  and
  g463
  (
    n443,
    n312,
    n229,
    n253,
    n436
  );


  or
  g464
  (
    n513,
    n299,
    n302,
    n158,
    n430
  );


  xor
  g465
  (
    n529,
    n194,
    n420,
    n285,
    n290
  );


  and
  g466
  (
    n526,
    n296,
    n434,
    n414,
    n221
  );


  xnor
  g467
  (
    n500,
    n162,
    n170,
    n429,
    n255
  );


  nand
  g468
  (
    n490,
    n281,
    n245,
    n231,
    n220
  );


  xnor
  g469
  (
    n456,
    n218,
    n174,
    n277,
    n424
  );


  xor
  g470
  (
    n491,
    n231,
    n259,
    n238,
    n290
  );


  xor
  g471
  (
    n447,
    n181,
    n175,
    n255,
    n429
  );


  xnor
  g472
  (
    n485,
    n297,
    n268,
    n422,
    n307
  );


  or
  g473
  (
    n475,
    n300,
    n213,
    n421,
    n227
  );


  nor
  g474
  (
    n454,
    n292,
    n311,
    n258,
    n165
  );


  nand
  g475
  (
    n517,
    n226,
    n263,
    n415,
    n168
  );


  xor
  g476
  (
    n522,
    n177,
    n414,
    n423,
    n313
  );


  nor
  g477
  (
    n487,
    n438,
    n430,
    n188,
    n160
  );


  nand
  g478
  (
    n458,
    n201,
    n243,
    n195,
    n313
  );


  xor
  g479
  (
    n510,
    n416,
    n439,
    n274,
    n437
  );


  or
  g480
  (
    n468,
    n295,
    n420,
    n426,
    n173
  );


  xor
  g481
  (
    n534,
    n310,
    n285,
    n276,
    n258
  );


  nand
  g482
  (
    n446,
    n179,
    n437,
    n436,
    n259
  );


  nand
  g483
  (
    n481,
    n287,
    n232,
    n432,
    n204
  );


  xor
  g484
  (
    n538,
    n305,
    n430,
    n190,
    n423
  );


  xor
  g485
  (
    KeyWire_0_8,
    n217,
    n176,
    n433,
    n419
  );


  xnor
  g486
  (
    n465,
    n193,
    n222,
    n435,
    n307
  );


  xnor
  g487
  (
    n469,
    n171,
    n247,
    n206,
    n438
  );


  nand
  g488
  (
    n441,
    n209,
    n215,
    n252,
    n235
  );


  xnor
  g489
  (
    n450,
    n236,
    n182,
    n187,
    n197
  );


  xor
  g490
  (
    n525,
    n233,
    n280,
    n225
  );


  xnor
  g491
  (
    n512,
    n270,
    n200,
    n427,
    n168
  );


  nand
  g492
  (
    KeyWire_0_63,
    n248,
    n419,
    n428,
    n427
  );


  xnor
  g493
  (
    n516,
    n418,
    n265,
    n254,
    n220
  );


  and
  g494
  (
    n461,
    n207,
    n263,
    n281,
    n415
  );


  xor
  g495
  (
    n483,
    n432,
    n433,
    n426,
    n173
  );


  nor
  g496
  (
    n508,
    n200,
    n432,
    n277,
    n227
  );


  nand
  g497
  (
    n530,
    n279,
    n417,
    n264,
    n433
  );


  nor
  g498
  (
    n531,
    n416,
    n273,
    n304,
    n237
  );


  nor
  g499
  (
    n496,
    n415,
    n216,
    n223,
    n178
  );


  nand
  g500
  (
    n521,
    n316,
    n426,
    n170,
    n254
  );


  nand
  g501
  (
    n541,
    n288,
    n202,
    n182,
    n436
  );


  xnor
  g502
  (
    n467,
    n279,
    n178,
    n291,
    n191
  );


  nor
  g503
  (
    n542,
    n269,
    n210,
    n169,
    n153
  );


  or
  g504
  (
    n470,
    n274,
    n439,
    n431,
    n230
  );


  nand
  g505
  (
    n518,
    n418,
    n262,
    n250,
    n306
  );


  nor
  g506
  (
    n543,
    n205,
    n213,
    n293,
    n241
  );


  xnor
  g507
  (
    KeyWire_0_37,
    n431,
    n266,
    n293,
    n245
  );


  xor
  g508
  (
    n466,
    n242,
    n176,
    n191,
    n435
  );


  nand
  g509
  (
    n495,
    n172,
    n232,
    n315,
    n159
  );


  nand
  g510
  (
    n445,
    n183,
    n246,
    n278,
    n425
  );


  xor
  g511
  (
    n476,
    n434,
    n179,
    n196,
    n240
  );


  nor
  g512
  (
    KeyWire_0_43,
    n203,
    n186,
    n234,
    n167
  );


  xor
  g513
  (
    n536,
    n423,
    n428,
    n185,
    n166
  );


  nor
  g514
  (
    n509,
    n210,
    n421,
    n422,
    n301
  );


  xor
  g515
  (
    n502,
    n276,
    n294,
    n228,
    n169
  );


  xnor
  g516
  (
    n555,
    n354,
    n352,
    n344,
    n391
  );


  nor
  g517
  (
    n582,
    n354,
    n515,
    n377,
    n364
  );


  or
  g518
  (
    n561,
    n376,
    n383,
    n351,
    n346
  );


  nor
  g519
  (
    n571,
    n368,
    n106,
    n350,
    n324
  );


  xor
  g520
  (
    n605,
    n497,
    n319,
    n512,
    n378
  );


  and
  g521
  (
    n576,
    n443,
    n375,
    n385,
    n387
  );


  xor
  g522
  (
    n595,
    n485,
    n363,
    n110,
    n530
  );


  xor
  g523
  (
    n622,
    n338,
    n471,
    n362,
    n389
  );


  nand
  g524
  (
    n577,
    n379,
    n331,
    n455,
    n366
  );


  nand
  g525
  (
    KeyWire_0_61,
    n382,
    n101,
    n339,
    n104
  );


  xnor
  g526
  (
    n628,
    n349,
    n518,
    n331,
    n453
  );


  xnor
  g527
  (
    n592,
    n357,
    n488,
    n379,
    n343
  );


  xnor
  g528
  (
    n560,
    n344,
    n531,
    n350,
    n353
  );


  xnor
  g529
  (
    n544,
    n441,
    n475,
    n109,
    n354
  );


  nand
  g530
  (
    n631,
    n384,
    n360,
    n377,
    n380
  );


  and
  g531
  (
    n606,
    n342,
    n377,
    n393,
    n379
  );


  xor
  g532
  (
    n642,
    n395,
    n338,
    n348,
    n26
  );


  xnor
  g533
  (
    n565,
    n365,
    n322,
    n492,
    n347
  );


  xnor
  g534
  (
    n645,
    n348,
    n371,
    n355,
    n326
  );


  xor
  g535
  (
    KeyWire_0_58,
    n364,
    n371,
    n365,
    n388
  );


  nor
  g536
  (
    n640,
    n496,
    n318,
    n105,
    n389
  );


  or
  g537
  (
    n545,
    n337,
    n337,
    n26,
    n528
  );


  nor
  g538
  (
    n619,
    n508,
    n370,
    n527,
    n449
  );


  nor
  g539
  (
    n617,
    n447,
    n369,
    n103,
    n363
  );


  or
  g540
  (
    n648,
    n457,
    n330,
    n339,
    n483
  );


  nand
  g541
  (
    n625,
    n371,
    n387,
    n341,
    n110
  );


  and
  g542
  (
    n610,
    n394,
    n327,
    n108,
    n516
  );


  nand
  g543
  (
    n553,
    n395,
    n359,
    n342
  );


  xor
  g544
  (
    n623,
    n456,
    n459,
    n26,
    n350
  );


  xnor
  g545
  (
    n575,
    n392,
    n340,
    n376,
    n393
  );


  xnor
  g546
  (
    n566,
    n516,
    n349,
    n332,
    n345
  );


  xnor
  g547
  (
    n594,
    n355,
    n355,
    n372,
    n526
  );


  or
  g548
  (
    n638,
    n329,
    n317,
    n476,
    n370
  );


  xnor
  g549
  (
    KeyWire_0_9,
    n506,
    n386,
    n390,
    n323
  );


  xor
  g550
  (
    n643,
    n364,
    n382,
    n336,
    n387
  );


  xor
  g551
  (
    KeyWire_0_28,
    n366,
    n332,
    n358,
    n464
  );


  nand
  g552
  (
    KeyWire_0_55,
    n369,
    n329,
    n375,
    n491
  );


  xor
  g553
  (
    n651,
    n100,
    n463,
    n384,
    n520
  );


  nand
  g554
  (
    n599,
    n367,
    n525,
    n379,
    n460
  );


  nand
  g555
  (
    KeyWire_0_23,
    n360,
    n102,
    n372,
    n345
  );


  xnor
  g556
  (
    KeyWire_0_10,
    n451,
    n502,
    n360,
    n322
  );


  nand
  g557
  (
    n564,
    n361,
    n321,
    n27,
    n100
  );


  or
  g558
  (
    n615,
    n111,
    n509,
    n360,
    n378
  );


  xor
  g559
  (
    n548,
    n477,
    n347,
    n353,
    n361
  );


  and
  g560
  (
    n621,
    n388,
    n524,
    n325,
    n101
  );


  nor
  g561
  (
    KeyWire_0_2,
    n388,
    n376,
    n389,
    n366
  );


  nor
  g562
  (
    n629,
    n381,
    n103,
    n521,
    n442
  );


  and
  g563
  (
    n585,
    n380,
    n383,
    n320,
    n343
  );


  xor
  g564
  (
    n587,
    n374,
    n378,
    n371,
    n394
  );


  nor
  g565
  (
    n637,
    n351,
    n501,
    n390,
    n367
  );


  or
  g566
  (
    n641,
    n481,
    n390,
    n363,
    n366
  );


  xor
  g567
  (
    n616,
    n529,
    n107,
    n462,
    n368
  );


  and
  g568
  (
    n611,
    n106,
    n469,
    n356,
    n522
  );


  nor
  g569
  (
    KeyWire_0_48,
    n498,
    n350,
    n394,
    n367
  );


  nor
  g570
  (
    n633,
    n385,
    n383,
    n382,
    n102
  );


  xor
  g571
  (
    n563,
    n334,
    n104,
    n386,
    n482
  );


  nand
  g572
  (
    n613,
    n520,
    n103,
    n359,
    n109
  );


  nand
  g573
  (
    n546,
    n103,
    n369,
    n109,
    n110
  );


  or
  g574
  (
    KeyWire_0_40,
    n357,
    n487,
    n110,
    n356
  );


  and
  g575
  (
    n632,
    n364,
    n474,
    n374,
    n381
  );


  nor
  g576
  (
    n549,
    n368,
    n374,
    n479,
    n104
  );


  and
  g577
  (
    n644,
    n107,
    n109,
    n522,
    n333
  );


  xnor
  g578
  (
    n590,
    n383,
    n388,
    n466,
    n344
  );


  xor
  g579
  (
    n574,
    n510,
    n27,
    n472,
    n377
  );


  or
  g580
  (
    n552,
    n486,
    n100,
    n105,
    n529
  );


  xnor
  g581
  (
    n607,
    n374,
    n448,
    n523,
    n384
  );


  xnor
  g582
  (
    n551,
    n393,
    n357,
    n367,
    n362
  );


  and
  g583
  (
    KeyWire_0_39,
    n27,
    n323,
    n320,
    n339
  );


  and
  g584
  (
    KeyWire_0_18,
    n351,
    n505,
    n528,
    n499
  );


  xor
  g585
  (
    n646,
    n369,
    n445,
    n342,
    n348
  );


  and
  g586
  (
    n593,
    n381,
    n467,
    n99,
    n25
  );


  or
  g587
  (
    n559,
    n345,
    n317,
    n513,
    n484
  );


  nor
  g588
  (
    n627,
    n465,
    n111,
    n328,
    n341
  );


  nand
  g589
  (
    n649,
    n444,
    n100,
    n343,
    n346
  );


  or
  g590
  (
    n626,
    n385,
    n517,
    n380,
    n500
  );


  nand
  g591
  (
    n580,
    n382,
    n511,
    n515,
    n346
  );


  xnor
  g592
  (
    n608,
    n328,
    n391,
    n346,
    n375
  );


  and
  g593
  (
    n579,
    n373,
    n358,
    n504,
    n490
  );


  and
  g594
  (
    n618,
    n394,
    n321,
    n334,
    n513
  );


  xnor
  g595
  (
    n654,
    n461,
    n108,
    n386,
    n530
  );


  xnor
  g596
  (
    n567,
    n356,
    n495,
    n335,
    n378
  );


  nand
  g597
  (
    n647,
    n519,
    n106,
    n478,
    n503
  );


  and
  g598
  (
    n630,
    n392,
    n108,
    n390,
    n352
  );


  and
  g599
  (
    n554,
    n395,
    n348,
    n393,
    n102
  );


  and
  g600
  (
    n558,
    n341,
    n343,
    n26,
    n318
  );


  xnor
  g601
  (
    n550,
    n362,
    n365,
    n470,
    n458
  );


  nor
  g602
  (
    n609,
    n356,
    n27,
    n353,
    n384
  );


  nor
  g603
  (
    n584,
    n494,
    n370,
    n440
  );


  and
  g604
  (
    KeyWire_0_56,
    n101,
    n373,
    n518,
    n514
  );


  and
  g605
  (
    n603,
    n352,
    n396,
    n480,
    n108
  );


  xor
  g606
  (
    n588,
    n392,
    n351,
    n361,
    n347
  );


  nor
  g607
  (
    n547,
    n523,
    n316,
    n368,
    n373
  );


  and
  g608
  (
    n573,
    n473,
    n330,
    n358,
    n333
  );


  or
  g609
  (
    n568,
    n362,
    n335,
    n373,
    n391
  );


  nand
  g610
  (
    n602,
    n326,
    n372,
    n489,
    n386
  );


  nand
  g611
  (
    n639,
    n358,
    n363,
    n340,
    n519
  );


  nand
  g612
  (
    n570,
    n454,
    n507,
    n359,
    n396
  );


  xnor
  g613
  (
    n598,
    n352,
    n353,
    n385,
    n517
  );


  xnor
  g614
  (
    n589,
    n340,
    n375,
    n395,
    n355
  );


  and
  g615
  (
    n652,
    n327,
    n349,
    n340,
    n101
  );


  xor
  g616
  (
    n578,
    n372,
    n347,
    n102,
    n106
  );


  xor
  g617
  (
    n557,
    n514,
    n446,
    n392,
    n338
  );


  and
  g618
  (
    n601,
    n468,
    n349,
    n380,
    n341
  );


  xor
  g619
  (
    n597,
    n105,
    n450,
    n339,
    n493
  );


  nor
  g620
  (
    n569,
    n357,
    n521,
    n525,
    n107
  );


  nor
  g621
  (
    n612,
    n381,
    n361,
    n526,
    n325
  );


  xnor
  g622
  (
    n596,
    n512,
    n345,
    n111,
    n365
  );


  xor
  g623
  (
    n572,
    n376,
    n319,
    n391,
    n336
  );


  xnor
  g624
  (
    n634,
    n387,
    n105,
    n524,
    n104
  );


  xnor
  g625
  (
    n624,
    n107,
    n359,
    n324,
    n354
  );


  or
  g626
  (
    n635,
    n344,
    n452,
    n389,
    n527
  );


  not
  g627
  (
    n658,
    n531
  );


  not
  g628
  (
    n661,
    n548
  );


  buf
  g629
  (
    n657,
    n546
  );


  buf
  g630
  (
    n656,
    n549
  );


  buf
  g631
  (
    n660,
    n532
  );


  not
  g632
  (
    n659,
    n547
  );


  nand
  g633
  (
    n655,
    n550,
    n545,
    n544
  );


  and
  g634
  (
    n681,
    n597,
    n556,
    n575,
    n587
  );


  or
  g635
  (
    n679,
    n631,
    n623,
    n574,
    n657
  );


  or
  g636
  (
    n676,
    n613,
    n571,
    n581,
    n582
  );


  xnor
  g637
  (
    n684,
    n660,
    n658,
    n661,
    n553
  );


  nor
  g638
  (
    n685,
    n551,
    n660,
    n594,
    n656
  );


  nor
  g639
  (
    n678,
    n656,
    n555,
    n657,
    n585
  );


  nor
  g640
  (
    n675,
    n554,
    n628,
    n611,
    n626
  );


  xnor
  g641
  (
    n669,
    n624,
    n655,
    n615,
    n608
  );


  or
  g642
  (
    n677,
    n593,
    n614,
    n592,
    n603
  );


  xnor
  g643
  (
    n687,
    n604,
    n589,
    n620,
    n625
  );


  nor
  g644
  (
    n664,
    n655,
    n606,
    n661,
    n612
  );


  nor
  g645
  (
    n667,
    n568,
    n569,
    n618,
    n591
  );


  nor
  g646
  (
    n672,
    n610,
    n605,
    n659,
    n599
  );


  nand
  g647
  (
    n662,
    n588,
    n561,
    n564,
    n590
  );


  nor
  g648
  (
    n673,
    n629,
    n570,
    n661,
    n659
  );


  nor
  g649
  (
    n682,
    n622,
    n660,
    n563,
    n627
  );


  nor
  g650
  (
    n668,
    n562,
    n572,
    n578,
    n558
  );


  nor
  g651
  (
    n674,
    n583,
    n657,
    n566,
    n658
  );


  nor
  g652
  (
    n671,
    n621,
    n576,
    n602,
    n586
  );


  nor
  g653
  (
    n688,
    n661,
    n552,
    n658,
    n573
  );


  nor
  g654
  (
    n680,
    n656,
    n560,
    n617,
    n616
  );


  nor
  g655
  (
    n666,
    n565,
    n658,
    n584,
    n656
  );


  or
  g656
  (
    n670,
    n657,
    n601,
    n659,
    n579
  );


  xor
  g657
  (
    n686,
    n609,
    n596,
    n580,
    n660
  );


  xnor
  g658
  (
    n663,
    n655,
    n607,
    n577,
    n630
  );


  and
  g659
  (
    n665,
    n595,
    n619,
    n600,
    n598
  );


  nand
  g660
  (
    n683,
    n559,
    n557,
    n659,
    n567
  );


  or
  g661
  (
    n692,
    n119,
    n121,
    n115,
    n117
  );


  or
  g662
  (
    n707,
    n113,
    n116,
    n124,
    n125
  );


  nor
  g663
  (
    n703,
    n663,
    n117,
    n673,
    n675
  );


  and
  g664
  (
    n701,
    n664,
    n118,
    n122
  );


  or
  g665
  (
    n697,
    n114,
    n669,
    n119,
    n112
  );


  or
  g666
  (
    n696,
    n114,
    n668,
    n676,
    n124
  );


  nand
  g667
  (
    n689,
    n121,
    n125,
    n117,
    n111
  );


  or
  g668
  (
    KeyWire_0_53,
    n676,
    n120,
    n118
  );


  nor
  g669
  (
    n690,
    n676,
    n113,
    n122,
    n123
  );


  xnor
  g670
  (
    KeyWire_0_47,
    n674,
    n119,
    n662,
    n123
  );


  or
  g671
  (
    n704,
    n121,
    n671,
    n675,
    n126
  );


  and
  g672
  (
    n693,
    n123,
    n118,
    n121,
    n122
  );


  nand
  g673
  (
    n705,
    n115,
    n113,
    n125
  );


  nor
  g674
  (
    n691,
    n124,
    n114,
    n675,
    n115
  );


  xor
  g675
  (
    n702,
    n120,
    n113,
    n666,
    n124
  );


  nor
  g676
  (
    n708,
    n118,
    n114,
    n119,
    n672
  );


  and
  g677
  (
    n694,
    n670,
    n675,
    n126,
    n120
  );


  or
  g678
  (
    n699,
    n123,
    n116,
    n665,
    n112
  );


  nand
  g679
  (
    n706,
    n117,
    n116,
    n115
  );


  xor
  g680
  (
    KeyWire_0_19,
    n667,
    n126,
    n112
  );


  xor
  g681
  (
    n721,
    n397,
    n402,
    n406,
    n696
  );


  xor
  g682
  (
    n722,
    n404,
    n407,
    n400,
    n697
  );


  xor
  g683
  (
    n710,
    n399,
    n397,
    n404,
    n401
  );


  nand
  g684
  (
    n718,
    n703,
    n398,
    n400
  );


  or
  g685
  (
    n712,
    n405,
    n396,
    n403,
    n401
  );


  or
  g686
  (
    n717,
    n702,
    n397,
    n407,
    n398
  );


  nor
  g687
  (
    n719,
    n399,
    n706,
    n701,
    n407
  );


  nand
  g688
  (
    n711,
    n406,
    n707,
    n705,
    n397
  );


  and
  g689
  (
    n724,
    n400,
    n398,
    n403
  );


  or
  g690
  (
    n723,
    n694,
    n399,
    n396,
    n402
  );


  nor
  g691
  (
    n716,
    n402,
    n693,
    n403,
    n404
  );


  nand
  g692
  (
    n713,
    n708,
    n408,
    n699
  );


  xor
  g693
  (
    n714,
    n399,
    n401,
    n406,
    n700
  );


  xor
  g694
  (
    n720,
    n406,
    n698,
    n405
  );


  and
  g695
  (
    KeyWire_0_45,
    n407,
    n404,
    n402,
    n405
  );


  xor
  g696
  (
    n715,
    n695,
    n401,
    n704,
    n403
  );


  nor
  g697
  (
    n726,
    n649,
    n648,
    n640,
    n652
  );


  nor
  g698
  (
    n725,
    n635,
    n710,
    n643
  );


  nor
  g699
  (
    n727,
    n642,
    n710,
    n709
  );


  nand
  g700
  (
    n729,
    n632,
    n650,
    n637,
    n647
  );


  or
  g701
  (
    n728,
    n645,
    n646,
    n641,
    n638
  );


  or
  g702
  (
    n730,
    n636,
    n644,
    n709
  );


  nand
  g703
  (
    n731,
    n634,
    n651,
    n633,
    n639
  );


  nand
  g704
  (
    n741,
    n717,
    n718,
    n728,
    n713
  );


  xnor
  g705
  (
    n742,
    n713,
    n716,
    n711,
    n712
  );


  nand
  g706
  (
    n733,
    n717,
    n716,
    n729,
    n712
  );


  nand
  g707
  (
    n734,
    n717,
    n711,
    n712,
    n728
  );


  xnor
  g708
  (
    n732,
    n714,
    n717,
    n715,
    n716
  );


  xor
  g709
  (
    n737,
    n718,
    n714,
    n729
  );


  nand
  g710
  (
    n735,
    n718,
    n713,
    n719,
    n726
  );


  nand
  g711
  (
    n739,
    n715,
    n725,
    n727,
    n714
  );


  nand
  g712
  (
    n738,
    n712,
    n715,
    n711,
    n718
  );


  nor
  g713
  (
    KeyWire_0_25,
    n711,
    n727,
    n728
  );


  nand
  g714
  (
    n736,
    n713,
    n715,
    n728,
    n716
  );


  and
  g715
  (
    n743,
    n680,
    n409,
    n734,
    n679
  );


  xor
  g716
  (
    n749,
    n680,
    n678,
    n677
  );


  nand
  g717
  (
    n748,
    n678,
    n408,
    n679
  );


  xnor
  g718
  (
    n747,
    n737,
    n680,
    n677
  );


  and
  g719
  (
    n745,
    n735,
    n678,
    n733,
    n732
  );


  xor
  g720
  (
    n746,
    n677,
    n681,
    n676,
    n738
  );


  or
  g721
  (
    n744,
    n736,
    n679,
    n408,
    n680
  );


  nand
  g722
  (
    n753,
    n744,
    n739,
    n748,
    n533
  );


  xnor
  g723
  (
    n752,
    n742,
    n721,
    n740,
    n720
  );


  xnor
  g724
  (
    n751,
    n746,
    n719,
    n721
  );


  xnor
  g725
  (
    n750,
    n533,
    n743,
    n720,
    n719
  );


  xnor
  g726
  (
    n755,
    n741,
    n720,
    n745,
    n747
  );


  and
  g727
  (
    n754,
    n721,
    n719,
    n720,
    n532
  );


  xor
  g728
  (
    KeyWire_0_34,
    n681,
    n682,
    n752
  );


  nor
  g729
  (
    n756,
    n750,
    n681,
    n722
  );


  nand
  g730
  (
    n757,
    n683,
    n751,
    n682
  );


  and
  g731
  (
    n760,
    n757,
    n730
  );


  xnor
  g732
  (
    n759,
    n729,
    n729,
    n730,
    n756
  );


  xnor
  g733
  (
    n762,
    n723,
    n723,
    n760,
    n722
  );


  nor
  g734
  (
    n761,
    n722,
    n759,
    n760,
    n723
  );


  nor
  g735
  (
    n763,
    n722,
    n724,
    n723
  );


  buf
  g736
  (
    n770,
    n761
  );


  not
  g737
  (
    n766,
    n731
  );


  not
  g738
  (
    n764,
    n762
  );


  buf
  g739
  (
    n769,
    n731
  );


  buf
  g740
  (
    n768,
    n731
  );


  buf
  g741
  (
    n773,
    n762
  );


  not
  g742
  (
    n772,
    n749
  );


  and
  g743
  (
    n765,
    n683,
    n763,
    n731
  );


  xnor
  g744
  (
    n767,
    n763,
    n761,
    n762
  );


  nor
  g745
  (
    n771,
    n762,
    n763
  );


  not
  g746
  (
    n775,
    n764
  );


  not
  g747
  (
    n774,
    n764
  );


  xnor
  g748
  (
    n779,
    n774,
    n765,
    n764,
    n769
  );


  xnor
  g749
  (
    n776,
    n766,
    n766,
    n775,
    n768
  );


  or
  g750
  (
    n783,
    n768,
    n766,
    n765,
    n774
  );


  nor
  g751
  (
    KeyWire_0_31,
    n765,
    n766,
    n768,
    n764
  );


  xnor
  g752
  (
    n780,
    n774,
    n724,
    n767,
    n775
  );


  nand
  g753
  (
    n781,
    n767,
    n767,
    n768,
    n774
  );


  or
  g754
  (
    n782,
    n775,
    n769,
    n767
  );


  nor
  g755
  (
    n777,
    n769,
    n765,
    n775,
    n724
  );


  not
  g756
  (
    n791,
    n410
  );


  not
  g757
  (
    KeyWire_0_42,
    n410
  );


  not
  g758
  (
    n786,
    n412
  );


  buf
  g759
  (
    n790,
    n779
  );


  nand
  g760
  (
    n785,
    n778,
    n776,
    n409,
    n410
  );


  or
  g761
  (
    n788,
    n412,
    n411,
    n780,
    n409
  );


  or
  g762
  (
    n789,
    n781,
    n411,
    n779
  );


  nand
  g763
  (
    n787,
    n778,
    n410,
    n412,
    n777
  );


  nand
  g764
  (
    n784,
    n780,
    n409,
    n412,
    n411
  );


  buf
  g765
  (
    n793,
    n784
  );


  not
  g766
  (
    n794,
    n784
  );


  or
  g767
  (
    n795,
    n794,
    n413
  );


  xnor
  g768
  (
    n796,
    n755,
    n654,
    n795,
    n753
  );


  nor
  g769
  (
    n797,
    n653,
    n795,
    n758,
    n754
  );


  xnor
  g770
  (
    n798,
    n796,
    n770
  );


  or
  g771
  (
    n799,
    n798,
    n786,
    n787
  );


  xnor
  g772
  (
    n801,
    n787,
    n788,
    n798,
    n786
  );


  nand
  g773
  (
    n800,
    n787,
    n786,
    n785
  );


  nor
  g774
  (
    n802,
    n797,
    n798,
    n788
  );


  or
  g775
  (
    n816,
    n536,
    n802,
    n535,
    n543
  );


  nand
  g776
  (
    n803,
    n540,
    n771,
    n537,
    n782
  );


  and
  g777
  (
    n813,
    n538,
    n772,
    n801
  );


  nand
  g778
  (
    n804,
    n802,
    n773,
    n684,
    n800
  );


  xor
  g779
  (
    n814,
    n772,
    n799,
    n800
  );


  and
  g780
  (
    n818,
    n537,
    n536,
    n540,
    n800
  );


  nand
  g781
  (
    n805,
    n541,
    n773,
    n126,
    n535
  );


  nor
  g782
  (
    n808,
    n801,
    n685,
    n772,
    n534
  );


  nand
  g783
  (
    n812,
    n771,
    n802,
    n801,
    n799
  );


  nand
  g784
  (
    n806,
    n771,
    n538,
    n683,
    n782
  );


  xor
  g785
  (
    KeyWire_0_36,
    n781,
    n542,
    n771
  );


  xor
  g786
  (
    n815,
    n772,
    n543,
    n539,
    n773
  );


  or
  g787
  (
    n817,
    n413,
    n684
  );


  xor
  g788
  (
    n810,
    n683,
    n800,
    n799,
    n770
  );


  and
  g789
  (
    KeyWire_0_54,
    n534,
    n802,
    n685,
    n539
  );


  xnor
  g790
  (
    n811,
    n685,
    n541,
    n783
  );


  or
  g791
  (
    KeyWire_0_59,
    n810,
    n773,
    n807,
    n804
  );


  and
  g792
  (
    n819,
    n811,
    n791,
    n688,
    n790
  );


  nor
  g793
  (
    n826,
    n688,
    n685,
    n791,
    n818
  );


  nand
  g794
  (
    n821,
    n803,
    n790,
    n686,
    n687
  );


  xnor
  g795
  (
    n829,
    n792,
    n687,
    n791
  );


  xnor
  g796
  (
    KeyWire_0_51,
    n815,
    n817,
    n788,
    n790
  );


  or
  g797
  (
    n822,
    n790,
    n688,
    n687,
    n792
  );


  xnor
  g798
  (
    n830,
    n805,
    n816,
    n789,
    n791
  );


  nor
  g799
  (
    n827,
    n808,
    n686,
    n789,
    n792
  );


  or
  g800
  (
    n824,
    n792,
    n813,
    n812,
    n789
  );


  or
  g801
  (
    n823,
    n688,
    n788,
    n789,
    n809
  );


  nand
  g802
  (
    n825,
    n686,
    n686,
    n814,
    n806
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n334,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n111,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n583,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n434,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n245,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n196,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n104,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n404,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n507,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n562,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n591,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n250,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n511,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n29,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n258,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n112,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n92,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n114,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n600,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n695,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n63,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n93,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n110,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n586,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n182,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n740,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n121,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n285,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n614,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n383,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n439,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n778,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n71,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n335,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n758,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n161,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n809,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n492,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n49,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n650,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n653,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n251,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n792,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n499,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n177,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n709,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n87,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n698,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n581,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n238,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n311,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n828,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n120,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n700,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n807,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n556,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n604,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n307,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n636,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n820,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n153,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n620,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n78,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n449,
    KeyNOTWire_0_63
  );


endmodule


