// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1120_14_8 written by SynthGen on 2021/05/24 19:42:17
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1120_14_8 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25,
 n1108, n1097, n1103, n1098, n1104, n1099, n1100, n1086,
 n1101, n1089, n1106, n1091, n1134, n1136, n1140, n1142,
 n1141, n1143, n1144, n1145, n1139);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25;

output n1108, n1097, n1103, n1098, n1104, n1099, n1100, n1086,
 n1101, n1089, n1106, n1091, n1134, n1136, n1140, n1142,
 n1141, n1143, n1144, n1145, n1139;

wire n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
 n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
 n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
 n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
 n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
 n1082, n1083, n1084, n1085, n1087, n1088, n1090, n1092,
 n1093, n1094, n1095, n1096, n1102, n1105, n1107, n1109,
 n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
 n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
 n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
 n1135, n1137, n1138;

buf  g0 (n28, n2);
not  g1 (n27, n3);
not  g2 (n34, n7);
not  g3 (n33, n3);
not  g4 (n30, n1);
buf  g5 (n36, n8);
not  g6 (n35, n2);
buf  g7 (n32, n5);
buf  g8 (n29, n6);
not  g9 (n37, n2);
not  g10 (n31, n4);
or   g11 (n39, n6, n4, n7, n5);
xor  g12 (n38, n3, n7, n6, n4);
xnor g13 (n26, n5, n8, n1);
not  g14 (n43, n32);
buf  g15 (n40, n27);
not  g16 (n49, n28);
buf  g17 (n51, n31);
buf  g18 (n41, n34);
buf  g19 (n52, n28);
buf  g20 (n53, n37);
buf  g21 (n57, n29);
nand g22 (n42, n26, n30);
and  g23 (n47, n33, n32, n29);
and  g24 (n55, n36, n26, n27);
and  g25 (n54, n34, n36, n30, n33);
and  g26 (n44, n32, n28, n35, n31);
or   g27 (n58, n28, n36, n35);
nand g28 (n48, n34, n27, n30, n35);
nor  g29 (n46, n30, n35, n27, n31);
or   g30 (n45, n33, n31, n26, n37);
or   g31 (n50, n34, n29, n32, n33);
nor  g32 (n56, n37, n38);
or   g33 (n64, n42, n50, n55, n56);
xnor g34 (n62, n40, n53, n54, n49);
nor  g35 (n61, n51, n50, n53, n41);
or   g36 (n63, n43, n48, n54, n44);
xor  g37 (n60, n47, n55, n51);
xor  g38 (n59, n45, n52, n46);
buf  g39 (n74, n59);
not  g40 (n73, n38);
not  g41 (n67, n38);
buf  g42 (n70, n64);
buf  g43 (n65, n9);
not  g44 (n72, n9);
buf  g45 (n71, n8);
not  g46 (n68, n63);
not  g47 (n66, n63);
not  g48 (n79, n60);
buf  g49 (n77, n62);
buf  g50 (n69, n59);
and  g51 (n75, n62, n64, n9, n63);
nand g52 (n76, n62, n61, n64, n9);
nand g53 (n78, n63, n60, n10, n59);
or   g54 (n80, n60, n61, n64);
not  g55 (n90, n70);
buf  g56 (n100, n13);
not  g57 (n82, n73);
not  g58 (n86, n56);
buf  g59 (n102, n13);
buf  g60 (n91, n68);
xor  g61 (n96, n14, n77);
or   g62 (n95, n71, n78);
nand g63 (n83, n78, n77);
nand g64 (n110, n76, n11);
nand g65 (n101, n14, n11);
xnor g66 (n87, n75, n77);
or   g67 (n93, n65, n74);
and  g68 (n92, n80, n14);
and  g69 (n107, n15, n72);
xnor g70 (n85, n79, n76);
xor  g71 (n109, n12, n73);
and  g72 (n111, n10, n66);
and  g73 (n89, n15, n67);
or   g74 (n97, n11, n12);
buf  g75 (n104, n79);
and  g76 (n112, n16, n80);
nor  g77 (n81, n13, n16);
nand g78 (n84, n69, n75);
nor  g79 (n98, n15, n12);
and  g80 (n88, n75, n74);
and  g81 (n106, n78, n73);
xor  g82 (n105, n14, n13);
or   g83 (n108, n12, n15);
or   g84 (n94, n10, n74);
or   g85 (n103, n10, n11);
nand g86 (n99, n80, n76);
not  g87 (n117, n81);
not  g88 (n205, n92);
buf  g89 (n148, n87);
buf  g90 (n214, n106);
buf  g91 (n139, n97);
not  g92 (n136, n101);
buf  g93 (n125, n101);
not  g94 (n113, n93);
not  g95 (n239, n88);
buf  g96 (n198, n90);
not  g97 (n114, n104);
buf  g98 (n206, n98);
buf  g99 (n119, n111);
buf  g100 (n210, n112);
not  g101 (n132, n102);
buf  g102 (n202, n83);
buf  g103 (n207, n93);
not  g104 (n153, n82);
not  g105 (n219, n102);
not  g106 (n134, n88);
buf  g107 (n116, n89);
not  g108 (n222, n112);
buf  g109 (n124, n107);
not  g110 (n221, n103);
buf  g111 (n179, n101);
not  g112 (n181, n104);
not  g113 (n204, n85);
not  g114 (n176, n81);
buf  g115 (n175, n103);
not  g116 (n232, n106);
buf  g117 (n201, n95);
buf  g118 (n229, n89);
buf  g119 (n190, n94);
not  g120 (n140, n89);
buf  g121 (n200, n111);
not  g122 (n189, n110);
buf  g123 (n171, n99);
buf  g124 (n185, n89);
not  g125 (n195, n97);
buf  g126 (n180, n82);
not  g127 (n162, n90);
not  g128 (n143, n85);
not  g129 (n122, n86);
not  g130 (n235, n100);
buf  g131 (n147, n109);
buf  g132 (n127, n108);
buf  g133 (n126, n99);
not  g134 (n160, n102);
buf  g135 (n217, n106);
buf  g136 (n178, n97);
not  g137 (n224, n86);
buf  g138 (n120, n97);
buf  g139 (n118, n81);
not  g140 (n166, n94);
not  g141 (n233, n90);
buf  g142 (n177, n110);
not  g143 (n228, n96);
buf  g144 (n142, n95);
buf  g145 (n129, n84);
buf  g146 (n169, n95);
not  g147 (n155, n92);
buf  g148 (n216, n83);
not  g149 (n208, n87);
not  g150 (n130, n81);
buf  g151 (n141, n95);
buf  g152 (n227, n107);
not  g153 (n193, n84);
not  g154 (n240, n108);
not  g155 (n225, n92);
not  g156 (n203, n93);
not  g157 (n196, n99);
buf  g158 (n123, n98);
buf  g159 (n150, n82);
buf  g160 (n213, n106);
buf  g161 (n223, n87);
not  g162 (n212, n105);
not  g163 (n154, n98);
not  g164 (n194, n109);
not  g165 (n236, n105);
buf  g166 (n135, n93);
not  g167 (n220, n108);
buf  g168 (n133, n107);
not  g169 (n173, n96);
buf  g170 (n174, n92);
buf  g171 (n215, n85);
not  g172 (n164, n100);
not  g173 (n152, n111);
not  g174 (n238, n91);
not  g175 (n234, n82);
buf  g176 (n159, n100);
not  g177 (n158, n112);
buf  g178 (n151, n101);
not  g179 (n167, n84);
buf  g180 (n209, n98);
buf  g181 (n161, n102);
buf  g182 (n156, n85);
buf  g183 (n168, n105);
not  g184 (n226, n91);
not  g185 (n192, n90);
not  g186 (n163, n87);
buf  g187 (n186, n91);
not  g188 (n231, n86);
buf  g189 (n211, n111);
not  g190 (n237, n100);
buf  g191 (n182, n88);
buf  g192 (n157, n103);
not  g193 (n137, n96);
not  g194 (n165, n96);
not  g195 (n115, n83);
buf  g196 (n146, n110);
not  g197 (n183, n104);
buf  g198 (n184, n112);
not  g199 (n149, n84);
buf  g200 (n121, n94);
not  g201 (n170, n109);
buf  g202 (n138, n91);
buf  g203 (n230, n103);
buf  g204 (n197, n94);
buf  g205 (n128, n86);
buf  g206 (n187, n99);
buf  g207 (n218, n110);
buf  g208 (n144, n83);
not  g209 (n131, n88);
not  g210 (n172, n108);
buf  g211 (n188, n109);
buf  g212 (n199, n107);
not  g213 (n145, n104);
buf  g214 (n191, n105);
not  g215 (n406, n116);
buf  g216 (n452, n120);
buf  g217 (n372, n220);
not  g218 (n414, n236);
buf  g219 (n428, n196);
not  g220 (n367, n127);
not  g221 (n479, n173);
not  g222 (n285, n189);
not  g223 (n358, n228);
buf  g224 (n312, n213);
buf  g225 (n346, n184);
not  g226 (n331, n214);
buf  g227 (n337, n151);
not  g228 (n326, n208);
not  g229 (n419, n157);
buf  g230 (n482, n154);
buf  g231 (n332, n178);
not  g232 (n304, n178);
not  g233 (n311, n207);
buf  g234 (n274, n224);
buf  g235 (n437, n220);
not  g236 (n261, n202);
buf  g237 (n328, n228);
buf  g238 (n383, n179);
not  g239 (n499, n206);
not  g240 (n457, n134);
buf  g241 (n402, n176);
not  g242 (n266, n227);
buf  g243 (n315, n178);
not  g244 (n434, n197);
buf  g245 (n345, n157);
buf  g246 (n470, n238);
not  g247 (n291, n126);
buf  g248 (n405, n181);
not  g249 (n483, n144);
buf  g250 (n333, n143);
not  g251 (n458, n183);
buf  g252 (n469, n125);
not  g253 (n427, n163);
buf  g254 (n282, n179);
buf  g255 (n362, n159);
not  g256 (n490, n155);
buf  g257 (n276, n153);
not  g258 (n454, n129);
buf  g259 (n410, n117);
buf  g260 (n342, n122);
not  g261 (n415, n233);
buf  g262 (n356, n132);
not  g263 (n330, n174);
not  g264 (n303, n195);
buf  g265 (n322, n215);
not  g266 (n382, n135);
not  g267 (n387, n161);
not  g268 (n253, n158);
not  g269 (n249, n177);
not  g270 (n471, n169);
buf  g271 (n307, n227);
not  g272 (n497, n161);
not  g273 (n246, n128);
buf  g274 (n318, n212);
not  g275 (n306, n133);
buf  g276 (n302, n211);
buf  g277 (n334, n149);
buf  g278 (n280, n237);
buf  g279 (n338, n193);
buf  g280 (n461, n177);
buf  g281 (n329, n149);
not  g282 (n412, n199);
buf  g283 (n289, n148);
buf  g284 (n449, n223);
buf  g285 (n409, n131);
buf  g286 (n258, n184);
buf  g287 (n354, n231);
not  g288 (n250, n176);
not  g289 (n324, n176);
not  g290 (n456, n234);
buf  g291 (n448, n130);
not  g292 (n468, n118);
buf  g293 (n502, n156);
not  g294 (n259, n207);
buf  g295 (n496, n178);
not  g296 (n385, n129);
buf  g297 (n264, n194);
not  g298 (n283, n204);
not  g299 (n263, n222);
not  g300 (n341, n237);
not  g301 (n284, n209);
buf  g302 (n265, n132);
not  g303 (n391, n234);
buf  g304 (n316, n126);
buf  g305 (n420, n196);
not  g306 (n435, n199);
not  g307 (n487, n228);
not  g308 (n492, n233);
buf  g309 (n393, n201);
not  g310 (n270, n200);
not  g311 (n277, n159);
buf  g312 (n422, n56);
buf  g313 (n371, n215);
buf  g314 (n272, n168);
not  g315 (n464, n197);
buf  g316 (n401, n136);
buf  g317 (n426, n164);
buf  g318 (n295, n239);
not  g319 (n474, n161);
not  g320 (n369, n196);
buf  g321 (n467, n114);
buf  g322 (n475, n140);
not  g323 (n488, n156);
buf  g324 (n460, n122);
not  g325 (n248, n159);
not  g326 (n439, n115);
not  g327 (n299, n218);
not  g328 (n273, n170);
not  g329 (n494, n164);
buf  g330 (n376, n165);
not  g331 (n363, n136);
buf  g332 (n357, n172);
buf  g333 (n486, n156);
buf  g334 (n404, n236);
not  g335 (n374, n216);
not  g336 (n390, n212);
not  g337 (n394, n149);
buf  g338 (n375, n157);
not  g339 (n498, n234);
not  g340 (n466, n217);
buf  g341 (n472, n132);
not  g342 (n365, n167);
buf  g343 (n313, n165);
not  g344 (n429, n152);
buf  g345 (n335, n174);
not  g346 (n484, n145);
not  g347 (n290, n166);
not  g348 (n396, n153);
buf  g349 (n244, n240);
buf  g350 (n389, n150);
not  g351 (n267, n113);
buf  g352 (n325, n116);
buf  g353 (n453, n123);
buf  g354 (n241, n120);
buf  g355 (n355, n181);
not  g356 (n441, n163);
not  g357 (n403, n128);
buf  g358 (n443, n195);
not  g359 (n243, n232);
buf  g360 (n408, n240);
buf  g361 (n268, n193);
buf  g362 (n336, n224);
not  g363 (n378, n138);
buf  g364 (n432, n206);
buf  g365 (n257, n122);
buf  g366 (n278, n118);
buf  g367 (n339, n186);
buf  g368 (n296, n177);
not  g369 (n310, n172);
buf  g370 (n353, n188);
buf  g371 (n301, n130);
not  g372 (n397, n138);
not  g373 (n424, n141);
not  g374 (n478, n230);
not  g375 (n379, n224);
buf  g376 (n352, n233);
buf  g377 (n314, n187);
buf  g378 (n481, n114);
buf  g379 (n451, n223);
not  g380 (n377, n182);
buf  g381 (n392, n123);
buf  g382 (n317, n142);
buf  g383 (n308, n230);
not  g384 (n400, n135);
not  g385 (n254, n129);
buf  g386 (n431, n162);
not  g387 (n319, n222);
not  g388 (n373, n224);
not  g389 (n347, n191);
buf  g390 (n288, n125);
buf  g391 (n349, n239);
buf  g392 (n294, n238);
and  g393 (n361, n182, n127, n218);
nor  g394 (n269, n194, n133, n236, n128);
xnor g395 (n298, n157, n193, n137, n139);
and  g396 (n255, n232, n126, n217, n196);
xnor g397 (n446, n183, n148, n180, n121);
nor  g398 (n380, n197, n225, n173, n162);
xnor g399 (n245, n201, n211, n210, n161);
xor  g400 (n501, n189, n226, n152, n160);
or   g401 (n242, n173, n205, n235, n127);
xnor g402 (n351, n229, n135, n190, n221);
xor  g403 (n275, n165, n212, n185, n215);
and  g404 (n251, n183, n206, n154, n150);
xnor g405 (n411, n131, n141, n119, n221);
xor  g406 (n309, n166, n210, n174, n170);
or   g407 (n416, n147, n147, n159, n152);
xor  g408 (n366, n185, n203, n115, n163);
and  g409 (n381, n235, n188, n184, n216);
or   g410 (n413, n191, n232, n210, n144);
nor  g411 (n386, n203, n167, n143, n151);
and  g412 (n297, n134, n208, n204, n215);
nor  g413 (n440, n237, n198, n131, n136);
nand g414 (n340, n194, n170, n190, n216);
or   g415 (n477, n184, n119, n221, n118);
or   g416 (n485, n164, n199, n183, n181);
or   g417 (n450, n192, n238, n171, n239);
xor  g418 (n463, n218, n162, n202, n131);
xor  g419 (n252, n180, n129, n229, n182);
or   g420 (n465, n137, n237, n192, n115);
or   g421 (n287, n190, n197, n121, n217);
nand g422 (n292, n122, n226, n181, n177);
and  g423 (n407, n195, n113, n185, n182);
and  g424 (n370, n227, n154, n155, n124);
nand g425 (n430, n160, n155, n192, n240);
or   g426 (n442, n146, n142, n164, n219);
or   g427 (n279, n175, n175, n231, n128);
or   g428 (n271, n198, n230, n186, n225);
nand g429 (n438, n141, n145, n125, n205);
nor  g430 (n359, n123, n124, n216, n205);
and  g431 (n348, n133, n141, n226, n235);
and  g432 (n462, n179, n170, n140, n199);
and  g433 (n360, n174, n117, n234, n213);
xnor g434 (n398, n211, n120, n143, n166);
xor  g435 (n491, n180, n139, n144);
and  g436 (n480, n114, n185, n162, n207);
nor  g437 (n489, n145, n172, n168, n142);
nand g438 (n495, n232, n190, n225, n220);
nor  g439 (n321, n201, n228, n203, n167);
nor  g440 (n445, n125, n186, n147, n146);
xor  g441 (n327, n113, n158, n222, n203);
xor  g442 (n305, n124, n238, n139, n116);
and  g443 (n473, n193, n113, n172, n192);
and  g444 (n395, n213, n117, n223, n187);
or   g445 (n323, n163, n188, n155, n239);
xor  g446 (n476, n175, n133, n200, n209);
or   g447 (n417, n219, n143, n189, n168);
and  g448 (n350, n117, n227, n231, n142);
or   g449 (n344, n119, n160, n231, n114);
and  g450 (n455, n158, n145, n147, n171);
or   g451 (n384, n194, n121, n201, n195);
xor  g452 (n256, n209, n212, n167, n225);
xnor g453 (n320, n189, n153, n198, n148);
nor  g454 (n459, n138, n148, n134, n136);
xnor g455 (n444, n205, n169, n208, n175);
or   g456 (n500, n149, n176, n200, n150);
nand g457 (n364, n121, n130, n191, n187);
and  g458 (n433, n156, n119, n166, n168);
or   g459 (n493, n206, n204, n217, n137);
or   g460 (n293, n218, n140, n132, n207);
or   g461 (n447, n229, n219, n151, n126);
xnor g462 (n423, n116, n169, n230, n118);
and  g463 (n247, n115, n214, n135, n236);
xnor g464 (n388, n139, n233, n208, n153);
xnor g465 (n300, n179, n140, n214, n165);
nor  g466 (n425, n180, n200, n123, n198);
nand g467 (n418, n146, n226, n187, n210);
and  g468 (n421, n150, n219, n154, n146);
or   g469 (n260, n169, n120, n202, n173);
xor  g470 (n343, n188, n152, n240, n221);
xnor g471 (n281, n171, n151, n204, n186);
nand g472 (n436, n211, n220, n158, n127);
or   g473 (n399, n222, n137, n130, n171);
or   g474 (n368, n191, n214, n202, n124);
xor  g475 (n262, n138, n213, n229, n209);
or   g476 (n286, n134, n223, n160, n235);
not  g477 (n762, n337);
buf  g478 (n673, n402);
buf  g479 (n682, n456);
not  g480 (n534, n279);
not  g481 (n845, n348);
buf  g482 (n590, n299);
not  g483 (n528, n344);
buf  g484 (n747, n18);
not  g485 (n823, n320);
not  g486 (n776, n483);
not  g487 (n899, n374);
not  g488 (n721, n477);
not  g489 (n654, n259);
buf  g490 (n798, n303);
buf  g491 (n792, n312);
buf  g492 (n810, n374);
not  g493 (n584, n376);
buf  g494 (n724, n345);
buf  g495 (n917, n403);
buf  g496 (n913, n323);
not  g497 (n729, n273);
buf  g498 (n872, n441);
buf  g499 (n780, n461);
buf  g500 (n625, n475);
not  g501 (n617, n389);
buf  g502 (n740, n409);
buf  g503 (n681, n57);
not  g504 (n831, n482);
not  g505 (n766, n337);
not  g506 (n954, n390);
buf  g507 (n842, n411);
not  g508 (n542, n360);
not  g509 (n609, n417);
not  g510 (n870, n443);
buf  g511 (n518, n18);
not  g512 (n647, n417);
not  g513 (n770, n446);
not  g514 (n697, n329);
not  g515 (n962, n245);
buf  g516 (n613, n485);
buf  g517 (n541, n469);
not  g518 (n514, n281);
buf  g519 (n895, n495);
not  g520 (n704, n476);
not  g521 (n649, n283);
not  g522 (n614, n344);
not  g523 (n522, n272);
buf  g524 (n765, n267);
buf  g525 (n841, n452);
not  g526 (n540, n296);
buf  g527 (n879, n423);
not  g528 (n675, n300);
not  g529 (n888, n302);
not  g530 (n859, n299);
not  g531 (n858, n368);
not  g532 (n607, n380);
not  g533 (n904, n342);
not  g534 (n964, n458);
buf  g535 (n887, n471);
not  g536 (n662, n472);
not  g537 (n652, n341);
buf  g538 (n574, n248);
not  g539 (n703, n250);
buf  g540 (n644, n248);
buf  g541 (n808, n479);
buf  g542 (n637, n411);
buf  g543 (n725, n277);
not  g544 (n559, n313);
not  g545 (n728, n413);
not  g546 (n757, n400);
buf  g547 (n715, n367);
buf  g548 (n612, n251);
not  g549 (n633, n382);
buf  g550 (n796, n308);
buf  g551 (n783, n241);
buf  g552 (n691, n488);
not  g553 (n670, n408);
not  g554 (n549, n312);
not  g555 (n521, n338);
not  g556 (n961, n397);
buf  g557 (n722, n498);
buf  g558 (n925, n421);
not  g559 (n854, n317);
not  g560 (n733, n454);
buf  g561 (n579, n419);
buf  g562 (n587, n363);
buf  g563 (n867, n265);
not  g564 (n717, n430);
not  g565 (n640, n461);
buf  g566 (n832, n454);
buf  g567 (n865, n311);
buf  g568 (n892, n308);
buf  g569 (n509, n362);
buf  g570 (n695, n296);
not  g571 (n781, n490);
not  g572 (n850, n387);
buf  g573 (n575, n365);
buf  g574 (n567, n279);
not  g575 (n642, n325);
not  g576 (n802, n354);
buf  g577 (n804, n260);
buf  g578 (n536, n267);
not  g579 (n545, n326);
not  g580 (n539, n251);
buf  g581 (n576, n491);
not  g582 (n566, n426);
buf  g583 (n631, n334);
buf  g584 (n634, n481);
buf  g585 (n864, n289);
not  g586 (n732, n310);
buf  g587 (n905, n385);
not  g588 (n799, n380);
not  g589 (n684, n379);
not  g590 (n818, n442);
not  g591 (n583, n289);
buf  g592 (n839, n318);
not  g593 (n746, n365);
not  g594 (n943, n338);
not  g595 (n803, n280);
buf  g596 (n606, n308);
buf  g597 (n742, n364);
not  g598 (n581, n375);
not  g599 (n713, n348);
buf  g600 (n585, n271);
buf  g601 (n743, n413);
buf  g602 (n779, n297);
not  g603 (n761, n328);
not  g604 (n886, n375);
buf  g605 (n772, n309);
not  g606 (n941, n464);
not  g607 (n608, n266);
not  g608 (n690, n389);
not  g609 (n664, n279);
buf  g610 (n526, n378);
not  g611 (n699, n335);
buf  g612 (n786, n374);
not  g613 (n828, n306);
not  g614 (n829, n255);
not  g615 (n693, n488);
buf  g616 (n598, n485);
buf  g617 (n955, n502);
buf  g618 (n951, n482);
buf  g619 (n530, n309);
buf  g620 (n689, n323);
buf  g621 (n914, n487);
buf  g622 (n911, n491);
not  g623 (n705, n383);
buf  g624 (n618, n398);
not  g625 (n718, n308);
buf  g626 (n927, n276);
buf  g627 (n727, n295);
buf  g628 (n547, n254);
buf  g629 (n548, n307);
buf  g630 (n702, n492);
buf  g631 (n696, n435);
not  g632 (n550, n344);
not  g633 (n855, n315);
buf  g634 (n869, n18);
not  g635 (n593, n379);
buf  g636 (n834, n17);
not  g637 (n745, n270);
buf  g638 (n931, n268);
buf  g639 (n853, n386);
buf  g640 (n674, n252);
not  g641 (n785, n340);
not  g642 (n846, n16);
not  g643 (n656, n356);
buf  g644 (n592, n322);
buf  g645 (n885, n249);
not  g646 (n738, n254);
buf  g647 (n830, n405);
buf  g648 (n597, n391);
buf  g649 (n601, n356);
buf  g650 (n908, n263);
buf  g651 (n963, n282);
buf  g652 (n833, n478);
buf  g653 (n760, n404);
buf  g654 (n815, n492);
not  g655 (n852, n345);
not  g656 (n525, n378);
buf  g657 (n700, n355);
buf  g658 (n944, n399);
not  g659 (n657, n294);
not  g660 (n929, n442);
buf  g661 (n671, n242);
not  g662 (n650, n464);
buf  g663 (n873, n290);
not  g664 (n685, n304);
not  g665 (n714, n17);
not  g666 (n755, n459);
not  g667 (n897, n440);
buf  g668 (n767, n441);
not  g669 (n805, n388);
buf  g670 (n558, n264);
not  g671 (n701, n422);
not  g672 (n748, n352);
buf  g673 (n641, n365);
not  g674 (n546, n448);
not  g675 (n946, n478);
buf  g676 (n639, n288);
buf  g677 (n953, n325);
not  g678 (n898, n17);
not  g679 (n847, n447);
buf  g680 (n512, n309);
buf  g681 (n933, n463);
buf  g682 (n555, n405);
buf  g683 (n591, n306);
not  g684 (n775, n459);
buf  g685 (n744, n498);
not  g686 (n942, n323);
buf  g687 (n794, n463);
buf  g688 (n616, n450);
buf  g689 (n874, n39);
buf  g690 (n809, n347);
not  g691 (n688, n352);
buf  g692 (n615, n462);
not  g693 (n825, n320);
not  g694 (n720, n442);
not  g695 (n707, n295);
not  g696 (n737, n256);
not  g697 (n503, n350);
not  g698 (n920, n246);
buf  g699 (n838, n317);
not  g700 (n570, n294);
not  g701 (n533, n386);
buf  g702 (n921, n476);
buf  g703 (n891, n294);
not  g704 (n800, n304);
not  g705 (n948, n396);
not  g706 (n824, n490);
buf  g707 (n513, n423);
not  g708 (n749, n293);
not  g709 (n949, n450);
buf  g710 (n679, n355);
buf  g711 (n940, n458);
not  g712 (n790, n292);
not  g713 (n677, n413);
buf  g714 (n843, n415);
not  g715 (n645, n385);
buf  g716 (n739, n333);
buf  g717 (n643, n331);
not  g718 (n698, n362);
not  g719 (n814, n499);
not  g720 (n706, n18);
buf  g721 (n894, n282);
not  g722 (n939, n492);
not  g723 (n906, n493);
not  g724 (n777, n342);
buf  g725 (n801, n452);
buf  g726 (n900, n490);
buf  g727 (n957, n501);
not  g728 (n840, n19);
not  g729 (n519, n432);
buf  g730 (n544, n290);
buf  g731 (n543, n253);
buf  g732 (n537, n377);
buf  g733 (n508, n343);
buf  g734 (n907, n486);
buf  g735 (n789, n332);
buf  g736 (n924, n324);
not  g737 (n646, n484);
buf  g738 (n569, n367);
not  g739 (n915, n431);
not  g740 (n868, n323);
not  g741 (n588, n443);
xnor g742 (n596, n298, n348);
nand g743 (n936, n368, n357, n341, n356);
nand g744 (n602, n410, n493, n370, n325);
xor  g745 (n626, n400, n366, n363, n359);
nor  g746 (n932, n424, n435, n247, n482);
and  g747 (n827, n425, n281, n346, n242);
nand g748 (n667, n331, n366, n336, n496);
xor  g749 (n551, n262, n457, n388, n479);
nor  g750 (n883, n350, n421, n414, n392);
xnor g751 (n938, n259, n422, n429, n257);
and  g752 (n826, n375, n270, n420, n429);
and  g753 (n912, n415, n500, n361, n377);
xnor g754 (n511, n438, n405, n39, n428);
and  g755 (n945, n336, n486, n360, n418);
nor  g756 (n532, n351, n291, n253, n274);
and  g757 (n935, n301, n276, n395, n488);
and  g758 (n764, n440, n387, n343, n363);
xnor g759 (n716, n257, n466, n480, n370);
and  g760 (n788, n305, n320, n424, n278);
and  g761 (n622, n380, n252, n495, n17);
and  g762 (n758, n272, n430, n368, n392);
nor  g763 (n750, n342, n357, n437, n355);
nand g764 (n564, n439, n241, n484, n483);
and  g765 (n510, n401, n502, n305, n416);
xnor g766 (n910, n371, n433, n243, n400);
or   g767 (n821, n427, n299, n485, n278);
xor  g768 (n861, n307, n384, n321, n427);
or   g769 (n571, n429, n493, n398);
or   g770 (n604, n295, n340, n302, n258);
nand g771 (n605, n291, n487, n277, n501);
or   g772 (n552, n334, n329, n371, n495);
nand g773 (n860, n440, n263, n393, n500);
nor  g774 (n603, n290, n252, n269, n258);
nand g775 (n623, n412, n428, n335, n367);
nor  g776 (n556, n359, n245, n447, n329);
nand g777 (n934, n286, n462, n403, n371);
nand g778 (n782, n353, n465, n268, n285);
nand g779 (n730, n407, n305, n446, n462);
nand g780 (n735, n474, n354, n477, n351);
and  g781 (n531, n445, n258, n491, n343);
or   g782 (n620, n465, n401, n427, n246);
xor  g783 (n902, n319, n341, n387, n490);
nor  g784 (n573, n473, n481, n393, n461);
and  g785 (n947, n451, n367, n352, n260);
and  g786 (n527, n322, n395, n423, n460);
nand g787 (n769, n409, n424, n410, n342);
xnor g788 (n928, n251, n261, n466, n285);
and  g789 (n816, n287, n281, n494, n316);
xnor g790 (n712, n498, n425, n386, n369);
xor  g791 (n635, n482, n468, n285, n280);
nor  g792 (n572, n262, n309, n340, n440);
xor  g793 (n889, n284, n287, n419, n426);
xnor g794 (n880, n477, n385, n283, n404);
and  g795 (n683, n286, n481, n349, n288);
and  g796 (n965, n393, n480, n477, n470);
nand g797 (n669, n273, n409, n394, n470);
xor  g798 (n568, n306, n354, n313, n345);
nand g799 (n580, n288, n470, n417, n497);
nand g800 (n844, n288, n303, n439, n275);
xor  g801 (n771, n337, n273, n326, n500);
xor  g802 (n866, n412, n311, n262, n270);
or   g803 (n565, n435, n411, n473, n331);
and  g804 (n751, n461, n349, n329, n366);
xor  g805 (n586, n349, n416, n265, n418);
nand g806 (n563, n394, n256, n258, n415);
xnor g807 (n875, n424, n491, n352, n414);
or   g808 (n589, n468, n460, n343, n313);
or   g809 (n708, n406, n405, n332, n336);
or   g810 (n863, n416, n437, n403, n419);
nor  g811 (n922, n330, n327, n277, n339);
nand g812 (n950, n271, n346, n318, n410);
or   g813 (n797, n267, n396, n334, n353);
and  g814 (n515, n437, n472, n257, n391);
or   g815 (n806, n250, n486, n398, n358);
nand g816 (n817, n255, n331, n303, n423);
nor  g817 (n595, n407, n264, n313, n426);
nor  g818 (n926, n260, n397, n243, n422);
xnor g819 (n791, n292, n328, n448, n314);
xor  g820 (n877, n251, n254, n249, n322);
xor  g821 (n960, n432, n357, n389, n449);
nor  g822 (n636, n381, n341, n407, n496);
nor  g823 (n600, n421, n446, n346, n403);
or   g824 (n582, n397, n452, n484, n383);
nor  g825 (n516, n457, n319, n434, n360);
nand g826 (n837, n500, n428, n442, n411);
xor  g827 (n561, n391, n453, n378, n298);
and  g828 (n666, n377, n454, n374, n381);
nand g829 (n710, n362, n335, n372, n497);
nand g830 (n878, n373, n274, n291, n471);
or   g831 (n711, n269, n456, n262, n266);
and  g832 (n752, n447, n276, n271, n468);
xnor g833 (n857, n432, n253, n324, n314);
nor  g834 (n517, n315, n321, n299, n479);
xnor g835 (n958, n282, n419, n346, n370);
and  g836 (n773, n416, n466, n301, n383);
or   g837 (n807, n363, n489, n360, n268);
nand g838 (n651, n383, n320, n418, n420);
nor  g839 (n734, n255, n364, n347, n289);
nand g840 (n520, n297, n449, n314, n379);
or   g841 (n668, n487, n441, n443, n369);
nand g842 (n630, n316, n380, n353, n399);
or   g843 (n754, n444, n270, n430, n389);
xnor g844 (n655, n499, n387, n324, n275);
xnor g845 (n903, n265, n437, n469, n285);
and  g846 (n632, n420, n464, n485, n399);
nor  g847 (n909, n354, n489, n396, n317);
xor  g848 (n562, n470, n496, n349, n361);
or   g849 (n741, n439, n263, n372, n394);
xor  g850 (n918, n444, n487, n295, n368);
xor  g851 (n660, n376, n286, n254, n492);
and  g852 (n884, n384, n333, n350, n361);
nand g853 (n610, n330, n404, n436, n336);
nand g854 (n836, n460, n372, n392, n248);
or   g855 (n624, n444, n333, n496, n322);
nor  g856 (n694, n16, n358, n244, n401);
nand g857 (n901, n473, n307, n373, n406);
and  g858 (n768, n436, n431, n330, n402);
xor  g859 (n523, n245, n266, n296, n450);
and  g860 (n553, n438, n364, n479, n388);
or   g861 (n505, n339, n465, n247, n451);
xnor g862 (n822, n328, n445, n427, n391);
and  g863 (n628, n327, n364, n301, n247);
or   g864 (n952, n356, n351, n337, n481);
xor  g865 (n648, n425, n256, n414, n249);
and  g866 (n611, n319, n422, n438, n358);
nand g867 (n956, n292, n448, n269, n497);
xor  g868 (n638, n373, n501, n311, n280);
xnor g869 (n529, n328, n456, n399, n256);
xnor g870 (n930, n426, n494, n264, n448);
xnor g871 (n778, n459, n303, n434, n339);
or   g872 (n507, n296, n402, n287, n289);
nand g873 (n723, n472, n272, n277, n244);
xor  g874 (n524, n483, n369, n480, n283);
nand g875 (n663, n443, n459, n316, n445);
xor  g876 (n557, n460, n259, n395, n474);
nor  g877 (n937, n458, n347, n281, n400);
or   g878 (n919, n455, n408, n465, n499);
or   g879 (n848, n304, n351, n392, n488);
xnor g880 (n882, n318, n259, n269, n475);
nand g881 (n759, n475, n39, n406, n489);
nand g882 (n820, n338, n432, n433, n483);
nor  g883 (n627, n287, n311, n332, n330);
nor  g884 (n813, n434, n494, n464, n446);
or   g885 (n736, n453, n271, n457, n340);
xor  g886 (n812, n292, n257, n324, n314);
xor  g887 (n659, n407, n293, n390, n333);
nor  g888 (n916, n300, n347, n406, n371);
or   g889 (n680, n434, n325, n372, n267);
xnor g890 (n658, n307, n458, n462, n265);
xor  g891 (n896, n456, n286, n431, n344);
xnor g892 (n763, n421, n498, n19, n469);
xnor g893 (n795, n410, n495, n381, n279);
xor  g894 (n678, n348, n291, n260, n390);
and  g895 (n774, n476, n316, n359, n350);
nor  g896 (n560, n429, n358, n420, n390);
nand g897 (n692, n384, n318, n275, n430);
nand g898 (n811, n317, n357, n474, n370);
nor  g899 (n506, n475, n376, n339, n402);
xor  g900 (n793, n353, n297, n451, n369);
xor  g901 (n881, n293, n282, n396, n244);
xnor g902 (n726, n393, n398, n304, n335);
or   g903 (n687, n274, n438, n253, n453);
nand g904 (n535, n376, n327, n263, n284);
nand g905 (n672, n241, n417, n382, n455);
xnor g906 (n835, n468, n312, n294, n321);
and  g907 (n893, n319, n455, n290, n471);
nand g908 (n621, n467, n473, n478, n302);
xor  g909 (n577, n261, n457, n409, n441);
xor  g910 (n686, n243, n361, n272, n449);
nand g911 (n862, n486, n408, n268);
nor  g912 (n661, n480, n433, n418, n300);
nor  g913 (n890, n315, n401, n366, n502);
xnor g914 (n876, n332, n280, n278, n467);
or   g915 (n554, n474, n450, n255, n246);
nand g916 (n578, n453, n306, n463, n394);
xor  g917 (n665, n471, n310, n447, n428);
and  g918 (n784, n365, n415, n355, n466);
xor  g919 (n849, n362, n375, n382, n435);
nor  g920 (n619, n454, n312, n39, n310);
xor  g921 (n871, n359, n274, n300, n242);
xnor g922 (n504, n463, n382, n297, n439);
nand g923 (n851, n378, n326, n452, n436);
nor  g924 (n959, n326, n472, n388, n444);
and  g925 (n787, n315, n502, n455, n478);
and  g926 (n923, n467, n449, n381, n278);
or   g927 (n856, n275, n250, n264, n298);
xor  g928 (n753, n377, n501, n436, n397);
xnor g929 (n538, n261, n425, n445, n284);
xor  g930 (n819, n412, n476, n384, n413);
nand g931 (n599, n284, n433, n310, n261);
xor  g932 (n731, n489, n385, n414, n494);
xnor g933 (n719, n252, n412, n386, n298);
xnor g934 (n676, n404, n302, n334, n338);
nor  g935 (n653, n379, n266, n345, n431);
or   g936 (n629, n321, n373, n467, n283);
or   g937 (n756, n293, n276, n484, n273);
nor  g938 (n709, n497, n499, n327, n469);
xnor g939 (n594, n395, n305, n451, n301);
xnor g940 (n1065, n964, n676, n796, n761);
xnor g941 (n1015, n520, n632, n963, n829);
xnor g942 (n1011, n954, n755, n546, n771);
or   g943 (n966, n673, n619, n898, n798);
nand g944 (n1071, n887, n958, n665, n578);
xnor g945 (n1080, n651, n772, n835, n960);
nor  g946 (n1035, n884, n911, n720, n633);
xor  g947 (n1009, n932, n569, n856, n737);
xor  g948 (n1068, n740, n641, n852, n838);
xnor g949 (n1063, n751, n645, n853, n843);
and  g950 (n1000, n913, n867, n515, n945);
or   g951 (n986, n809, n621, n612, n953);
nor  g952 (n968, n734, n817, n943, n821);
nand g953 (n1029, n560, n675, n758, n618);
xor  g954 (n970, n699, n568, n797, n636);
nor  g955 (n1053, n875, n625, n775, n731);
xor  g956 (n1008, n959, n929, n643, n690);
nor  g957 (n1023, n837, n869, n537, n539);
xnor g958 (n1039, n600, n886, n890, n799);
or   g959 (n1042, n519, n629, n790, n933);
nand g960 (n1046, n710, n698, n759, n601);
or   g961 (n1083, n942, n963, n711, n514);
or   g962 (n1005, n536, n604, n779, n727);
xnor g963 (n1075, n679, n575, n635, n952);
and  g964 (n1062, n693, n926, n548, n683);
xor  g965 (n1041, n812, n895, n824, n791);
xnor g966 (n1051, n879, n605, n940, n802);
xor  g967 (n1048, n844, n863, n777, n792);
nand g968 (n981, n544, n707, n960, n881);
and  g969 (n1001, n672, n860, n505, n961);
nor  g970 (n1074, n834, n658, n778, n573);
and  g971 (n1076, n677, n717, n756, n745);
nor  g972 (n1081, n598, n811, n893, n752);
nand g973 (n1037, n694, n614, n748, n735);
nand g974 (n987, n814, n706, n764, n511);
xor  g975 (n974, n905, n956, n729, n701);
and  g976 (n980, n522, n868, n800, n883);
xnor g977 (n994, n577, n934, n552, n957);
xnor g978 (n998, n921, n611, n521, n682);
xnor g979 (n1034, n718, n902, n785, n702);
or   g980 (n1020, n556, n565, n857, n832);
nand g981 (n989, n557, n849, n616, n951);
xor  g982 (n1047, n649, n958, n674, n566);
and  g983 (n977, n874, n916, n952, n613);
xnor g984 (n1066, n754, n965, n610, n789);
xnor g985 (n1018, n864, n634, n862, n527);
nand g986 (n973, n769, n762, n508, n586);
nor  g987 (n991, n558, n816, n554, n861);
xnor g988 (n1033, n736, n591, n647, n846);
nand g989 (n1030, n813, n962, n786, n865);
or   g990 (n992, n845, n903, n750, n631);
nand g991 (n1043, n794, n908, n526, n739);
or   g992 (n978, n741, n842, n815, n776);
xnor g993 (n1010, n553, n551, n766, n582);
xnor g994 (n1038, n770, n581, n545, n685);
nor  g995 (n995, n839, n939, n567, n744);
xor  g996 (n1070, n584, n650, n697, n946);
xnor g997 (n1024, n962, n877, n858, n657);
or   g998 (n997, n836, n851, n607, n914);
nand g999 (n1077, n524, n894, n725, n507);
nand g1000 (n1028, n630, n904, n572, n746);
nor  g1001 (n975, n749, n826, n922, n543);
or   g1002 (n976, n724, n555, n599, n804);
xnor g1003 (n1002, n823, n620, n708, n907);
xnor g1004 (n999, n892, n660, n924, n954);
nand g1005 (n1049, n533, n955, n885, n589);
xnor g1006 (n1016, n595, n623, n918, n965);
or   g1007 (n1055, n678, n882, n803, n901);
nand g1008 (n1058, n726, n959, n593, n767);
nor  g1009 (n1012, n615, n663, n847, n506);
or   g1010 (n1027, n805, n587, n897, n841);
and  g1011 (n1054, n850, n757, n919, n900);
xor  g1012 (n1013, n656, n781, n912, n585);
or   g1013 (n1006, n529, n733, n662, n906);
and  g1014 (n1064, n518, n563, n872, n655);
nor  g1015 (n1079, n628, n878, n760, n590);
xor  g1016 (n1044, n580, n542, n525, n915);
or   g1017 (n1007, n592, n859, n899, n774);
and  g1018 (n1014, n602, n531, n541, n828);
xor  g1019 (n1040, n889, n719, n747, n638);
xor  g1020 (n1073, n583, n920, n876, n936);
or   g1021 (n1082, n705, n830, n788, n855);
and  g1022 (n1022, n848, n709, n671, n571);
xor  g1023 (n988, n528, n696, n576, n550);
xor  g1024 (n1067, n715, n941, n810, n742);
nor  g1025 (n1069, n603, n723, n646, n949);
nor  g1026 (n1057, n637, n819, n686, n820);
xor  g1027 (n971, n961, n948, n609, n784);
xnor g1028 (n996, n668, n654, n714, n669);
or   g1029 (n1031, n753, n938, n713, n688);
nor  g1030 (n1004, n953, n806, n680, n574);
xnor g1031 (n1050, n763, n930, n866, n523);
nor  g1032 (n993, n666, n642, n597, n831);
nand g1033 (n1036, n570, n712, n782, n854);
xnor g1034 (n1017, n716, n738, n684, n722);
and  g1035 (n1072, n562, n691, n925, n703);
or   g1036 (n984, n670, n534, n937, n549);
or   g1037 (n967, n957, n822, n639, n773);
and  g1038 (n990, n840, n516, n743, n538);
xnor g1039 (n985, n730, n692, n644, n765);
xor  g1040 (n1003, n659, n917, n513, n579);
xor  g1041 (n1026, n624, n667, n808, n928);
nor  g1042 (n983, n880, n964, n653, n947);
and  g1043 (n972, n732, n594, n910, n956);
nand g1044 (n969, n931, n768, n535, n661);
or   g1045 (n979, n721, n695, n681, n728);
nor  g1046 (n1032, n873, n532, n807, n588);
and  g1047 (n982, n564, n617, n783, n793);
xor  g1048 (n1045, n935, n627, n704, n801);
xor  g1049 (n1060, n606, n825, n795, n559);
xor  g1050 (n1056, n787, n504, n871, n512);
or   g1051 (n1021, n664, n944, n780, n626);
nor  g1052 (n1084, n608, n888, n510, n540);
nand g1053 (n1052, n640, n833, n909, n517);
or   g1054 (n1078, n891, n927, n870, n530);
xnor g1055 (n1061, n955, n827, n547, n596);
nor  g1056 (n1059, n509, n622, n648, n923);
xnor g1057 (n1025, n818, n689, n896, n561);
or   g1058 (n1019, n950, n700, n652, n687);
nand g1059 (n1111, n990, n1051, n1079, n1015);
xnor g1060 (n1110, n1040, n1034, n1035, n974);
xor  g1061 (n1091, n1066, n1064, n1020, n1014);
nand g1062 (n1101, n1003, n1000, n1036, n1056);
or   g1063 (n1106, n1065, n1010, n1026, n1002);
or   g1064 (n1100, n994, n1012, n979, n1021);
nand g1065 (n1094, n1080, n1068, n1075, n1022);
nor  g1066 (n1109, n1057, n1071, n1006, n986);
xor  g1067 (n1112, n969, n995, n1031, n1039);
or   g1068 (n1095, n968, n981, n1044, n1053);
or   g1069 (n1087, n1050, n989, n996, n966);
xor  g1070 (n1108, n1063, n1058, n1009, n988);
xor  g1071 (n1104, n1073, n1016, n1025, n1052);
and  g1072 (n1092, n978, n997, n1061, n1028);
xor  g1073 (n1088, n1024, n980, n1011, n1019);
nor  g1074 (n1090, n973, n1005, n1042, n971);
nand g1075 (n1085, n1017, n972, n1033, n1077);
nor  g1076 (n1089, n998, n1037, n1008, n967);
xnor g1077 (n1096, n1067, n1004, n991, n1018);
nor  g1078 (n1093, n1007, n1046, n985, n1001);
nand g1079 (n1097, n1072, n970, n1029, n1070);
xnor g1080 (n1105, n1043, n1060, n987, n1048);
xnor g1081 (n1103, n983, n1013, n993, n984);
xnor g1082 (n1102, n992, n1059, n1030, n976);
xor  g1083 (n1113, n1081, n1078, n1049, n975);
and  g1084 (n1107, n1076, n977, n1027, n1069);
nor  g1085 (n1099, n1045, n1047, n1032, n1062);
nor  g1086 (n1086, n999, n1023, n982, n1041);
nand g1087 (n1098, n1054, n1038, n1055, n1074);
xor  g1088 (n1123, n24, n58, n25, n1111);
or   g1089 (n1121, n21, n21, n25, n20);
and  g1090 (n1125, n23, n22, n57);
nor  g1091 (n1122, n1110, n23, n20, n24);
xor  g1092 (n1119, n1097, n1102, n1107, n19);
nand g1093 (n1118, n1105, n58, n1104, n1098);
nand g1094 (n1117, n1100, n23, n19);
nand g1095 (n1115, n1103, n22, n57);
nand g1096 (n1120, n25, n20, n58, n1099);
xnor g1097 (n1116, n21, n1112, n1108, n25);
xnor g1098 (n1124, n1106, n1109, n24, n1101);
xnor g1099 (n1114, n21, n20, n1113, n24);
buf  g1100 (n1129, n1114);
not  g1101 (n1127, n1115);
or   g1102 (n1128, n1118, n1117, n1115, n1114);
xnor g1103 (n1130, n1118, n1115, n1116, n1117);
xor  g1104 (n1126, n1114, n1116, n1117);
and  g1105 (n1132, n1119, n1127, n1118);
and  g1106 (n1138, n1128, n1127, n1084, n1126);
xnor g1107 (n1136, n1130, n1126, n1129, n1127);
nor  g1108 (n1133, n1126, n1128, n1129, n1118);
nor  g1109 (n1135, n1120, n1129, n1130);
nor  g1110 (n1131, n1128, n1119, n1083);
xor  g1111 (n1137, n1120, n1119, n1082, n1126);
or   g1112 (n1134, n1130, n1129, n1120, n1128);
xor  g1113 (n1139, n1120, n1123, n1122, n1121);
xor  g1114 (n1141, n1123, n1122, n1121);
or   g1115 (n1142, n1121, n1122, n1137, n1125);
xor  g1116 (n1144, n1121, n1124, n1125);
or   g1117 (n1140, n1123, n1134, n1125, n1133);
nor  g1118 (n1145, n1125, n1136, n1124, n1123);
and  g1119 (n1143, n1135, n1132, n1138, n1124);
endmodule
