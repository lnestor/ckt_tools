

module Stat_2000_224
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1188,
  n1172,
  n1175,
  n1185,
  n1170,
  n1183,
  n1181,
  n1171,
  n1182,
  n1189,
  n1190,
  n1213,
  n1215,
  n1221,
  n1250,
  n1246,
  n1243,
  n1249,
  n1238,
  n1257,
  n1236,
  n1237,
  n1248,
  n1244,
  n1256,
  n1254,
  n1245,
  n1247,
  n1240,
  n1242,
  n2031,
  n2032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n1188;
  output n1172;
  output n1175;
  output n1185;
  output n1170;
  output n1183;
  output n1181;
  output n1171;
  output n1182;
  output n1189;
  output n1190;
  output n1213;
  output n1215;
  output n1221;
  output n1250;
  output n1246;
  output n1243;
  output n1249;
  output n1238;
  output n1257;
  output n1236;
  output n1237;
  output n1248;
  output n1244;
  output n1256;
  output n1254;
  output n1245;
  output n1247;
  output n1240;
  output n1242;
  output n2031;
  output n2032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1173;
  wire n1174;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1184;
  wire n1186;
  wire n1187;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1214;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1239;
  wire n1241;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1255;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    n112,
    n14
  );


  not
  g1
  (
    n148,
    n23
  );


  buf
  g2
  (
    n81,
    n12
  );


  not
  g3
  (
    n83,
    n26
  );


  not
  g4
  (
    n58,
    n27
  );


  not
  g5
  (
    n119,
    n20
  );


  buf
  g6
  (
    n107,
    n19
  );


  buf
  g7
  (
    n137,
    n4
  );


  not
  g8
  (
    n141,
    n27
  );


  not
  g9
  (
    n86,
    n9
  );


  buf
  g10
  (
    n149,
    n7
  );


  buf
  g11
  (
    n48,
    n18
  );


  buf
  g12
  (
    n153,
    n28
  );


  not
  g13
  (
    n96,
    n24
  );


  not
  g14
  (
    n90,
    n28
  );


  buf
  g15
  (
    n37,
    n16
  );


  buf
  g16
  (
    n118,
    n7
  );


  buf
  g17
  (
    n70,
    n14
  );


  not
  g18
  (
    n139,
    n21
  );


  buf
  g19
  (
    n125,
    n8
  );


  not
  g20
  (
    n134,
    n31
  );


  buf
  g21
  (
    n129,
    n29
  );


  not
  g22
  (
    n72,
    n21
  );


  not
  g23
  (
    n79,
    n24
  );


  buf
  g24
  (
    KeyWire_0_31,
    n23
  );


  buf
  g25
  (
    n126,
    n16
  );


  not
  g26
  (
    n66,
    n10
  );


  not
  g27
  (
    n136,
    n19
  );


  buf
  g28
  (
    n142,
    n1
  );


  not
  g29
  (
    n65,
    n28
  );


  buf
  g30
  (
    n52,
    n25
  );


  buf
  g31
  (
    n111,
    n29
  );


  not
  g32
  (
    n133,
    n32
  );


  buf
  g33
  (
    n150,
    n22
  );


  not
  g34
  (
    n109,
    n20
  );


  buf
  g35
  (
    n120,
    n30
  );


  buf
  g36
  (
    n108,
    n23
  );


  not
  g37
  (
    n44,
    n20
  );


  buf
  g38
  (
    n53,
    n12
  );


  buf
  g39
  (
    n97,
    n32
  );


  buf
  g40
  (
    n159,
    n8
  );


  buf
  g41
  (
    n75,
    n5
  );


  buf
  g42
  (
    n144,
    n2
  );


  buf
  g43
  (
    n87,
    n26
  );


  not
  g44
  (
    n45,
    n28
  );


  buf
  g45
  (
    n122,
    n19
  );


  buf
  g46
  (
    n95,
    n18
  );


  not
  g47
  (
    n131,
    n10
  );


  not
  g48
  (
    n84,
    n25
  );


  not
  g49
  (
    n101,
    n16
  );


  buf
  g50
  (
    n41,
    n2
  );


  not
  g51
  (
    n33,
    n6
  );


  not
  g52
  (
    n39,
    n9
  );


  buf
  g53
  (
    n103,
    n18
  );


  buf
  g54
  (
    n82,
    n19
  );


  buf
  g55
  (
    n35,
    n15
  );


  buf
  g56
  (
    n110,
    n5
  );


  buf
  g57
  (
    n123,
    n16
  );


  not
  g58
  (
    n38,
    n24
  );


  buf
  g59
  (
    n61,
    n27
  );


  not
  g60
  (
    n68,
    n4
  );


  not
  g61
  (
    n105,
    n3
  );


  not
  g62
  (
    n124,
    n26
  );


  buf
  g63
  (
    n130,
    n11
  );


  not
  g64
  (
    n56,
    n29
  );


  buf
  g65
  (
    n73,
    n13
  );


  not
  g66
  (
    n51,
    n13
  );


  not
  g67
  (
    n47,
    n24
  );


  not
  g68
  (
    n115,
    n14
  );


  buf
  g69
  (
    n100,
    n17
  );


  buf
  g70
  (
    n76,
    n25
  );


  not
  g71
  (
    n121,
    n31
  );


  buf
  g72
  (
    n155,
    n17
  );


  buf
  g73
  (
    n55,
    n30
  );


  buf
  g74
  (
    n102,
    n9
  );


  buf
  g75
  (
    n98,
    n1
  );


  not
  g76
  (
    n138,
    n9
  );


  not
  g77
  (
    n40,
    n17
  );


  buf
  g78
  (
    n154,
    n11
  );


  not
  g79
  (
    n117,
    n10
  );


  buf
  g80
  (
    n34,
    n1
  );


  not
  g81
  (
    n157,
    n32
  );


  buf
  g82
  (
    n89,
    n6
  );


  not
  g83
  (
    n160,
    n6
  );


  not
  g84
  (
    n74,
    n32
  );


  buf
  g85
  (
    n146,
    n12
  );


  buf
  g86
  (
    n104,
    n26
  );


  buf
  g87
  (
    n88,
    n17
  );


  buf
  g88
  (
    n85,
    n8
  );


  not
  g89
  (
    n60,
    n30
  );


  buf
  g90
  (
    n94,
    n10
  );


  buf
  g91
  (
    n106,
    n21
  );


  not
  g92
  (
    n127,
    n13
  );


  buf
  g93
  (
    n140,
    n22
  );


  not
  g94
  (
    n49,
    n4
  );


  buf
  g95
  (
    n63,
    n22
  );


  not
  g96
  (
    n69,
    n8
  );


  not
  g97
  (
    n147,
    n5
  );


  not
  g98
  (
    n77,
    n5
  );


  buf
  g99
  (
    n92,
    n15
  );


  buf
  g100
  (
    n59,
    n31
  );


  buf
  g101
  (
    n151,
    n18
  );


  buf
  g102
  (
    n152,
    n25
  );


  not
  g103
  (
    n116,
    n20
  );


  buf
  g104
  (
    n64,
    n7
  );


  not
  g105
  (
    n54,
    n31
  );


  not
  g106
  (
    n93,
    n23
  );


  not
  g107
  (
    n50,
    n15
  );


  not
  g108
  (
    n71,
    n14
  );


  buf
  g109
  (
    n158,
    n30
  );


  not
  g110
  (
    KeyWire_0_22,
    n21
  );


  not
  g111
  (
    n62,
    n2
  );


  not
  g112
  (
    n67,
    n22
  );


  buf
  g113
  (
    n57,
    n3
  );


  buf
  g114
  (
    n113,
    n11
  );


  buf
  g115
  (
    n80,
    n12
  );


  buf
  g116
  (
    n46,
    n13
  );


  buf
  g117
  (
    n143,
    n11
  );


  buf
  g118
  (
    n114,
    n1
  );


  not
  g119
  (
    n145,
    n27
  );


  buf
  g120
  (
    n99,
    n4
  );


  not
  g121
  (
    n42,
    n3
  );


  not
  g122
  (
    n128,
    n29
  );


  buf
  g123
  (
    n135,
    n15
  );


  buf
  g124
  (
    n78,
    n3
  );


  buf
  g125
  (
    n43,
    n2
  );


  buf
  g126
  (
    n156,
    n6
  );


  not
  g127
  (
    n36,
    n7
  );


  buf
  g128
  (
    n295,
    n37
  );


  buf
  g129
  (
    n243,
    n136
  );


  not
  g130
  (
    n375,
    n129
  );


  not
  g131
  (
    n248,
    n70
  );


  buf
  g132
  (
    n489,
    n45
  );


  buf
  g133
  (
    n550,
    n84
  );


  buf
  g134
  (
    n214,
    n127
  );


  not
  g135
  (
    n250,
    n48
  );


  buf
  g136
  (
    n434,
    n100
  );


  not
  g137
  (
    n176,
    n58
  );


  buf
  g138
  (
    n168,
    n131
  );


  not
  g139
  (
    n480,
    n137
  );


  not
  g140
  (
    n535,
    n44
  );


  buf
  g141
  (
    n445,
    n115
  );


  not
  g142
  (
    n408,
    n111
  );


  buf
  g143
  (
    n513,
    n87
  );


  buf
  g144
  (
    n310,
    n66
  );


  buf
  g145
  (
    KeyWire_0_3,
    n108
  );


  buf
  g146
  (
    n567,
    n74
  );


  not
  g147
  (
    n163,
    n58
  );


  buf
  g148
  (
    n554,
    n47
  );


  buf
  g149
  (
    n350,
    n125
  );


  not
  g150
  (
    n270,
    n117
  );


  buf
  g151
  (
    n274,
    n135
  );


  buf
  g152
  (
    n210,
    n35
  );


  not
  g153
  (
    n212,
    n102
  );


  buf
  g154
  (
    n558,
    n55
  );


  not
  g155
  (
    n297,
    n51
  );


  not
  g156
  (
    n486,
    n42
  );


  not
  g157
  (
    n429,
    n40
  );


  buf
  g158
  (
    n303,
    n101
  );


  buf
  g159
  (
    n583,
    n69
  );


  not
  g160
  (
    n230,
    n89
  );


  buf
  g161
  (
    n478,
    n84
  );


  not
  g162
  (
    n406,
    n98
  );


  buf
  g163
  (
    n271,
    n56
  );


  buf
  g164
  (
    n544,
    n67
  );


  buf
  g165
  (
    n484,
    n92
  );


  buf
  g166
  (
    n397,
    n65
  );


  not
  g167
  (
    n525,
    n112
  );


  buf
  g168
  (
    n213,
    n37
  );


  buf
  g169
  (
    n342,
    n117
  );


  not
  g170
  (
    n263,
    n110
  );


  buf
  g171
  (
    n341,
    n127
  );


  buf
  g172
  (
    n343,
    n46
  );


  buf
  g173
  (
    n430,
    n61
  );


  not
  g174
  (
    n469,
    n136
  );


  buf
  g175
  (
    n379,
    n94
  );


  not
  g176
  (
    n336,
    n113
  );


  not
  g177
  (
    n215,
    n39
  );


  buf
  g178
  (
    n587,
    n44
  );


  buf
  g179
  (
    n333,
    n70
  );


  buf
  g180
  (
    n165,
    n38
  );


  not
  g181
  (
    n519,
    n54
  );


  buf
  g182
  (
    n338,
    n129
  );


  not
  g183
  (
    n348,
    n141
  );


  buf
  g184
  (
    n461,
    n60
  );


  not
  g185
  (
    n533,
    n64
  );


  buf
  g186
  (
    n334,
    n87
  );


  not
  g187
  (
    n296,
    n45
  );


  not
  g188
  (
    n439,
    n83
  );


  buf
  g189
  (
    n288,
    n137
  );


  buf
  g190
  (
    n417,
    n130
  );


  not
  g191
  (
    n547,
    n128
  );


  buf
  g192
  (
    n565,
    n49
  );


  not
  g193
  (
    n265,
    n115
  );


  not
  g194
  (
    n532,
    n95
  );


  buf
  g195
  (
    n398,
    n119
  );


  not
  g196
  (
    n409,
    n81
  );


  buf
  g197
  (
    n233,
    n76
  );


  buf
  g198
  (
    n352,
    n95
  );


  not
  g199
  (
    n185,
    n108
  );


  buf
  g200
  (
    n292,
    n101
  );


  not
  g201
  (
    n568,
    n51
  );


  buf
  g202
  (
    n247,
    n111
  );


  not
  g203
  (
    n449,
    n76
  );


  not
  g204
  (
    n440,
    n38
  );


  not
  g205
  (
    n290,
    n79
  );


  buf
  g206
  (
    n471,
    n125
  );


  not
  g207
  (
    n563,
    n35
  );


  not
  g208
  (
    n592,
    n52
  );


  buf
  g209
  (
    n476,
    n130
  );


  not
  g210
  (
    n171,
    n133
  );


  not
  g211
  (
    n238,
    n133
  );


  not
  g212
  (
    n386,
    n57
  );


  not
  g213
  (
    n252,
    n132
  );


  buf
  g214
  (
    n428,
    n35
  );


  buf
  g215
  (
    n380,
    n114
  );


  buf
  g216
  (
    KeyWire_0_2,
    n121
  );


  not
  g217
  (
    n289,
    n93
  );


  buf
  g218
  (
    n578,
    n131
  );


  buf
  g219
  (
    n531,
    n106
  );


  not
  g220
  (
    n528,
    n118
  );


  not
  g221
  (
    n359,
    n122
  );


  not
  g222
  (
    n282,
    n80
  );


  buf
  g223
  (
    n521,
    n93
  );


  buf
  g224
  (
    n382,
    n127
  );


  buf
  g225
  (
    n421,
    n42
  );


  not
  g226
  (
    n574,
    n75
  );


  not
  g227
  (
    n362,
    n139
  );


  not
  g228
  (
    n317,
    n102
  );


  buf
  g229
  (
    n518,
    n86
  );


  not
  g230
  (
    n340,
    n99
  );


  not
  g231
  (
    n401,
    n33
  );


  not
  g232
  (
    n197,
    n135
  );


  buf
  g233
  (
    n299,
    n108
  );


  buf
  g234
  (
    n335,
    n135
  );


  not
  g235
  (
    n387,
    n97
  );


  buf
  g236
  (
    n242,
    n39
  );


  buf
  g237
  (
    n451,
    n56
  );


  not
  g238
  (
    n351,
    n139
  );


  not
  g239
  (
    n400,
    n103
  );


  buf
  g240
  (
    n231,
    n41
  );


  buf
  g241
  (
    n321,
    n36
  );


  buf
  g242
  (
    n306,
    n69
  );


  buf
  g243
  (
    n177,
    n88
  );


  not
  g244
  (
    n552,
    n86
  );


  buf
  g245
  (
    n260,
    n122
  );


  not
  g246
  (
    n229,
    n49
  );


  buf
  g247
  (
    KeyWire_0_27,
    n126
  );


  buf
  g248
  (
    n376,
    n72
  );


  buf
  g249
  (
    n286,
    n66
  );


  not
  g250
  (
    n576,
    n61
  );


  buf
  g251
  (
    n183,
    n94
  );


  not
  g252
  (
    n508,
    n88
  );


  not
  g253
  (
    n354,
    n90
  );


  not
  g254
  (
    n259,
    n59
  );


  buf
  g255
  (
    n545,
    n116
  );


  buf
  g256
  (
    n371,
    n116
  );


  not
  g257
  (
    n251,
    n36
  );


  buf
  g258
  (
    n581,
    n87
  );


  buf
  g259
  (
    n236,
    n78
  );


  buf
  g260
  (
    n169,
    n36
  );


  not
  g261
  (
    n447,
    n137
  );


  buf
  g262
  (
    n542,
    n69
  );


  not
  g263
  (
    n302,
    n119
  );


  buf
  g264
  (
    KeyWire_0_23,
    n127
  );


  not
  g265
  (
    n590,
    n100
  );


  not
  g266
  (
    n173,
    n34
  );


  not
  g267
  (
    n355,
    n139
  );


  not
  g268
  (
    n249,
    n93
  );


  not
  g269
  (
    n194,
    n48
  );


  buf
  g270
  (
    n239,
    n140
  );


  buf
  g271
  (
    n524,
    n86
  );


  buf
  g272
  (
    n497,
    n43
  );


  not
  g273
  (
    n534,
    n107
  );


  buf
  g274
  (
    n457,
    n78
  );


  buf
  g275
  (
    n232,
    n105
  );


  buf
  g276
  (
    n298,
    n134
  );


  not
  g277
  (
    n385,
    n50
  );


  not
  g278
  (
    n283,
    n124
  );


  not
  g279
  (
    n422,
    n47
  );


  buf
  g280
  (
    n224,
    n93
  );


  buf
  g281
  (
    n276,
    n126
  );


  buf
  g282
  (
    n418,
    n107
  );


  not
  g283
  (
    n312,
    n64
  );


  buf
  g284
  (
    n579,
    n65
  );


  not
  g285
  (
    n218,
    n83
  );


  not
  g286
  (
    n394,
    n106
  );


  buf
  g287
  (
    n227,
    n85
  );


  not
  g288
  (
    n483,
    n51
  );


  buf
  g289
  (
    n217,
    n66
  );


  buf
  g290
  (
    n284,
    n57
  );


  buf
  g291
  (
    n506,
    n52
  );


  not
  g292
  (
    n204,
    n59
  );


  not
  g293
  (
    n589,
    n59
  );


  not
  g294
  (
    n586,
    n75
  );


  not
  g295
  (
    n569,
    n84
  );


  not
  g296
  (
    n555,
    n34
  );


  buf
  g297
  (
    n370,
    n133
  );


  not
  g298
  (
    n221,
    n34
  );


  buf
  g299
  (
    n501,
    n130
  );


  buf
  g300
  (
    n455,
    n74
  );


  buf
  g301
  (
    n209,
    n112
  );


  buf
  g302
  (
    n211,
    n41
  );


  not
  g303
  (
    n245,
    n54
  );


  not
  g304
  (
    n325,
    n46
  );


  not
  g305
  (
    n487,
    n117
  );


  not
  g306
  (
    n454,
    n47
  );


  buf
  g307
  (
    n395,
    n134
  );


  not
  g308
  (
    n237,
    n107
  );


  buf
  g309
  (
    n553,
    n47
  );


  buf
  g310
  (
    n437,
    n115
  );


  buf
  g311
  (
    n328,
    n82
  );


  buf
  g312
  (
    n548,
    n79
  );


  buf
  g313
  (
    n320,
    n109
  );


  not
  g314
  (
    n186,
    n36
  );


  not
  g315
  (
    n369,
    n75
  );


  buf
  g316
  (
    n361,
    n106
  );


  not
  g317
  (
    n436,
    n50
  );


  buf
  g318
  (
    n322,
    n120
  );


  not
  g319
  (
    n588,
    n89
  );


  not
  g320
  (
    n427,
    n43
  );


  buf
  g321
  (
    n470,
    n98
  );


  not
  g322
  (
    n393,
    n40
  );


  buf
  g323
  (
    n384,
    n111
  );


  not
  g324
  (
    n278,
    n132
  );


  buf
  g325
  (
    n256,
    n90
  );


  not
  g326
  (
    n346,
    n39
  );


  buf
  g327
  (
    n420,
    n96
  );


  buf
  g328
  (
    n526,
    n81
  );


  buf
  g329
  (
    n192,
    n91
  );


  not
  g330
  (
    n515,
    n121
  );


  buf
  g331
  (
    n268,
    n99
  );


  not
  g332
  (
    n507,
    n89
  );


  not
  g333
  (
    n490,
    n121
  );


  buf
  g334
  (
    n316,
    n38
  );


  not
  g335
  (
    n414,
    n81
  );


  buf
  g336
  (
    n195,
    n119
  );


  not
  g337
  (
    n413,
    n49
  );


  buf
  g338
  (
    n572,
    n109
  );


  not
  g339
  (
    n344,
    n77
  );


  not
  g340
  (
    n466,
    n108
  );


  not
  g341
  (
    n330,
    n137
  );


  buf
  g342
  (
    n562,
    n125
  );


  not
  g343
  (
    n477,
    n88
  );


  buf
  g344
  (
    n407,
    n77
  );


  not
  g345
  (
    n191,
    n65
  );


  not
  g346
  (
    n304,
    n38
  );


  not
  g347
  (
    n255,
    n124
  );


  not
  g348
  (
    n225,
    n99
  );


  not
  g349
  (
    n582,
    n90
  );


  not
  g350
  (
    n326,
    n40
  );


  not
  g351
  (
    n530,
    n138
  );


  not
  g352
  (
    n426,
    n44
  );


  not
  g353
  (
    n488,
    n33
  );


  buf
  g354
  (
    n235,
    n87
  );


  buf
  g355
  (
    n491,
    n64
  );


  not
  g356
  (
    n162,
    n55
  );


  not
  g357
  (
    KeyWire_0_12,
    n141
  );


  buf
  g358
  (
    n216,
    n104
  );


  buf
  g359
  (
    n473,
    n52
  );


  not
  g360
  (
    n402,
    n48
  );


  not
  g361
  (
    n253,
    n81
  );


  not
  g362
  (
    n580,
    n128
  );


  not
  g363
  (
    n411,
    n119
  );


  buf
  g364
  (
    n465,
    n135
  );


  buf
  g365
  (
    n234,
    n88
  );


  not
  g366
  (
    n546,
    n68
  );


  buf
  g367
  (
    n442,
    n72
  );


  not
  g368
  (
    n285,
    n80
  );


  not
  g369
  (
    n479,
    n51
  );


  buf
  g370
  (
    n468,
    n110
  );


  buf
  g371
  (
    n509,
    n133
  );


  buf
  g372
  (
    n403,
    n37
  );


  not
  g373
  (
    n458,
    n71
  );


  not
  g374
  (
    n349,
    n95
  );


  buf
  g375
  (
    n360,
    n82
  );


  buf
  g376
  (
    n161,
    n52
  );


  buf
  g377
  (
    n199,
    n96
  );


  buf
  g378
  (
    n485,
    n136
  );


  buf
  g379
  (
    n228,
    n79
  );


  not
  g380
  (
    n594,
    n129
  );


  not
  g381
  (
    n517,
    n44
  );


  buf
  g382
  (
    n511,
    n120
  );


  not
  g383
  (
    n241,
    n126
  );


  not
  g384
  (
    n551,
    n80
  );


  buf
  g385
  (
    n331,
    n91
  );


  buf
  g386
  (
    n172,
    n50
  );


  not
  g387
  (
    n499,
    n138
  );


  not
  g388
  (
    n573,
    n63
  );


  not
  g389
  (
    n358,
    n138
  );


  not
  g390
  (
    n196,
    n65
  );


  buf
  g391
  (
    n311,
    n41
  );


  not
  g392
  (
    n366,
    n94
  );


  not
  g393
  (
    n182,
    n104
  );


  buf
  g394
  (
    n564,
    n79
  );


  not
  g395
  (
    n281,
    n92
  );


  buf
  g396
  (
    n577,
    n107
  );


  not
  g397
  (
    n464,
    n121
  );


  not
  g398
  (
    n512,
    n85
  );


  buf
  g399
  (
    n319,
    n103
  );


  buf
  g400
  (
    n424,
    n136
  );


  buf
  g401
  (
    n264,
    n125
  );


  buf
  g402
  (
    n500,
    n130
  );


  buf
  g403
  (
    n452,
    n114
  );


  buf
  g404
  (
    n166,
    n120
  );


  not
  g405
  (
    n543,
    n75
  );


  buf
  g406
  (
    n262,
    n91
  );


  not
  g407
  (
    n257,
    n94
  );


  buf
  g408
  (
    n433,
    n54
  );


  buf
  g409
  (
    n431,
    n71
  );


  not
  g410
  (
    n584,
    n102
  );


  not
  g411
  (
    n324,
    n83
  );


  buf
  g412
  (
    n462,
    n134
  );


  buf
  g413
  (
    n223,
    n110
  );


  buf
  g414
  (
    n448,
    n104
  );


  not
  g415
  (
    n367,
    n68
  );


  buf
  g416
  (
    n323,
    n63
  );


  not
  g417
  (
    n307,
    n126
  );


  not
  g418
  (
    n453,
    n103
  );


  not
  g419
  (
    n178,
    n131
  );


  buf
  g420
  (
    n301,
    n33
  );


  buf
  g421
  (
    n293,
    n123
  );


  buf
  g422
  (
    n273,
    n90
  );


  buf
  g423
  (
    n503,
    n73
  );


  buf
  g424
  (
    n443,
    n77
  );


  buf
  g425
  (
    n520,
    n85
  );


  not
  g426
  (
    n167,
    n74
  );


  not
  g427
  (
    n363,
    n113
  );


  buf
  g428
  (
    n450,
    n115
  );


  not
  g429
  (
    n593,
    n131
  );


  not
  g430
  (
    n475,
    n78
  );


  not
  g431
  (
    n537,
    n76
  );


  buf
  g432
  (
    n536,
    n62
  );


  buf
  g433
  (
    n189,
    n109
  );


  buf
  g434
  (
    n365,
    n43
  );


  buf
  g435
  (
    n498,
    n113
  );


  buf
  g436
  (
    n246,
    n98
  );


  not
  g437
  (
    n309,
    n49
  );


  not
  g438
  (
    n514,
    n118
  );


  buf
  g439
  (
    n180,
    n96
  );


  buf
  g440
  (
    n294,
    n67
  );


  not
  g441
  (
    n318,
    n110
  );


  buf
  g442
  (
    n493,
    n129
  );


  buf
  g443
  (
    n392,
    n97
  );


  not
  g444
  (
    n164,
    n70
  );


  buf
  g445
  (
    n527,
    n91
  );


  buf
  g446
  (
    n388,
    n140
  );


  buf
  g447
  (
    n492,
    n123
  );


  not
  g448
  (
    n200,
    n138
  );


  not
  g449
  (
    n313,
    n57
  );


  buf
  g450
  (
    n441,
    n61
  );


  not
  g451
  (
    n353,
    n53
  );


  buf
  g452
  (
    n383,
    n66
  );


  not
  g453
  (
    n337,
    n134
  );


  not
  g454
  (
    n372,
    n105
  );


  not
  g455
  (
    n300,
    n100
  );


  not
  g456
  (
    n315,
    n102
  );


  not
  g457
  (
    n205,
    n54
  );


  not
  g458
  (
    n279,
    n76
  );


  not
  g459
  (
    n444,
    n132
  );


  not
  g460
  (
    n280,
    n71
  );


  buf
  g461
  (
    n415,
    n34
  );


  not
  g462
  (
    n538,
    n53
  );


  not
  g463
  (
    n561,
    n122
  );


  buf
  g464
  (
    n396,
    n82
  );


  buf
  g465
  (
    n381,
    n60
  );


  buf
  g466
  (
    n174,
    n59
  );


  buf
  g467
  (
    n539,
    n39
  );


  buf
  g468
  (
    n347,
    n105
  );


  not
  g469
  (
    n275,
    n120
  );


  buf
  g470
  (
    KeyWire_0_24,
    n101
  );


  buf
  g471
  (
    n220,
    n117
  );


  buf
  g472
  (
    n472,
    n40
  );


  buf
  g473
  (
    KeyWire_0_17,
    n55
  );


  not
  g474
  (
    n585,
    n78
  );


  buf
  g475
  (
    n556,
    n72
  );


  not
  g476
  (
    n244,
    n86
  );


  not
  g477
  (
    n198,
    n55
  );


  buf
  g478
  (
    n287,
    n95
  );


  not
  g479
  (
    n240,
    n73
  );


  not
  g480
  (
    n460,
    n48
  );


  not
  g481
  (
    n368,
    n46
  );


  buf
  g482
  (
    n570,
    n140
  );


  not
  g483
  (
    n208,
    n71
  );


  not
  g484
  (
    n481,
    n124
  );


  not
  g485
  (
    n446,
    n62
  );


  buf
  g486
  (
    n571,
    n46
  );


  not
  g487
  (
    n378,
    n33
  );


  not
  g488
  (
    n467,
    n122
  );


  not
  g489
  (
    n356,
    n100
  );


  not
  g490
  (
    n314,
    n61
  );


  buf
  g491
  (
    n181,
    n63
  );


  buf
  g492
  (
    n389,
    n113
  );


  not
  g493
  (
    n474,
    n111
  );


  not
  g494
  (
    n494,
    n43
  );


  not
  g495
  (
    n184,
    n97
  );


  not
  g496
  (
    n254,
    n105
  );


  not
  g497
  (
    n291,
    n123
  );


  buf
  g498
  (
    n502,
    n92
  );


  buf
  g499
  (
    n364,
    n112
  );


  not
  g500
  (
    n591,
    n60
  );


  buf
  g501
  (
    n496,
    n67
  );


  buf
  g502
  (
    n269,
    n112
  );


  buf
  g503
  (
    n305,
    n72
  );


  buf
  g504
  (
    n559,
    n116
  );


  not
  g505
  (
    KeyWire_0_11,
    n101
  );


  not
  g506
  (
    n226,
    n84
  );


  buf
  g507
  (
    n391,
    n58
  );


  buf
  g508
  (
    n405,
    n92
  );


  buf
  g509
  (
    n175,
    n118
  );


  not
  g510
  (
    n438,
    n73
  );


  not
  g511
  (
    n190,
    n37
  );


  not
  g512
  (
    n377,
    n70
  );


  not
  g513
  (
    n201,
    n41
  );


  buf
  g514
  (
    n329,
    n116
  );


  not
  g515
  (
    n435,
    n74
  );


  buf
  g516
  (
    n459,
    n56
  );


  buf
  g517
  (
    KeyWire_0_29,
    n67
  );


  buf
  g518
  (
    n258,
    n42
  );


  buf
  g519
  (
    n456,
    n58
  );


  not
  g520
  (
    n202,
    n68
  );


  buf
  g521
  (
    n193,
    n57
  );


  not
  g522
  (
    n272,
    n69
  );


  not
  g523
  (
    n412,
    n68
  );


  buf
  g524
  (
    n541,
    n53
  );


  buf
  g525
  (
    n261,
    n42
  );


  buf
  g526
  (
    n170,
    n109
  );


  not
  g527
  (
    n425,
    n128
  );


  buf
  g528
  (
    n187,
    n45
  );


  not
  g529
  (
    n423,
    n45
  );


  buf
  g530
  (
    n266,
    n98
  );


  not
  g531
  (
    n523,
    n60
  );


  buf
  g532
  (
    n505,
    n114
  );


  buf
  g533
  (
    n566,
    n64
  );


  buf
  g534
  (
    n374,
    n140
  );


  buf
  g535
  (
    n404,
    n77
  );


  not
  g536
  (
    n332,
    n53
  );


  not
  g537
  (
    n416,
    n106
  );


  buf
  g538
  (
    n549,
    n80
  );


  not
  g539
  (
    n357,
    n83
  );


  not
  g540
  (
    n529,
    n128
  );


  buf
  g541
  (
    n222,
    n62
  );


  buf
  g542
  (
    n504,
    n73
  );


  not
  g543
  (
    n327,
    n96
  );


  buf
  g544
  (
    n516,
    n124
  );


  not
  g545
  (
    n463,
    n89
  );


  buf
  g546
  (
    n399,
    n97
  );


  buf
  g547
  (
    n522,
    n103
  );


  buf
  g548
  (
    n419,
    n99
  );


  not
  g549
  (
    n277,
    n123
  );


  not
  g550
  (
    n206,
    n118
  );


  not
  g551
  (
    n203,
    n35
  );


  buf
  g552
  (
    n179,
    n63
  );


  not
  g553
  (
    n188,
    n139
  );


  not
  g554
  (
    n267,
    n104
  );


  buf
  g555
  (
    n410,
    n62
  );


  buf
  g556
  (
    n345,
    n56
  );


  not
  g557
  (
    n308,
    n114
  );


  not
  g558
  (
    n575,
    n50
  );


  buf
  g559
  (
    n219,
    n82
  );


  not
  g560
  (
    n339,
    n132
  );


  buf
  g561
  (
    n557,
    n85
  );


  buf
  g562
  (
    n714,
    n177
  );


  buf
  g563
  (
    n724,
    n240
  );


  buf
  g564
  (
    n716,
    n234
  );


  not
  g565
  (
    n713,
    n303
  );


  not
  g566
  (
    n694,
    n321
  );


  not
  g567
  (
    n672,
    n275
  );


  buf
  g568
  (
    n605,
    n170
  );


  not
  g569
  (
    n637,
    n256
  );


  buf
  g570
  (
    n621,
    n179
  );


  not
  g571
  (
    n718,
    n314
  );


  buf
  g572
  (
    n810,
    n226
  );


  not
  g573
  (
    n653,
    n333
  );


  not
  g574
  (
    n812,
    n191
  );


  not
  g575
  (
    n646,
    n297
  );


  not
  g576
  (
    n680,
    n263
  );


  not
  g577
  (
    n811,
    n185
  );


  not
  g578
  (
    n667,
    n165
  );


  not
  g579
  (
    n691,
    n339
  );


  not
  g580
  (
    n739,
    n172
  );


  not
  g581
  (
    n725,
    n231
  );


  buf
  g582
  (
    n727,
    n363
  );


  buf
  g583
  (
    n731,
    n326
  );


  not
  g584
  (
    n651,
    n194
  );


  buf
  g585
  (
    n729,
    n341
  );


  not
  g586
  (
    KeyWire_0_13,
    n306
  );


  buf
  g587
  (
    n793,
    n262
  );


  not
  g588
  (
    n632,
    n355
  );


  buf
  g589
  (
    n604,
    n218
  );


  not
  g590
  (
    n626,
    n344
  );


  not
  g591
  (
    n698,
    n203
  );


  buf
  g592
  (
    n740,
    n184
  );


  not
  g593
  (
    n790,
    n270
  );


  not
  g594
  (
    n797,
    n276
  );


  buf
  g595
  (
    n623,
    n290
  );


  not
  g596
  (
    n615,
    n332
  );


  buf
  g597
  (
    n663,
    n244
  );


  not
  g598
  (
    n678,
    n351
  );


  not
  g599
  (
    n655,
    n318
  );


  not
  g600
  (
    n597,
    n247
  );


  buf
  g601
  (
    n649,
    n374
  );


  not
  g602
  (
    n730,
    n282
  );


  not
  g603
  (
    n699,
    n222
  );


  not
  g604
  (
    n695,
    n175
  );


  buf
  g605
  (
    n654,
    n214
  );


  not
  g606
  (
    n643,
    n242
  );


  buf
  g607
  (
    n669,
    n252
  );


  not
  g608
  (
    n755,
    n274
  );


  not
  g609
  (
    n747,
    n310
  );


  not
  g610
  (
    n738,
    n239
  );


  buf
  g611
  (
    n690,
    n192
  );


  buf
  g612
  (
    n765,
    n198
  );


  buf
  g613
  (
    n737,
    n292
  );


  buf
  g614
  (
    n757,
    n280
  );


  buf
  g615
  (
    n754,
    n383
  );


  not
  g616
  (
    n786,
    n215
  );


  buf
  g617
  (
    n816,
    n385
  );


  not
  g618
  (
    n750,
    n250
  );


  buf
  g619
  (
    n610,
    n291
  );


  buf
  g620
  (
    n785,
    n277
  );


  not
  g621
  (
    n783,
    n271
  );


  buf
  g622
  (
    n728,
    n173
  );


  buf
  g623
  (
    n760,
    n230
  );


  not
  g624
  (
    n802,
    n354
  );


  buf
  g625
  (
    KeyWire_0_10,
    n286
  );


  buf
  g626
  (
    n676,
    n387
  );


  not
  g627
  (
    n787,
    n300
  );


  not
  g628
  (
    n666,
    n377
  );


  not
  g629
  (
    n636,
    n375
  );


  not
  g630
  (
    n608,
    n302
  );


  not
  g631
  (
    n659,
    n201
  );


  not
  g632
  (
    n813,
    n287
  );


  buf
  g633
  (
    n689,
    n273
  );


  not
  g634
  (
    n683,
    n269
  );


  buf
  g635
  (
    n687,
    n255
  );


  buf
  g636
  (
    n741,
    n164
  );


  buf
  g637
  (
    n796,
    n307
  );


  not
  g638
  (
    n657,
    n206
  );


  not
  g639
  (
    n688,
    n216
  );


  buf
  g640
  (
    n821,
    n340
  );


  buf
  g641
  (
    n719,
    n338
  );


  not
  g642
  (
    n662,
    n245
  );


  not
  g643
  (
    n707,
    n268
  );


  buf
  g644
  (
    n817,
    n220
  );


  buf
  g645
  (
    n625,
    n254
  );


  not
  g646
  (
    n697,
    n359
  );


  buf
  g647
  (
    n661,
    n352
  );


  buf
  g648
  (
    n778,
    n362
  );


  not
  g649
  (
    n733,
    n209
  );


  not
  g650
  (
    n723,
    n248
  );


  buf
  g651
  (
    n686,
    n370
  );


  buf
  g652
  (
    n700,
    n295
  );


  not
  g653
  (
    n619,
    n217
  );


  not
  g654
  (
    n819,
    n337
  );


  not
  g655
  (
    n709,
    n238
  );


  buf
  g656
  (
    n761,
    n180
  );


  not
  g657
  (
    n758,
    n371
  );


  buf
  g658
  (
    n684,
    n304
  );


  not
  g659
  (
    n638,
    n350
  );


  not
  g660
  (
    n614,
    n233
  );


  not
  g661
  (
    n631,
    n284
  );


  not
  g662
  (
    n806,
    n211
  );


  buf
  g663
  (
    n627,
    n357
  );


  buf
  g664
  (
    n808,
    n246
  );


  buf
  g665
  (
    n599,
    n278
  );


  buf
  g666
  (
    n650,
    n166
  );


  not
  g667
  (
    n799,
    n182
  );


  not
  g668
  (
    n679,
    n241
  );


  buf
  g669
  (
    n722,
    n235
  );


  not
  g670
  (
    n762,
    n336
  );


  buf
  g671
  (
    n671,
    n379
  );


  not
  g672
  (
    n617,
    n348
  );


  not
  g673
  (
    n682,
    n213
  );


  not
  g674
  (
    n668,
    n260
  );


  not
  g675
  (
    n780,
    n312
  );


  buf
  g676
  (
    n658,
    n199
  );


  not
  g677
  (
    n732,
    n174
  );


  buf
  g678
  (
    n721,
    n257
  );


  buf
  g679
  (
    n702,
    n261
  );


  buf
  g680
  (
    n814,
    n187
  );


  buf
  g681
  (
    n807,
    n294
  );


  not
  g682
  (
    n748,
    n353
  );


  buf
  g683
  (
    n751,
    n358
  );


  not
  g684
  (
    n715,
    n168
  );


  not
  g685
  (
    n600,
    n361
  );


  not
  g686
  (
    n753,
    n299
  );


  not
  g687
  (
    n805,
    n328
  );


  not
  g688
  (
    n711,
    n259
  );


  not
  g689
  (
    n763,
    n369
  );


  buf
  g690
  (
    n804,
    n335
  );


  not
  g691
  (
    n673,
    n204
  );


  buf
  g692
  (
    n598,
    n202
  );


  buf
  g693
  (
    n781,
    n372
  );


  not
  g694
  (
    n693,
    n221
  );


  buf
  g695
  (
    n611,
    n176
  );


  buf
  g696
  (
    n792,
    n356
  );


  buf
  g697
  (
    n639,
    n193
  );


  buf
  g698
  (
    n717,
    n283
  );


  not
  g699
  (
    n624,
    n183
  );


  not
  g700
  (
    n784,
    n229
  );


  not
  g701
  (
    n656,
    n197
  );


  not
  g702
  (
    n675,
    n330
  );


  not
  g703
  (
    n776,
    n305
  );


  not
  g704
  (
    n681,
    n293
  );


  not
  g705
  (
    n633,
    n232
  );


  not
  g706
  (
    n759,
    n320
  );


  not
  g707
  (
    n767,
    n200
  );


  not
  g708
  (
    n710,
    n342
  );


  buf
  g709
  (
    n641,
    n360
  );


  not
  g710
  (
    n798,
    n324
  );


  not
  g711
  (
    n774,
    n207
  );


  buf
  g712
  (
    n685,
    n272
  );


  buf
  g713
  (
    n772,
    n329
  );


  buf
  g714
  (
    n602,
    n210
  );


  buf
  g715
  (
    n764,
    n169
  );


  not
  g716
  (
    n674,
    n162
  );


  not
  g717
  (
    n742,
    n381
  );


  not
  g718
  (
    n794,
    n224
  );


  buf
  g719
  (
    n795,
    n311
  );


  not
  g720
  (
    n736,
    n279
  );


  buf
  g721
  (
    n712,
    n258
  );


  buf
  g722
  (
    n703,
    n315
  );


  buf
  g723
  (
    n818,
    n378
  );


  buf
  g724
  (
    n803,
    n237
  );


  not
  g725
  (
    n642,
    n253
  );


  buf
  g726
  (
    n601,
    n322
  );


  buf
  g727
  (
    n769,
    n345
  );


  buf
  g728
  (
    n670,
    n316
  );


  buf
  g729
  (
    n768,
    n265
  );


  not
  g730
  (
    n647,
    n346
  );


  not
  g731
  (
    n815,
    n181
  );


  buf
  g732
  (
    n612,
    n288
  );


  not
  g733
  (
    n644,
    n386
  );


  buf
  g734
  (
    n596,
    n325
  );


  buf
  g735
  (
    n696,
    n349
  );


  buf
  g736
  (
    n820,
    n189
  );


  not
  g737
  (
    n752,
    n266
  );


  not
  g738
  (
    n620,
    n368
  );


  buf
  g739
  (
    n791,
    n367
  );


  buf
  g740
  (
    n609,
    n347
  );


  buf
  g741
  (
    n734,
    n285
  );


  not
  g742
  (
    n630,
    n301
  );


  buf
  g743
  (
    n745,
    n308
  );


  buf
  g744
  (
    n616,
    n227
  );


  buf
  g745
  (
    n749,
    n251
  );


  not
  g746
  (
    n634,
    n319
  );


  buf
  g747
  (
    n788,
    n208
  );


  not
  g748
  (
    n701,
    n190
  );


  buf
  g749
  (
    n606,
    n366
  );


  not
  g750
  (
    n622,
    n196
  );


  buf
  g751
  (
    n660,
    n298
  );


  not
  g752
  (
    n595,
    n289
  );


  buf
  g753
  (
    n708,
    n188
  );


  not
  g754
  (
    n770,
    n331
  );


  buf
  g755
  (
    n665,
    n323
  );


  not
  g756
  (
    n771,
    n212
  );


  not
  g757
  (
    n705,
    n219
  );


  buf
  g758
  (
    n628,
    n161
  );


  not
  g759
  (
    n692,
    n313
  );


  buf
  g760
  (
    n726,
    n373
  );


  not
  g761
  (
    n704,
    n327
  );


  buf
  g762
  (
    n744,
    n334
  );


  not
  g763
  (
    n746,
    n380
  );


  not
  g764
  (
    n607,
    n382
  );


  buf
  g765
  (
    n652,
    n167
  );


  not
  g766
  (
    n629,
    n186
  );


  not
  g767
  (
    n735,
    n171
  );


  not
  g768
  (
    n648,
    n364
  );


  not
  g769
  (
    n800,
    n267
  );


  not
  g770
  (
    n789,
    n249
  );


  not
  g771
  (
    n756,
    n223
  );


  buf
  g772
  (
    n603,
    n195
  );


  not
  g773
  (
    n640,
    n317
  );


  not
  g774
  (
    n677,
    n205
  );


  buf
  g775
  (
    n743,
    n228
  );


  buf
  g776
  (
    n706,
    n264
  );


  buf
  g777
  (
    n782,
    n365
  );


  buf
  g778
  (
    n779,
    n309
  );


  buf
  g779
  (
    n635,
    n281
  );


  not
  g780
  (
    n801,
    n376
  );


  buf
  g781
  (
    n773,
    n384
  );


  not
  g782
  (
    n809,
    n343
  );


  not
  g783
  (
    n766,
    n163
  );


  not
  g784
  (
    n613,
    n296
  );


  buf
  g785
  (
    n775,
    n225
  );


  not
  g786
  (
    n618,
    n236
  );


  not
  g787
  (
    n720,
    n243
  );


  buf
  g788
  (
    n777,
    n178
  );


  or
  g789
  (
    n826,
    n481,
    n652,
    n146,
    n557
  );


  xor
  g790
  (
    n867,
    n788,
    n455,
    n147,
    n602
  );


  nand
  g791
  (
    n834,
    n471,
    n656,
    n469,
    n555
  );


  and
  g792
  (
    n1026,
    n745,
    n806,
    n617,
    n535
  );


  or
  g793
  (
    n944,
    n488,
    n498,
    n701,
    n423
  );


  and
  g794
  (
    n901,
    n507,
    n467,
    n489,
    n571
  );


  nand
  g795
  (
    n940,
    n160,
    n412,
    n451,
    n157
  );


  or
  g796
  (
    n1039,
    n523,
    n720,
    n474,
    n537
  );


  or
  g797
  (
    n926,
    n550,
    n684,
    n539,
    n538
  );


  and
  g798
  (
    n905,
    n728,
    n808,
    n467,
    n679
  );


  nor
  g799
  (
    n951,
    n520,
    n751,
    n508,
    n525
  );


  nand
  g800
  (
    n849,
    n550,
    n472,
    n763,
    n146
  );


  or
  g801
  (
    n921,
    n390,
    n621,
    n556,
    n157
  );


  nor
  g802
  (
    n900,
    n634,
    n618,
    n419,
    n563
  );


  nand
  g803
  (
    n1033,
    n502,
    n155,
    n399,
    n710
  );


  xnor
  g804
  (
    n1030,
    n538,
    n802,
    n774,
    n567
  );


  or
  g805
  (
    n842,
    n665,
    n424,
    n468,
    n519
  );


  xor
  g806
  (
    n927,
    n541,
    n469,
    n493,
    n509
  );


  nand
  g807
  (
    n1017,
    n405,
    n452,
    n553,
    n516
  );


  or
  g808
  (
    n994,
    n719,
    n156,
    n532,
    n449
  );


  xor
  g809
  (
    n966,
    n635,
    n804,
    n655,
    n455
  );


  or
  g810
  (
    n967,
    n748,
    n533,
    n680,
    n657
  );


  nand
  g811
  (
    n1021,
    n468,
    n506,
    n663,
    n512
  );


  nand
  g812
  (
    n832,
    n555,
    n553,
    n693,
    n156
  );


  and
  g813
  (
    n862,
    n527,
    n803,
    n159,
    n487
  );


  xnor
  g814
  (
    n989,
    n158,
    n542,
    n544,
    n744
  );


  and
  g815
  (
    n870,
    n575,
    n461,
    n791,
    n146
  );


  or
  g816
  (
    n863,
    n767,
    n451,
    n612,
    n782
  );


  and
  g817
  (
    n1045,
    n155,
    n443,
    n631,
    n568
  );


  xnor
  g818
  (
    n1001,
    n444,
    n649,
    n486,
    n482
  );


  or
  g819
  (
    n960,
    n638,
    n503,
    n526,
    n493
  );


  or
  g820
  (
    n840,
    n765,
    n559,
    n445,
    n542
  );


  or
  g821
  (
    n1022,
    n648,
    n644,
    n489,
    n508
  );


  xor
  g822
  (
    n824,
    n601,
    n558,
    n536,
    n153
  );


  xor
  g823
  (
    n933,
    n520,
    n805,
    n819,
    n504
  );


  xor
  g824
  (
    n873,
    n151,
    n490,
    n526,
    n674
  );


  xnor
  g825
  (
    n886,
    n658,
    n515,
    n713,
    n535
  );


  nor
  g826
  (
    KeyWire_0_14,
    n773,
    n524,
    n470,
    n462
  );


  xor
  g827
  (
    n854,
    n152,
    n450,
    n496,
    n148
  );


  and
  g828
  (
    n1019,
    n514,
    n464,
    n510,
    n483
  );


  and
  g829
  (
    n918,
    n458,
    n467,
    n457,
    n555
  );


  xnor
  g830
  (
    n916,
    n687,
    n526,
    n513,
    n486
  );


  xnor
  g831
  (
    n880,
    n550,
    n577,
    n724,
    n480
  );


  xnor
  g832
  (
    n1004,
    n651,
    n472,
    n682,
    n444
  );


  nand
  g833
  (
    n985,
    n549,
    n500,
    n757,
    n566
  );


  xnor
  g834
  (
    n974,
    n731,
    n558,
    n503,
    n517
  );


  xnor
  g835
  (
    n860,
    n686,
    n540,
    n572,
    n158
  );


  xnor
  g836
  (
    n848,
    n460,
    n509,
    n754,
    n442
  );


  nor
  g837
  (
    n1010,
    n487,
    n495,
    n596,
    n548
  );


  or
  g838
  (
    n1042,
    n570,
    n495,
    n471,
    n456
  );


  or
  g839
  (
    n1028,
    n703,
    n490,
    n159,
    n677
  );


  xor
  g840
  (
    n984,
    n552,
    n570,
    n454,
    n145
  );


  or
  g841
  (
    KeyWire_0_5,
    n143,
    n747,
    n396,
    n554
  );


  or
  g842
  (
    n1034,
    n455,
    n546,
    n454,
    n467
  );


  xor
  g843
  (
    n1005,
    n565,
    n154,
    n578,
    n784
  );


  xor
  g844
  (
    n1007,
    n416,
    n560,
    n510,
    n499
  );


  nand
  g845
  (
    n1043,
    n150,
    n534,
    n453,
    n741
  );


  nand
  g846
  (
    n908,
    n502,
    n530,
    n477
  );


  nand
  g847
  (
    n979,
    n800,
    n551,
    n492,
    n641
  );


  nor
  g848
  (
    n879,
    n155,
    n603,
    n477,
    n694
  );


  nor
  g849
  (
    n1046,
    n450,
    n515,
    n469,
    n573
  );


  and
  g850
  (
    n953,
    n495,
    n604,
    n511,
    n153
  );


  xor
  g851
  (
    n858,
    n398,
    n531,
    n484,
    n551
  );


  or
  g852
  (
    n935,
    n470,
    n525,
    n569,
    n639
  );


  nand
  g853
  (
    n844,
    n466,
    n623,
    n810,
    n538
  );


  xor
  g854
  (
    n833,
    n462,
    n705,
    n444,
    n556
  );


  nor
  g855
  (
    n947,
    n445,
    n446,
    n477,
    n654
  );


  or
  g856
  (
    n871,
    n572,
    n547,
    n555,
    n493
  );


  or
  g857
  (
    n845,
    n561,
    n492,
    n550,
    n480
  );


  nand
  g858
  (
    n991,
    n458,
    n160,
    n568,
    n737
  );


  nand
  g859
  (
    n825,
    n636,
    n653,
    n154,
    n799
  );


  and
  g860
  (
    n1031,
    n501,
    n786,
    n395,
    n559
  );


  or
  g861
  (
    n949,
    n552,
    n485,
    n643,
    n557
  );


  and
  g862
  (
    n856,
    n570,
    n464,
    n615,
    n690
  );


  nor
  g863
  (
    n1024,
    n413,
    n498,
    n716,
    n708
  );


  xnor
  g864
  (
    n883,
    n483,
    n438,
    n146,
    n414
  );


  and
  g865
  (
    n983,
    n459,
    n609,
    n457,
    n557
  );


  nand
  g866
  (
    n830,
    n537,
    n752,
    n521,
    n702
  );


  xor
  g867
  (
    n982,
    n536,
    n760,
    n448,
    n787
  );


  or
  g868
  (
    n847,
    n697,
    n556,
    n598,
    n431
  );


  xnor
  g869
  (
    n978,
    n500,
    n496,
    n567,
    n151
  );


  and
  g870
  (
    n972,
    n507,
    n496,
    n154,
    n820
  );


  and
  g871
  (
    KeyWire_0_0,
    n148,
    n485,
    n498,
    n563
  );


  nor
  g872
  (
    n923,
    n145,
    n441,
    n149,
    n778
  );


  nor
  g873
  (
    n975,
    n501,
    n143,
    n676,
    n528
  );


  xor
  g874
  (
    n997,
    n552,
    n528,
    n474,
    n484
  );


  or
  g875
  (
    n1029,
    n633,
    n487,
    n515,
    n394
  );


  nand
  g876
  (
    n861,
    n459,
    n489,
    n508,
    n789
  );


  or
  g877
  (
    n981,
    n521,
    n670,
    n545,
    n527
  );


  xnor
  g878
  (
    n934,
    n462,
    n532,
    n447,
    n474
  );


  nand
  g879
  (
    n930,
    n482,
    n699,
    n451,
    n759
  );


  or
  g880
  (
    n1040,
    n573,
    n775,
    n479,
    n420
  );


  nand
  g881
  (
    n1041,
    n564,
    n523,
    n700,
    n527
  );


  or
  g882
  (
    n995,
    n475,
    n522,
    n148,
    n459
  );


  nand
  g883
  (
    n1002,
    n611,
    n544,
    n529,
    n500
  );


  nand
  g884
  (
    n961,
    n410,
    n147,
    n797,
    n764
  );


  and
  g885
  (
    n998,
    n573,
    n738,
    n465,
    n145
  );


  or
  g886
  (
    n885,
    n566,
    n486,
    n688,
    n732
  );


  xnor
  g887
  (
    n906,
    n560,
    n464,
    n511,
    n407
  );


  xor
  g888
  (
    n1027,
    n567,
    n534,
    n517,
    n449
  );


  nand
  g889
  (
    n1032,
    n411,
    n450,
    n562,
    n722
  );


  xor
  g890
  (
    n846,
    n489,
    n622,
    n572,
    n531
  );


  xnor
  g891
  (
    n1047,
    n574,
    n526,
    n463,
    n152
  );


  nor
  g892
  (
    n868,
    n566,
    n532,
    n678,
    n492
  );


  or
  g893
  (
    n941,
    n696,
    n536,
    n561,
    n491
  );


  xnor
  g894
  (
    n877,
    n669,
    n559,
    n798,
    n403
  );


  or
  g895
  (
    n1025,
    n664,
    n547,
    n402,
    n608
  );


  or
  g896
  (
    n999,
    n453,
    n578,
    n430,
    n736
  );


  or
  g897
  (
    n922,
    n562,
    n541,
    n454,
    n406
  );


  and
  g898
  (
    n936,
    n480,
    n553,
    n507,
    n554
  );


  or
  g899
  (
    n881,
    n514,
    n563,
    n450,
    n479
  );


  nand
  g900
  (
    n915,
    n575,
    n546,
    n533,
    n513
  );


  xor
  g901
  (
    n907,
    n448,
    n474,
    n465,
    n142
  );


  nand
  g902
  (
    n896,
    n642,
    n510,
    n478,
    n575
  );


  xnor
  g903
  (
    n950,
    n597,
    n795,
    n691,
    n614
  );


  xor
  g904
  (
    n986,
    n408,
    n432,
    n498,
    n717
  );


  xnor
  g905
  (
    n822,
    n613,
    n445,
    n516,
    n721
  );


  and
  g906
  (
    n973,
    n466,
    n630,
    n558,
    n443
  );


  nand
  g907
  (
    n962,
    n478,
    n535,
    n729,
    n490
  );


  or
  g908
  (
    n823,
    n625,
    n454,
    n397,
    n516
  );


  and
  g909
  (
    n874,
    n154,
    n447,
    n725
  );


  xnor
  g910
  (
    n990,
    n768,
    n451,
    n607,
    n476
  );


  and
  g911
  (
    n892,
    n542,
    n142,
    n425,
    n756
  );


  or
  g912
  (
    n945,
    n776,
    n755,
    n461,
    n624
  );


  and
  g913
  (
    n852,
    n508,
    n545,
    n144,
    n466
  );


  xnor
  g914
  (
    n836,
    n574,
    n758,
    n783,
    n535
  );


  nor
  g915
  (
    n831,
    n560,
    n689,
    n541,
    n479
  );


  xor
  g916
  (
    n889,
    n496,
    n683,
    n505,
    n675
  );


  and
  g917
  (
    n893,
    n158,
    n544,
    n156,
    n494
  );


  and
  g918
  (
    n993,
    n141,
    n551,
    n792,
    n509
  );


  nor
  g919
  (
    n1003,
    n743,
    n472,
    n147,
    n742
  );


  xor
  g920
  (
    n903,
    n149,
    n531,
    n506
  );


  xnor
  g921
  (
    n894,
    n541,
    n620,
    n692,
    n750
  );


  and
  g922
  (
    n955,
    n746,
    n548,
    n524,
    n433
  );


  nor
  g923
  (
    n920,
    n497,
    n718,
    n473,
    n151
  );


  and
  g924
  (
    n948,
    n527,
    n561,
    n150,
    n143
  );


  and
  g925
  (
    n865,
    n144,
    n505,
    n152,
    n150
  );


  or
  g926
  (
    n876,
    n565,
    n574,
    n142,
    n532
  );


  nor
  g927
  (
    n943,
    n512,
    n576,
    n446,
    n707
  );


  xor
  g928
  (
    n864,
    n494,
    n521,
    n488,
    n761
  );


  and
  g929
  (
    n954,
    n463,
    n517,
    n492,
    n730
  );


  xnor
  g930
  (
    n931,
    n540,
    n785,
    n144,
    n577
  );


  nor
  g931
  (
    n1016,
    n435,
    n497,
    n506,
    n427
  );


  nand
  g932
  (
    n942,
    n519,
    n514,
    n463,
    n734
  );


  or
  g933
  (
    n913,
    n816,
    n681,
    n156,
    n605
  );


  nor
  g934
  (
    n932,
    n512,
    n557,
    n507,
    n502
  );


  or
  g935
  (
    n977,
    n448,
    n434,
    n545,
    n400
  );


  and
  g936
  (
    n859,
    n452,
    n571,
    n476,
    n461
  );


  nand
  g937
  (
    n956,
    n712,
    n632,
    n469,
    n520
  );


  nand
  g938
  (
    n875,
    n447,
    n491,
    n142,
    n659
  );


  xor
  g939
  (
    n855,
    n662,
    n452,
    n568,
    n484
  );


  and
  g940
  (
    n992,
    n567,
    n436,
    n158,
    n462
  );


  xor
  g941
  (
    n1035,
    n539,
    n704,
    n530,
    n749
  );


  nand
  g942
  (
    n851,
    n511,
    n569,
    n388,
    n453
  );


  xnor
  g943
  (
    n971,
    n506,
    n155,
    n514,
    n569
  );


  xor
  g944
  (
    n888,
    n576,
    n473,
    n543,
    n525
  );


  xor
  g945
  (
    n839,
    n619,
    n437,
    n781,
    n706
  );


  and
  g946
  (
    n988,
    n637,
    n772,
    n486,
    n159
  );


  nand
  g947
  (
    n980,
    n534,
    n475,
    n524,
    n770
  );


  and
  g948
  (
    n869,
    n476,
    n160,
    n666
  );


  nand
  g949
  (
    n1009,
    n534,
    n460,
    n672,
    n472
  );


  or
  g950
  (
    n964,
    n487,
    n504,
    n546,
    n443
  );


  and
  g951
  (
    n976,
    n537,
    n522,
    n449,
    n153
  );


  and
  g952
  (
    n968,
    n446,
    n739,
    n726,
    n539
  );


  xor
  g953
  (
    n1006,
    n811,
    n524,
    n471,
    n610
  );


  nand
  g954
  (
    n828,
    n495,
    n480,
    n482,
    n548
  );


  or
  g955
  (
    n1018,
    n478,
    n518,
    n391,
    n576
  );


  nor
  g956
  (
    n970,
    n497,
    n442,
    n818,
    n460
  );


  or
  g957
  (
    n919,
    n505,
    n456,
    n417,
    n484
  );


  xnor
  g958
  (
    n965,
    n551,
    n481,
    n468,
    n512
  );


  and
  g959
  (
    n939,
    n481,
    n521,
    n698,
    n599
  );


  xnor
  g960
  (
    n895,
    n491,
    n456,
    n418,
    n577
  );


  and
  g961
  (
    n917,
    n566,
    n501,
    n545,
    n564
  );


  or
  g962
  (
    n872,
    n149,
    n536,
    n723,
    n539
  );


  or
  g963
  (
    n1023,
    n459,
    n504,
    n460,
    n563
  );


  and
  g964
  (
    n853,
    n715,
    n777,
    n485,
    n452
  );


  nor
  g965
  (
    n843,
    n516,
    n667,
    n145,
    n404
  );


  or
  g966
  (
    n891,
    n509,
    n503,
    n499,
    n533
  );


  and
  g967
  (
    n1036,
    n528,
    n479,
    n695,
    n470
  );


  nand
  g968
  (
    n1015,
    n466,
    n513,
    n790,
    n529
  );


  and
  g969
  (
    n996,
    n150,
    n780,
    n809,
    n570
  );


  xnor
  g970
  (
    n866,
    n483,
    n428,
    n422,
    n626
  );


  xnor
  g971
  (
    n884,
    n762,
    n538,
    n488,
    n540
  );


  xnor
  g972
  (
    n946,
    n457,
    n569,
    n794,
    n389
  );


  xor
  g973
  (
    n1013,
    n673,
    n456,
    n812,
    n628
  );


  nor
  g974
  (
    n882,
    n548,
    n709,
    n801,
    n616
  );


  nor
  g975
  (
    n912,
    n499,
    n711,
    n813,
    n473
  );


  or
  g976
  (
    n1044,
    n529,
    n473,
    n515,
    n769
  );


  nand
  g977
  (
    n898,
    n753,
    n556,
    n650,
    n144
  );


  xnor
  g978
  (
    n924,
    n445,
    n494,
    n574,
    n568
  );


  nand
  g979
  (
    n959,
    n564,
    n401,
    n500,
    n595
  );


  or
  g980
  (
    n838,
    n523,
    n547,
    n733,
    n627
  );


  nor
  g981
  (
    n952,
    n558,
    n537,
    n494,
    n511
  );


  nor
  g982
  (
    n938,
    n468,
    n529,
    n552,
    n807
  );


  and
  g983
  (
    n841,
    n577,
    n544,
    n528,
    n540
  );


  nand
  g984
  (
    n899,
    n571,
    n393,
    n448,
    n546
  );


  and
  g985
  (
    n958,
    n685,
    n564,
    n485,
    n470
  );


  xnor
  g986
  (
    n914,
    n542,
    n793,
    n549,
    n449
  );


  and
  g987
  (
    n904,
    n645,
    n554,
    n153,
    n159
  );


  and
  g988
  (
    n850,
    n565,
    n522,
    n465,
    n562
  );


  or
  g989
  (
    n878,
    n409,
    n475,
    n415,
    n518
  );


  xnor
  g990
  (
    n837,
    n796,
    n525,
    n392,
    n157
  );


  xor
  g991
  (
    n937,
    n553,
    n562,
    n533,
    n483
  );


  nand
  g992
  (
    n969,
    n714,
    n573,
    n561,
    n148
  );


  xor
  g993
  (
    n835,
    n455,
    n510,
    n149,
    n476
  );


  nand
  g994
  (
    n909,
    n458,
    n458,
    n439,
    n499
  );


  xnor
  g995
  (
    n963,
    n143,
    n578,
    n727,
    n446
  );


  xnor
  g996
  (
    n890,
    n543,
    n629,
    n661,
    n481
  );


  nand
  g997
  (
    n1037,
    n475,
    n464,
    n501,
    n817
  );


  and
  g998
  (
    n911,
    n523,
    n490,
    n543,
    n488
  );


  xor
  g999
  (
    n1038,
    n766,
    n668,
    n493,
    n554
  );


  nand
  g1000
  (
    n1012,
    n565,
    n571,
    n157,
    n513
  );


  nand
  g1001
  (
    n910,
    n530,
    n600,
    n478,
    n660
  );


  or
  g1002
  (
    n928,
    n606,
    n444,
    n771,
    n547
  );


  xor
  g1003
  (
    n857,
    n578,
    n740,
    n814,
    n504
  );


  nor
  g1004
  (
    n929,
    n522,
    n517,
    n646,
    n457
  );


  and
  g1005
  (
    n902,
    n518,
    n440,
    n549,
    n421
  );


  nor
  g1006
  (
    n897,
    n560,
    n465,
    n502,
    n482
  );


  xnor
  g1007
  (
    n1014,
    n443,
    n576,
    n503,
    n152
  );


  nor
  g1008
  (
    n1020,
    n147,
    n151,
    n549,
    n735
  );


  nor
  g1009
  (
    n925,
    n429,
    n815,
    n497,
    n491
  );


  xnor
  g1010
  (
    n987,
    n471,
    n671,
    n575,
    n426
  );


  xor
  g1011
  (
    n957,
    n518,
    n572,
    n779,
    n477
  );


  xnor
  g1012
  (
    n1008,
    n141,
    n519,
    n520,
    n461
  );


  nor
  g1013
  (
    n887,
    n519,
    n640,
    n505,
    n543
  );


  nor
  g1014
  (
    n827,
    n559,
    n453,
    n463,
    n647
  );


  not
  g1015
  (
    n1049,
    n823
  );


  buf
  g1016
  (
    n1048,
    n824
  );


  or
  g1017
  (
    n1053,
    n579,
    n582,
    n581,
    n580
  );


  nand
  g1018
  (
    n1056,
    n582,
    n581,
    n583,
    n579
  );


  nand
  g1019
  (
    n1055,
    n582,
    n580,
    n579,
    n1049
  );


  xor
  g1020
  (
    n1054,
    n580,
    n584,
    n1048
  );


  xor
  g1021
  (
    n1052,
    n583,
    n584,
    n579
  );


  nand
  g1022
  (
    n1057,
    n580,
    n1049
  );


  and
  g1023
  (
    n1050,
    n583,
    n581,
    n1048,
    n582
  );


  and
  g1024
  (
    n1051,
    n583,
    n1048,
    n581,
    n584
  );


  not
  g1025
  (
    n1065,
    n825
  );


  buf
  g1026
  (
    n1063,
    n1053
  );


  buf
  g1027
  (
    n1076,
    n589
  );


  buf
  g1028
  (
    n1082,
    n1052
  );


  buf
  g1029
  (
    n1072,
    n1055
  );


  not
  g1030
  (
    n1075,
    n591
  );


  not
  g1031
  (
    n1078,
    n832
  );


  not
  g1032
  (
    n1062,
    n587
  );


  not
  g1033
  (
    n1073,
    n585
  );


  not
  g1034
  (
    n1058,
    n587
  );


  not
  g1035
  (
    n1084,
    n590
  );


  xor
  g1036
  (
    n1068,
    n588,
    n1054,
    n1052
  );


  nand
  g1037
  (
    n1079,
    n588,
    n1055,
    n833
  );


  or
  g1038
  (
    n1080,
    n588,
    n1053,
    n838,
    n586
  );


  nor
  g1039
  (
    n1059,
    n1051,
    n831,
    n586,
    n837
  );


  and
  g1040
  (
    n1071,
    n1055,
    n591,
    n586,
    n834
  );


  xnor
  g1041
  (
    n1067,
    n1054,
    n1057,
    n839,
    n589
  );


  or
  g1042
  (
    n1081,
    n826,
    n1056,
    n590,
    n835
  );


  xor
  g1043
  (
    n1077,
    n1053,
    n1056,
    n590,
    n1057
  );


  and
  g1044
  (
    n1074,
    n1056,
    n828,
    n842,
    n1052
  );


  xnor
  g1045
  (
    n1060,
    n585,
    n836,
    n588,
    n591
  );


  nand
  g1046
  (
    n1069,
    n589,
    n1057,
    n587,
    n1053
  );


  and
  g1047
  (
    n1083,
    n1050,
    n589,
    n585,
    n587
  );


  nor
  g1048
  (
    n1064,
    n1056,
    n590,
    n829,
    n840
  );


  xor
  g1049
  (
    n1061,
    n830,
    n585,
    n1054,
    n827
  );


  or
  g1050
  (
    n1066,
    n841,
    n586,
    n591,
    n1057
  );


  or
  g1051
  (
    n1070,
    n592,
    n1051,
    n1052,
    n1054
  );


  not
  g1052
  (
    n1097,
    n1071
  );


  not
  g1053
  (
    n1102,
    n881
  );


  buf
  g1054
  (
    n1115,
    n1075
  );


  buf
  g1055
  (
    n1146,
    n1072
  );


  not
  g1056
  (
    n1134,
    n849
  );


  buf
  g1057
  (
    n1149,
    n865
  );


  not
  g1058
  (
    n1159,
    n1076
  );


  not
  g1059
  (
    n1104,
    n1067
  );


  buf
  g1060
  (
    n1151,
    n1062
  );


  not
  g1061
  (
    n1091,
    n1058
  );


  buf
  g1062
  (
    n1128,
    n1064
  );


  buf
  g1063
  (
    n1136,
    n1063
  );


  buf
  g1064
  (
    n1099,
    n1069
  );


  not
  g1065
  (
    n1129,
    n853
  );


  not
  g1066
  (
    n1142,
    n877
  );


  buf
  g1067
  (
    n1092,
    n1075
  );


  buf
  g1068
  (
    n1095,
    n1071
  );


  buf
  g1069
  (
    n1126,
    n1074
  );


  buf
  g1070
  (
    n1137,
    n863
  );


  buf
  g1071
  (
    n1087,
    n880
  );


  not
  g1072
  (
    n1140,
    n1065
  );


  not
  g1073
  (
    n1130,
    n851
  );


  buf
  g1074
  (
    n1119,
    n1058
  );


  buf
  g1075
  (
    n1162,
    n848
  );


  not
  g1076
  (
    n1112,
    n1069
  );


  buf
  g1077
  (
    n1135,
    n1068
  );


  not
  g1078
  (
    n1131,
    n1061
  );


  buf
  g1079
  (
    n1085,
    n1069
  );


  buf
  g1080
  (
    n1153,
    n1065
  );


  not
  g1081
  (
    n1163,
    n847
  );


  not
  g1082
  (
    n1096,
    n1060
  );


  buf
  g1083
  (
    n1148,
    n1068
  );


  buf
  g1084
  (
    n1094,
    n1065
  );


  buf
  g1085
  (
    KeyWire_0_6,
    n1076
  );


  not
  g1086
  (
    n1088,
    n1067
  );


  not
  g1087
  (
    n1143,
    n846
  );


  not
  g1088
  (
    n1121,
    n1070
  );


  not
  g1089
  (
    n1164,
    n1070
  );


  buf
  g1090
  (
    n1093,
    n1058
  );


  not
  g1091
  (
    n1105,
    n856
  );


  not
  g1092
  (
    n1132,
    n1064
  );


  buf
  g1093
  (
    KeyWire_0_28,
    n845
  );


  buf
  g1094
  (
    n1114,
    n1060
  );


  not
  g1095
  (
    n1113,
    n860
  );


  buf
  g1096
  (
    n1124,
    n1058
  );


  not
  g1097
  (
    n1133,
    n1061
  );


  buf
  g1098
  (
    n1127,
    n858
  );


  not
  g1099
  (
    n1161,
    n1069
  );


  buf
  g1100
  (
    n1141,
    n1073
  );


  not
  g1101
  (
    n1160,
    n1060
  );


  not
  g1102
  (
    n1090,
    n1059
  );


  not
  g1103
  (
    n1109,
    n864
  );


  buf
  g1104
  (
    n1125,
    n1071
  );


  not
  g1105
  (
    n1157,
    n876
  );


  buf
  g1106
  (
    n1111,
    n1076
  );


  buf
  g1107
  (
    n1158,
    n875
  );


  not
  g1108
  (
    n1106,
    n1068
  );


  not
  g1109
  (
    n1118,
    n862
  );


  not
  g1110
  (
    n1144,
    n1062
  );


  buf
  g1111
  (
    n1110,
    n1066
  );


  and
  g1112
  (
    n1145,
    n1062,
    n874,
    n1073
  );


  nand
  g1113
  (
    n1138,
    n1059,
    n867,
    n854
  );


  xnor
  g1114
  (
    n1139,
    n1074,
    n1064,
    n1066
  );


  and
  g1115
  (
    n1150,
    n1072,
    n1070,
    n844
  );


  xor
  g1116
  (
    n1103,
    n882,
    n1073,
    n868
  );


  or
  g1117
  (
    n1089,
    n843,
    n852,
    n1061
  );


  xnor
  g1118
  (
    n1101,
    n1072,
    n1075,
    n1073
  );


  or
  g1119
  (
    n1154,
    n1068,
    n1063,
    n1071
  );


  nor
  g1120
  (
    n1123,
    n850,
    n1067,
    n866
  );


  nor
  g1121
  (
    n1117,
    n1077,
    n1075,
    n1074
  );


  nor
  g1122
  (
    n1147,
    n855,
    n1063,
    n1070
  );


  nand
  g1123
  (
    n1155,
    n1059,
    n1077,
    n1074
  );


  xnor
  g1124
  (
    KeyWire_0_4,
    n1060,
    n1059,
    n871
  );


  xor
  g1125
  (
    n1156,
    n879,
    n1065,
    n1077
  );


  nand
  g1126
  (
    n1122,
    n1061,
    n1066,
    n859
  );


  xnor
  g1127
  (
    n1100,
    n1072,
    n1067,
    n861
  );


  nor
  g1128
  (
    n1108,
    n1064,
    n1076,
    n869
  );


  nor
  g1129
  (
    n1152,
    n873,
    n1066,
    n1062
  );


  and
  g1130
  (
    n1116,
    n857,
    n872,
    n1077
  );


  nor
  g1131
  (
    n1098,
    n878,
    n870,
    n1063
  );


  or
  g1132
  (
    n1166,
    n891,
    n899,
    n951,
    n929
  );


  xnor
  g1133
  (
    n1190,
    n1086,
    n906,
    n890,
    n1090
  );


  or
  g1134
  (
    n1174,
    n932,
    n927,
    n963,
    n898
  );


  xor
  g1135
  (
    n1165,
    n1088,
    n948,
    n946,
    n940
  );


  and
  g1136
  (
    n1183,
    n1086,
    n907,
    n1085,
    n926
  );


  and
  g1137
  (
    n1169,
    n888,
    n908,
    n894,
    n945
  );


  and
  g1138
  (
    n1178,
    n900,
    n955,
    n883,
    n942
  );


  nor
  g1139
  (
    n1168,
    n887,
    n1087,
    n950
  );


  nand
  g1140
  (
    n1188,
    n1087,
    n904,
    n1088,
    n1089
  );


  nor
  g1141
  (
    n1185,
    n1091,
    n917,
    n923,
    n941
  );


  xor
  g1142
  (
    n1167,
    n1090,
    n919,
    n1085,
    n962
  );


  xnor
  g1143
  (
    KeyWire_0_21,
    n952,
    n924,
    n914,
    n1087
  );


  and
  g1144
  (
    n1181,
    n1089,
    n1090,
    n910,
    n897
  );


  or
  g1145
  (
    n1170,
    n934,
    n889,
    n960,
    n901
  );


  and
  g1146
  (
    n1173,
    n956,
    n925,
    n896,
    n892
  );


  xnor
  g1147
  (
    n1191,
    n922,
    n953,
    n1086,
    n886
  );


  xnor
  g1148
  (
    n1187,
    n1088,
    n916,
    n1089,
    n913
  );


  nor
  g1149
  (
    n1179,
    n935,
    n909,
    n1086,
    n928
  );


  xor
  g1150
  (
    n1171,
    n958,
    n1091,
    n893,
    n954
  );


  xnor
  g1151
  (
    n1172,
    n905,
    n961,
    n947,
    n911
  );


  xnor
  g1152
  (
    n1175,
    n944,
    n1090,
    n912,
    n918
  );


  and
  g1153
  (
    n1184,
    n930,
    n1085,
    n957,
    n937
  );


  xor
  g1154
  (
    n1186,
    n895,
    n938,
    n936,
    n903
  );


  and
  g1155
  (
    n1180,
    n920,
    n1091,
    n939,
    n885
  );


  xor
  g1156
  (
    n1176,
    n1085,
    n1089,
    n884,
    n931
  );


  nor
  g1157
  (
    n1177,
    n959,
    n949,
    n1088,
    n933
  );


  and
  g1158
  (
    n1182,
    n943,
    n902,
    n915,
    n921
  );


  xnor
  g1159
  (
    n1195,
    n1079,
    n1189,
    n1186,
    n975
  );


  or
  g1160
  (
    n1204,
    n977,
    n1082,
    n1177
  );


  and
  g1161
  (
    n1197,
    n593,
    n1080,
    n1083,
    n592
  );


  or
  g1162
  (
    n1196,
    n1185,
    n1084,
    n1178,
    n1078
  );


  nand
  g1163
  (
    n1199,
    n1079,
    n1079,
    n1084,
    n967
  );


  and
  g1164
  (
    n1200,
    n1080,
    n1182,
    n974,
    n821
  );


  nand
  g1165
  (
    n1198,
    n972,
    n1183,
    n1083
  );


  nand
  g1166
  (
    n1202,
    n976,
    n1081,
    n1082,
    n1078
  );


  xor
  g1167
  (
    n1206,
    n1188,
    n1191,
    n592,
    n979
  );


  and
  g1168
  (
    n1207,
    n1184,
    n965,
    n966,
    n1176
  );


  xnor
  g1169
  (
    n1205,
    n1083,
    n971,
    n1081,
    n1080
  );


  xnor
  g1170
  (
    n1194,
    n964,
    n1187,
    n969,
    n1082
  );


  or
  g1171
  (
    KeyWire_0_15,
    n1078,
    n968,
    n1181,
    n1081
  );


  nor
  g1172
  (
    n1201,
    n1081,
    n593,
    n970,
    n1079
  );


  or
  g1173
  (
    n1203,
    n1179,
    n1078,
    n1190,
    n1180
  );


  nor
  g1174
  (
    n1192,
    n1080,
    n978,
    n592,
    n973
  );


  xnor
  g1175
  (
    n1221,
    n1084,
    n1205,
    n1095,
    n1092
  );


  xnor
  g1176
  (
    n1211,
    n1098,
    n987,
    n1206,
    n993
  );


  xnor
  g1177
  (
    n1214,
    n982,
    n986,
    n1204,
    n1093
  );


  xnor
  g1178
  (
    n1217,
    n992,
    n1097,
    n1093,
    n1202
  );


  xor
  g1179
  (
    n1212,
    n1203,
    n1096,
    n988,
    n1097
  );


  nand
  g1180
  (
    n1216,
    n1094,
    n980,
    n985,
    n1096
  );


  xnor
  g1181
  (
    n1218,
    n1199,
    n990,
    n1200,
    n1198
  );


  or
  g1182
  (
    n1220,
    n991,
    n1092,
    n1093
  );


  xnor
  g1183
  (
    n1213,
    n1196,
    n983,
    n1094
  );


  xnor
  g1184
  (
    n1215,
    n1193,
    n1092,
    n1098,
    n1195
  );


  and
  g1185
  (
    n1208,
    n1201,
    n1095,
    n1096,
    n1197
  );


  nor
  g1186
  (
    n1209,
    n994,
    n1095,
    n1096,
    n1094
  );


  xor
  g1187
  (
    n1210,
    n1097,
    n984,
    n1084,
    n1091
  );


  and
  g1188
  (
    n1219,
    n1095,
    n981,
    n1194,
    n1192
  );


  xor
  g1189
  (
    n1222,
    n989,
    n1098,
    n1093,
    n1097
  );


  nor
  g1190
  (
    n1231,
    n1100,
    n1104,
    n1103
  );


  and
  g1191
  (
    n1226,
    n1215,
    n1101,
    n1213,
    n1211
  );


  xnor
  g1192
  (
    n1230,
    n1106,
    n1106,
    n1105,
    n1099
  );


  nand
  g1193
  (
    n1227,
    n1222,
    n1105,
    n1217,
    n1218
  );


  and
  g1194
  (
    n1224,
    n1221,
    n1101,
    n1220
  );


  or
  g1195
  (
    n1232,
    n1106,
    n1098,
    n1102,
    n1104
  );


  or
  g1196
  (
    n1223,
    n1100,
    n1105,
    n1102
  );


  xor
  g1197
  (
    n1229,
    n1102,
    n1100,
    n1103,
    n1216
  );


  or
  g1198
  (
    n1233,
    n1107,
    n1100,
    n1104,
    n1101
  );


  nor
  g1199
  (
    n1225,
    n1106,
    n1107,
    n1104,
    n1214
  );


  nand
  g1200
  (
    n1228,
    n1103,
    n1102,
    n1099,
    n1219
  );


  and
  g1201
  (
    n1234,
    n1212,
    n1107,
    n1099
  );


  not
  g1202
  (
    n1248,
    n1223
  );


  buf
  g1203
  (
    n1251,
    n1224
  );


  buf
  g1204
  (
    n1235,
    n1223
  );


  not
  g1205
  (
    n1253,
    n1228
  );


  buf
  g1206
  (
    n1238,
    n1107
  );


  not
  g1207
  (
    n1256,
    n1227
  );


  buf
  g1208
  (
    n1237,
    n1224
  );


  not
  g1209
  (
    n1254,
    n1228
  );


  not
  g1210
  (
    n1240,
    n1226
  );


  buf
  g1211
  (
    n1239,
    n1225
  );


  not
  g1212
  (
    n1255,
    n1227
  );


  buf
  g1213
  (
    n1247,
    n1225
  );


  buf
  g1214
  (
    n1242,
    n1108
  );


  buf
  g1215
  (
    n1245,
    n1227
  );


  not
  g1216
  (
    n1243,
    n1224
  );


  not
  g1217
  (
    n1249,
    n1226
  );


  buf
  g1218
  (
    n1236,
    n1225
  );


  buf
  g1219
  (
    n1241,
    n1108
  );


  buf
  g1220
  (
    n1246,
    n1108
  );


  buf
  g1221
  (
    n1244,
    n1226
  );


  nand
  g1222
  (
    n1257,
    n1227,
    n1226
  );


  xor
  g1223
  (
    n1250,
    n1225,
    n1224,
    n1108,
    n1109
  );


  xnor
  g1224
  (
    n1258,
    n1109,
    n1223,
    n1228
  );


  nand
  g1225
  (
    n1252,
    n1110,
    n1109,
    n1223
  );


  not
  g1226
  (
    n1259,
    n1238
  );


  not
  g1227
  (
    n1266,
    n1241
  );


  not
  g1228
  (
    n1262,
    n1240
  );


  not
  g1229
  (
    n1263,
    n1239
  );


  buf
  g1230
  (
    n1260,
    n1241
  );


  not
  g1231
  (
    n1265,
    n1236
  );


  buf
  g1232
  (
    n1264,
    n1239
  );


  not
  g1233
  (
    n1268,
    n1240
  );


  buf
  g1234
  (
    n1261,
    n1235
  );


  buf
  g1235
  (
    n1267,
    n1237
  );


  buf
  g1236
  (
    n1269,
    n1261
  );


  not
  g1237
  (
    n1280,
    n1259
  );


  buf
  g1238
  (
    n1271,
    n1262
  );


  buf
  g1239
  (
    n1278,
    n1259
  );


  not
  g1240
  (
    n1284,
    n1262
  );


  not
  g1241
  (
    n1283,
    n1260
  );


  buf
  g1242
  (
    n1273,
    n1262
  );


  buf
  g1243
  (
    n1275,
    n1261
  );


  buf
  g1244
  (
    n1286,
    n1261
  );


  not
  g1245
  (
    n1285,
    n1259
  );


  buf
  g1246
  (
    n1272,
    n1260
  );


  not
  g1247
  (
    n1270,
    n1262
  );


  buf
  g1248
  (
    n1274,
    n1259
  );


  buf
  g1249
  (
    n1282,
    n1260
  );


  buf
  g1250
  (
    n1277,
    n1260
  );


  buf
  g1251
  (
    n1276,
    n1261
  );


  not
  g1252
  (
    n1279,
    n1263
  );


  buf
  g1253
  (
    n1281,
    n1263
  );


  buf
  g1254
  (
    n1291,
    n1278
  );


  buf
  g1255
  (
    n1315,
    n1112
  );


  buf
  g1256
  (
    n1344,
    n1273
  );


  buf
  g1257
  (
    n1325,
    n1285
  );


  not
  g1258
  (
    n1326,
    n1269
  );


  not
  g1259
  (
    n1314,
    n1280
  );


  buf
  g1260
  (
    n1331,
    n1286
  );


  not
  g1261
  (
    n1335,
    n1270
  );


  not
  g1262
  (
    n1310,
    n1278
  );


  not
  g1263
  (
    n1312,
    n1283
  );


  not
  g1264
  (
    n1334,
    n1277
  );


  buf
  g1265
  (
    n1336,
    n1284
  );


  buf
  g1266
  (
    n1309,
    n1277
  );


  not
  g1267
  (
    n1339,
    n1271
  );


  not
  g1268
  (
    KeyWire_0_30,
    n1286
  );


  buf
  g1269
  (
    n1332,
    n1279
  );


  buf
  g1270
  (
    n1296,
    n1001
  );


  buf
  g1271
  (
    n1289,
    n1269
  );


  buf
  g1272
  (
    n1323,
    n1280
  );


  buf
  g1273
  (
    n1316,
    n1274
  );


  not
  g1274
  (
    n1299,
    n1277
  );


  not
  g1275
  (
    n1292,
    n996
  );


  not
  g1276
  (
    n1295,
    n1000
  );


  buf
  g1277
  (
    n1294,
    n1276
  );


  not
  g1278
  (
    n1357,
    n1271
  );


  buf
  g1279
  (
    n1288,
    n1270
  );


  buf
  g1280
  (
    n1307,
    n1275
  );


  not
  g1281
  (
    n1303,
    n1284
  );


  buf
  g1282
  (
    n1293,
    n1112
  );


  not
  g1283
  (
    n1356,
    n1271
  );


  buf
  g1284
  (
    n1321,
    n1282
  );


  not
  g1285
  (
    n1329,
    n1276
  );


  buf
  g1286
  (
    n1300,
    n1269
  );


  buf
  g1287
  (
    n1298,
    n1275
  );


  not
  g1288
  (
    KeyWire_0_9,
    n1285
  );


  buf
  g1289
  (
    n1330,
    n1286
  );


  not
  g1290
  (
    n1345,
    n1272
  );


  buf
  g1291
  (
    n1318,
    n1112
  );


  buf
  g1292
  (
    n1317,
    n1274
  );


  not
  g1293
  (
    n1324,
    n1281
  );


  not
  g1294
  (
    n1343,
    n1276
  );


  buf
  g1295
  (
    n1352,
    n1283
  );


  buf
  g1296
  (
    n1354,
    n1275
  );


  buf
  g1297
  (
    n1311,
    n1279
  );


  buf
  g1298
  (
    n1320,
    n1110
  );


  not
  g1299
  (
    n1328,
    n1283
  );


  not
  g1300
  (
    n1340,
    n998
  );


  buf
  g1301
  (
    n1327,
    n1111
  );


  buf
  g1302
  (
    n1301,
    n1273
  );


  not
  g1303
  (
    n1337,
    n1282
  );


  buf
  g1304
  (
    KeyWire_0_7,
    n1280
  );


  not
  g1305
  (
    n1358,
    n1270
  );


  buf
  g1306
  (
    n1350,
    n1273
  );


  not
  g1307
  (
    n1304,
    n1283
  );


  buf
  g1308
  (
    n1347,
    n1284
  );


  not
  g1309
  (
    n1319,
    n1284
  );


  not
  g1310
  (
    n1351,
    n1271
  );


  not
  g1311
  (
    n1308,
    n1281
  );


  not
  g1312
  (
    n1302,
    n1272
  );


  not
  g1313
  (
    n1341,
    n1285
  );


  buf
  g1314
  (
    n1305,
    n1003
  );


  not
  g1315
  (
    n1313,
    n1281
  );


  not
  g1316
  (
    n1342,
    n997
  );


  buf
  g1317
  (
    n1306,
    n1280
  );


  buf
  g1318
  (
    n1287,
    n1111
  );


  nand
  g1319
  (
    n1353,
    n1278,
    n1002,
    n1279
  );


  xnor
  g1320
  (
    n1333,
    n1275,
    n1110,
    n1277,
    n1285
  );


  xor
  g1321
  (
    n1355,
    n1270,
    n1286,
    n1273,
    n1274
  );


  xor
  g1322
  (
    n1322,
    n1269,
    n1281,
    n1278,
    n999
  );


  and
  g1323
  (
    n1338,
    n1110,
    n1272,
    n1276
  );


  nand
  g1324
  (
    n1297,
    n995,
    n1274,
    n1111
  );


  xnor
  g1325
  (
    n1290,
    n1279,
    n1282,
    n1112
  );


  buf
  g1326
  (
    n1586,
    n1251
  );


  buf
  g1327
  (
    n1415,
    n1324
  );


  buf
  g1328
  (
    n1469,
    n1007
  );


  buf
  g1329
  (
    n1587,
    n1325
  );


  buf
  g1330
  (
    n1392,
    n1328
  );


  not
  g1331
  (
    n1515,
    n1321
  );


  not
  g1332
  (
    n1424,
    n1231
  );


  buf
  g1333
  (
    n1579,
    n1301
  );


  buf
  g1334
  (
    n1481,
    n1249
  );


  not
  g1335
  (
    n1466,
    n1253
  );


  not
  g1336
  (
    n1482,
    n1116
  );


  buf
  g1337
  (
    n1369,
    n1344
  );


  not
  g1338
  (
    n1542,
    n1113
  );


  not
  g1339
  (
    n1370,
    n1339
  );


  not
  g1340
  (
    n1366,
    n1306
  );


  not
  g1341
  (
    n1551,
    n1241
  );


  buf
  g1342
  (
    n1390,
    n1231
  );


  buf
  g1343
  (
    n1381,
    n1254
  );


  not
  g1344
  (
    n1589,
    n1297
  );


  not
  g1345
  (
    n1590,
    n1328
  );


  buf
  g1346
  (
    n1486,
    n1329
  );


  not
  g1347
  (
    n1436,
    n1242
  );


  not
  g1348
  (
    n1537,
    n1329
  );


  buf
  g1349
  (
    n1489,
    n1297
  );


  not
  g1350
  (
    n1360,
    n1251
  );


  not
  g1351
  (
    n1536,
    n1250
  );


  not
  g1352
  (
    n1543,
    n1319
  );


  not
  g1353
  (
    n1437,
    n1334
  );


  buf
  g1354
  (
    n1376,
    n1250
  );


  buf
  g1355
  (
    n1566,
    n1289
  );


  not
  g1356
  (
    n1539,
    n1344
  );


  not
  g1357
  (
    n1457,
    n1343
  );


  not
  g1358
  (
    n1364,
    n1232
  );


  not
  g1359
  (
    n1528,
    n1231
  );


  not
  g1360
  (
    n1388,
    n1312
  );


  not
  g1361
  (
    n1496,
    n1334
  );


  buf
  g1362
  (
    n1491,
    n1332
  );


  buf
  g1363
  (
    n1545,
    n1333
  );


  not
  g1364
  (
    n1401,
    n1250
  );


  not
  g1365
  (
    n1488,
    n1296
  );


  buf
  g1366
  (
    n1588,
    n1255
  );


  buf
  g1367
  (
    n1581,
    n1253
  );


  not
  g1368
  (
    n1474,
    n1318
  );


  not
  g1369
  (
    n1449,
    n1312
  );


  buf
  g1370
  (
    n1386,
    n1307
  );


  not
  g1371
  (
    n1414,
    n1320
  );


  buf
  g1372
  (
    KeyWire_0_19,
    n1330
  );


  not
  g1373
  (
    n1442,
    n1336
  );


  not
  g1374
  (
    n1490,
    n1115
  );


  buf
  g1375
  (
    n1406,
    n1316
  );


  buf
  g1376
  (
    n1432,
    n1342
  );


  not
  g1377
  (
    n1361,
    n1335
  );


  not
  g1378
  (
    n1402,
    n1004
  );


  buf
  g1379
  (
    n1571,
    n1306
  );


  buf
  g1380
  (
    n1529,
    n1315
  );


  buf
  g1381
  (
    n1525,
    n1243
  );


  not
  g1382
  (
    n1384,
    n1254
  );


  not
  g1383
  (
    n1371,
    n1230
  );


  not
  g1384
  (
    n1487,
    n1317
  );


  buf
  g1385
  (
    n1417,
    n1249
  );


  not
  g1386
  (
    n1577,
    n1293
  );


  buf
  g1387
  (
    n1429,
    n1305
  );


  buf
  g1388
  (
    n1404,
    n1299
  );


  buf
  g1389
  (
    n1483,
    n1255
  );


  buf
  g1390
  (
    n1391,
    n1247
  );


  buf
  g1391
  (
    n1430,
    n1295
  );


  not
  g1392
  (
    n1478,
    n1234
  );


  buf
  g1393
  (
    n1476,
    n1319
  );


  buf
  g1394
  (
    n1573,
    n1247
  );


  buf
  g1395
  (
    n1428,
    n1207
  );


  not
  g1396
  (
    n1544,
    n1321
  );


  buf
  g1397
  (
    n1484,
    n1243
  );


  not
  g1398
  (
    n1519,
    n1318
  );


  not
  g1399
  (
    n1568,
    n1320
  );


  buf
  g1400
  (
    n1574,
    n1315
  );


  buf
  g1401
  (
    n1421,
    n1012
  );


  buf
  g1402
  (
    n1452,
    n1324
  );


  not
  g1403
  (
    n1526,
    n1308
  );


  not
  g1404
  (
    n1368,
    n1305
  );


  not
  g1405
  (
    n1555,
    n1310
  );


  not
  g1406
  (
    n1565,
    n1331
  );


  not
  g1407
  (
    n1359,
    n1337
  );


  buf
  g1408
  (
    n1448,
    n1326
  );


  not
  g1409
  (
    n1471,
    n1009
  );


  not
  g1410
  (
    n1470,
    n1242
  );


  buf
  g1411
  (
    n1382,
    n1298
  );


  not
  g1412
  (
    n1434,
    n1244
  );


  not
  g1413
  (
    n1582,
    n1344
  );


  buf
  g1414
  (
    n1462,
    n1312
  );


  not
  g1415
  (
    n1441,
    n1304
  );


  not
  g1416
  (
    n1563,
    n1116
  );


  buf
  g1417
  (
    n1499,
    n1317
  );


  buf
  g1418
  (
    n1372,
    n1231
  );


  buf
  g1419
  (
    n1527,
    n1294
  );


  not
  g1420
  (
    n1497,
    n1315
  );


  not
  g1421
  (
    n1422,
    n1339
  );


  buf
  g1422
  (
    n1451,
    n1249
  );


  buf
  g1423
  (
    n1518,
    n1310
  );


  not
  g1424
  (
    n1559,
    n1323
  );


  not
  g1425
  (
    n1547,
    n1302
  );


  not
  g1426
  (
    n1400,
    n1323
  );


  not
  g1427
  (
    n1500,
    n1343
  );


  not
  g1428
  (
    n1458,
    n1319
  );


  not
  g1429
  (
    n1535,
    n1309
  );


  buf
  g1430
  (
    n1447,
    n1314
  );


  buf
  g1431
  (
    n1514,
    n1243
  );


  not
  g1432
  (
    n1585,
    n1250
  );


  not
  g1433
  (
    n1405,
    n1322
  );


  buf
  g1434
  (
    n1549,
    n1332
  );


  buf
  g1435
  (
    n1494,
    n1312
  );


  not
  g1436
  (
    n1572,
    n1287
  );


  buf
  g1437
  (
    n1367,
    n1311
  );


  buf
  g1438
  (
    n1440,
    n1115
  );


  buf
  g1439
  (
    n1377,
    n1243
  );


  buf
  g1440
  (
    n1517,
    n1317
  );


  buf
  g1441
  (
    n1465,
    n1332
  );


  buf
  g1442
  (
    n1455,
    n1323
  );


  buf
  g1443
  (
    n1420,
    n1251
  );


  not
  g1444
  (
    n1416,
    n1244
  );


  buf
  g1445
  (
    n1562,
    n1336
  );


  buf
  g1446
  (
    n1530,
    n1306
  );


  buf
  g1447
  (
    n1385,
    n1330
  );


  buf
  g1448
  (
    n1433,
    n1320
  );


  not
  g1449
  (
    n1495,
    n1308
  );


  not
  g1450
  (
    n1459,
    n1233
  );


  buf
  g1451
  (
    n1550,
    n1326
  );


  not
  g1452
  (
    n1541,
    n1256
  );


  not
  g1453
  (
    n1375,
    n1249
  );


  buf
  g1454
  (
    n1521,
    n1295
  );


  buf
  g1455
  (
    n1560,
    n1289
  );


  buf
  g1456
  (
    n1473,
    n1296
  );


  buf
  g1457
  (
    n1576,
    n1340
  );


  buf
  g1458
  (
    n1389,
    n1311
  );


  buf
  g1459
  (
    n1511,
    n1248
  );


  buf
  g1460
  (
    n1394,
    n1337
  );


  not
  g1461
  (
    n1443,
    n1335
  );


  not
  g1462
  (
    n1399,
    n1298
  );


  not
  g1463
  (
    n1524,
    n1294
  );


  buf
  g1464
  (
    n1591,
    n1313
  );


  buf
  g1465
  (
    n1533,
    n1328
  );


  buf
  g1466
  (
    n1523,
    n1234
  );


  buf
  g1467
  (
    n1395,
    n1245
  );


  buf
  g1468
  (
    n1554,
    n1293
  );


  buf
  g1469
  (
    n1463,
    n1006
  );


  buf
  g1470
  (
    n1507,
    n1345
  );


  not
  g1471
  (
    n1410,
    n1327
  );


  buf
  g1472
  (
    n1584,
    n1229
  );


  buf
  g1473
  (
    n1431,
    n1242
  );


  not
  g1474
  (
    n1540,
    n1317
  );


  buf
  g1475
  (
    n1553,
    n1338
  );


  not
  g1476
  (
    n1479,
    n1335
  );


  buf
  g1477
  (
    n1504,
    n1335
  );


  not
  g1478
  (
    n1467,
    n1301
  );


  not
  g1479
  (
    n1450,
    n1326
  );


  buf
  g1480
  (
    n1509,
    n1114
  );


  not
  g1481
  (
    n1387,
    n1288
  );


  not
  g1482
  (
    n1461,
    n1114
  );


  not
  g1483
  (
    n1444,
    n1113
  );


  buf
  g1484
  (
    n1580,
    n1328
  );


  not
  g1485
  (
    n1446,
    n1305
  );


  buf
  g1486
  (
    n1561,
    n1322
  );


  not
  g1487
  (
    n1439,
    n1309
  );


  not
  g1488
  (
    n1583,
    n1255
  );


  buf
  g1489
  (
    n1556,
    n1301
  );


  buf
  g1490
  (
    n1508,
    n1301
  );


  not
  g1491
  (
    n1454,
    n1307
  );


  buf
  g1492
  (
    n1485,
    n1232
  );


  not
  g1493
  (
    n1503,
    n1315
  );


  buf
  g1494
  (
    n1522,
    n1252
  );


  not
  g1495
  (
    n1492,
    n1232
  );


  not
  g1496
  (
    n1569,
    n1332
  );


  buf
  g1497
  (
    n1567,
    n1309
  );


  not
  g1498
  (
    n1426,
    n1337
  );


  buf
  g1499
  (
    n1380,
    n1234
  );


  buf
  g1500
  (
    n1501,
    n1008
  );


  buf
  g1501
  (
    n1412,
    n1336
  );


  buf
  g1502
  (
    n1397,
    n1252
  );


  buf
  g1503
  (
    n1411,
    n1229
  );


  buf
  g1504
  (
    n1513,
    n1230
  );


  buf
  g1505
  (
    n1413,
    n1343
  );


  not
  g1506
  (
    n1468,
    n1253
  );


  buf
  g1507
  (
    n1419,
    n1329
  );


  buf
  g1508
  (
    n1538,
    n1339
  );


  buf
  g1509
  (
    n1578,
    n1341
  );


  not
  g1510
  (
    n1365,
    n1246
  );


  not
  g1511
  (
    n1362,
    n1302
  );


  buf
  g1512
  (
    n1464,
    n1297
  );


  not
  g1513
  (
    n1534,
    n1313
  );


  not
  g1514
  (
    n1456,
    n1256
  );


  buf
  g1515
  (
    n1408,
    n1327
  );


  not
  g1516
  (
    n1558,
    n1304
  );


  not
  g1517
  (
    n1512,
    n1307
  );


  buf
  g1518
  (
    n1546,
    n1254
  );


  not
  g1519
  (
    n1418,
    n1321
  );


  buf
  g1520
  (
    n1373,
    n1314
  );


  buf
  g1521
  (
    n1407,
    n1340
  );


  nand
  g1522
  (
    n1435,
    n1295,
    n1341,
    n1302,
    n1290
  );


  xnor
  g1523
  (
    n1532,
    n1011,
    n1293,
    n1324,
    n1287
  );


  xor
  g1524
  (
    n1363,
    n1311,
    n1305,
    n1318,
    n1233
  );


  nand
  g1525
  (
    n1548,
    n1327,
    n1287,
    n1322,
    n1207
  );


  xnor
  g1526
  (
    n1506,
    n1336,
    n1248,
    n1114,
    n1232
  );


  xor
  g1527
  (
    n1505,
    n1116,
    n1299,
    n1292,
    n1115
  );


  nand
  g1528
  (
    n1472,
    n1290,
    n1338,
    n1316,
    n1255
  );


  xnor
  g1529
  (
    n1423,
    n1291,
    n1291,
    n1244,
    n1241
  );


  nor
  g1530
  (
    n1564,
    n1251,
    n1246,
    n1327,
    n1290
  );


  and
  g1531
  (
    n1557,
    n1324,
    n1247,
    n1010,
    n1242
  );


  xnor
  g1532
  (
    n1425,
    n1321,
    n1325,
    n1331,
    n1248
  );


  or
  g1533
  (
    n1383,
    n1331,
    n1294,
    n1303
  );


  and
  g1534
  (
    n1531,
    n1341,
    n1340,
    n1297,
    n1306
  );


  and
  g1535
  (
    n1409,
    n1308,
    n1333,
    n1298,
    n1233
  );


  and
  g1536
  (
    n1438,
    n1294,
    n1309,
    n1325,
    n1342
  );


  and
  g1537
  (
    n1393,
    n1303,
    n1322,
    n1245,
    n1295
  );


  or
  g1538
  (
    n1445,
    n1314,
    n1288,
    n1310,
    n1292
  );


  and
  g1539
  (
    n1480,
    n1310,
    n1288,
    n1114,
    n1290
  );


  xnor
  g1540
  (
    n1374,
    n1246,
    n1244,
    n1230,
    n1229
  );


  xnor
  g1541
  (
    n1510,
    n1343,
    n1113,
    n1246,
    n1230
  );


  or
  g1542
  (
    n1453,
    n1325,
    n1233,
    n1291,
    n1299
  );


  xor
  g1543
  (
    n1427,
    n1245,
    n1115,
    n1314,
    n1300
  );


  nor
  g1544
  (
    n1379,
    n1299,
    n1326,
    n1331,
    n1245
  );


  and
  g1545
  (
    n1396,
    n1330,
    n1288,
    n1316,
    n1344
  );


  xnor
  g1546
  (
    n1516,
    n1320,
    n1293,
    n1340,
    n1338
  );


  nand
  g1547
  (
    n1378,
    n1318,
    n1113,
    n1333,
    n1298
  );


  xnor
  g1548
  (
    n1520,
    n1287,
    n1289,
    n1292,
    n1334
  );


  xnor
  g1549
  (
    n1477,
    n1316,
    n1248,
    n1308,
    n1254
  );


  xnor
  g1550
  (
    n1502,
    n1300,
    n1116,
    n1252,
    n1342
  );


  or
  g1551
  (
    n1570,
    n1296,
    n1252,
    n1292,
    n1330
  );


  and
  g1552
  (
    n1398,
    n1339,
    n1329,
    n1307,
    n1338
  );


  xnor
  g1553
  (
    n1460,
    n1005,
    n1303,
    n1319,
    n1289
  );


  xnor
  g1554
  (
    n1575,
    n1304,
    n1341,
    n1247,
    n1300
  );


  or
  g1555
  (
    n1403,
    n1342,
    n1323,
    n1304,
    n1291
  );


  xor
  g1556
  (
    n1552,
    n1311,
    n1300,
    n1229,
    n1337
  );


  nor
  g1557
  (
    KeyWire_0_18,
    n1333,
    n1253,
    n1334,
    n1296
  );


  and
  g1558
  (
    n1498,
    n1234,
    n1313,
    n1302
  );


  buf
  g1559
  (
    n1597,
    n1131
  );


  buf
  g1560
  (
    KeyWire_0_20,
    n1533
  );


  not
  g1561
  (
    n1601,
    n1427
  );


  buf
  g1562
  (
    n1799,
    n1137
  );


  buf
  g1563
  (
    n1810,
    n1539
  );


  not
  g1564
  (
    n1802,
    n1510
  );


  not
  g1565
  (
    n1788,
    n1533
  );


  not
  g1566
  (
    n1605,
    n593
  );


  not
  g1567
  (
    n1742,
    n1537
  );


  not
  g1568
  (
    n1855,
    n1542
  );


  not
  g1569
  (
    n1781,
    n1121
  );


  buf
  g1570
  (
    n1666,
    n1523
  );


  buf
  g1571
  (
    n1770,
    n1372
  );


  not
  g1572
  (
    n1661,
    n1021
  );


  not
  g1573
  (
    n1740,
    n1485
  );


  not
  g1574
  (
    n1596,
    n1122
  );


  buf
  g1575
  (
    n1704,
    n1418
  );


  buf
  g1576
  (
    n1752,
    n1542
  );


  buf
  g1577
  (
    n1638,
    n1152
  );


  buf
  g1578
  (
    n1845,
    n1495
  );


  not
  g1579
  (
    n1634,
    n1122
  );


  buf
  g1580
  (
    n1633,
    n1144
  );


  buf
  g1581
  (
    n1644,
    n1121
  );


  buf
  g1582
  (
    n1827,
    n1142
  );


  buf
  g1583
  (
    n1785,
    n1136
  );


  buf
  g1584
  (
    n1631,
    n1267
  );


  buf
  g1585
  (
    n1860,
    n1406
  );


  not
  g1586
  (
    n1805,
    n1256
  );


  buf
  g1587
  (
    n1608,
    n1151
  );


  buf
  g1588
  (
    n1739,
    n1435
  );


  buf
  g1589
  (
    n1617,
    n1548
  );


  not
  g1590
  (
    n1690,
    n1517
  );


  buf
  g1591
  (
    n1843,
    n1526
  );


  not
  g1592
  (
    n1763,
    n1531
  );


  buf
  g1593
  (
    n1736,
    n1144
  );


  buf
  g1594
  (
    n1602,
    n1521
  );


  not
  g1595
  (
    n1754,
    n1135
  );


  not
  g1596
  (
    n1723,
    n1424
  );


  not
  g1597
  (
    n1636,
    n1157
  );


  buf
  g1598
  (
    n1741,
    n1517
  );


  buf
  g1599
  (
    n1794,
    n1510
  );


  not
  g1600
  (
    n1701,
    n1361
  );


  buf
  g1601
  (
    n1751,
    n1547
  );


  not
  g1602
  (
    n1619,
    n1023
  );


  buf
  g1603
  (
    n1700,
    n1267
  );


  not
  g1604
  (
    n1643,
    n1131
  );


  buf
  g1605
  (
    n1696,
    n1502
  );


  buf
  g1606
  (
    n1773,
    n1155
  );


  buf
  g1607
  (
    n1728,
    n1134
  );


  not
  g1608
  (
    n1823,
    n1151
  );


  buf
  g1609
  (
    n1651,
    n1154
  );


  buf
  g1610
  (
    n1657,
    n1436
  );


  buf
  g1611
  (
    n1642,
    n1442
  );


  not
  g1612
  (
    n1618,
    n1535
  );


  not
  g1613
  (
    n1777,
    n1536
  );


  not
  g1614
  (
    n1613,
    n1461
  );


  not
  g1615
  (
    n1746,
    n1028
  );


  buf
  g1616
  (
    n1796,
    n1540
  );


  buf
  g1617
  (
    n1852,
    n1519
  );


  buf
  g1618
  (
    n1635,
    n1141
  );


  not
  g1619
  (
    n1820,
    n1524
  );


  not
  g1620
  (
    n1665,
    n1146
  );


  buf
  g1621
  (
    n1699,
    n1135
  );


  buf
  g1622
  (
    n1679,
    n1537
  );


  buf
  g1623
  (
    n1790,
    n1473
  );


  not
  g1624
  (
    n1615,
    n1503
  );


  buf
  g1625
  (
    n1705,
    n1129
  );


  not
  g1626
  (
    n1603,
    n1149
  );


  buf
  g1627
  (
    n1767,
    n1482
  );


  buf
  g1628
  (
    n1819,
    n1153
  );


  not
  g1629
  (
    n1744,
    n1462
  );


  not
  g1630
  (
    n1821,
    n1149
  );


  buf
  g1631
  (
    n1832,
    n1123
  );


  buf
  g1632
  (
    n1667,
    n1526
  );


  buf
  g1633
  (
    n1645,
    n1145
  );


  not
  g1634
  (
    n1656,
    n1530
  );


  buf
  g1635
  (
    n1851,
    n1438
  );


  not
  g1636
  (
    n1839,
    n1016
  );


  buf
  g1637
  (
    n1726,
    n1120
  );


  not
  g1638
  (
    n1753,
    n1513
  );


  buf
  g1639
  (
    n1664,
    n1147
  );


  not
  g1640
  (
    n1652,
    n1382
  );


  not
  g1641
  (
    n1857,
    n1128
  );


  buf
  g1642
  (
    n1594,
    n1159
  );


  buf
  g1643
  (
    n1717,
    n1157
  );


  not
  g1644
  (
    n1674,
    n1540
  );


  not
  g1645
  (
    n1778,
    n1134
  );


  not
  g1646
  (
    n1691,
    n1139
  );


  not
  g1647
  (
    n1765,
    n1147
  );


  not
  g1648
  (
    n1648,
    n1394
  );


  not
  g1649
  (
    n1818,
    n1143
  );


  buf
  g1650
  (
    n1621,
    n1143
  );


  not
  g1651
  (
    n1609,
    n1504
  );


  buf
  g1652
  (
    n1676,
    n1534
  );


  not
  g1653
  (
    n1620,
    n1265
  );


  buf
  g1654
  (
    n1738,
    n1157
  );


  buf
  g1655
  (
    n1853,
    n1152
  );


  buf
  g1656
  (
    n1858,
    n1160
  );


  buf
  g1657
  (
    n1693,
    n1430
  );


  buf
  g1658
  (
    n1782,
    n1022
  );


  buf
  g1659
  (
    n1737,
    n1156
  );


  buf
  g1660
  (
    n1817,
    n1138
  );


  not
  g1661
  (
    n1718,
    n1264
  );


  buf
  g1662
  (
    n1686,
    n1266
  );


  not
  g1663
  (
    n1842,
    n1128
  );


  not
  g1664
  (
    n1775,
    n1157
  );


  not
  g1665
  (
    n1724,
    n1416
  );


  not
  g1666
  (
    n1716,
    n1136
  );


  not
  g1667
  (
    n1720,
    n1547
  );


  buf
  g1668
  (
    n1806,
    n1523
  );


  not
  g1669
  (
    n1703,
    n1525
  );


  buf
  g1670
  (
    n1761,
    n1145
  );


  buf
  g1671
  (
    n1830,
    n1548
  );


  not
  g1672
  (
    n1797,
    n1405
  );


  buf
  g1673
  (
    n1684,
    n1486
  );


  buf
  g1674
  (
    n1706,
    n1545
  );


  buf
  g1675
  (
    KeyWire_0_25,
    n1506
  );


  buf
  g1676
  (
    n1688,
    n1444
  );


  buf
  g1677
  (
    n1721,
    n1428
  );


  not
  g1678
  (
    n1628,
    n1540
  );


  buf
  g1679
  (
    n1829,
    n1265
  );


  buf
  g1680
  (
    n1697,
    n1371
  );


  buf
  g1681
  (
    n1756,
    n1409
  );


  buf
  g1682
  (
    n1670,
    n1162
  );


  not
  g1683
  (
    n1623,
    n1266
  );


  buf
  g1684
  (
    n1814,
    n1142
  );


  not
  g1685
  (
    n1774,
    n1150
  );


  buf
  g1686
  (
    n1807,
    n1120
  );


  buf
  g1687
  (
    n1825,
    n1396
  );


  not
  g1688
  (
    n1840,
    n1496
  );


  not
  g1689
  (
    n1816,
    n1538
  );


  not
  g1690
  (
    n1592,
    n1376
  );


  buf
  g1691
  (
    n1713,
    n1147
  );


  buf
  g1692
  (
    n1624,
    n1136
  );


  buf
  g1693
  (
    n1764,
    n1121
  );


  not
  g1694
  (
    n1727,
    n1160
  );


  not
  g1695
  (
    n1714,
    n1470
  );


  not
  g1696
  (
    KeyWire_0_26,
    n1159
  );


  buf
  g1697
  (
    n1598,
    n1528
  );


  buf
  g1698
  (
    n1672,
    n1378
  );


  not
  g1699
  (
    n1712,
    n1489
  );


  not
  g1700
  (
    n1847,
    n1119
  );


  buf
  g1701
  (
    n1707,
    n1540
  );


  buf
  g1702
  (
    n1834,
    n1163
  );


  buf
  g1703
  (
    n1689,
    n1464
  );


  buf
  g1704
  (
    n1828,
    n1164
  );


  buf
  g1705
  (
    n1692,
    n1137
  );


  not
  g1706
  (
    n1604,
    n1515
  );


  buf
  g1707
  (
    n1622,
    n1431
  );


  not
  g1708
  (
    n1732,
    n594
  );


  not
  g1709
  (
    n1812,
    n1119
  );


  not
  g1710
  (
    n1607,
    n1161
  );


  buf
  g1711
  (
    n1715,
    n1541
  );


  not
  g1712
  (
    n1861,
    n1144
  );


  buf
  g1713
  (
    n1668,
    n1140
  );


  not
  g1714
  (
    n1722,
    n1129
  );


  buf
  g1715
  (
    n1698,
    n1440
  );


  buf
  g1716
  (
    n1862,
    n1392
  );


  buf
  g1717
  (
    n1610,
    n1487
  );


  not
  g1718
  (
    n1757,
    n1393
  );


  not
  g1719
  (
    n1729,
    n1366
  );


  not
  g1720
  (
    n1629,
    n1256
  );


  not
  g1721
  (
    n1687,
    n1151
  );


  buf
  g1722
  (
    n1683,
    n1538
  );


  buf
  g1723
  (
    n1606,
    n1447
  );


  not
  g1724
  (
    n1616,
    n1140
  );


  buf
  g1725
  (
    n1694,
    n1529
  );


  buf
  g1726
  (
    n1653,
    n1544
  );


  not
  g1727
  (
    n1748,
    n1018
  );


  not
  g1728
  (
    n1760,
    n1119
  );


  buf
  g1729
  (
    n1669,
    n1535
  );


  buf
  g1730
  (
    n1789,
    n1377
  );


  buf
  g1731
  (
    n1640,
    n1543
  );


  buf
  g1732
  (
    n1836,
    n1130
  );


  buf
  g1733
  (
    n1734,
    n1125
  );


  buf
  g1734
  (
    n1646,
    n1415
  );


  buf
  g1735
  (
    n1848,
    n1155
  );


  buf
  g1736
  (
    n1815,
    n1128
  );


  buf
  g1737
  (
    n1822,
    n1543
  );


  buf
  g1738
  (
    n1671,
    n1448
  );


  not
  g1739
  (
    n1659,
    n1451
  );


  not
  g1740
  (
    n1747,
    n1511
  );


  buf
  g1741
  (
    n1673,
    n1395
  );


  buf
  g1742
  (
    n1745,
    n1375
  );


  not
  g1743
  (
    n1680,
    n1268
  );


  buf
  g1744
  (
    n1725,
    n1544
  );


  not
  g1745
  (
    n1844,
    n1155
  );


  buf
  g1746
  (
    n1771,
    n1534
  );


  nor
  g1747
  (
    n1682,
    n1145,
    n1452,
    n1480
  );


  nor
  g1748
  (
    n1813,
    n1432,
    n1494,
    n1434,
    n1437
  );


  xnor
  g1749
  (
    n1731,
    n1031,
    n1460,
    n1118,
    n1541
  );


  and
  g1750
  (
    n1735,
    n1514,
    n1155,
    n1501,
    n1373
  );


  xnor
  g1751
  (
    n1709,
    n1403,
    n1158,
    n1163,
    n1265
  );


  nand
  g1752
  (
    n1826,
    n1387,
    n1381,
    n1140,
    n1433
  );


  and
  g1753
  (
    n1637,
    n1507,
    n1493,
    n1439,
    n1401
  );


  and
  g1754
  (
    n1685,
    n1399,
    n1502,
    n1388,
    n1535
  );


  and
  g1755
  (
    n1758,
    n1263,
    n1449,
    n1126,
    n1386
  );


  nor
  g1756
  (
    n1647,
    n1459,
    n1118,
    n1360,
    n1142
  );


  nor
  g1757
  (
    KeyWire_0_1,
    n1152,
    n1530,
    n1404,
    n1129
  );


  nor
  g1758
  (
    n1800,
    n1455,
    n1127,
    n1120
  );


  and
  g1759
  (
    n1791,
    n1423,
    n1137,
    n1521,
    n1505
  );


  nor
  g1760
  (
    n1654,
    n1363,
    n1429,
    n1153,
    n1425
  );


  nand
  g1761
  (
    n1824,
    n1258,
    n1144,
    n1441,
    n1549
  );


  nor
  g1762
  (
    n1600,
    n1466,
    n1390,
    n1125,
    n1148
  );


  nor
  g1763
  (
    n1837,
    n1546,
    n1463,
    n1267,
    n1499
  );


  nor
  g1764
  (
    n1663,
    n1407,
    n1529,
    n1141,
    n1126
  );


  and
  g1765
  (
    n1801,
    n1478,
    n1422,
    n1158,
    n1149
  );


  and
  g1766
  (
    n1662,
    n1545,
    n1139,
    n1148,
    n1514
  );


  nor
  g1767
  (
    n1776,
    n1136,
    n1491,
    n1135,
    n1267
  );


  nor
  g1768
  (
    n1750,
    n1015,
    n1543,
    n1148,
    n1151
  );


  xnor
  g1769
  (
    n1841,
    n1156,
    n1268,
    n1125,
    n1522
  );


  nand
  g1770
  (
    n1831,
    n1152,
    n1124,
    n1369,
    n1402
  );


  xnor
  g1771
  (
    n1749,
    n1146,
    n1468,
    n1539,
    n1408
  );


  xnor
  g1772
  (
    n1838,
    n1413,
    n1483,
    n1127,
    n1522
  );


  xnor
  g1773
  (
    n1733,
    n1374,
    n1501,
    n1146,
    n1268
  );


  and
  g1774
  (
    n1599,
    n1411,
    n1503,
    n1532,
    n1257
  );


  nand
  g1775
  (
    n1803,
    n1549,
    n1266,
    n1511,
    n1117
  );


  xnor
  g1776
  (
    n1678,
    n1135,
    n1539,
    n1027,
    n1124
  );


  xor
  g1777
  (
    n1792,
    n1128,
    n1161,
    n1160,
    n1454
  );


  xor
  g1778
  (
    n1649,
    n1154,
    n1457,
    n1537,
    n1126
  );


  xnor
  g1779
  (
    n1675,
    n1162,
    n1426,
    n1159,
    n1528
  );


  or
  g1780
  (
    n1632,
    n1545,
    n1117,
    n1547,
    n1158
  );


  nand
  g1781
  (
    n1658,
    n1453,
    n1398,
    n1516,
    n1532
  );


  or
  g1782
  (
    n1854,
    n1158,
    n1024,
    n1133,
    n1500
  );


  xnor
  g1783
  (
    n1787,
    n1017,
    n1362,
    n1153,
    n1263
  );


  xor
  g1784
  (
    n1625,
    n1476,
    n1154,
    n1264,
    n1465
  );


  xor
  g1785
  (
    n1762,
    n1484,
    n1549,
    n1132,
    n1159
  );


  nand
  g1786
  (
    n1595,
    n1509,
    n1518,
    n1467,
    n1124
  );


  or
  g1787
  (
    n1780,
    n593,
    n1014,
    n1025,
    n1456
  );


  nor
  g1788
  (
    n1759,
    n1548,
    n1120,
    n1264,
    n1153
  );


  nand
  g1789
  (
    n1835,
    n1458,
    n1515,
    n1013,
    n1469
  );


  and
  g1790
  (
    n1626,
    n1020,
    n1141,
    n1477,
    n1118
  );


  xnor
  g1791
  (
    n1630,
    n1368,
    n1029,
    n1512,
    n1531
  );


  xnor
  g1792
  (
    n1798,
    n1367,
    n1132,
    n1545,
    n1140
  );


  nand
  g1793
  (
    n1772,
    n1266,
    n1257,
    n1536,
    n1410
  );


  xnor
  g1794
  (
    n1859,
    n1542,
    n1479,
    n1117,
    n1139
  );


  or
  g1795
  (
    n1655,
    n1133,
    n1492,
    n1417,
    n1524
  );


  and
  g1796
  (
    n1639,
    n1546,
    n1384,
    n1019,
    n1033
  );


  xnor
  g1797
  (
    n1833,
    n1475,
    n1268,
    n1138,
    n1541
  );


  xnor
  g1798
  (
    n1710,
    n1129,
    n1516,
    n1504,
    n1130
  );


  xnor
  g1799
  (
    n1795,
    n1414,
    n1364,
    n1162,
    n1512
  );


  xor
  g1800
  (
    KeyWire_0_16,
    n1161,
    n1519,
    n1122,
    n1118
  );


  xor
  g1801
  (
    n1702,
    n1536,
    n1123,
    n1125,
    n1538
  );


  xor
  g1802
  (
    n1711,
    n1490,
    n1472,
    n1421,
    n1123
  );


  xor
  g1803
  (
    n1849,
    n1412,
    n1520,
    n1507,
    n1154
  );


  xnor
  g1804
  (
    n1784,
    n1420,
    n1132,
    n1359,
    n1537
  );


  or
  g1805
  (
    n1809,
    n1149,
    n1258,
    n1123,
    n1257
  );


  xor
  g1806
  (
    n1850,
    n1163,
    n1471,
    n1546,
    n1142
  );


  or
  g1807
  (
    n1804,
    n1538,
    n1509,
    n1150
  );


  xnor
  g1808
  (
    n1611,
    n1132,
    n1163,
    n1548,
    n1370
  );


  xnor
  g1809
  (
    n1768,
    n1379,
    n1400,
    n1397,
    n1481
  );


  and
  g1810
  (
    n1641,
    n1544,
    n1122,
    n1541,
    n1445
  );


  xnor
  g1811
  (
    n1769,
    n1543,
    n1498,
    n1147,
    n1138
  );


  xnor
  g1812
  (
    n1593,
    n1130,
    n1419,
    n1139,
    n1391
  );


  nor
  g1813
  (
    n1612,
    n1143,
    n1446,
    n1488,
    n1138
  );


  or
  g1814
  (
    n1730,
    n1518,
    n1544,
    n1257,
    n1450
  );


  nand
  g1815
  (
    n1614,
    n1145,
    n1474,
    n1525,
    n1542
  );


  or
  g1816
  (
    n1695,
    n1143,
    n1026,
    n1133,
    n1161
  );


  nand
  g1817
  (
    n1660,
    n1264,
    n1539,
    n1148,
    n1508
  );


  xnor
  g1818
  (
    n1743,
    n1505,
    n1385,
    n1547,
    n1119
  );


  nand
  g1819
  (
    n1811,
    n1500,
    n1383,
    n1131,
    n1156
  );


  nor
  g1820
  (
    n1793,
    n1032,
    n1506,
    n1162,
    n1443
  );


  nand
  g1821
  (
    n1719,
    n1121,
    n1380,
    n1535,
    n1160
  );


  and
  g1822
  (
    n1779,
    n1164,
    n1150,
    n1124,
    n1527
  );


  nand
  g1823
  (
    n1766,
    n594,
    n1133,
    n1130,
    n1258
  );


  xor
  g1824
  (
    n1786,
    n1365,
    n1030,
    n1134,
    n1549
  );


  and
  g1825
  (
    n1856,
    n1513,
    n1126,
    n1520,
    n1146
  );


  xnor
  g1826
  (
    n1677,
    n1389,
    n1536,
    n1258,
    n594
  );


  nor
  g1827
  (
    n1846,
    n1497,
    n1508,
    n1546,
    n1156
  );


  xor
  g1828
  (
    n1708,
    n1134,
    n1131,
    n1141,
    n1527
  );


  nor
  g1829
  (
    n1681,
    n1117,
    n1265,
    n1127,
    n1137
  );


  xor
  g1830
  (
    n1934,
    n1696,
    n1553,
    n1783,
    n1571
  );


  xor
  g1831
  (
    n1958,
    n1353,
    n1570,
    n1636,
    n1807
  );


  nor
  g1832
  (
    n1867,
    n1625,
    n1643,
    n1588,
    n1558
  );


  nor
  g1833
  (
    n1897,
    n1688,
    n1782,
    n1565,
    n1358
  );


  and
  g1834
  (
    n1988,
    n1582,
    n1814,
    n1792,
    n1571
  );


  xnor
  g1835
  (
    n1953,
    n1701,
    n1621,
    n1853,
    n1638
  );


  nand
  g1836
  (
    n1937,
    n1580,
    n1606,
    n1756,
    n1347
  );


  nor
  g1837
  (
    n1914,
    n1042,
    n1349,
    n1711,
    n1572
  );


  nand
  g1838
  (
    n1903,
    n1553,
    n1558,
    n1713,
    n1641
  );


  xor
  g1839
  (
    n1881,
    n1345,
    n1589,
    n1786,
    n1582
  );


  xnor
  g1840
  (
    n1892,
    n1795,
    n1854,
    n1607,
    n1700
  );


  xor
  g1841
  (
    n1922,
    n1768,
    n1770,
    n1590,
    n1806
  );


  nor
  g1842
  (
    n1879,
    n1860,
    n1578,
    n1798,
    n1629
  );


  nor
  g1843
  (
    n1933,
    n1743,
    n1704,
    n1813,
    n1559
  );


  xnor
  g1844
  (
    n1886,
    n1594,
    n1345,
    n1829,
    n1824
  );


  nand
  g1845
  (
    n1906,
    n1679,
    n1618,
    n1586,
    n1851
  );


  and
  g1846
  (
    n1901,
    n1821,
    n1666,
    n1573,
    n1748
  );


  or
  g1847
  (
    n1912,
    n1772,
    n1758,
    n1352,
    n1619
  );


  nand
  g1848
  (
    n1951,
    n1550,
    n1751,
    n1562,
    n1569
  );


  xnor
  g1849
  (
    n1908,
    n1357,
    n1047,
    n1551,
    n1567
  );


  or
  g1850
  (
    n1938,
    n1582,
    n1586,
    n1348,
    n1574
  );


  nand
  g1851
  (
    n1925,
    n1555,
    n1587,
    n1797,
    n1830
  );


  or
  g1852
  (
    n1963,
    n1678,
    n1556,
    n1587,
    n1707
  );


  or
  g1853
  (
    n1913,
    n1579,
    n1767,
    n1581,
    n1759
  );


  nor
  g1854
  (
    n1907,
    n1708,
    n1551,
    n1835,
    n1753
  );


  xnor
  g1855
  (
    n1889,
    n1691,
    n1761,
    n1723,
    n1351
  );


  xor
  g1856
  (
    n1982,
    n1356,
    n1802,
    n1568,
    n1724
  );


  and
  g1857
  (
    n1987,
    n1844,
    n1794,
    n1584,
    n1664
  );


  xnor
  g1858
  (
    n1921,
    n1750,
    n1354,
    n1356,
    n1826
  );


  or
  g1859
  (
    n1874,
    n1601,
    n1557,
    n594,
    n1591
  );


  nand
  g1860
  (
    n1928,
    n1648,
    n1039,
    n1034,
    n1634
  );


  or
  g1861
  (
    n1919,
    n1357,
    n1551,
    n1580,
    n1552
  );


  xnor
  g1862
  (
    n1971,
    n1843,
    n1769,
    n1347,
    n1043
  );


  nor
  g1863
  (
    n1976,
    n1347,
    n1575,
    n1846,
    n1612
  );


  xnor
  g1864
  (
    n1936,
    n1694,
    n1561,
    n1659,
    n1693
  );


  nor
  g1865
  (
    n1966,
    n1728,
    n1576,
    n1584,
    n1702
  );


  nor
  g1866
  (
    n1872,
    n1726,
    n1668,
    n1567,
    n1583
  );


  and
  g1867
  (
    n1989,
    n1706,
    n1699,
    n1345,
    n1858
  );


  nand
  g1868
  (
    n1969,
    n1632,
    n1552,
    n1350,
    n1720
  );


  and
  g1869
  (
    n1948,
    n1599,
    n1838,
    n1589,
    n1732
  );


  xor
  g1870
  (
    n1876,
    n1849,
    n1604,
    n1808,
    n1555
  );


  xnor
  g1871
  (
    n1985,
    n1689,
    n1627,
    n1595,
    n1605
  );


  nor
  g1872
  (
    n1893,
    n1577,
    n1556,
    n1590,
    n1038
  );


  nor
  g1873
  (
    n1970,
    n1622,
    n1587,
    n1557,
    n1036
  );


  xnor
  g1874
  (
    n1972,
    n1351,
    n1040,
    n1785,
    n1573
  );


  xnor
  g1875
  (
    n1968,
    n1561,
    n1349,
    n1352,
    n1690
  );


  and
  g1876
  (
    n1931,
    n1581,
    n1817,
    n1347,
    n1661
  );


  nor
  g1877
  (
    n1870,
    n1593,
    n1739,
    n1353,
    n1575
  );


  and
  g1878
  (
    n1957,
    n1552,
    n1553,
    n1041,
    n1771
  );


  xor
  g1879
  (
    n1900,
    n1586,
    n1667,
    n1583,
    n1568
  );


  nor
  g1880
  (
    n1965,
    n1778,
    n1764,
    n1585,
    n1616
  );


  nor
  g1881
  (
    n1949,
    n1681,
    n1850,
    n1554,
    n1749
  );


  or
  g1882
  (
    n1871,
    n1788,
    n1358,
    n1714,
    n1855
  );


  nor
  g1883
  (
    n1909,
    n1579,
    n1355,
    n1351,
    n1755
  );


  xnor
  g1884
  (
    n1961,
    n1591,
    n1765,
    n1164,
    n1563
  );


  nand
  g1885
  (
    n1939,
    n1662,
    n1737,
    n1566,
    n1349
  );


  and
  g1886
  (
    n1896,
    n1719,
    n1572,
    n1839,
    n1776
  );


  nand
  g1887
  (
    n1910,
    n1774,
    n1804,
    n1669,
    n1356
  );


  or
  g1888
  (
    n1975,
    n1831,
    n1561,
    n1348,
    n1574
  );


  and
  g1889
  (
    n1944,
    n1550,
    n1845,
    n1346,
    n1567
  );


  xnor
  g1890
  (
    n1866,
    n1164,
    n1568,
    n1609,
    n1672
  );


  xnor
  g1891
  (
    n1895,
    n1712,
    n1583,
    n1563
  );


  and
  g1892
  (
    n1979,
    n1775,
    n1551,
    n1591,
    n1566
  );


  nor
  g1893
  (
    n1902,
    n1640,
    n1357,
    n1354,
    n1762
  );


  nand
  g1894
  (
    n1918,
    n1044,
    n1574,
    n1350,
    n1822
  );


  nand
  g1895
  (
    n1915,
    n1573,
    n1564,
    n1588,
    n1677
  );


  and
  g1896
  (
    n1920,
    n1574,
    n1570,
    n1705,
    n1742
  );


  xor
  g1897
  (
    n1983,
    n1709,
    n1703,
    n1348,
    n1833
  );


  nor
  g1898
  (
    n1865,
    n1611,
    n1684,
    n1576,
    n1564
  );


  and
  g1899
  (
    n1932,
    n1559,
    n1591,
    n1354,
    n1575
  );


  or
  g1900
  (
    n1887,
    n1576,
    n1746,
    n1583,
    n1578
  );


  nor
  g1901
  (
    n1898,
    n1654,
    n1856,
    n1560,
    n1572
  );


  xnor
  g1902
  (
    n1899,
    n1587,
    n1727,
    n1686,
    n1613
  );


  and
  g1903
  (
    n1990,
    n1562,
    n1645,
    n1358,
    n1581
  );


  xor
  g1904
  (
    n1880,
    n1784,
    n1692,
    n1675,
    n1862
  );


  and
  g1905
  (
    n1924,
    n1584,
    n1556,
    n1550,
    n1557
  );


  xor
  g1906
  (
    n1977,
    n1738,
    n1823,
    n1578,
    n1810
  );


  and
  g1907
  (
    n1927,
    n1564,
    n1576,
    n1584,
    n1631
  );


  and
  g1908
  (
    n1978,
    n1791,
    n1354,
    n1796,
    n1570
  );


  and
  g1909
  (
    n1904,
    n1716,
    n1592,
    n1585,
    n1803
  );


  xnor
  g1910
  (
    n1917,
    n1734,
    n1600,
    n1580,
    n1577
  );


  and
  g1911
  (
    n1878,
    n1801,
    n1680,
    n1671,
    n1790
  );


  and
  g1912
  (
    n1923,
    n1842,
    n1588,
    n1799,
    n1346
  );


  xor
  g1913
  (
    n1926,
    n1682,
    n1837,
    n1861,
    n1752
  );


  nor
  g1914
  (
    n1980,
    n1626,
    n1566,
    n1663,
    n1683
  );


  nand
  g1915
  (
    n1929,
    n1349,
    n1745,
    n1554,
    n1590
  );


  and
  g1916
  (
    n1888,
    n1560,
    n1565,
    n1685,
    n1623
  );


  nand
  g1917
  (
    n1905,
    n1588,
    n1670,
    n1565,
    n1655
  );


  or
  g1918
  (
    n1868,
    n1353,
    n1773,
    n1718,
    n1741
  );


  xnor
  g1919
  (
    n1950,
    n1346,
    n1565,
    n1562,
    n1351
  );


  xor
  g1920
  (
    n1941,
    n1614,
    n1589,
    n1780,
    n1649
  );


  and
  g1921
  (
    n1935,
    n1602,
    n1781,
    n1633,
    n1352
  );


  nor
  g1922
  (
    n1959,
    n1725,
    n1564,
    n1350,
    n1571
  );


  xor
  g1923
  (
    n1891,
    n1766,
    n1763,
    n1555,
    n1819
  );


  xor
  g1924
  (
    n1940,
    n1847,
    n1554,
    n1793,
    n1779
  );


  nor
  g1925
  (
    n1945,
    n1848,
    n1590,
    n1721,
    n1715
  );


  nor
  g1926
  (
    n1873,
    n1355,
    n1577,
    n1656,
    n1673
  );


  nand
  g1927
  (
    n1863,
    n1859,
    n1836,
    n1757,
    n1575
  );


  and
  g1928
  (
    n1885,
    n1580,
    n1740,
    n1566,
    n1550
  );


  and
  g1929
  (
    KeyWire_0_8,
    n1560,
    n1852,
    n1577,
    n1617
  );


  xor
  g1930
  (
    n1974,
    n1809,
    n1815,
    n1350,
    n1811
  );


  nor
  g1931
  (
    n1967,
    n1573,
    n1585,
    n1832,
    n1571
  );


  nand
  g1932
  (
    n1960,
    n1559,
    n1820,
    n1596,
    n1597
  );


  xnor
  g1933
  (
    n1946,
    n1559,
    n1658,
    n1754,
    n1642
  );


  xnor
  g1934
  (
    n1973,
    n1805,
    n1676,
    n1818,
    n1615
  );


  nor
  g1935
  (
    n1864,
    n1787,
    n1777,
    n1834,
    n1825
  );


  xor
  g1936
  (
    n1916,
    n1035,
    n1731,
    n1624,
    n1047
  );


  nor
  g1937
  (
    n1954,
    n1660,
    n1582,
    n1046,
    n1572
  );


  nand
  g1938
  (
    n1875,
    n1552,
    n1579,
    n1603,
    n1567
  );


  and
  g1939
  (
    n1882,
    n1717,
    n1562,
    n1828,
    n1665
  );


  or
  g1940
  (
    n1952,
    n1729,
    n1569,
    n1744,
    n1557
  );


  or
  g1941
  (
    n1883,
    n1355,
    n1747,
    n1553,
    n1598
  );


  nor
  g1942
  (
    n1981,
    n1789,
    n1352,
    n1346,
    n1644
  );


  xnor
  g1943
  (
    n1943,
    n1348,
    n1730,
    n1647,
    n1635
  );


  nand
  g1944
  (
    n1877,
    n1646,
    n1736,
    n1695,
    n1637
  );


  or
  g1945
  (
    n1962,
    n1650,
    n1356,
    n1556,
    n1037
  );


  nor
  g1946
  (
    n1890,
    n1840,
    n1586,
    n1841,
    n1651
  );


  xor
  g1947
  (
    n1894,
    n1561,
    n1674,
    n1563,
    n1687
  );


  xnor
  g1948
  (
    n1947,
    n1639,
    n1710,
    n1800,
    n1857
  );


  nand
  g1949
  (
    n1911,
    n1697,
    n1579,
    n1760,
    n1560
  );


  nand
  g1950
  (
    n1884,
    n1558,
    n1628,
    n1652,
    n1816
  );


  xor
  g1951
  (
    n1955,
    n1353,
    n1558,
    n1630,
    n1733
  );


  nor
  g1952
  (
    n1869,
    n1355,
    n1620,
    n1735,
    n1610
  );


  nand
  g1953
  (
    n1942,
    n1827,
    n1570,
    n1578,
    n1555
  );


  and
  g1954
  (
    n1986,
    n1698,
    n1657,
    n1589,
    n1608
  );


  nand
  g1955
  (
    n1964,
    n1653,
    n1358,
    n1569,
    n1812
  );


  and
  g1956
  (
    n1956,
    n1585,
    n1568,
    n1569,
    n1581
  );


  nand
  g1957
  (
    n1984,
    n1554,
    n1045,
    n1357,
    n1722
  );


  and
  g1958
  (
    n2007,
    n1880,
    n1922,
    n1885,
    n1952
  );


  nor
  g1959
  (
    n2009,
    n1863,
    n1927,
    n1987,
    n1982
  );


  xor
  g1960
  (
    n1999,
    n1873,
    n1884,
    n1970,
    n1864
  );


  nand
  g1961
  (
    n2008,
    n1871,
    n1954,
    n1946,
    n1938
  );


  nand
  g1962
  (
    n2017,
    n1915,
    n1974,
    n1920,
    n1900
  );


  nor
  g1963
  (
    n1996,
    n1909,
    n1950,
    n1988,
    n1957
  );


  xnor
  g1964
  (
    n2004,
    n1866,
    n1961,
    n1872,
    n1969
  );


  nand
  g1965
  (
    n2014,
    n1980,
    n1942,
    n1895,
    n1870
  );


  and
  g1966
  (
    n1993,
    n1965,
    n1892,
    n1935,
    n1887
  );


  xnor
  g1967
  (
    n2012,
    n1914,
    n1888,
    n1986,
    n1874
  );


  xnor
  g1968
  (
    n2016,
    n1877,
    n1929,
    n1931,
    n1905
  );


  xor
  g1969
  (
    n1991,
    n1985,
    n1930,
    n1959,
    n1875
  );


  xor
  g1970
  (
    n2019,
    n1923,
    n1926,
    n1968,
    n1912
  );


  xnor
  g1971
  (
    n1995,
    n1889,
    n1886,
    n1940,
    n1917
  );


  nor
  g1972
  (
    n1997,
    n1924,
    n1962,
    n1971,
    n1967
  );


  nand
  g1973
  (
    n2022,
    n1983,
    n1941,
    n1936,
    n1964
  );


  and
  g1974
  (
    n2021,
    n1893,
    n1984,
    n1911,
    n1953
  );


  nand
  g1975
  (
    n1994,
    n1896,
    n1975,
    n1960,
    n1868
  );


  xnor
  g1976
  (
    n2003,
    n1949,
    n1955,
    n1990,
    n1865
  );


  and
  g1977
  (
    n2013,
    n1972,
    n1944,
    n1881,
    n1907
  );


  xnor
  g1978
  (
    n2010,
    n1921,
    n1978,
    n1883,
    n1878
  );


  xor
  g1979
  (
    n2015,
    n1876,
    n1901,
    n1908,
    n1904
  );


  xor
  g1980
  (
    n1998,
    n1976,
    n1947,
    n1897,
    n1966
  );


  nand
  g1981
  (
    n2000,
    n1943,
    n1948,
    n1899,
    n1937
  );


  xnor
  g1982
  (
    n2005,
    n1903,
    n1891,
    n1989,
    n1934
  );


  xor
  g1983
  (
    n1992,
    n1906,
    n1918,
    n1902,
    n1933
  );


  and
  g1984
  (
    n2011,
    n1932,
    n1977,
    n1939,
    n1879
  );


  or
  g1985
  (
    n2002,
    n1898,
    n1869,
    n1919,
    n1979
  );


  and
  g1986
  (
    n2001,
    n1951,
    n1981,
    n1913,
    n1867
  );


  nor
  g1987
  (
    n2020,
    n1882,
    n1925,
    n1958,
    n1963
  );


  nand
  g1988
  (
    n2006,
    n1894,
    n1916,
    n1928,
    n1910
  );


  and
  g1989
  (
    n2018,
    n1890,
    n1973,
    n1945,
    n1956
  );


  nand
  g1990
  (
    n2027,
    n2019,
    n2016,
    n2017,
    n1996
  );


  xnor
  g1991
  (
    n2026,
    n1992,
    n2009,
    n1997,
    n1999
  );


  xor
  g1992
  (
    n2028,
    n1993,
    n2003,
    n2011,
    n2014
  );


  and
  g1993
  (
    n2024,
    n1994,
    n2004,
    n2010,
    n2015
  );


  xnor
  g1994
  (
    n2030,
    n1998,
    n2006,
    n2020,
    n2018
  );


  or
  g1995
  (
    n2023,
    n2008,
    n2005,
    n2021,
    n2002
  );


  xor
  g1996
  (
    n2025,
    n1991,
    n1995,
    n2000,
    n2001
  );


  xnor
  g1997
  (
    n2029,
    n2012,
    n2007,
    n2013,
    n2022
  );


  nand
  g1998
  (
    n2031,
    n2029,
    n2030,
    n2026,
    n2025
  );


  nand
  g1999
  (
    n2032,
    n2028,
    n2024,
    n2027,
    n2023
  );


  xnor
  KeyGate_0_0
  (
    n1000,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1808,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n373,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n560,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1107,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n829,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1086,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1346,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1930,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1349,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n645,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n390,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n495,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n664,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1011,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1193,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1783,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n510,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1475,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n1493,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1755,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1189,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n91,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n432,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n540,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1627,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1650,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n207,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1120,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n482,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1348,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n132,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

