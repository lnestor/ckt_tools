

module Stat_1363_31_10
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n45,
  n46,
  n47,
  n48,
  n1117,
  n1123,
  n1116,
  n1121,
  n1110,
  n1124,
  n1122,
  n1119,
  n1118,
  n1128,
  n1409,
  n1407,
  n1403,
  n1401,
  n1410,
  n1408,
  n1405,
  n1411,
  n1402,
  n1406,
  n1404,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63,
  keyIn_0_64,
  keyIn_0_65,
  keyIn_0_66,
  keyIn_0_67,
  keyIn_0_68,
  keyIn_0_69,
  keyIn_0_70,
  keyIn_0_71,
  keyIn_0_72,
  keyIn_0_73,
  keyIn_0_74,
  keyIn_0_75,
  keyIn_0_76,
  keyIn_0_77,
  keyIn_0_78,
  keyIn_0_79,
  keyIn_0_80,
  keyIn_0_81,
  keyIn_0_82,
  keyIn_0_83,
  keyIn_0_84,
  keyIn_0_85,
  keyIn_0_86,
  keyIn_0_87,
  keyIn_0_88,
  keyIn_0_89,
  keyIn_0_90,
  keyIn_0_91,
  keyIn_0_92,
  keyIn_0_93,
  keyIn_0_94,
  keyIn_0_95
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input n40;input n41;input n42;input n43;input n44;input n45;input n46;input n47;input n48;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;input keyIn_0_64;input keyIn_0_65;input keyIn_0_66;input keyIn_0_67;input keyIn_0_68;input keyIn_0_69;input keyIn_0_70;input keyIn_0_71;input keyIn_0_72;input keyIn_0_73;input keyIn_0_74;input keyIn_0_75;input keyIn_0_76;input keyIn_0_77;input keyIn_0_78;input keyIn_0_79;input keyIn_0_80;input keyIn_0_81;input keyIn_0_82;input keyIn_0_83;input keyIn_0_84;input keyIn_0_85;input keyIn_0_86;input keyIn_0_87;input keyIn_0_88;input keyIn_0_89;input keyIn_0_90;input keyIn_0_91;input keyIn_0_92;input keyIn_0_93;input keyIn_0_94;input keyIn_0_95;
  output n1117;output n1123;output n1116;output n1121;output n1110;output n1124;output n1122;output n1119;output n1118;output n1128;output n1409;output n1407;output n1403;output n1401;output n1410;output n1408;output n1405;output n1411;output n1402;output n1406;output n1404;
  wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1120;wire n1125;wire n1126;wire n1127;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire g_input_0_32;wire gbar_input_0_32;wire g_input_0_33;wire gbar_input_0_33;wire g_input_0_34;wire gbar_input_0_34;wire g_input_0_35;wire gbar_input_0_35;wire g_input_0_36;wire gbar_input_0_36;wire g_input_0_37;wire gbar_input_0_37;wire g_input_0_38;wire gbar_input_0_38;wire g_input_0_39;wire gbar_input_0_39;wire g_input_0_40;wire gbar_input_0_40;wire g_input_0_41;wire gbar_input_0_41;wire g_input_0_42;wire gbar_input_0_42;wire g_input_0_43;wire gbar_input_0_43;wire g_input_0_44;wire gbar_input_0_44;wire g_input_0_45;wire gbar_input_0_45;wire g_input_0_46;wire gbar_input_0_46;wire g_input_0_47;wire gbar_input_0_47;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n178,
    n3
  );


  buf
  g1
  (
    n58,
    n36
  );


  buf
  g2
  (
    n196,
    n24
  );


  buf
  g3
  (
    n208,
    n42
  );


  not
  g4
  (
    n189,
    n1
  );


  buf
  g5
  (
    n110,
    n4
  );


  not
  g6
  (
    n120,
    n10
  );


  buf
  g7
  (
    n215,
    n11
  );


  not
  g8
  (
    n154,
    n9
  );


  buf
  g9
  (
    n116,
    n36
  );


  not
  g10
  (
    n114,
    n28
  );


  not
  g11
  (
    n81,
    n24
  );


  not
  g12
  (
    n49,
    n37
  );


  buf
  g13
  (
    n216,
    n8
  );


  buf
  g14
  (
    n129,
    n16
  );


  not
  g15
  (
    n157,
    n21
  );


  not
  g16
  (
    n199,
    n5
  );


  not
  g17
  (
    n64,
    n41
  );


  not
  g18
  (
    n94,
    n28
  );


  buf
  g19
  (
    n193,
    n6
  );


  buf
  g20
  (
    n141,
    n10
  );


  buf
  g21
  (
    n174,
    n32
  );


  buf
  g22
  (
    n133,
    n33
  );


  buf
  g23
  (
    n186,
    n7
  );


  buf
  g24
  (
    n105,
    n18
  );


  buf
  g25
  (
    n102,
    n5
  );


  not
  g26
  (
    n77,
    n8
  );


  not
  g27
  (
    n175,
    n41
  );


  not
  g28
  (
    n52,
    n2
  );


  not
  g29
  (
    n185,
    n25
  );


  buf
  g30
  (
    n167,
    n7
  );


  not
  g31
  (
    n112,
    n23
  );


  not
  g32
  (
    n184,
    n15
  );


  buf
  g33
  (
    n214,
    n8
  );


  not
  g34
  (
    n176,
    n14
  );


  buf
  g35
  (
    n180,
    n26
  );


  buf
  g36
  (
    n88,
    n4
  );


  not
  g37
  (
    n137,
    n27
  );


  not
  g38
  (
    n128,
    n6
  );


  not
  g39
  (
    n104,
    n29
  );


  buf
  g40
  (
    n205,
    n31
  );


  buf
  g41
  (
    n50,
    n9
  );


  not
  g42
  (
    n73,
    n33
  );


  buf
  g43
  (
    n90,
    n29
  );


  not
  g44
  (
    n107,
    n30
  );


  buf
  g45
  (
    n111,
    n37
  );


  buf
  g46
  (
    n158,
    n17
  );


  buf
  g47
  (
    n192,
    n6
  );


  not
  g48
  (
    n132,
    n13
  );


  not
  g49
  (
    n86,
    n41
  );


  buf
  g50
  (
    n82,
    n26
  );


  not
  g51
  (
    n68,
    n17
  );


  buf
  g52
  (
    n163,
    n33
  );


  buf
  g53
  (
    n188,
    n23
  );


  not
  g54
  (
    n70,
    n13
  );


  not
  g55
  (
    n209,
    n29
  );


  buf
  g56
  (
    n206,
    n12
  );


  not
  g57
  (
    n170,
    n3
  );


  not
  g58
  (
    n63,
    n41
  );


  buf
  g59
  (
    n172,
    n24
  );


  not
  g60
  (
    n165,
    n35
  );


  buf
  g61
  (
    n67,
    n42
  );


  buf
  g62
  (
    n181,
    n13
  );


  not
  g63
  (
    n156,
    n7
  );


  buf
  g64
  (
    n54,
    n10
  );


  not
  g65
  (
    n144,
    n4
  );


  not
  g66
  (
    n62,
    n2
  );


  buf
  g67
  (
    n93,
    n15
  );


  buf
  g68
  (
    n169,
    n20
  );


  buf
  g69
  (
    n65,
    n25
  );


  not
  g70
  (
    n145,
    n42
  );


  buf
  g71
  (
    n113,
    n19
  );


  buf
  g72
  (
    n127,
    n40
  );


  not
  g73
  (
    n147,
    n23
  );


  buf
  g74
  (
    n194,
    n20
  );


  buf
  g75
  (
    n166,
    n10
  );


  buf
  g76
  (
    n213,
    n34
  );


  buf
  g77
  (
    n103,
    n28
  );


  not
  g78
  (
    n123,
    n9
  );


  buf
  g79
  (
    n210,
    n19
  );


  buf
  g80
  (
    n198,
    n29
  );


  not
  g81
  (
    n131,
    n22
  );


  buf
  g82
  (
    n142,
    n17
  );


  not
  g83
  (
    n191,
    n21
  );


  buf
  g84
  (
    n56,
    n22
  );


  buf
  g85
  (
    n152,
    n34
  );


  not
  g86
  (
    n177,
    n11
  );


  not
  g87
  (
    n97,
    n3
  );


  buf
  g88
  (
    n190,
    n28
  );


  buf
  g89
  (
    n161,
    n9
  );


  buf
  g90
  (
    n99,
    n38
  );


  buf
  g91
  (
    n117,
    n16
  );


  buf
  g92
  (
    n160,
    n42
  );


  not
  g93
  (
    n53,
    n30
  );


  not
  g94
  (
    n85,
    n18
  );


  not
  g95
  (
    n173,
    n35
  );


  buf
  g96
  (
    n101,
    n34
  );


  not
  g97
  (
    n149,
    n4
  );


  not
  g98
  (
    n168,
    n35
  );


  not
  g99
  (
    n211,
    n8
  );


  not
  g100
  (
    n98,
    n20
  );


  not
  g101
  (
    n138,
    n40
  );


  buf
  g102
  (
    n153,
    n27
  );


  buf
  g103
  (
    n202,
    n38
  );


  buf
  g104
  (
    n92,
    n12
  );


  buf
  g105
  (
    n79,
    n31
  );


  buf
  g106
  (
    n171,
    n32
  );


  not
  g107
  (
    n151,
    n14
  );


  not
  g108
  (
    n162,
    n31
  );


  not
  g109
  (
    n207,
    n21
  );


  buf
  g110
  (
    n96,
    n5
  );


  not
  g111
  (
    n115,
    n6
  );


  not
  g112
  (
    n84,
    n24
  );


  buf
  g113
  (
    n126,
    n26
  );


  not
  g114
  (
    n95,
    n40
  );


  not
  g115
  (
    n135,
    n30
  );


  buf
  g116
  (
    n71,
    n19
  );


  not
  g117
  (
    n91,
    n18
  );


  not
  g118
  (
    n197,
    n16
  );


  not
  g119
  (
    n183,
    n40
  );


  not
  g120
  (
    n89,
    n12
  );


  buf
  g121
  (
    n87,
    n2
  );


  buf
  g122
  (
    n136,
    n37
  );


  not
  g123
  (
    n143,
    n31
  );


  buf
  g124
  (
    n80,
    n39
  );


  buf
  g125
  (
    n130,
    n38
  );


  buf
  g126
  (
    n60,
    n15
  );


  not
  g127
  (
    n51,
    n27
  );


  not
  g128
  (
    n134,
    n32
  );


  not
  g129
  (
    n182,
    n32
  );


  not
  g130
  (
    n108,
    n15
  );


  not
  g131
  (
    n148,
    n27
  );


  buf
  g132
  (
    n203,
    n14
  );


  buf
  g133
  (
    n204,
    n25
  );


  buf
  g134
  (
    n75,
    n5
  );


  buf
  g135
  (
    n100,
    n21
  );


  buf
  g136
  (
    n187,
    n22
  );


  not
  g137
  (
    n72,
    n16
  );


  not
  g138
  (
    n146,
    n13
  );


  not
  g139
  (
    n109,
    n1
  );


  buf
  g140
  (
    n125,
    n38
  );


  not
  g141
  (
    n200,
    n1
  );


  not
  g142
  (
    n179,
    n3
  );


  not
  g143
  (
    n159,
    n36
  );


  not
  g144
  (
    n106,
    n11
  );


  not
  g145
  (
    n61,
    n20
  );


  not
  g146
  (
    n124,
    n17
  );


  not
  g147
  (
    n201,
    n26
  );


  not
  g148
  (
    n212,
    n36
  );


  not
  g149
  (
    n121,
    n35
  );


  buf
  g150
  (
    n83,
    n39
  );


  not
  g151
  (
    n155,
    n12
  );


  not
  g152
  (
    n66,
    n1
  );


  buf
  g153
  (
    n195,
    n33
  );


  not
  g154
  (
    n139,
    n14
  );


  buf
  g155
  (
    n164,
    n2
  );


  not
  g156
  (
    n55,
    n34
  );


  not
  g157
  (
    n78,
    n18
  );


  not
  g158
  (
    n57,
    n25
  );


  buf
  g159
  (
    n59,
    n11
  );


  buf
  g160
  (
    n150,
    n39
  );


  not
  g161
  (
    n74,
    n19
  );


  not
  g162
  (
    n76,
    n39
  );


  not
  g163
  (
    n118,
    n23
  );


  not
  g164
  (
    n140,
    n22
  );


  not
  g165
  (
    n119,
    n37
  );


  not
  g166
  (
    n69,
    n30
  );


  not
  g167
  (
    n122,
    n7
  );


  not
  g168
  (
    n653,
    n137
  );


  buf
  g169
  (
    n818,
    n125
  );


  buf
  g170
  (
    n353,
    n178
  );


  buf
  g171
  (
    n566,
    n150
  );


  buf
  g172
  (
    n227,
    n135
  );


  not
  g173
  (
    n218,
    n161
  );


  buf
  g174
  (
    n248,
    n115
  );


  not
  g175
  (
    n692,
    n131
  );


  buf
  g176
  (
    n501,
    n125
  );


  not
  g177
  (
    n698,
    n162
  );


  buf
  g178
  (
    n365,
    n69
  );


  not
  g179
  (
    n799,
    n115
  );


  not
  g180
  (
    n350,
    n79
  );


  buf
  g181
  (
    n622,
    n142
  );


  buf
  g182
  (
    n803,
    n88
  );


  not
  g183
  (
    n774,
    n143
  );


  buf
  g184
  (
    n487,
    n187
  );


  buf
  g185
  (
    n656,
    n112
  );


  buf
  g186
  (
    n759,
    n153
  );


  buf
  g187
  (
    n328,
    n167
  );


  not
  g188
  (
    n804,
    n191
  );


  not
  g189
  (
    n513,
    n137
  );


  not
  g190
  (
    n287,
    n163
  );


  not
  g191
  (
    n447,
    n112
  );


  not
  g192
  (
    n289,
    n124
  );


  buf
  g193
  (
    n363,
    n142
  );


  not
  g194
  (
    n712,
    n189
  );


  buf
  g195
  (
    n702,
    n192
  );


  buf
  g196
  (
    n628,
    n100
  );


  not
  g197
  (
    n836,
    n93
  );


  not
  g198
  (
    n709,
    n147
  );


  not
  g199
  (
    n681,
    n188
  );


  not
  g200
  (
    n730,
    n87
  );


  not
  g201
  (
    n242,
    n63
  );


  not
  g202
  (
    n834,
    n73
  );


  not
  g203
  (
    n543,
    n104
  );


  not
  g204
  (
    n255,
    n121
  );


  buf
  g205
  (
    n846,
    n91
  );


  not
  g206
  (
    n439,
    n59
  );


  buf
  g207
  (
    n641,
    n181
  );


  not
  g208
  (
    n294,
    n191
  );


  buf
  g209
  (
    n415,
    n84
  );


  not
  g210
  (
    n408,
    n112
  );


  not
  g211
  (
    n547,
    n115
  );


  not
  g212
  (
    n637,
    n151
  );


  not
  g213
  (
    n824,
    n68
  );


  not
  g214
  (
    n463,
    n169
  );


  buf
  g215
  (
    n417,
    n170
  );


  buf
  g216
  (
    n428,
    n85
  );


  not
  g217
  (
    n288,
    n128
  );


  buf
  g218
  (
    n636,
    n64
  );


  not
  g219
  (
    n310,
    n55
  );


  not
  g220
  (
    n564,
    n145
  );


  not
  g221
  (
    n259,
    n202
  );


  not
  g222
  (
    n714,
    n50
  );


  not
  g223
  (
    n745,
    n175
  );


  buf
  g224
  (
    n652,
    n188
  );


  not
  g225
  (
    n555,
    n65
  );


  not
  g226
  (
    n472,
    n101
  );


  not
  g227
  (
    n507,
    n175
  );


  not
  g228
  (
    n768,
    n152
  );


  buf
  g229
  (
    n512,
    n133
  );


  not
  g230
  (
    n706,
    n132
  );


  buf
  g231
  (
    n783,
    n148
  );


  buf
  g232
  (
    n696,
    n75
  );


  not
  g233
  (
    n635,
    n204
  );


  not
  g234
  (
    n378,
    n112
  );


  buf
  g235
  (
    n701,
    n66
  );


  buf
  g236
  (
    n356,
    n49
  );


  not
  g237
  (
    n568,
    n55
  );


  not
  g238
  (
    n320,
    n120
  );


  not
  g239
  (
    n838,
    n205
  );


  not
  g240
  (
    n506,
    n104
  );


  buf
  g241
  (
    n740,
    n127
  );


  not
  g242
  (
    n282,
    n127
  );


  not
  g243
  (
    n674,
    n66
  );


  buf
  g244
  (
    n737,
    n113
  );


  buf
  g245
  (
    n226,
    n127
  );


  not
  g246
  (
    n843,
    n158
  );


  buf
  g247
  (
    n492,
    n100
  );


  not
  g248
  (
    n615,
    n92
  );


  buf
  g249
  (
    n784,
    n106
  );


  buf
  g250
  (
    n708,
    n180
  );


  buf
  g251
  (
    n241,
    n160
  );


  buf
  g252
  (
    n497,
    n85
  );


  not
  g253
  (
    n291,
    n100
  );


  buf
  g254
  (
    n546,
    n70
  );


  buf
  g255
  (
    n277,
    n182
  );


  not
  g256
  (
    n519,
    n173
  );


  buf
  g257
  (
    n584,
    n113
  );


  not
  g258
  (
    n822,
    n76
  );


  buf
  g259
  (
    n461,
    n111
  );


  buf
  g260
  (
    n411,
    n132
  );


  buf
  g261
  (
    n613,
    n143
  );


  buf
  g262
  (
    n420,
    n86
  );


  buf
  g263
  (
    n359,
    n79
  );


  buf
  g264
  (
    n658,
    n150
  );


  buf
  g265
  (
    n526,
    n108
  );


  buf
  g266
  (
    n751,
    n168
  );


  buf
  g267
  (
    n357,
    n117
  );


  buf
  g268
  (
    n471,
    n49
  );


  buf
  g269
  (
    n811,
    n123
  );


  not
  g270
  (
    n223,
    n180
  );


  buf
  g271
  (
    n764,
    n76
  );


  not
  g272
  (
    n738,
    n197
  );


  not
  g273
  (
    n433,
    n207
  );


  buf
  g274
  (
    n625,
    n124
  );


  buf
  g275
  (
    n258,
    n155
  );


  buf
  g276
  (
    n781,
    n152
  );


  not
  g277
  (
    n264,
    n83
  );


  not
  g278
  (
    n581,
    n169
  );


  not
  g279
  (
    n779,
    n190
  );


  not
  g280
  (
    n565,
    n109
  );


  not
  g281
  (
    n302,
    n147
  );


  not
  g282
  (
    n343,
    n199
  );


  not
  g283
  (
    n261,
    n188
  );


  not
  g284
  (
    n377,
    n164
  );


  buf
  g285
  (
    n413,
    n107
  );


  buf
  g286
  (
    n587,
    n206
  );


  not
  g287
  (
    n435,
    n92
  );


  buf
  g288
  (
    n247,
    n147
  );


  buf
  g289
  (
    n621,
    n140
  );


  buf
  g290
  (
    n796,
    n126
  );


  not
  g291
  (
    n484,
    n137
  );


  not
  g292
  (
    n713,
    n190
  );


  not
  g293
  (
    n347,
    n80
  );


  not
  g294
  (
    n369,
    n165
  );


  buf
  g295
  (
    n711,
    n150
  );


  buf
  g296
  (
    n485,
    n110
  );


  buf
  g297
  (
    n829,
    n72
  );


  not
  g298
  (
    n772,
    n122
  );


  not
  g299
  (
    n493,
    n58
  );


  buf
  g300
  (
    n807,
    n128
  );


  not
  g301
  (
    n296,
    n188
  );


  not
  g302
  (
    n518,
    n173
  );


  buf
  g303
  (
    n601,
    n60
  );


  not
  g304
  (
    n585,
    n171
  );


  buf
  g305
  (
    n429,
    n183
  );


  buf
  g306
  (
    n573,
    n161
  );


  not
  g307
  (
    n780,
    n174
  );


  buf
  g308
  (
    n797,
    n164
  );


  not
  g309
  (
    n747,
    n50
  );


  not
  g310
  (
    n726,
    n96
  );


  not
  g311
  (
    n577,
    n49
  );


  buf
  g312
  (
    n321,
    n62
  );


  buf
  g313
  (
    n578,
    n126
  );


  buf
  g314
  (
    n776,
    n88
  );


  buf
  g315
  (
    n399,
    n72
  );


  buf
  g316
  (
    n785,
    n189
  );


  not
  g317
  (
    n693,
    n129
  );


  buf
  g318
  (
    n596,
    n82
  );


  buf
  g319
  (
    n643,
    n160
  );


  buf
  g320
  (
    n603,
    n67
  );


  buf
  g321
  (
    n375,
    n156
  );


  not
  g322
  (
    n449,
    n167
  );


  buf
  g323
  (
    n600,
    n176
  );


  not
  g324
  (
    n389,
    n96
  );


  not
  g325
  (
    n539,
    n114
  );


  not
  g326
  (
    n246,
    n73
  );


  buf
  g327
  (
    n267,
    n119
  );


  buf
  g328
  (
    n406,
    n56
  );


  buf
  g329
  (
    n346,
    n78
  );


  buf
  g330
  (
    n669,
    n133
  );


  not
  g331
  (
    n753,
    n63
  );


  buf
  g332
  (
    n544,
    n76
  );


  not
  g333
  (
    n503,
    n98
  );


  buf
  g334
  (
    n739,
    n179
  );


  buf
  g335
  (
    n680,
    n197
  );


  buf
  g336
  (
    n474,
    n85
  );


  buf
  g337
  (
    n450,
    n79
  );


  buf
  g338
  (
    n252,
    n157
  );


  buf
  g339
  (
    n763,
    n98
  );


  not
  g340
  (
    n383,
    n133
  );


  buf
  g341
  (
    n397,
    n138
  );


  buf
  g342
  (
    n524,
    n96
  );


  buf
  g343
  (
    n612,
    n107
  );


  buf
  g344
  (
    n238,
    n197
  );


  buf
  g345
  (
    n283,
    n168
  );


  buf
  g346
  (
    n367,
    n142
  );


  buf
  g347
  (
    n823,
    n158
  );


  not
  g348
  (
    n298,
    n153
  );


  not
  g349
  (
    n672,
    n194
  );


  not
  g350
  (
    n315,
    n152
  );


  not
  g351
  (
    n541,
    n151
  );


  buf
  g352
  (
    n480,
    n174
  );


  not
  g353
  (
    n830,
    n102
  );


  buf
  g354
  (
    n390,
    n165
  );


  not
  g355
  (
    n814,
    n85
  );


  not
  g356
  (
    n683,
    n72
  );


  not
  g357
  (
    n793,
    n93
  );


  buf
  g358
  (
    n662,
    n87
  );


  buf
  g359
  (
    n618,
    n67
  );


  not
  g360
  (
    n736,
    n80
  );


  not
  g361
  (
    n454,
    n199
  );


  buf
  g362
  (
    n704,
    n154
  );


  not
  g363
  (
    n778,
    n68
  );


  buf
  g364
  (
    n404,
    n191
  );


  not
  g365
  (
    n278,
    n65
  );


  not
  g366
  (
    n393,
    n91
  );


  not
  g367
  (
    n733,
    n167
  );


  not
  g368
  (
    n514,
    n196
  );


  buf
  g369
  (
    n465,
    n132
  );


  not
  g370
  (
    n611,
    n157
  );


  not
  g371
  (
    n540,
    n54
  );


  not
  g372
  (
    n767,
    n139
  );


  buf
  g373
  (
    n219,
    n68
  );


  buf
  g374
  (
    n322,
    n156
  );


  not
  g375
  (
    n668,
    n132
  );


  buf
  g376
  (
    n409,
    n125
  );


  not
  g377
  (
    n243,
    n149
  );


  not
  g378
  (
    n607,
    n175
  );


  buf
  g379
  (
    n624,
    n121
  );


  buf
  g380
  (
    n281,
    n190
  );


  buf
  g381
  (
    n634,
    n131
  );


  not
  g382
  (
    n629,
    n53
  );


  not
  g383
  (
    n679,
    n166
  );


  not
  g384
  (
    n372,
    n51
  );


  buf
  g385
  (
    n262,
    n93
  );


  buf
  g386
  (
    n617,
    n69
  );


  buf
  g387
  (
    n231,
    n179
  );


  buf
  g388
  (
    n609,
    n141
  );


  buf
  g389
  (
    n269,
    n69
  );


  not
  g390
  (
    n334,
    n113
  );


  buf
  g391
  (
    n639,
    n151
  );


  not
  g392
  (
    n667,
    n199
  );


  not
  g393
  (
    n659,
    n198
  );


  not
  g394
  (
    n791,
    n111
  );


  not
  g395
  (
    n813,
    n129
  );


  not
  g396
  (
    n542,
    n110
  );


  buf
  g397
  (
    n309,
    n90
  );


  buf
  g398
  (
    n305,
    n162
  );


  not
  g399
  (
    n469,
    n166
  );


  buf
  g400
  (
    n695,
    n206
  );


  not
  g401
  (
    n268,
    n193
  );


  not
  g402
  (
    n563,
    n78
  );


  buf
  g403
  (
    n230,
    n59
  );


  buf
  g404
  (
    n689,
    n198
  );


  not
  g405
  (
    n478,
    n121
  );


  not
  g406
  (
    n479,
    n185
  );


  not
  g407
  (
    n810,
    n144
  );


  buf
  g408
  (
    n462,
    n52
  );


  not
  g409
  (
    n286,
    n195
  );


  buf
  g410
  (
    n528,
    n77
  );


  buf
  g411
  (
    n339,
    n155
  );


  buf
  g412
  (
    n762,
    n164
  );


  not
  g413
  (
    n582,
    n56
  );


  buf
  g414
  (
    n551,
    n116
  );


  not
  g415
  (
    n424,
    n56
  );


  not
  g416
  (
    n645,
    n205
  );


  buf
  g417
  (
    n646,
    n148
  );


  not
  g418
  (
    n591,
    n115
  );


  not
  g419
  (
    n398,
    n58
  );


  buf
  g420
  (
    n414,
    n200
  );


  not
  g421
  (
    n719,
    n136
  );


  not
  g422
  (
    n240,
    n134
  );


  buf
  g423
  (
    n533,
    n189
  );


  buf
  g424
  (
    n847,
    n99
  );


  buf
  g425
  (
    n827,
    n67
  );


  buf
  g426
  (
    n604,
    n172
  );


  not
  g427
  (
    n486,
    n190
  );


  not
  g428
  (
    n279,
    n136
  );


  buf
  g429
  (
    n387,
    n106
  );


  not
  g430
  (
    n438,
    n52
  );


  not
  g431
  (
    n351,
    n140
  );


  buf
  g432
  (
    n718,
    n95
  );


  buf
  g433
  (
    n532,
    n203
  );


  not
  g434
  (
    n329,
    n207
  );


  buf
  g435
  (
    n537,
    n146
  );


  not
  g436
  (
    n456,
    n70
  );


  buf
  g437
  (
    n556,
    n160
  );


  buf
  g438
  (
    n312,
    n50
  );


  buf
  g439
  (
    n703,
    n186
  );


  buf
  g440
  (
    n395,
    n170
  );


  buf
  g441
  (
    n481,
    n87
  );


  buf
  g442
  (
    n815,
    n80
  );


  not
  g443
  (
    n729,
    n77
  );


  buf
  g444
  (
    n642,
    n51
  );


  not
  g445
  (
    n446,
    n89
  );


  not
  g446
  (
    n835,
    n121
  );


  buf
  g447
  (
    n598,
    n59
  );


  not
  g448
  (
    n427,
    n74
  );


  not
  g449
  (
    n345,
    n183
  );


  not
  g450
  (
    n444,
    n184
  );


  not
  g451
  (
    n661,
    n172
  );


  not
  g452
  (
    n274,
    n177
  );


  buf
  g453
  (
    n304,
    n136
  );


  not
  g454
  (
    n549,
    n158
  );


  buf
  g455
  (
    n579,
    n150
  );


  not
  g456
  (
    n798,
    n134
  );


  not
  g457
  (
    n314,
    n111
  );


  not
  g458
  (
    n839,
    n106
  );


  buf
  g459
  (
    n782,
    n145
  );


  buf
  g460
  (
    n690,
    n154
  );


  not
  g461
  (
    n233,
    n128
  );


  buf
  g462
  (
    n300,
    n157
  );


  not
  g463
  (
    n496,
    n80
  );


  buf
  g464
  (
    n225,
    n141
  );


  not
  g465
  (
    n816,
    n145
  );


  buf
  g466
  (
    n728,
    n60
  );


  not
  g467
  (
    n741,
    n193
  );


  buf
  g468
  (
    n786,
    n181
  );


  not
  g469
  (
    n384,
    n99
  );


  buf
  g470
  (
    n284,
    n56
  );


  not
  g471
  (
    n498,
    n167
  );


  buf
  g472
  (
    n236,
    n202
  );


  buf
  g473
  (
    n545,
    n77
  );


  not
  g474
  (
    n657,
    n194
  );


  not
  g475
  (
    n337,
    n94
  );


  not
  g476
  (
    n280,
    n185
  );


  not
  g477
  (
    n371,
    n53
  );


  not
  g478
  (
    n531,
    n65
  );


  buf
  g479
  (
    n677,
    n105
  );


  not
  g480
  (
    n760,
    n170
  );


  buf
  g481
  (
    n648,
    n164
  );


  buf
  g482
  (
    n234,
    n181
  );


  not
  g483
  (
    n841,
    n141
  );


  buf
  g484
  (
    n299,
    n71
  );


  buf
  g485
  (
    n732,
    n81
  );


  buf
  g486
  (
    n473,
    n72
  );


  not
  g487
  (
    n735,
    n124
  );


  not
  g488
  (
    n567,
    n171
  );


  buf
  g489
  (
    n686,
    n101
  );


  not
  g490
  (
    n228,
    n182
  );


  buf
  g491
  (
    n673,
    n61
  );


  not
  g492
  (
    n602,
    n146
  );


  not
  g493
  (
    n301,
    n109
  );


  not
  g494
  (
    n335,
    n95
  );


  not
  g495
  (
    n499,
    n86
  );


  not
  g496
  (
    n491,
    n178
  );


  buf
  g497
  (
    n220,
    n110
  );


  not
  g498
  (
    n405,
    n204
  );


  not
  g499
  (
    n520,
    n136
  );


  buf
  g500
  (
    n434,
    n103
  );


  not
  g501
  (
    n442,
    n198
  );


  not
  g502
  (
    n569,
    n203
  );


  not
  g503
  (
    n421,
    n103
  );


  not
  g504
  (
    n235,
    n75
  );


  not
  g505
  (
    n694,
    n159
  );


  buf
  g506
  (
    n316,
    n172
  );


  not
  g507
  (
    n410,
    n144
  );


  buf
  g508
  (
    n344,
    n113
  );


  buf
  g509
  (
    n597,
    n71
  );


  not
  g510
  (
    n794,
    n192
  );


  buf
  g511
  (
    n515,
    n91
  );


  buf
  g512
  (
    n401,
    n195
  );


  not
  g513
  (
    n251,
    n123
  );


  buf
  g514
  (
    n423,
    n105
  );


  not
  g515
  (
    n826,
    n97
  );


  buf
  g516
  (
    n580,
    n123
  );


  not
  g517
  (
    n670,
    n159
  );


  buf
  g518
  (
    n821,
    n169
  );


  buf
  g519
  (
    n691,
    n205
  );


  buf
  g520
  (
    n654,
    n120
  );


  not
  g521
  (
    n403,
    n96
  );


  not
  g522
  (
    n361,
    n57
  );


  buf
  g523
  (
    n490,
    n74
  );


  buf
  g524
  (
    n769,
    n129
  );


  buf
  g525
  (
    n483,
    n148
  );


  buf
  g526
  (
    n400,
    n60
  );


  not
  g527
  (
    n808,
    n205
  );


  not
  g528
  (
    n529,
    n90
  );


  buf
  g529
  (
    n755,
    n98
  );


  not
  g530
  (
    n336,
    n82
  );


  not
  g531
  (
    n527,
    n183
  );


  not
  g532
  (
    n502,
    n201
  );


  buf
  g533
  (
    n592,
    n62
  );


  not
  g534
  (
    n352,
    n51
  );


  not
  g535
  (
    n276,
    n97
  );


  not
  g536
  (
    n575,
    n75
  );


  not
  g537
  (
    n459,
    n54
  );


  not
  g538
  (
    n599,
    n57
  );


  buf
  g539
  (
    n222,
    n53
  );


  buf
  g540
  (
    n663,
    n147
  );


  buf
  g541
  (
    n746,
    n177
  );


  not
  g542
  (
    n576,
    n58
  );


  buf
  g543
  (
    n530,
    n71
  );


  not
  g544
  (
    n623,
    n81
  );


  buf
  g545
  (
    n265,
    n61
  );


  buf
  g546
  (
    n303,
    n171
  );


  not
  g547
  (
    n716,
    n186
  );


  not
  g548
  (
    n705,
    n101
  );


  buf
  g549
  (
    n844,
    n143
  );


  buf
  g550
  (
    n470,
    n123
  );


  not
  g551
  (
    n426,
    n66
  );


  buf
  g552
  (
    n809,
    n182
  );


  not
  g553
  (
    n761,
    n166
  );


  not
  g554
  (
    n536,
    n117
  );


  buf
  g555
  (
    n293,
    n204
  );


  buf
  g556
  (
    n270,
    n187
  );


  buf
  g557
  (
    n789,
    n81
  );


  not
  g558
  (
    n458,
    n139
  );


  not
  g559
  (
    n550,
    n206
  );


  not
  g560
  (
    n752,
    n84
  );


  buf
  g561
  (
    n845,
    n161
  );


  buf
  g562
  (
    n440,
    n163
  );


  not
  g563
  (
    n717,
    n77
  );


  buf
  g564
  (
    n848,
    n78
  );


  buf
  g565
  (
    n317,
    n53
  );


  not
  g566
  (
    n833,
    n145
  );


  buf
  g567
  (
    n297,
    n92
  );


  buf
  g568
  (
    n432,
    n153
  );


  buf
  g569
  (
    n430,
    n65
  );


  buf
  g570
  (
    n385,
    n161
  );


  not
  g571
  (
    n700,
    n75
  );


  buf
  g572
  (
    n237,
    n49
  );


  not
  g573
  (
    n801,
    n149
  );


  buf
  g574
  (
    n720,
    n88
  );


  buf
  g575
  (
    n460,
    n122
  );


  buf
  g576
  (
    n381,
    n120
  );


  buf
  g577
  (
    n368,
    n54
  );


  buf
  g578
  (
    n306,
    n142
  );


  buf
  g579
  (
    n311,
    n197
  );


  not
  g580
  (
    n684,
    n172
  );


  buf
  g581
  (
    n805,
    n187
  );


  not
  g582
  (
    n825,
    n144
  );


  buf
  g583
  (
    n562,
    n169
  );


  buf
  g584
  (
    n790,
    n138
  );


  not
  g585
  (
    n224,
    n168
  );


  not
  g586
  (
    n425,
    n162
  );


  buf
  g587
  (
    n715,
    n81
  );


  not
  g588
  (
    n254,
    n203
  );


  buf
  g589
  (
    n849,
    n98
  );


  buf
  g590
  (
    n295,
    n195
  );


  not
  g591
  (
    n837,
    n187
  );


  not
  g592
  (
    n245,
    n126
  );


  not
  g593
  (
    n391,
    n97
  );


  not
  g594
  (
    n676,
    n183
  );


  buf
  g595
  (
    n457,
    n118
  );


  buf
  g596
  (
    n374,
    n66
  );


  buf
  g597
  (
    n558,
    n107
  );


  not
  g598
  (
    n724,
    n202
  );


  buf
  g599
  (
    n557,
    n178
  );


  buf
  g600
  (
    n734,
    n156
  );


  not
  g601
  (
    n710,
    n149
  );


  not
  g602
  (
    n272,
    n110
  );


  not
  g603
  (
    n475,
    n69
  );


  not
  g604
  (
    n436,
    n195
  );


  buf
  g605
  (
    n742,
    n107
  );


  buf
  g606
  (
    n770,
    n86
  );


  not
  g607
  (
    n342,
    n118
  );


  buf
  g608
  (
    n614,
    n73
  );


  not
  g609
  (
    n416,
    n117
  );


  buf
  g610
  (
    n412,
    n76
  );


  buf
  g611
  (
    n232,
    n109
  );


  not
  g612
  (
    n758,
    n191
  );


  buf
  g613
  (
    n806,
    n63
  );


  not
  g614
  (
    n535,
    n60
  );


  not
  g615
  (
    n504,
    n201
  );


  not
  g616
  (
    n360,
    n61
  );


  buf
  g617
  (
    n553,
    n83
  );


  buf
  g618
  (
    n508,
    n138
  );


  buf
  g619
  (
    n370,
    n116
  );


  not
  g620
  (
    n419,
    n189
  );


  not
  g621
  (
    n627,
    n200
  );


  buf
  g622
  (
    n616,
    n61
  );


  not
  g623
  (
    n330,
    n87
  );


  not
  g624
  (
    n355,
    n119
  );


  not
  g625
  (
    n650,
    n140
  );


  not
  g626
  (
    n548,
    n159
  );


  not
  g627
  (
    n257,
    n184
  );


  not
  g628
  (
    n271,
    n70
  );


  buf
  g629
  (
    n748,
    n71
  );


  buf
  g630
  (
    n773,
    n184
  );


  buf
  g631
  (
    n244,
    n95
  );


  buf
  g632
  (
    n586,
    n109
  );


  buf
  g633
  (
    n757,
    n86
  );


  buf
  g634
  (
    n831,
    n163
  );


  buf
  g635
  (
    n338,
    n67
  );


  buf
  g636
  (
    n756,
    n204
  );


  not
  g637
  (
    n638,
    n151
  );


  buf
  g638
  (
    n510,
    n58
  );


  buf
  g639
  (
    n445,
    n54
  );


  not
  g640
  (
    n290,
    n83
  );


  buf
  g641
  (
    n500,
    n193
  );


  buf
  g642
  (
    n792,
    n84
  );


  buf
  g643
  (
    n422,
    n198
  );


  not
  g644
  (
    n840,
    n180
  );


  buf
  g645
  (
    n340,
    n146
  );


  buf
  g646
  (
    n448,
    n68
  );


  not
  g647
  (
    n590,
    n70
  );


  buf
  g648
  (
    n464,
    n130
  );


  not
  g649
  (
    n788,
    n148
  );


  not
  g650
  (
    n812,
    n138
  );


  not
  g651
  (
    n678,
    n114
  );


  buf
  g652
  (
    n358,
    n128
  );


  buf
  g653
  (
    n509,
    n55
  );


  not
  g654
  (
    n292,
    n108
  );


  not
  g655
  (
    n800,
    n141
  );


  buf
  g656
  (
    n256,
    n120
  );


  buf
  g657
  (
    n707,
    n158
  );


  not
  g658
  (
    n561,
    n51
  );


  not
  g659
  (
    n610,
    n135
  );


  not
  g660
  (
    n386,
    n114
  );


  not
  g661
  (
    n229,
    n140
  );


  not
  g662
  (
    n402,
    n201
  );


  buf
  g663
  (
    n495,
    n186
  );


  buf
  g664
  (
    n766,
    n144
  );


  not
  g665
  (
    n828,
    n192
  );


  not
  g666
  (
    n333,
    n74
  );


  buf
  g667
  (
    n332,
    n64
  );


  buf
  g668
  (
    n494,
    n152
  );


  not
  g669
  (
    n249,
    n101
  );


  buf
  g670
  (
    n593,
    n196
  );


  buf
  g671
  (
    n572,
    n179
  );


  not
  g672
  (
    n687,
    n180
  );


  not
  g673
  (
    n559,
    n55
  );


  buf
  g674
  (
    n407,
    n117
  );


  not
  g675
  (
    n731,
    n63
  );


  not
  g676
  (
    n647,
    n94
  );


  buf
  g677
  (
    n534,
    n124
  );


  not
  g678
  (
    n795,
    n57
  );


  buf
  g679
  (
    n285,
    n134
  );


  buf
  g680
  (
    n476,
    n82
  );


  buf
  g681
  (
    n632,
    n173
  );


  not
  g682
  (
    n606,
    n83
  );


  buf
  g683
  (
    n787,
    n199
  );


  buf
  g684
  (
    n671,
    n116
  );


  not
  g685
  (
    n522,
    n130
  );


  not
  g686
  (
    n665,
    n182
  );


  buf
  g687
  (
    n313,
    n89
  );


  not
  g688
  (
    n777,
    n73
  );


  not
  g689
  (
    n376,
    n122
  );


  not
  g690
  (
    n239,
    n177
  );


  buf
  g691
  (
    n323,
    n139
  );


  not
  g692
  (
    n832,
    n106
  );


  buf
  g693
  (
    n666,
    n157
  );


  buf
  g694
  (
    n554,
    n59
  );


  buf
  g695
  (
    n331,
    n185
  );


  not
  g696
  (
    n688,
    n118
  );


  buf
  g697
  (
    n754,
    n57
  );


  not
  g698
  (
    n324,
    n166
  );


  not
  g699
  (
    n517,
    n79
  );


  buf
  g700
  (
    n588,
    n52
  );


  buf
  g701
  (
    n660,
    n155
  );


  not
  g702
  (
    n675,
    n91
  );


  buf
  g703
  (
    n725,
    n181
  );


  buf
  g704
  (
    n488,
    n194
  );


  not
  g705
  (
    n468,
    n165
  );


  not
  g706
  (
    n620,
    n162
  );


  not
  g707
  (
    n765,
    n122
  );


  not
  g708
  (
    n221,
    n108
  );


  buf
  g709
  (
    n341,
    n130
  );


  buf
  g710
  (
    n307,
    n89
  );


  not
  g711
  (
    n354,
    n94
  );


  not
  g712
  (
    n589,
    n116
  );


  not
  g713
  (
    n552,
    n88
  );


  not
  g714
  (
    n366,
    n108
  );


  not
  g715
  (
    n452,
    n50
  );


  buf
  g716
  (
    n364,
    n104
  );


  buf
  g717
  (
    n253,
    n90
  );


  buf
  g718
  (
    n505,
    n103
  );


  buf
  g719
  (
    n318,
    n129
  );


  not
  g720
  (
    n743,
    n104
  );


  buf
  g721
  (
    n727,
    n168
  );


  not
  g722
  (
    n392,
    n105
  );


  buf
  g723
  (
    n583,
    n163
  );


  not
  g724
  (
    n273,
    n103
  );


  not
  g725
  (
    n850,
    n93
  );


  not
  g726
  (
    n349,
    n178
  );


  buf
  g727
  (
    n651,
    n194
  );


  buf
  g728
  (
    n373,
    n64
  );


  not
  g729
  (
    n466,
    n89
  );


  buf
  g730
  (
    n560,
    n102
  );


  not
  g731
  (
    n451,
    n196
  );


  not
  g732
  (
    n489,
    n170
  );


  buf
  g733
  (
    n266,
    n175
  );


  buf
  g734
  (
    n594,
    n137
  );


  buf
  g735
  (
    n263,
    n185
  );


  buf
  g736
  (
    n388,
    n90
  );


  not
  g737
  (
    n699,
    n154
  );


  buf
  g738
  (
    n467,
    n62
  );


  not
  g739
  (
    n644,
    n97
  );


  not
  g740
  (
    n664,
    n203
  );


  not
  g741
  (
    n626,
    n174
  );


  buf
  g742
  (
    n308,
    n171
  );


  not
  g743
  (
    n362,
    n119
  );


  buf
  g744
  (
    n655,
    n206
  );


  not
  g745
  (
    n418,
    n100
  );


  buf
  g746
  (
    n453,
    n82
  );


  not
  g747
  (
    n477,
    n94
  );


  buf
  g748
  (
    n574,
    n102
  );


  not
  g749
  (
    n379,
    n131
  );


  not
  g750
  (
    n685,
    n186
  );


  not
  g751
  (
    n721,
    n176
  );


  not
  g752
  (
    n538,
    n99
  );


  not
  g753
  (
    n217,
    n176
  );


  buf
  g754
  (
    n851,
    n105
  );


  buf
  g755
  (
    n749,
    n102
  );


  buf
  g756
  (
    n608,
    n99
  );


  not
  g757
  (
    n771,
    n92
  );


  not
  g758
  (
    n649,
    n133
  );


  buf
  g759
  (
    n441,
    n139
  );


  buf
  g760
  (
    n640,
    n125
  );


  not
  g761
  (
    n571,
    n78
  );


  buf
  g762
  (
    n744,
    n177
  );


  not
  g763
  (
    n380,
    n64
  );


  not
  g764
  (
    n820,
    n179
  );


  not
  g765
  (
    n443,
    n193
  );


  not
  g766
  (
    n523,
    n160
  );


  buf
  g767
  (
    n842,
    n149
  );


  buf
  g768
  (
    n697,
    n84
  );


  not
  g769
  (
    n817,
    n184
  );


  not
  g770
  (
    n437,
    n156
  );


  buf
  g771
  (
    n630,
    n207
  );


  not
  g772
  (
    n605,
    n135
  );


  buf
  g773
  (
    n631,
    n146
  );


  buf
  g774
  (
    n802,
    n154
  );


  buf
  g775
  (
    n525,
    n200
  );


  not
  g776
  (
    n516,
    n131
  );


  buf
  g777
  (
    n723,
    n134
  );


  not
  g778
  (
    n250,
    n196
  );


  not
  g779
  (
    n327,
    n62
  );


  buf
  g780
  (
    n431,
    n95
  );


  not
  g781
  (
    n750,
    n155
  );


  buf
  g782
  (
    n260,
    n114
  );


  buf
  g783
  (
    n325,
    n143
  );


  buf
  g784
  (
    n396,
    n135
  );


  buf
  g785
  (
    n382,
    n130
  );


  not
  g786
  (
    n722,
    n118
  );


  buf
  g787
  (
    n511,
    n127
  );


  not
  g788
  (
    n570,
    n202
  );


  not
  g789
  (
    n775,
    n165
  );


  buf
  g790
  (
    n455,
    n74
  );


  buf
  g791
  (
    n326,
    n119
  );


  buf
  g792
  (
    n682,
    n153
  );


  not
  g793
  (
    n275,
    n111
  );


  not
  g794
  (
    n595,
    n159
  );


  not
  g795
  (
    n319,
    n201
  );


  not
  g796
  (
    n619,
    n176
  );


  buf
  g797
  (
    n394,
    n173
  );


  not
  g798
  (
    n482,
    n52
  );


  not
  g799
  (
    n633,
    n200
  );


  buf
  g800
  (
    n819,
    n192
  );


  not
  g801
  (
    n521,
    n126
  );


  buf
  g802
  (
    n348,
    n174
  );


  xnor
  g803
  (
    n949,
    n470,
    n290,
    n447,
    n420
  );


  or
  g804
  (
    n948,
    n429,
    n387,
    n418,
    n445
  );


  xor
  g805
  (
    n916,
    n441,
    n348,
    n584,
    n334
  );


  or
  g806
  (
    n895,
    n656,
    n306,
    n323,
    n281
  );


  or
  g807
  (
    n961,
    n226,
    n384,
    n315,
    n502
  );


  nand
  g808
  (
    n974,
    n625,
    n528,
    n375,
    n642
  );


  nand
  g809
  (
    n893,
    n761,
    n769,
    n771,
    n788
  );


  and
  g810
  (
    n859,
    n758,
    n358,
    n262,
    n609
  );


  nor
  g811
  (
    n878,
    n593,
    n278,
    n512,
    n777
  );


  nor
  g812
  (
    n892,
    n643,
    n551,
    n293,
    n605
  );


  nor
  g813
  (
    n942,
    n751,
    n602,
    n288,
    n545
  );


  and
  g814
  (
    n889,
    n530,
    n667,
    n572,
    n564
  );


  xnor
  g815
  (
    n988,
    n388,
    n608,
    n604,
    n475
  );


  and
  g816
  (
    n955,
    n220,
    n600,
    n424,
    n238
  );


  xor
  g817
  (
    n900,
    n207,
    n535,
    n689,
    n465
  );


  and
  g818
  (
    n968,
    n736,
    n303,
    n340,
    n362
  );


  nor
  g819
  (
    n917,
    n663,
    n491,
    n742,
    n794
  );


  xor
  g820
  (
    n918,
    n623,
    n639,
    n416,
    n511
  );


  or
  g821
  (
    n959,
    n489,
    n628,
    n529,
    n498
  );


  xor
  g822
  (
    n899,
    n360,
    n371,
    n433,
    n658
  );


  nand
  g823
  (
    n962,
    n403,
    n251,
    n611,
    n641
  );


  or
  g824
  (
    n911,
    n634,
    n727,
    n257,
    n504
  );


  xnor
  g825
  (
    n934,
    n563,
    n582,
    n693,
    n601
  );


  nor
  g826
  (
    n935,
    n701,
    n411,
    n263,
    n542
  );


  or
  g827
  (
    n932,
    n786,
    n382,
    n485,
    n302
  );


  nor
  g828
  (
    n869,
    n676,
    n330,
    n749,
    n737
  );


  xnor
  g829
  (
    n923,
    n482,
    n533,
    n432,
    n380
  );


  or
  g830
  (
    n868,
    n633,
    n785,
    n274,
    n754
  );


  xor
  g831
  (
    n958,
    n299,
    n507,
    n265,
    n366
  );


  nor
  g832
  (
    n910,
    n450,
    n493,
    n280,
    n479
  );


  nand
  g833
  (
    n969,
    n789,
    n264,
    n253,
    n589
  );


  xor
  g834
  (
    n896,
    n685,
    n467,
    n648,
    n506
  );


  xnor
  g835
  (
    n865,
    n614,
    n588,
    n461,
    n774
  );


  xor
  g836
  (
    n928,
    n409,
    n252,
    n421,
    n718
  );


  nand
  g837
  (
    n936,
    n228,
    n569,
    n795,
    n574
  );


  and
  g838
  (
    n901,
    n790,
    n462,
    n399,
    n760
  );


  and
  g839
  (
    n913,
    n456,
    n515,
    n679,
    n219
  );


  nand
  g840
  (
    n960,
    n463,
    n596,
    n617,
    n494
  );


  or
  g841
  (
    n938,
    n578,
    n223,
    n250,
    n546
  );


  or
  g842
  (
    n866,
    n446,
    n335,
    n301,
    n757
  );


  and
  g843
  (
    n951,
    n495,
    n417,
    n552,
    n367
  );


  and
  g844
  (
    n920,
    n240,
    n540,
    n464,
    n566
  );


  nor
  g845
  (
    n886,
    n733,
    n695,
    n653,
    n230
  );


  nor
  g846
  (
    n981,
    n428,
    n256,
    n621,
    n324
  );


  and
  g847
  (
    n941,
    n555,
    n597,
    n710,
    n668
  );


  xnor
  g848
  (
    n864,
    n361,
    n513,
    n332,
    n694
  );


  nor
  g849
  (
    n979,
    n644,
    n365,
    n592,
    n452
  );


  nor
  g850
  (
    n984,
    n556,
    n675,
    n791,
    n692
  );


  nor
  g851
  (
    n929,
    n357,
    n442,
    n624,
    n469
  );


  nand
  g852
  (
    n983,
    n747,
    n410,
    n313,
    n570
  );


  xor
  g853
  (
    n858,
    n729,
    n275,
    n440,
    n618
  );


  nor
  g854
  (
    n905,
    n686,
    n327,
    n590,
    n347
  );


  or
  g855
  (
    n952,
    n354,
    n460,
    n717,
    n522
  );


  xor
  g856
  (
    n973,
    n339,
    n286,
    n239,
    n364
  );


  xnor
  g857
  (
    n922,
    n708,
    n343,
    n647,
    n294
  );


  xor
  g858
  (
    n943,
    n422,
    n431,
    n224,
    n547
  );


  and
  g859
  (
    n933,
    n383,
    n688,
    n379,
    n586
  );


  xnor
  g860
  (
    n867,
    n650,
    n743,
    n374,
    n405
  );


  xor
  g861
  (
    n915,
    n439,
    n319,
    n603,
    n594
  );


  xor
  g862
  (
    n987,
    n386,
    n671,
    n407,
    n517
  );


  nor
  g863
  (
    n919,
    n395,
    n630,
    n300,
    n539
  );


  xor
  g864
  (
    n975,
    n350,
    n778,
    n244,
    n304
  );


  or
  g865
  (
    n853,
    n363,
    n497,
    n712,
    n328
  );


  xor
  g866
  (
    n931,
    n599,
    n553,
    n295,
    n659
  );


  or
  g867
  (
    n991,
    n261,
    n268,
    n472,
    n401
  );


  or
  g868
  (
    n950,
    n558,
    n776,
    n466,
    n732
  );


  xnor
  g869
  (
    n921,
    n784,
    n780,
    n753,
    n707
  );


  xnor
  g870
  (
    n937,
    n703,
    n237,
    n698,
    n673
  );


  nand
  g871
  (
    n906,
    n412,
    n458,
    n247,
    n490
  );


  xnor
  g872
  (
    n927,
    n745,
    n266,
    n705,
    n775
  );


  or
  g873
  (
    n926,
    n505,
    n400,
    n322,
    n437
  );


  nand
  g874
  (
    n863,
    n598,
    n550,
    n538,
    n503
  );


  nand
  g875
  (
    n884,
    n393,
    n724,
    n520,
    n782
  );


  nand
  g876
  (
    n872,
    n738,
    n474,
    n662,
    n516
  );


  xor
  g877
  (
    n874,
    n756,
    n235,
    n255,
    n351
  );


  xor
  g878
  (
    n857,
    n748,
    n763,
    n765,
    n344
  );


  and
  g879
  (
    n982,
    n402,
    n587,
    n620,
    n514
  );


  or
  g880
  (
    n940,
    n532,
    n459,
    n276,
    n660
  );


  xor
  g881
  (
    n904,
    n414,
    n372,
    n764,
    n585
  );


  xnor
  g882
  (
    n887,
    n779,
    n486,
    n273,
    n355
  );


  xor
  g883
  (
    n870,
    n752,
    n792,
    n687,
    n426
  );


  xor
  g884
  (
    n956,
    n267,
    n483,
    n534,
    n787
  );


  nor
  g885
  (
    n976,
    n723,
    n218,
    n557,
    n320
  );


  xor
  g886
  (
    n971,
    n562,
    n269,
    n652,
    n773
  );


  or
  g887
  (
    n882,
    n560,
    n317,
    n622,
    n312
  );


  nand
  g888
  (
    n989,
    n651,
    n677,
    n318,
    n523
  );


  xor
  g889
  (
    n890,
    n443,
    n510,
    n316,
    n755
  );


  and
  g890
  (
    n902,
    n481,
    n279,
    n619,
    n683
  );


  and
  g891
  (
    n912,
    n283,
    n715,
    n739,
    n271
  );


  xor
  g892
  (
    n860,
    n478,
    n666,
    n720,
    n356
  );


  xor
  g893
  (
    n925,
    n419,
    n436,
    n455,
    n616
  );


  nor
  g894
  (
    n966,
    n728,
    n338,
    n245,
    n635
  );


  nand
  g895
  (
    n992,
    n243,
    n607,
    n632,
    n438
  );


  nor
  g896
  (
    n894,
    n649,
    n242,
    n711,
    n772
  );


  xnor
  g897
  (
    n881,
    n484,
    n285,
    n615,
    n329
  );


  nand
  g898
  (
    n862,
    n249,
    n565,
    n413,
    n548
  );


  and
  g899
  (
    n970,
    n398,
    n561,
    n337,
    n292
  );


  xor
  g900
  (
    n898,
    n770,
    n640,
    n581,
    n225
  );


  nor
  g901
  (
    n963,
    n744,
    n352,
    n654,
    n699
  );


  and
  g902
  (
    n897,
    n759,
    n377,
    n521,
    n314
  );


  xor
  g903
  (
    n994,
    n310,
    n369,
    n353,
    n696
  );


  or
  g904
  (
    n891,
    n454,
    n722,
    n719,
    n378
  );


  and
  g905
  (
    n930,
    n227,
    n576,
    n451,
    n298
  );


  xnor
  g906
  (
    n875,
    n783,
    n746,
    n396,
    n741
  );


  nand
  g907
  (
    n985,
    n704,
    n793,
    n571,
    n691
  );


  xnor
  g908
  (
    n965,
    n473,
    n305,
    n277,
    n735
  );


  nand
  g909
  (
    n852,
    n331,
    n381,
    n270,
    n664
  );


  or
  g910
  (
    n888,
    n716,
    n449,
    n488,
    n246
  );


  or
  g911
  (
    n996,
    n681,
    n341,
    n531,
    n453
  );


  xnor
  g912
  (
    n856,
    n536,
    n404,
    n713,
    n579
  );


  nor
  g913
  (
    n972,
    n518,
    n231,
    n731,
    n389
  );


  xnor
  g914
  (
    n967,
    n645,
    n448,
    n241,
    n670
  );


  xnor
  g915
  (
    n903,
    n349,
    n415,
    n333,
    n346
  );


  and
  g916
  (
    n855,
    n629,
    n359,
    n509,
    n408
  );


  nand
  g917
  (
    n964,
    n549,
    n610,
    n222,
    n326
  );


  nor
  g918
  (
    n879,
    n457,
    n730,
    n311,
    n248
  );


  and
  g919
  (
    n873,
    n373,
    n376,
    n740,
    n684
  );


  or
  g920
  (
    n990,
    n568,
    n697,
    n307,
    n537
  );


  xor
  g921
  (
    n885,
    n613,
    n674,
    n526,
    n544
  );


  nor
  g922
  (
    n947,
    n406,
    n519,
    n287,
    n527
  );


  and
  g923
  (
    n907,
    n427,
    n236,
    n390,
    n525
  );


  xor
  g924
  (
    n908,
    n444,
    n471,
    n233,
    n750
  );


  and
  g925
  (
    n909,
    n487,
    n342,
    n725,
    n655
  );


  xor
  g926
  (
    n861,
    n309,
    n259,
    n700,
    n591
  );


  or
  g927
  (
    n953,
    n284,
    n612,
    n595,
    n260
  );


  xor
  g928
  (
    n939,
    n657,
    n682,
    n468,
    n661
  );


  xnor
  g929
  (
    n978,
    n709,
    n423,
    n606,
    n234
  );


  and
  g930
  (
    n986,
    n706,
    n480,
    n714,
    n282
  );


  nand
  g931
  (
    n944,
    n325,
    n781,
    n258,
    n434
  );


  or
  g932
  (
    n924,
    n768,
    n678,
    n492,
    n627
  );


  and
  g933
  (
    n946,
    n345,
    n541,
    n336,
    n680
  );


  or
  g934
  (
    n954,
    n577,
    n297,
    n291,
    n477
  );


  nor
  g935
  (
    n854,
    n394,
    n646,
    n500,
    n573
  );


  xor
  g936
  (
    n876,
    n397,
    n499,
    n496,
    n554
  );


  or
  g937
  (
    n883,
    n232,
    n626,
    n476,
    n721
  );


  xnor
  g938
  (
    n880,
    n669,
    n665,
    n289,
    n726
  );


  or
  g939
  (
    n993,
    n229,
    n767,
    n690,
    n296
  );


  nor
  g940
  (
    n877,
    n580,
    n430,
    n524,
    n637
  );


  and
  g941
  (
    n957,
    n559,
    n308,
    n501,
    n391
  );


  and
  g942
  (
    n914,
    n370,
    n272,
    n385,
    n368
  );


  and
  g943
  (
    n945,
    n636,
    n567,
    n435,
    n702
  );


  xor
  g944
  (
    n995,
    n254,
    n672,
    n221,
    n321
  );


  or
  g945
  (
    n980,
    n631,
    n508,
    n762,
    n217
  );


  and
  g946
  (
    n871,
    n425,
    n734,
    n543,
    n583
  );


  xor
  g947
  (
    n977,
    n766,
    n638,
    n575,
    n392
  );


  xnor
  g948
  (
    n1001,
    n852,
    n864
  );


  nor
  g949
  (
    n1004,
    n869,
    n874
  );


  xnor
  g950
  (
    n1003,
    n879,
    n881
  );


  nor
  g951
  (
    n1005,
    n878,
    n883
  );


  or
  g952
  (
    n999,
    n872,
    n859
  );


  xor
  g953
  (
    n1007,
    n871,
    n876
  );


  xor
  g954
  (
    n1002,
    n863,
    n868
  );


  nand
  g955
  (
    n1008,
    n877,
    n856
  );


  or
  g956
  (
    n1009,
    n882,
    n860
  );


  xnor
  g957
  (
    n1000,
    n853,
    n854
  );


  nor
  g958
  (
    n997,
    n867,
    n865
  );


  nand
  g959
  (
    n998,
    n857,
    n873
  );


  and
  g960
  (
    n1011,
    n858,
    n862
  );


  xor
  g961
  (
    n1006,
    n866,
    n880
  );


  and
  g962
  (
    n1012,
    n855,
    n875
  );


  and
  g963
  (
    n1010,
    n870,
    n861
  );


  buf
  g964
  (
    n1013,
    n998
  );


  buf
  g965
  (
    n1014,
    n997
  );


  buf
  g966
  (
    n1018,
    n1013
  );


  not
  g967
  (
    n1017,
    n1013
  );


  not
  g968
  (
    n1016,
    n1013
  );


  not
  g969
  (
    n1015,
    n1013
  );


  xor
  g970
  (
    n1019,
    n900,
    n1001,
    n1015,
    n1003
  );


  xor
  g971
  (
    n1025,
    n906,
    n1004,
    n887,
    n902
  );


  xnor
  g972
  (
    n1022,
    n1015,
    n1001,
    n911,
    n999
  );


  xnor
  g973
  (
    n1024,
    n1001,
    n1016,
    n897,
    n905
  );


  nand
  g974
  (
    n1021,
    n889,
    n1017,
    n899,
    n1002
  );


  and
  g975
  (
    n1020,
    n884,
    n891,
    n1015,
    n910
  );


  nor
  g976
  (
    n1027,
    n1016,
    n1000,
    n907,
    n901
  );


  nand
  g977
  (
    n1032,
    n1004,
    n1017,
    n1002,
    n898
  );


  nor
  g978
  (
    n1033,
    n1000,
    n894,
    n1017,
    n1016
  );


  nor
  g979
  (
    n1023,
    n1018,
    n1018,
    n890,
    n1001
  );


  or
  g980
  (
    n1031,
    n912,
    n904,
    n1018,
    n1015
  );


  xor
  g981
  (
    n1034,
    n903,
    n1017,
    n886,
    n1002
  );


  and
  g982
  (
    n1029,
    n1018,
    n888,
    n1003
  );


  nand
  g983
  (
    n1028,
    n1016,
    n1003,
    n885,
    n895
  );


  nor
  g984
  (
    n1030,
    n909,
    n893,
    n1004,
    n892
  );


  or
  g985
  (
    n1026,
    n896,
    n1000,
    n908,
    n1002
  );


  or
  g986
  (
    n1037,
    n46,
    n47,
    n48
  );


  xor
  g987
  (
    n1041,
    n43,
    n1023,
    n45,
    n44
  );


  xnor
  g988
  (
    n1042,
    n43,
    n1026,
    n48,
    n45
  );


  xor
  g989
  (
    n1040,
    n1022,
    n43,
    n47,
    n44
  );


  nand
  g990
  (
    n1038,
    n43,
    n46,
    n1020,
    n1025
  );


  nand
  g991
  (
    n1036,
    n44,
    n45,
    n48,
    n1021
  );


  nor
  g992
  (
    n1039,
    n45,
    n48,
    n1019,
    n46
  );


  or
  g993
  (
    n1035,
    n46,
    n47,
    n1024,
    n44
  );


  not
  g994
  (
    n1063,
    n1040
  );


  not
  g995
  (
    n1050,
    n210
  );


  buf
  g996
  (
    n1060,
    n1038
  );


  buf
  g997
  (
    n1052,
    n1039
  );


  not
  g998
  (
    n1051,
    n1037
  );


  buf
  g999
  (
    n1061,
    n210
  );


  not
  g1000
  (
    n1047,
    n209
  );


  not
  g1001
  (
    n1059,
    n209
  );


  buf
  g1002
  (
    n1057,
    n208
  );


  not
  g1003
  (
    n1043,
    n208
  );


  not
  g1004
  (
    n1056,
    n1042
  );


  buf
  g1005
  (
    n1046,
    n1036
  );


  buf
  g1006
  (
    n1048,
    n208
  );


  not
  g1007
  (
    n1044,
    n1035
  );


  buf
  g1008
  (
    n1058,
    n1042
  );


  not
  g1009
  (
    n1062,
    n1041
  );


  not
  g1010
  (
    n1045,
    n1036
  );


  xor
  g1011
  (
    n1053,
    n1037,
    n1041,
    n1038
  );


  or
  g1012
  (
    n1054,
    n1041,
    n210,
    n209,
    n1040
  );


  and
  g1013
  (
    n1049,
    n1039,
    n209,
    n1040,
    n1042
  );


  xor
  g1014
  (
    n1055,
    n1040,
    n1035,
    n208,
    n1041
  );


  not
  g1015
  (
    n1075,
    n1043
  );


  buf
  g1016
  (
    n1067,
    n1043
  );


  buf
  g1017
  (
    n1065,
    n1043
  );


  not
  g1018
  (
    n1074,
    n796
  );


  buf
  g1019
  (
    n1071,
    n1044
  );


  buf
  g1020
  (
    n1070,
    n1044
  );


  buf
  g1021
  (
    n1064,
    n1045
  );


  buf
  g1022
  (
    n1072,
    n1045
  );


  not
  g1023
  (
    n1066,
    n1044
  );


  buf
  g1024
  (
    n1073,
    n1044
  );


  and
  g1025
  (
    n1068,
    n1043,
    n798
  );


  and
  g1026
  (
    n1069,
    n797,
    n1045,
    n799
  );


  buf
  g1027
  (
    n1085,
    n1064
  );


  not
  g1028
  (
    n1077,
    n1066
  );


  not
  g1029
  (
    n1089,
    n1067
  );


  not
  g1030
  (
    n1081,
    n1067
  );


  not
  g1031
  (
    n1080,
    n1067
  );


  not
  g1032
  (
    n1087,
    n1067
  );


  buf
  g1033
  (
    n1079,
    n1064
  );


  not
  g1034
  (
    n1090,
    n1066
  );


  not
  g1035
  (
    n1082,
    n1065
  );


  buf
  g1036
  (
    n1088,
    n1064
  );


  buf
  g1037
  (
    n1076,
    n1066
  );


  not
  g1038
  (
    n1078,
    n1065
  );


  buf
  g1039
  (
    n1084,
    n1066
  );


  buf
  g1040
  (
    n1086,
    n1064
  );


  buf
  g1041
  (
    n1083,
    n1065
  );


  buf
  g1042
  (
    n1091,
    n1065
  );


  not
  g1043
  (
    n1105,
    n1079
  );


  not
  g1044
  (
    n1108,
    n1077
  );


  not
  g1045
  (
    n1107,
    n1076
  );


  not
  g1046
  (
    n1093,
    n1079
  );


  buf
  g1047
  (
    n1103,
    n1080
  );


  not
  g1048
  (
    n1095,
    n1078
  );


  buf
  g1049
  (
    n1106,
    n1079
  );


  buf
  g1050
  (
    n1098,
    n1077
  );


  not
  g1051
  (
    n1096,
    n1076
  );


  buf
  g1052
  (
    n1099,
    n1078
  );


  buf
  g1053
  (
    n1094,
    n1080
  );


  not
  g1054
  (
    n1100,
    n1077
  );


  buf
  g1055
  (
    n1104,
    n1078
  );


  buf
  g1056
  (
    n1109,
    n1077
  );


  not
  g1057
  (
    n1092,
    n1076
  );


  buf
  g1058
  (
    n1101,
    n1078
  );


  not
  g1059
  (
    n1097,
    n1076
  );


  not
  g1060
  (
    n1102,
    n1079
  );


  not
  g1061
  (
    n1115,
    n918
  );


  not
  g1062
  (
    n1119,
    n1094
  );


  buf
  g1063
  (
    n1117,
    n1092
  );


  not
  g1064
  (
    n1123,
    n914
  );


  not
  g1065
  (
    n1111,
    n1095
  );


  not
  g1066
  (
    n1126,
    n1094
  );


  not
  g1067
  (
    n1121,
    n1092
  );


  not
  g1068
  (
    n1127,
    n1014
  );


  not
  g1069
  (
    n1112,
    n1093
  );


  buf
  g1070
  (
    n1118,
    n1096
  );


  not
  g1071
  (
    n1122,
    n1014
  );


  not
  g1072
  (
    n1113,
    n1095
  );


  buf
  g1073
  (
    n1124,
    n1096
  );


  not
  g1074
  (
    n1116,
    n1014
  );


  buf
  g1075
  (
    n1110,
    n1095
  );


  xnor
  g1076
  (
    n1128,
    n915,
    n913
  );


  or
  g1077
  (
    n1114,
    n916,
    n917,
    n1093,
    n1096
  );


  and
  g1078
  (
    n1125,
    n1014,
    n1094,
    n1093
  );


  and
  g1079
  (
    n1120,
    n1094,
    n1092,
    n1095
  );


  xnor
  g1080
  (
    n1136,
    n214,
    n1122,
    n215
  );


  and
  g1081
  (
    n1131,
    n1121,
    n1120,
    n216,
    n210
  );


  nor
  g1082
  (
    n1137,
    n216,
    n1124,
    n919,
    n211
  );


  or
  g1083
  (
    n1129,
    n211,
    n214,
    n920,
    n1127
  );


  xnor
  g1084
  (
    n1130,
    n1125,
    n216,
    n212
  );


  xor
  g1085
  (
    n1132,
    n213,
    n213,
    n211,
    n1128
  );


  nor
  g1086
  (
    n1133,
    n211,
    n214,
    n212
  );


  and
  g1087
  (
    n1134,
    n1126,
    n213,
    n214
  );


  xnor
  g1088
  (
    n1135,
    n216,
    n215,
    n1123
  );


  nor
  g1089
  (
    n1149,
    n805,
    n808,
    n811,
    n801
  );


  xor
  g1090
  (
    n1144,
    n1028,
    n1031,
    n802,
    n1132
  );


  or
  g1091
  (
    n1145,
    n1132,
    n1133,
    n807,
    n814
  );


  xor
  g1092
  (
    n1146,
    n820,
    n804,
    n825,
    n824
  );


  xor
  g1093
  (
    n1147,
    n809,
    n1033,
    n1029,
    n1129
  );


  or
  g1094
  (
    n1141,
    n803,
    n812,
    n1133,
    n1131
  );


  nor
  g1095
  (
    n1148,
    n821,
    n1134,
    n1130,
    n1129
  );


  or
  g1096
  (
    n1140,
    n806,
    n1134,
    n819,
    n827
  );


  nor
  g1097
  (
    n1138,
    n813,
    n1130,
    n818,
    n1032
  );


  nor
  g1098
  (
    n1139,
    n816,
    n822,
    n817,
    n1131
  );


  nand
  g1099
  (
    n1143,
    n800,
    n810,
    n815,
    n1034
  );


  xnor
  g1100
  (
    n1142,
    n826,
    n1027,
    n1030,
    n823
  );


  not
  g1101
  (
    n1155,
    n1138
  );


  not
  g1102
  (
    n1150,
    n1138
  );


  not
  g1103
  (
    n1151,
    n1139
  );


  not
  g1104
  (
    n1154,
    n1139
  );


  not
  g1105
  (
    n1153,
    n1139
  );


  not
  g1106
  (
    n1152,
    n1139
  );


  nor
  g1107
  (
    n1158,
    n1057,
    n1152,
    n1062,
    n1054
  );


  nor
  g1108
  (
    n1175,
    n1058,
    n1153,
    n1055,
    n1061
  );


  and
  g1109
  (
    n1160,
    n1063,
    n1154,
    n1057
  );


  xor
  g1110
  (
    n1167,
    n1051,
    n1150,
    n1060,
    n1059
  );


  xor
  g1111
  (
    n1177,
    n1153,
    n1052,
    n1154,
    n1051
  );


  xor
  g1112
  (
    n1168,
    n1059,
    n1056,
    n1050,
    n1063
  );


  xor
  g1113
  (
    n1165,
    n1150,
    n1155,
    n1053
  );


  or
  g1114
  (
    n1171,
    n1063,
    n1152,
    n1047,
    n1051
  );


  and
  g1115
  (
    n1161,
    n1062,
    n1059,
    n1053,
    n1054
  );


  nor
  g1116
  (
    n1159,
    n1052,
    n1051,
    n1153,
    n1055
  );


  nor
  g1117
  (
    n1178,
    n1054,
    n1055,
    n1151,
    n1153
  );


  or
  g1118
  (
    n1173,
    n1154,
    n1049,
    n1152,
    n1050
  );


  nor
  g1119
  (
    n1170,
    n1060,
    n1060,
    n1049,
    n1055
  );


  nand
  g1120
  (
    n1156,
    n1151,
    n1048,
    n1047,
    n1046
  );


  nor
  g1121
  (
    n1176,
    n1155,
    n1151,
    n1054,
    n1058
  );


  or
  g1122
  (
    n1169,
    n1059,
    n1150,
    n1152,
    n1060
  );


  xor
  g1123
  (
    n1172,
    n1155,
    n1049,
    n1056
  );


  xor
  g1124
  (
    n1163,
    n1056,
    n1155,
    n1151,
    n1063
  );


  xor
  g1125
  (
    n1162,
    n1046,
    n1048,
    n1150
  );


  and
  g1126
  (
    n1164,
    n1047,
    n1053,
    n1046,
    n1061
  );


  and
  g1127
  (
    n1166,
    n1047,
    n1062,
    n1061
  );


  xnor
  g1128
  (
    n1174,
    n1050,
    n1057,
    n1052,
    n1049
  );


  nor
  g1129
  (
    n1157,
    n1154,
    n1058,
    n1061,
    n1050
  );


  nor
  g1130
  (
    n1179,
    n1058,
    n1052,
    n1046,
    n1048
  );


  buf
  g1131
  (
    n1183,
    n1156
  );


  buf
  g1132
  (
    n1181,
    n1158
  );


  not
  g1133
  (
    n1182,
    n1157
  );


  buf
  g1134
  (
    n1180,
    n1157
  );


  nand
  g1135
  (
    n1187,
    n1086,
    n1090,
    n1087,
    n1182
  );


  nand
  g1136
  (
    n1190,
    n1183,
    n1091,
    n1087,
    n1084
  );


  xor
  g1137
  (
    n1188,
    n1085,
    n1183,
    n1086,
    n1090
  );


  xnor
  g1138
  (
    n1186,
    n1089,
    n1088,
    n1083,
    n1082
  );


  or
  g1139
  (
    n1192,
    n1088,
    n1090,
    n1180,
    n1081
  );


  xor
  g1140
  (
    n1184,
    n1089,
    n1087,
    n1083,
    n1086
  );


  xnor
  g1141
  (
    n1185,
    n921,
    n1085,
    n1180,
    n1089
  );


  or
  g1142
  (
    n1197,
    n1182,
    n1181,
    n1088,
    n1080
  );


  xor
  g1143
  (
    n1198,
    n1084,
    n1086,
    n1091
  );


  nand
  g1144
  (
    n1193,
    n1088,
    n1084,
    n1083,
    n1180
  );


  or
  g1145
  (
    n1196,
    n1084,
    n1082,
    n1181
  );


  nor
  g1146
  (
    n1199,
    n1080,
    n1083,
    n1085,
    n1183
  );


  xnor
  g1147
  (
    n1195,
    n922,
    n1081,
    n1091
  );


  and
  g1148
  (
    n1194,
    n1180,
    n1181,
    n1085,
    n1090
  );


  and
  g1149
  (
    n1191,
    n1089,
    n1087,
    n1081,
    n1183
  );


  nor
  g1150
  (
    n1189,
    n1082,
    n1182,
    n1181
  );


  xor
  g1151
  (
    n1204,
    n1195,
    n1099,
    n1100,
    n1005
  );


  nand
  g1152
  (
    n1219,
    n1195,
    n1196,
    n1158,
    n1097
  );


  nand
  g1153
  (
    n1203,
    n1006,
    n1007,
    n1102,
    n1191
  );


  and
  g1154
  (
    n1221,
    n1196,
    n1159,
    n1107,
    n1008
  );


  xor
  g1155
  (
    n1208,
    n1103,
    n1187,
    n1098,
    n1188
  );


  xnor
  g1156
  (
    n1224,
    n1101,
    n1186,
    n1160,
    n1105
  );


  nor
  g1157
  (
    n1228,
    n1105,
    n1109,
    n1103,
    n1100
  );


  nand
  g1158
  (
    n1225,
    n1104,
    n1097,
    n1193,
    n1160
  );


  and
  g1159
  (
    n1220,
    n1190,
    n1161,
    n1109,
    n1007
  );


  nor
  g1160
  (
    n1216,
    n1195,
    n1134,
    n1161,
    n1106
  );


  or
  g1161
  (
    n1217,
    n1098,
    n1163,
    n1107,
    n1193
  );


  nor
  g1162
  (
    n1222,
    n1107,
    n1005,
    n1162,
    n1159
  );


  nand
  g1163
  (
    n1211,
    n1007,
    n1106,
    n1005
  );


  or
  g1164
  (
    n1213,
    n1194,
    n1004,
    n1105,
    n1187
  );


  nand
  g1165
  (
    n1212,
    n1100,
    n1190,
    n1105,
    n1108
  );


  or
  g1166
  (
    n1201,
    n1194,
    n1194,
    n1101,
    n1102
  );


  or
  g1167
  (
    n1200,
    n1163,
    n1096,
    n1101,
    n1109
  );


  or
  g1168
  (
    n1226,
    n1163,
    n1108,
    n1097
  );


  and
  g1169
  (
    n1206,
    n1104,
    n1102,
    n1160,
    n1101
  );


  nand
  g1170
  (
    n1209,
    n1008,
    n1108,
    n1007,
    n1005
  );


  and
  g1171
  (
    n1218,
    n1184,
    n1099,
    n1192,
    n1104
  );


  nor
  g1172
  (
    n1214,
    n1162,
    n1103,
    n1189,
    n1163
  );


  and
  g1173
  (
    n1210,
    n1189,
    n1109,
    n1191,
    n1162
  );


  or
  g1174
  (
    n1223,
    n1100,
    n1192,
    n1104,
    n1006
  );


  nand
  g1175
  (
    n1202,
    n1008,
    n1097,
    n1006,
    n1193
  );


  xnor
  g1176
  (
    n1229,
    n1161,
    n1188,
    n1103,
    n1099
  );


  nor
  g1177
  (
    n1215,
    n1102,
    n1160,
    n1194,
    n1186
  );


  xnor
  g1178
  (
    n1227,
    n1161,
    n1195,
    n1162,
    n1193
  );


  nand
  g1179
  (
    n1205,
    n1106,
    n1098,
    n1008,
    n1099
  );


  nand
  g1180
  (
    n1207,
    n1185,
    n1006,
    n1098,
    n1107
  );


  not
  g1181
  (
    n1230,
    n1212
  );


  buf
  g1182
  (
    n1234,
    n1211
  );


  not
  g1183
  (
    n1235,
    n1216
  );


  buf
  g1184
  (
    n1242,
    n1202
  );


  not
  g1185
  (
    n1233,
    n1214
  );


  buf
  g1186
  (
    n1245,
    n1207
  );


  buf
  g1187
  (
    n1244,
    n1203
  );


  not
  g1188
  (
    n1240,
    n1210
  );


  not
  g1189
  (
    n1243,
    n1204
  );


  buf
  g1190
  (
    n1237,
    n1200
  );


  buf
  g1191
  (
    n1247,
    n1205
  );


  buf
  g1192
  (
    n1239,
    n1208
  );


  not
  g1193
  (
    n1236,
    n1217
  );


  buf
  g1194
  (
    n1238,
    n1209
  );


  buf
  g1195
  (
    n1231,
    n1213
  );


  not
  g1196
  (
    n1246,
    n1206
  );


  not
  g1197
  (
    n1232,
    n1201
  );


  not
  g1198
  (
    n1241,
    n1215
  );


  not
  g1199
  (
    n1250,
    n1230
  );


  not
  g1200
  (
    n1249,
    n1230
  );


  not
  g1201
  (
    n1248,
    n1230
  );


  nand
  g1202
  (
    n1256,
    n1248,
    n1144,
    n1146,
    n1140
  );


  xor
  g1203
  (
    n1254,
    n1148,
    n1147,
    n1249,
    n1145
  );


  xnor
  g1204
  (
    n1259,
    n1147,
    n1144,
    n1145
  );


  or
  g1205
  (
    n1262,
    n1143,
    n1249,
    n1141,
    n1250
  );


  nor
  g1206
  (
    n1258,
    n1140,
    n1249,
    n1143
  );


  xor
  g1207
  (
    n1257,
    n1148,
    n1146,
    n1142
  );


  xnor
  g1208
  (
    n1253,
    n1147,
    n1248,
    n1141,
    n1146
  );


  nand
  g1209
  (
    n1251,
    n1144,
    n1143,
    n1248,
    n1145
  );


  xor
  g1210
  (
    n1260,
    n1148,
    n1145,
    n1248,
    n1140
  );


  or
  g1211
  (
    n1255,
    n1148,
    n1142,
    n1250
  );


  nand
  g1212
  (
    n1261,
    n1146,
    n1141,
    n1140
  );


  nor
  g1213
  (
    n1252,
    n1250,
    n1147,
    n1249,
    n1142
  );


  buf
  g1214
  (
    n1275,
    n1252
  );


  buf
  g1215
  (
    n1277,
    n956
  );


  not
  g1216
  (
    n1274,
    n933
  );


  nand
  g1217
  (
    n1278,
    n1254,
    n940,
    n936
  );


  or
  g1218
  (
    n1264,
    n1257,
    n953,
    n957,
    n1251
  );


  nand
  g1219
  (
    n1271,
    n951,
    n943,
    n925,
    n960
  );


  xor
  g1220
  (
    n1268,
    n1254,
    n934,
    n1252,
    n939
  );


  or
  g1221
  (
    n1266,
    n954,
    n944,
    n930,
    n937
  );


  or
  g1222
  (
    n1265,
    n927,
    n1257,
    n942,
    n1256
  );


  or
  g1223
  (
    n1276,
    n952,
    n1258,
    n924,
    n931
  );


  xnor
  g1224
  (
    n1269,
    n1253,
    n965,
    n947,
    n962
  );


  xnor
  g1225
  (
    n1280,
    n945,
    n932,
    n1251,
    n948
  );


  xnor
  g1226
  (
    n1267,
    n964,
    n1258,
    n941,
    n963
  );


  or
  g1227
  (
    n1263,
    n935,
    n926,
    n946,
    n1255
  );


  xnor
  g1228
  (
    n1272,
    n938,
    n961,
    n928,
    n949
  );


  and
  g1229
  (
    n1273,
    n923,
    n955,
    n1255,
    n1258
  );


  nor
  g1230
  (
    n1279,
    n966,
    n950,
    n929,
    n1259
  );


  or
  g1231
  (
    n1270,
    n1256,
    n1253,
    n958,
    n959
  );


  or
  g1232
  (
    n1282,
    n1263,
    n1166,
    n1164
  );


  or
  g1233
  (
    n1284,
    n1167,
    n1166,
    n1165,
    n1168
  );


  nor
  g1234
  (
    n1285,
    n1264,
    n1165
  );


  nor
  g1235
  (
    n1283,
    n1167,
    n1166,
    n1265,
    n1164
  );


  or
  g1236
  (
    n1286,
    n1167,
    n1267,
    n1268,
    n1168
  );


  nand
  g1237
  (
    n1281,
    n1266,
    n1167,
    n1164,
    n1166
  );


  buf
  g1238
  (
    n1287,
    n1281
  );


  buf
  g1239
  (
    n1288,
    n1283
  );


  not
  g1240
  (
    n1289,
    n1282
  );


  xor
  g1241
  (
    n1293,
    n1198,
    n1196,
    n1199,
    n1197
  );


  and
  g1242
  (
    n1291,
    n1197,
    n1198,
    n1289
  );


  or
  g1243
  (
    n1290,
    n1288,
    n1197,
    n1289,
    n1287
  );


  xnor
  g1244
  (
    n1292,
    n1199,
    n1199,
    n1269,
    n1288
  );


  or
  g1245
  (
    n1294,
    n1199,
    n1198,
    n1196,
    n1197
  );


  nand
  g1246
  (
    n1296,
    n1279,
    n1136,
    n1226,
    n1219
  );


  xor
  g1247
  (
    n1312,
    n1276,
    n1291,
    n1290,
    n1136
  );


  xnor
  g1248
  (
    n1310,
    n1277,
    n1226,
    n1224
  );


  and
  g1249
  (
    n1306,
    n1294,
    n1293,
    n1292
  );


  xnor
  g1250
  (
    n1299,
    n1135,
    n1229,
    n1222,
    n1225
  );


  xnor
  g1251
  (
    n1311,
    n1275,
    n1136,
    n1227
  );


  nand
  g1252
  (
    n1300,
    n1290,
    n1228,
    n1292,
    n1291
  );


  xor
  g1253
  (
    n1297,
    n1223,
    n1273,
    n1272,
    n1274
  );


  nor
  g1254
  (
    n1304,
    n1229,
    n1294,
    n1137,
    n1278
  );


  or
  g1255
  (
    n1303,
    n1278,
    n1291,
    n1273,
    n1226
  );


  and
  g1256
  (
    n1305,
    n1227,
    n1228,
    n1134,
    n1229
  );


  nor
  g1257
  (
    n1314,
    n1276,
    n1221,
    n1275,
    n1293
  );


  or
  g1258
  (
    n1298,
    n1277,
    n1270,
    n1220,
    n1135
  );


  and
  g1259
  (
    n1307,
    n1277,
    n1292,
    n1135,
    n1290
  );


  xnor
  g1260
  (
    n1295,
    n1218,
    n1225,
    n1293,
    n1229
  );


  nand
  g1261
  (
    n1301,
    n1225,
    n1277,
    n1227,
    n1224
  );


  nand
  g1262
  (
    n1309,
    n1135,
    n1223,
    n1271,
    n1292
  );


  nand
  g1263
  (
    n1308,
    n1228,
    n1272,
    n1290,
    n1278
  );


  or
  g1264
  (
    n1302,
    n1291,
    n1225,
    n1227,
    n1278
  );


  xnor
  g1265
  (
    n1313,
    n1228,
    n1294,
    n1274
  );


  and
  g1266
  (
    n1350,
    n842,
    n1245,
    n1313,
    n1312
  );


  xnor
  g1267
  (
    n1361,
    n1242,
    n1069,
    n844,
    n1238
  );


  or
  g1268
  (
    n1335,
    n829,
    n1011,
    n1238,
    n1074
  );


  nor
  g1269
  (
    n1318,
    n1010,
    n1285,
    n834,
    n1311
  );


  and
  g1270
  (
    n1322,
    n1300,
    n1233,
    n1231,
    n1235
  );


  or
  g1271
  (
    n1352,
    n1072,
    n848,
    n1240,
    n1010
  );


  or
  g1272
  (
    n1347,
    n1069,
    n1012,
    n1305,
    n1301
  );


  nor
  g1273
  (
    n1344,
    n1244,
    n1314,
    n1243,
    n1012
  );


  or
  g1274
  (
    n1328,
    n1241,
    n846,
    n1071,
    n828
  );


  nor
  g1275
  (
    n1343,
    n1069,
    n850,
    n1239
  );


  xor
  g1276
  (
    n1366,
    n1071,
    n1239,
    n847,
    n1074
  );


  or
  g1277
  (
    n1354,
    n1075,
    n839,
    n1302,
    n1073
  );


  and
  g1278
  (
    n1327,
    n1245,
    n830,
    n1242,
    n1244
  );


  nor
  g1279
  (
    n1333,
    n1073,
    n1259,
    n1075,
    n1307
  );


  xnor
  g1280
  (
    n1341,
    n1308,
    n1247,
    n1305,
    n1231
  );


  nor
  g1281
  (
    n1356,
    n1231,
    n1071,
    n1306,
    n1009
  );


  or
  g1282
  (
    n1359,
    n837,
    n1243,
    n840,
    n1070
  );


  xor
  g1283
  (
    n1321,
    n1236,
    n838,
    n831,
    n1012
  );


  xor
  g1284
  (
    n1357,
    n1240,
    n1235,
    n841,
    n1236
  );


  nand
  g1285
  (
    n1355,
    n1011,
    n1299,
    n1309,
    n1298
  );


  nand
  g1286
  (
    n1365,
    n1234,
    n1241,
    n1069,
    n845
  );


  nand
  g1287
  (
    n1362,
    n1149,
    n1279,
    n1313,
    n1247
  );


  nand
  g1288
  (
    n1358,
    n1075,
    n1305,
    n1149,
    n1231
  );


  or
  g1289
  (
    n1342,
    n843,
    n1308,
    n1299,
    n1071
  );


  and
  g1290
  (
    n1340,
    n967,
    n1074,
    n1312,
    n1313
  );


  xnor
  g1291
  (
    n1338,
    n1073,
    n1312,
    n1070,
    n1244
  );


  nor
  g1292
  (
    n1353,
    n1238,
    n1070,
    n1230,
    n1297
  );


  or
  g1293
  (
    n1316,
    n1072,
    n1297,
    n1240,
    n1241
  );


  and
  g1294
  (
    n1324,
    n1009,
    n1308,
    n1242,
    n1307
  );


  xor
  g1295
  (
    n1364,
    n1279,
    n1235,
    n1302,
    n1296
  );


  and
  g1296
  (
    n1351,
    n1068,
    n1243,
    n1244,
    n1234
  );


  or
  g1297
  (
    n1325,
    n1310,
    n1303,
    n1237,
    n1011
  );


  nand
  g1298
  (
    n1348,
    n1314,
    n1234,
    n1309,
    n1295
  );


  xor
  g1299
  (
    n1326,
    n1237,
    n1068,
    n1304,
    n836
  );


  xor
  g1300
  (
    n1329,
    n1070,
    n1072,
    n1296,
    n832
  );


  xnor
  g1301
  (
    n1363,
    n1068,
    n1236,
    n1075,
    n1072
  );


  and
  g1302
  (
    n1337,
    n968,
    n1284,
    n1246,
    n1237
  );


  xnor
  g1303
  (
    n1339,
    n1241,
    n1295,
    n1238,
    n1304
  );


  xnor
  g1304
  (
    n1319,
    n1242,
    n1012,
    n1232,
    n1313
  );


  nor
  g1305
  (
    n1345,
    n1237,
    n1246,
    n969,
    n1234
  );


  xnor
  g1306
  (
    n1317,
    n1309,
    n1232,
    n1042,
    n1233
  );


  or
  g1307
  (
    n1360,
    n1149,
    n851,
    n1009,
    n1010
  );


  nor
  g1308
  (
    n1346,
    n1235,
    n1286,
    n1314,
    n1307
  );


  or
  g1309
  (
    n1315,
    n1247,
    n1301,
    n1243,
    n1068
  );


  nor
  g1310
  (
    n1349,
    n1314,
    n835,
    n1310,
    n1233
  );


  xor
  g1311
  (
    n1331,
    n1311,
    n1011,
    n1310,
    n849
  );


  nor
  g1312
  (
    n1336,
    n1311,
    n1279,
    n1239,
    n1306
  );


  or
  g1313
  (
    n1334,
    n1009,
    n1246,
    n1010,
    n1232
  );


  or
  g1314
  (
    n1320,
    n1298,
    n1245,
    n1074,
    n1236
  );


  nand
  g1315
  (
    n1332,
    n1245,
    n1306,
    n1303,
    n1149
  );


  xnor
  g1316
  (
    n1323,
    n1233,
    n1232,
    n1300,
    n1246
  );


  xor
  g1317
  (
    n1330,
    n1247,
    n1073,
    n1240,
    n833
  );


  xor
  g1318
  (
    n1378,
    n1178,
    n1168,
    n1320,
    n1335
  );


  xor
  g1319
  (
    n1375,
    n1177,
    n1171,
    n992,
    n989
  );


  nor
  g1320
  (
    n1382,
    n1170,
    n1360,
    n1365,
    n1327
  );


  xnor
  g1321
  (
    n1385,
    n1329,
    n1179,
    n990,
    n1259
  );


  xnor
  g1322
  (
    n1389,
    n1325,
    n1352,
    n1350,
    n1174
  );


  and
  g1323
  (
    n1390,
    n1361,
    n1322,
    n1174,
    n1171
  );


  or
  g1324
  (
    n1371,
    n1176,
    n1179,
    n1362,
    n1354
  );


  xnor
  g1325
  (
    n1377,
    n1355,
    n1315,
    n1280,
    n974
  );


  xnor
  g1326
  (
    n1374,
    n1364,
    n1178,
    n1324,
    n1176
  );


  xnor
  g1327
  (
    n1397,
    n1363,
    n1340,
    n993,
    n1260
  );


  xor
  g1328
  (
    n1381,
    n1137,
    n1172,
    n1168
  );


  xnor
  g1329
  (
    n1391,
    n1280,
    n1323,
    n971,
    n1177
  );


  nor
  g1330
  (
    n1368,
    n1353,
    n1346,
    n1333,
    n1137
  );


  xnor
  g1331
  (
    n1370,
    n978,
    n1170,
    n1280,
    n1356
  );


  and
  g1332
  (
    n1398,
    n1172,
    n1345,
    n984,
    n982
  );


  nand
  g1333
  (
    n1379,
    n1169,
    n1177,
    n1171,
    n1178
  );


  xnor
  g1334
  (
    n1395,
    n1326,
    n979,
    n1173,
    n1316
  );


  xnor
  g1335
  (
    n1367,
    n1321,
    n1178,
    n1169,
    n1343
  );


  nor
  g1336
  (
    n1386,
    n1179,
    n994,
    n1170,
    n973
  );


  and
  g1337
  (
    n1388,
    n1338,
    n1179,
    n1357,
    n1366
  );


  nand
  g1338
  (
    n1394,
    n1334,
    n1331,
    n1342,
    n1344
  );


  xor
  g1339
  (
    n1369,
    n1259,
    n1349,
    n1339,
    n1359
  );


  nand
  g1340
  (
    n1396,
    n991,
    n983,
    n1319,
    n1170
  );


  xnor
  g1341
  (
    n1393,
    n986,
    n1348,
    n975,
    n1260
  );


  and
  g1342
  (
    n1383,
    n995,
    n1328,
    n976,
    n970
  );


  nand
  g1343
  (
    n1392,
    n1171,
    n1175,
    n987,
    n1358
  );


  and
  g1344
  (
    n1384,
    n1175,
    n1351,
    n1173,
    n1318
  );


  xor
  g1345
  (
    n1372,
    n977,
    n1169,
    n981,
    n1175
  );


  nand
  g1346
  (
    n1376,
    n1330,
    n1174,
    n1137,
    n972
  );


  xnor
  g1347
  (
    n1400,
    n1280,
    n1337,
    n1173,
    n985
  );


  and
  g1348
  (
    n1373,
    n996,
    n1177,
    n1317,
    n980
  );


  or
  g1349
  (
    n1387,
    n1174,
    n1332,
    n1169,
    n1172
  );


  nor
  g1350
  (
    n1380,
    n988,
    n1176,
    n1341
  );


  xnor
  g1351
  (
    n1399,
    n1336,
    n1175,
    n1173,
    n1347
  );


  or
  g1352
  (
    n1401,
    n1384,
    n1372,
    n1400,
    n1376
  );


  xor
  g1353
  (
    n1403,
    n1379,
    n1371,
    n1390,
    n1260
  );


  or
  g1354
  (
    n1405,
    n1262,
    n1388,
    n1398,
    n1374
  );


  and
  g1355
  (
    n1410,
    n1375,
    n1399,
    n1261,
    n1394
  );


  nand
  g1356
  (
    n1409,
    n1262,
    n1387,
    n1261,
    n1395
  );


  nor
  g1357
  (
    n1411,
    n1369,
    n1389,
    n1261,
    n1380
  );


  and
  g1358
  (
    n1402,
    n1377,
    n1370,
    n1397,
    n1383
  );


  xor
  g1359
  (
    n1406,
    n1373,
    n1378,
    n1260,
    n1381
  );


  nand
  g1360
  (
    n1404,
    n1367,
    n1393,
    n1368,
    n1386
  );


  nand
  g1361
  (
    n1407,
    n1382,
    n1261,
    n1392,
    n1391
  );


  xor
  g1362
  (
    AntiSAT_key_wire,
    n1385,
    n1396,
    n1262
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_0,
    keyIn_0_48,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_1,
    keyIn_0_49,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_2,
    keyIn_0_50,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_3,
    keyIn_0_51,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_4,
    keyIn_0_52,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_5,
    keyIn_0_53,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_6,
    keyIn_0_54,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_7,
    keyIn_0_55,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_8,
    keyIn_0_56,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_9,
    keyIn_0_57,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_10,
    keyIn_0_58,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_11,
    keyIn_0_59,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_12,
    keyIn_0_60,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_13,
    keyIn_0_61,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_14,
    keyIn_0_62,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_15,
    keyIn_0_63,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_64
  (
    gbar_input_0_16,
    keyIn_0_64,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_65
  (
    gbar_input_0_17,
    keyIn_0_65,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_66
  (
    gbar_input_0_18,
    keyIn_0_66,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_67
  (
    gbar_input_0_19,
    keyIn_0_67,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_68
  (
    gbar_input_0_20,
    keyIn_0_68,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_69
  (
    gbar_input_0_21,
    keyIn_0_69,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_70
  (
    gbar_input_0_22,
    keyIn_0_70,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_71
  (
    gbar_input_0_23,
    keyIn_0_71,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_72
  (
    gbar_input_0_24,
    keyIn_0_72,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_73
  (
    gbar_input_0_25,
    keyIn_0_73,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_74
  (
    gbar_input_0_26,
    keyIn_0_74,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_75
  (
    gbar_input_0_27,
    keyIn_0_75,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_76
  (
    gbar_input_0_28,
    keyIn_0_76,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_77
  (
    gbar_input_0_29,
    keyIn_0_77,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_78
  (
    gbar_input_0_30,
    keyIn_0_78,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_79
  (
    gbar_input_0_31,
    keyIn_0_79,
    n32
  );


  xor
  KeyPIGate_0_32
  (
    g_input_0_32,
    keyIn_0_32,
    n33
  );


  xor
  KeyPIGate_0_80
  (
    gbar_input_0_32,
    keyIn_0_80,
    n33
  );


  xor
  KeyPIGate_0_33
  (
    g_input_0_33,
    keyIn_0_33,
    n34
  );


  xor
  KeyPIGate_0_81
  (
    gbar_input_0_33,
    keyIn_0_81,
    n34
  );


  xor
  KeyPIGate_0_34
  (
    g_input_0_34,
    keyIn_0_34,
    n35
  );


  xor
  KeyPIGate_0_82
  (
    gbar_input_0_34,
    keyIn_0_82,
    n35
  );


  xor
  KeyPIGate_0_35
  (
    g_input_0_35,
    keyIn_0_35,
    n36
  );


  xor
  KeyPIGate_0_83
  (
    gbar_input_0_35,
    keyIn_0_83,
    n36
  );


  xor
  KeyPIGate_0_36
  (
    g_input_0_36,
    keyIn_0_36,
    n37
  );


  xor
  KeyPIGate_0_84
  (
    gbar_input_0_36,
    keyIn_0_84,
    n37
  );


  xor
  KeyPIGate_0_37
  (
    g_input_0_37,
    keyIn_0_37,
    n38
  );


  xor
  KeyPIGate_0_85
  (
    gbar_input_0_37,
    keyIn_0_85,
    n38
  );


  xor
  KeyPIGate_0_38
  (
    g_input_0_38,
    keyIn_0_38,
    n39
  );


  xor
  KeyPIGate_0_86
  (
    gbar_input_0_38,
    keyIn_0_86,
    n39
  );


  xor
  KeyPIGate_0_39
  (
    g_input_0_39,
    keyIn_0_39,
    n40
  );


  xor
  KeyPIGate_0_87
  (
    gbar_input_0_39,
    keyIn_0_87,
    n40
  );


  xor
  KeyPIGate_0_40
  (
    g_input_0_40,
    keyIn_0_40,
    n41
  );


  xor
  KeyPIGate_0_88
  (
    gbar_input_0_40,
    keyIn_0_88,
    n41
  );


  xor
  KeyPIGate_0_41
  (
    g_input_0_41,
    keyIn_0_41,
    n42
  );


  xor
  KeyPIGate_0_89
  (
    gbar_input_0_41,
    keyIn_0_89,
    n42
  );


  xor
  KeyPIGate_0_42
  (
    g_input_0_42,
    keyIn_0_42,
    n43
  );


  xor
  KeyPIGate_0_90
  (
    gbar_input_0_42,
    keyIn_0_90,
    n43
  );


  xor
  KeyPIGate_0_43
  (
    g_input_0_43,
    keyIn_0_43,
    n44
  );


  xor
  KeyPIGate_0_91
  (
    gbar_input_0_43,
    keyIn_0_91,
    n44
  );


  xor
  KeyPIGate_0_44
  (
    g_input_0_44,
    keyIn_0_44,
    n45
  );


  xor
  KeyPIGate_0_92
  (
    gbar_input_0_44,
    keyIn_0_92,
    n45
  );


  xor
  KeyPIGate_0_45
  (
    g_input_0_45,
    keyIn_0_45,
    n46
  );


  xor
  KeyPIGate_0_93
  (
    gbar_input_0_45,
    keyIn_0_93,
    n46
  );


  xor
  KeyPIGate_0_46
  (
    g_input_0_46,
    keyIn_0_46,
    n47
  );


  xor
  KeyPIGate_0_94
  (
    gbar_input_0_46,
    keyIn_0_94,
    n47
  );


  xor
  KeyPIGate_0_47
  (
    g_input_0_47,
    keyIn_0_47,
    n48
  );


  xor
  KeyPIGate_0_95
  (
    gbar_input_0_47,
    keyIn_0_95,
    n48
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31,
    g_input_0_32,
    g_input_0_33,
    g_input_0_34,
    g_input_0_35,
    g_input_0_36,
    g_input_0_37,
    g_input_0_38,
    g_input_0_39,
    g_input_0_40,
    g_input_0_41,
    g_input_0_42,
    g_input_0_43,
    g_input_0_44,
    g_input_0_45,
    g_input_0_46,
    g_input_0_47
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31,
    gbar_input_0_32,
    gbar_input_0_33,
    gbar_input_0_34,
    gbar_input_0_35,
    gbar_input_0_36,
    gbar_input_0_37,
    gbar_input_0_38,
    gbar_input_0_39,
    gbar_input_0_40,
    gbar_input_0_41,
    gbar_input_0_42,
    gbar_input_0_43,
    gbar_input_0_44,
    gbar_input_0_45,
    gbar_input_0_46,
    gbar_input_0_47
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n1408,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

