// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_147_624 written by SynthGen on 2021/05/24 19:45:40
module Stat_147_624( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18,
 n141, n149, n157, n162, n160, n165, n154, n151,
 n163, n158, n164, n150, n156, n161, n152, n153,
 n159, n155);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18;

output n141, n149, n157, n162, n160, n165, n154, n151,
 n163, n158, n164, n150, n156, n161, n152, n153,
 n159, n155;

wire n19, n20, n21, n22, n23, n24, n25, n26,
 n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n142, n143, n144, n145, n146, n147,
 n148;

not  g0 (n51, n2);
buf  g1 (n44, n6);
not  g2 (n59, n10);
not  g3 (n46, n12);
buf  g4 (n38, n1);
not  g5 (n39, n9);
buf  g6 (n32, n10);
buf  g7 (n58, n9);
not  g8 (n55, n7);
not  g9 (n31, n5);
not  g10 (n35, n8);
buf  g11 (n63, n8);
buf  g12 (n20, n11);
buf  g13 (n52, n6);
not  g14 (n56, n11);
not  g15 (n24, n7);
not  g16 (n50, n2);
not  g17 (n21, n12);
buf  g18 (n53, n3);
not  g19 (n49, n4);
not  g20 (n26, n5);
buf  g21 (n47, n5);
not  g22 (n28, n3);
buf  g23 (n43, n10);
buf  g24 (n64, n2);
buf  g25 (n19, n7);
buf  g26 (n34, n1);
not  g27 (n57, n5);
not  g28 (n62, n3);
buf  g29 (n29, n1);
not  g30 (n30, n2);
not  g31 (n33, n10);
buf  g32 (n22, n4);
not  g33 (n23, n8);
not  g34 (n40, n4);
not  g35 (n37, n6);
buf  g36 (n25, n9);
buf  g37 (n60, n9);
not  g38 (n45, n6);
not  g39 (n27, n3);
buf  g40 (n54, n11);
not  g41 (n48, n1);
not  g42 (n41, n8);
not  g43 (n42, n11);
not  g44 (n36, n4);
buf  g45 (n61, n7);
xor  g46 (n65, n19, n20);
xnor g47 (n66, n20, n19);
buf  g48 (n68, n66);
buf  g49 (n69, n66);
not  g50 (n67, n66);
not  g51 (n70, n66);
or   g52 (n83, n13, n17);
xnor g53 (n77, n15, n67);
xor  g54 (n84, n69, n15);
xor  g55 (n78, n70, n68);
nand g56 (n82, n70, n67);
xnor g57 (n71, n12, n17);
buf  g58 (n73, n18);
not  g59 (n85, n70);
xor  g60 (n74, n14, n69);
xnor g61 (n81, n16, n14);
buf  g62 (n76, n16);
nor  g63 (n72, n68, n13, n67);
and  g64 (n75, n16, n15, n69, n12);
or   g65 (n80, n68, n17, n69);
xor  g66 (n86, n18, n67, n68, n14);
nor  g67 (n79, n14, n13, n18, n15);
nand g68 (n147, n62, n22, n82);
xnor g69 (n109, n29, n76, n75);
nand g70 (n148, n21, n28, n55);
and  g71 (n125, n86, n30, n36);
xor  g72 (n126, n42, n72, n27);
and  g73 (n138, n42, n74, n40);
and  g74 (n95, n58, n86, n33);
and  g75 (n117, n22, n45, n30);
nand g76 (n141, n43, n76, n55, n72);
and  g77 (n142, n60, n77, n27, n85);
and  g78 (n100, n51, n86, n24, n71);
xor  g79 (n89, n82, n32, n37, n57);
and  g80 (n130, n51, n43, n40, n78);
nor  g81 (n110, n42, n46, n78, n44);
xor  g82 (n116, n40, n79, n53, n64);
or   g83 (n122, n82, n42, n83, n64);
xnor g84 (n129, n27, n39, n76, n37);
xnor g85 (n137, n35, n61, n62, n32);
and  g86 (n96, n34, n82, n25, n23);
and  g87 (n90, n72, n73, n21, n58);
nor  g88 (n91, n59, n21, n52, n74);
nand g89 (n88, n23, n60, n74, n56);
or   g90 (n120, n77, n33, n47, n61);
xor  g91 (n102, n79, n35, n45, n22);
xor  g92 (n139, n58, n56, n71, n85);
nor  g93 (n121, n38, n43, n75, n31);
or   g94 (n105, n60, n25, n52, n40);
xnor g95 (n104, n36, n44, n51, n85);
nand g96 (n144, n80, n52, n32, n61);
and  g97 (n101, n46, n83, n61, n76);
xor  g98 (n113, n28, n80, n72, n71);
nor  g99 (n115, n33, n74, n77, n50);
xor  g100 (n143, n63, n83, n28);
or   g101 (n106, n84, n36, n75, n30);
xor  g102 (n112, n73, n53, n41, n80);
nor  g103 (n107, n37, n59, n47, n45);
and  g104 (n99, n54, n85, n34, n59);
or   g105 (n140, n62, n59, n26, n57);
or   g106 (n93, n48, n39, n23, n45);
nor  g107 (n123, n47, n24, n64, n39);
nand g108 (n134, n63, n33, n56, n47);
xor  g109 (n128, n62, n30, n48, n37);
or   g110 (n124, n39, n26, n48);
xnor g111 (n132, n29, n31, n77, n35);
and  g112 (n111, n84, n79, n54, n28);
nand g113 (n87, n86, n48, n23, n29);
xnor g114 (n133, n53, n22, n51, n43);
or   g115 (n103, n53, n55, n56, n84);
nor  g116 (n94, n41, n50, n44, n46);
nand g117 (n127, n75, n49, n25, n81);
nor  g118 (n92, n29, n57, n21, n38);
or   g119 (n118, n81, n35, n80, n36);
and  g120 (n136, n54, n27, n73, n46);
nor  g121 (n145, n73, n38, n24);
nor  g122 (n146, n81, n50, n60, n79);
xnor g123 (n114, n34, n34, n50, n71);
or   g124 (n135, n49, n31, n38, n25);
xor  g125 (n131, n78, n49, n55);
xnor g126 (n97, n52, n81, n44, n54);
and  g127 (n98, n57, n31, n41, n63);
xor  g128 (n119, n78, n32, n84, n41);
nor  g129 (n108, n26, n64, n58, n63);
nand g130 (n152, n98, n131, n147, n113);
nor  g131 (n160, n90, n128, n144, n93);
xnor g132 (n163, n148, n147, n94, n140);
nand g133 (n158, n135, n147, n101, n141);
xnor g134 (n156, n121, n114, n89, n99);
nand g135 (n149, n136, n105, n110, n109);
nand g136 (n165, n104, n120, n118, n132);
nor  g137 (n162, n112, n87, n88, n108);
or   g138 (n161, n97, n129, n127, n96);
nand g139 (n155, n102, n148, n126, n125);
or   g140 (n159, n148, n146, n103, n119);
and  g141 (n164, n130, n91, n123, n106);
and  g142 (n150, n116, n107, n111, n95);
nand g143 (n151, n137, n100, n124, n122);
nor  g144 (n154, n117, n147, n92, n145);
xor  g145 (n153, n115, n138, n139, n134);
or   g146 (n157, n143, n148, n133, n142);
endmodule
