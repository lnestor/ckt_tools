

module Stat_1396_16_5
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n1289,
  n1271,
  n1274,
  n1262,
  n1291,
  n1283,
  n1290,
  n1261,
  n1268,
  n1266,
  n1264,
  n1265,
  n1278,
  n1286,
  n1270,
  n1277,
  n1276,
  n1263,
  n1287,
  n1285,
  n1281,
  n1273,
  n1415,
  n1418,
  n1413,
  n1410,
  n1411,
  n1416,
  n1417,
  n1412,
  n1409,
  n1414,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1289;output n1271;output n1274;output n1262;output n1291;output n1283;output n1290;output n1261;output n1268;output n1266;output n1264;output n1265;output n1278;output n1286;output n1270;output n1277;output n1276;output n1263;output n1287;output n1285;output n1281;output n1273;output n1415;output n1418;output n1413;output n1410;output n1411;output n1416;output n1417;output n1412;output n1409;output n1414;
  wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1267;wire n1269;wire n1272;wire n1275;wire n1279;wire n1280;wire n1282;wire n1284;wire n1288;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  buf
  g0
  (
    n90,
    n16
  );


  not
  g1
  (
    n77,
    n2
  );


  buf
  g2
  (
    n57,
    n17
  );


  not
  g3
  (
    n80,
    n5
  );


  buf
  g4
  (
    n88,
    n8
  );


  buf
  g5
  (
    n24,
    n19
  );


  buf
  g6
  (
    n38,
    n11
  );


  buf
  g7
  (
    n23,
    n16
  );


  buf
  g8
  (
    n69,
    n16
  );


  buf
  g9
  (
    n65,
    n19
  );


  buf
  g10
  (
    n58,
    n20
  );


  not
  g11
  (
    n78,
    n13
  );


  not
  g12
  (
    n76,
    n14
  );


  buf
  g13
  (
    n74,
    n10
  );


  not
  g14
  (
    n29,
    n11
  );


  not
  g15
  (
    n81,
    n1
  );


  buf
  g16
  (
    n85,
    n10
  );


  not
  g17
  (
    n39,
    n15
  );


  not
  g18
  (
    n89,
    n12
  );


  not
  g19
  (
    n97,
    n18
  );


  not
  g20
  (
    n67,
    n10
  );


  not
  g21
  (
    n36,
    n15
  );


  buf
  g22
  (
    n32,
    n10
  );


  not
  g23
  (
    n49,
    n5
  );


  buf
  g24
  (
    n75,
    n9
  );


  buf
  g25
  (
    n101,
    n6
  );


  buf
  g26
  (
    n42,
    n19
  );


  not
  g27
  (
    n99,
    n8
  );


  not
  g28
  (
    n95,
    n13
  );


  not
  g29
  (
    n51,
    n13
  );


  buf
  g30
  (
    n92,
    n7
  );


  buf
  g31
  (
    n61,
    n9
  );


  not
  g32
  (
    n55,
    n2
  );


  buf
  g33
  (
    n79,
    n3
  );


  buf
  g34
  (
    n64,
    n2
  );


  not
  g35
  (
    n83,
    n9
  );


  not
  g36
  (
    n53,
    n6
  );


  buf
  g37
  (
    n71,
    n3
  );


  buf
  g38
  (
    n44,
    n5
  );


  not
  g39
  (
    n28,
    n7
  );


  not
  g40
  (
    n93,
    n11
  );


  buf
  g41
  (
    n66,
    n5
  );


  not
  g42
  (
    n52,
    n17
  );


  buf
  g43
  (
    KeyWire_0_14,
    n1
  );


  buf
  g44
  (
    n86,
    n13
  );


  buf
  g45
  (
    n91,
    n8
  );


  buf
  g46
  (
    n33,
    n18
  );


  buf
  g47
  (
    n34,
    n7
  );


  not
  g48
  (
    n30,
    n6
  );


  not
  g49
  (
    n82,
    n4
  );


  not
  g50
  (
    n98,
    n19
  );


  not
  g51
  (
    n27,
    n12
  );


  not
  g52
  (
    n46,
    n17
  );


  not
  g53
  (
    KeyWire_0_31,
    n9
  );


  buf
  g54
  (
    n54,
    n1
  );


  not
  g55
  (
    n72,
    n16
  );


  not
  g56
  (
    n56,
    n20
  );


  not
  g57
  (
    n102,
    n12
  );


  not
  g58
  (
    n62,
    n3
  );


  not
  g59
  (
    n94,
    n6
  );


  not
  g60
  (
    n59,
    n11
  );


  buf
  g61
  (
    n37,
    n12
  );


  not
  g62
  (
    n40,
    n17
  );


  buf
  g63
  (
    n96,
    n14
  );


  not
  g64
  (
    n41,
    n3
  );


  buf
  g65
  (
    n60,
    n4
  );


  buf
  g66
  (
    n73,
    n14
  );


  buf
  g67
  (
    n31,
    n2
  );


  buf
  g68
  (
    n84,
    n20
  );


  buf
  g69
  (
    n35,
    n20
  );


  not
  g70
  (
    n100,
    n18
  );


  not
  g71
  (
    n68,
    n4
  );


  not
  g72
  (
    n50,
    n4
  );


  buf
  g73
  (
    n25,
    n15
  );


  buf
  g74
  (
    n26,
    n14
  );


  not
  g75
  (
    n48,
    n7
  );


  buf
  g76
  (
    n43,
    n1
  );


  buf
  g77
  (
    n47,
    n15
  );


  buf
  g78
  (
    n63,
    n8
  );


  buf
  g79
  (
    n87,
    n18
  );


  not
  g80
  (
    n343,
    n70
  );


  not
  g81
  (
    n355,
    n43
  );


  buf
  g82
  (
    n264,
    n76
  );


  not
  g83
  (
    n129,
    n31
  );


  buf
  g84
  (
    n244,
    n96
  );


  buf
  g85
  (
    n195,
    n100
  );


  buf
  g86
  (
    n358,
    n92
  );


  buf
  g87
  (
    n151,
    n95
  );


  not
  g88
  (
    n399,
    n50
  );


  not
  g89
  (
    n375,
    n24
  );


  not
  g90
  (
    n329,
    n70
  );


  buf
  g91
  (
    n156,
    n46
  );


  buf
  g92
  (
    n217,
    n67
  );


  buf
  g93
  (
    n376,
    n29
  );


  buf
  g94
  (
    n336,
    n71
  );


  not
  g95
  (
    n367,
    n61
  );


  not
  g96
  (
    n152,
    n82
  );


  buf
  g97
  (
    KeyWire_0_25,
    n68
  );


  not
  g98
  (
    n326,
    n39
  );


  not
  g99
  (
    n140,
    n56
  );


  buf
  g100
  (
    n397,
    n93
  );


  not
  g101
  (
    n110,
    n92
  );


  not
  g102
  (
    n351,
    n26
  );


  not
  g103
  (
    n126,
    n46
  );


  buf
  g104
  (
    n107,
    n28
  );


  buf
  g105
  (
    n414,
    n26
  );


  buf
  g106
  (
    n149,
    n79
  );


  buf
  g107
  (
    n410,
    n25
  );


  buf
  g108
  (
    n162,
    n48
  );


  not
  g109
  (
    n160,
    n55
  );


  buf
  g110
  (
    n188,
    n30
  );


  buf
  g111
  (
    n117,
    n82
  );


  buf
  g112
  (
    n280,
    n27
  );


  buf
  g113
  (
    n353,
    n88
  );


  not
  g114
  (
    n158,
    n29
  );


  buf
  g115
  (
    n384,
    n26
  );


  not
  g116
  (
    n252,
    n69
  );


  buf
  g117
  (
    n387,
    n30
  );


  buf
  g118
  (
    n164,
    n54
  );


  buf
  g119
  (
    n263,
    n92
  );


  not
  g120
  (
    n108,
    n78
  );


  buf
  g121
  (
    n148,
    n32
  );


  buf
  g122
  (
    n128,
    n33
  );


  buf
  g123
  (
    n334,
    n77
  );


  not
  g124
  (
    n119,
    n66
  );


  not
  g125
  (
    n255,
    n52
  );


  buf
  g126
  (
    n141,
    n67
  );


  buf
  g127
  (
    n193,
    n44
  );


  not
  g128
  (
    n390,
    n100
  );


  buf
  g129
  (
    n238,
    n83
  );


  buf
  g130
  (
    n190,
    n49
  );


  buf
  g131
  (
    n305,
    n23
  );


  not
  g132
  (
    n403,
    n23
  );


  not
  g133
  (
    n282,
    n77
  );


  not
  g134
  (
    n392,
    n45
  );


  buf
  g135
  (
    n401,
    n88
  );


  not
  g136
  (
    n239,
    n46
  );


  not
  g137
  (
    n216,
    n64
  );


  buf
  g138
  (
    n166,
    n85
  );


  buf
  g139
  (
    n237,
    n37
  );


  not
  g140
  (
    n249,
    n89
  );


  not
  g141
  (
    n223,
    n66
  );


  buf
  g142
  (
    n361,
    n96
  );


  not
  g143
  (
    n269,
    n91
  );


  not
  g144
  (
    n290,
    n41
  );


  buf
  g145
  (
    n114,
    n23
  );


  not
  g146
  (
    n192,
    n101
  );


  not
  g147
  (
    n243,
    n66
  );


  buf
  g148
  (
    n407,
    n85
  );


  buf
  g149
  (
    n327,
    n68
  );


  not
  g150
  (
    n364,
    n28
  );


  buf
  g151
  (
    n165,
    n53
  );


  not
  g152
  (
    n199,
    n40
  );


  buf
  g153
  (
    n250,
    n95
  );


  buf
  g154
  (
    n180,
    n45
  );


  not
  g155
  (
    n330,
    n75
  );


  not
  g156
  (
    n153,
    n62
  );


  buf
  g157
  (
    n159,
    n33
  );


  buf
  g158
  (
    n218,
    n77
  );


  not
  g159
  (
    n413,
    n89
  );


  not
  g160
  (
    n267,
    n90
  );


  buf
  g161
  (
    KeyWire_0_1,
    n55
  );


  buf
  g162
  (
    n396,
    n61
  );


  buf
  g163
  (
    n241,
    n28
  );


  not
  g164
  (
    n278,
    n32
  );


  buf
  g165
  (
    n229,
    n38
  );


  not
  g166
  (
    n279,
    n42
  );


  not
  g167
  (
    n275,
    n34
  );


  not
  g168
  (
    KeyWire_0_11,
    n65
  );


  not
  g169
  (
    n322,
    n96
  );


  buf
  g170
  (
    n183,
    n99
  );


  buf
  g171
  (
    n113,
    n43
  );


  buf
  g172
  (
    n260,
    n53
  );


  buf
  g173
  (
    n235,
    n99
  );


  not
  g174
  (
    n340,
    n41
  );


  not
  g175
  (
    n150,
    n87
  );


  buf
  g176
  (
    n104,
    n71
  );


  buf
  g177
  (
    n369,
    n36
  );


  buf
  g178
  (
    n171,
    n38
  );


  not
  g179
  (
    n179,
    n79
  );


  not
  g180
  (
    n311,
    n60
  );


  not
  g181
  (
    n385,
    n35
  );


  buf
  g182
  (
    n125,
    n48
  );


  not
  g183
  (
    n191,
    n63
  );


  not
  g184
  (
    n246,
    n26
  );


  not
  g185
  (
    n120,
    n62
  );


  buf
  g186
  (
    n176,
    n43
  );


  not
  g187
  (
    n291,
    n51
  );


  not
  g188
  (
    n394,
    n84
  );


  not
  g189
  (
    n258,
    n62
  );


  not
  g190
  (
    n337,
    n72
  );


  not
  g191
  (
    n389,
    n61
  );


  not
  g192
  (
    n286,
    n54
  );


  not
  g193
  (
    n167,
    n51
  );


  buf
  g194
  (
    n339,
    n91
  );


  not
  g195
  (
    n118,
    n84
  );


  not
  g196
  (
    n187,
    n51
  );


  buf
  g197
  (
    n319,
    n74
  );


  buf
  g198
  (
    n347,
    n25
  );


  buf
  g199
  (
    n111,
    n53
  );


  buf
  g200
  (
    n296,
    n93
  );


  buf
  g201
  (
    n200,
    n56
  );


  buf
  g202
  (
    n366,
    n63
  );


  buf
  g203
  (
    n324,
    n85
  );


  buf
  g204
  (
    n300,
    n33
  );


  buf
  g205
  (
    n298,
    n72
  );


  not
  g206
  (
    n133,
    n100
  );


  not
  g207
  (
    n228,
    n70
  );


  not
  g208
  (
    n220,
    n94
  );


  buf
  g209
  (
    KeyWire_0_21,
    n90
  );


  not
  g210
  (
    n372,
    n84
  );


  buf
  g211
  (
    n161,
    n33
  );


  not
  g212
  (
    n219,
    n46
  );


  buf
  g213
  (
    n147,
    n93
  );


  buf
  g214
  (
    n316,
    n86
  );


  buf
  g215
  (
    n380,
    n25
  );


  buf
  g216
  (
    n287,
    n75
  );


  buf
  g217
  (
    n234,
    n29
  );


  not
  g218
  (
    KeyWire_0_3,
    n38
  );


  buf
  g219
  (
    n175,
    n83
  );


  buf
  g220
  (
    n411,
    n71
  );


  not
  g221
  (
    n382,
    n49
  );


  not
  g222
  (
    n398,
    n78
  );


  not
  g223
  (
    n247,
    n47
  );


  buf
  g224
  (
    n360,
    n40
  );


  buf
  g225
  (
    n268,
    n91
  );


  not
  g226
  (
    n341,
    n81
  );


  buf
  g227
  (
    n145,
    n34
  );


  not
  g228
  (
    n371,
    n73
  );


  not
  g229
  (
    n121,
    n39
  );


  buf
  g230
  (
    n253,
    n45
  );


  buf
  g231
  (
    n373,
    n74
  );


  buf
  g232
  (
    n178,
    n29
  );


  buf
  g233
  (
    n314,
    n48
  );


  not
  g234
  (
    n211,
    n54
  );


  not
  g235
  (
    n132,
    n59
  );


  buf
  g236
  (
    n354,
    n58
  );


  not
  g237
  (
    n155,
    n97
  );


  not
  g238
  (
    n273,
    n86
  );


  buf
  g239
  (
    n185,
    n59
  );


  buf
  g240
  (
    n285,
    n60
  );


  buf
  g241
  (
    n400,
    n87
  );


  not
  g242
  (
    n402,
    n28
  );


  buf
  g243
  (
    n194,
    n68
  );


  not
  g244
  (
    n276,
    n95
  );


  buf
  g245
  (
    n144,
    n80
  );


  not
  g246
  (
    n310,
    n69
  );


  not
  g247
  (
    n124,
    n62
  );


  not
  g248
  (
    n302,
    n58
  );


  buf
  g249
  (
    n381,
    n35
  );


  buf
  g250
  (
    n204,
    n43
  );


  buf
  g251
  (
    n348,
    n31
  );


  buf
  g252
  (
    n198,
    n41
  );


  not
  g253
  (
    n123,
    n65
  );


  not
  g254
  (
    n309,
    n44
  );


  not
  g255
  (
    n307,
    n31
  );


  not
  g256
  (
    n405,
    n80
  );


  not
  g257
  (
    n303,
    n45
  );


  not
  g258
  (
    n212,
    n73
  );


  buf
  g259
  (
    n202,
    n81
  );


  not
  g260
  (
    n231,
    n39
  );


  buf
  g261
  (
    n257,
    n72
  );


  buf
  g262
  (
    n197,
    n64
  );


  buf
  g263
  (
    n168,
    n85
  );


  buf
  g264
  (
    n109,
    n97
  );


  buf
  g265
  (
    n295,
    n44
  );


  not
  g266
  (
    n226,
    n99
  );


  buf
  g267
  (
    n349,
    n93
  );


  buf
  g268
  (
    n272,
    n48
  );


  buf
  g269
  (
    n391,
    n63
  );


  buf
  g270
  (
    n404,
    n86
  );


  buf
  g271
  (
    n146,
    n25
  );


  not
  g272
  (
    n383,
    n23
  );


  buf
  g273
  (
    n271,
    n47
  );


  buf
  g274
  (
    n412,
    n86
  );


  buf
  g275
  (
    n352,
    n100
  );


  not
  g276
  (
    n288,
    n94
  );


  buf
  g277
  (
    n205,
    n41
  );


  buf
  g278
  (
    n363,
    n99
  );


  not
  g279
  (
    n379,
    n44
  );


  not
  g280
  (
    n186,
    n75
  );


  buf
  g281
  (
    n377,
    n36
  );


  buf
  g282
  (
    n338,
    n90
  );


  buf
  g283
  (
    n274,
    n50
  );


  not
  g284
  (
    n134,
    n60
  );


  not
  g285
  (
    n415,
    n37
  );


  not
  g286
  (
    n112,
    n56
  );


  not
  g287
  (
    n388,
    n54
  );


  buf
  g288
  (
    n306,
    n55
  );


  not
  g289
  (
    n143,
    n34
  );


  not
  g290
  (
    n251,
    n94
  );


  buf
  g291
  (
    n248,
    n55
  );


  buf
  g292
  (
    n131,
    n79
  );


  buf
  g293
  (
    n139,
    n75
  );


  not
  g294
  (
    n215,
    n34
  );


  buf
  g295
  (
    n362,
    n32
  );


  not
  g296
  (
    n262,
    n78
  );


  buf
  g297
  (
    n142,
    n52
  );


  buf
  g298
  (
    n332,
    n82
  );


  not
  g299
  (
    n173,
    n52
  );


  not
  g300
  (
    n224,
    n32
  );


  buf
  g301
  (
    n242,
    n87
  );


  not
  g302
  (
    n277,
    n73
  );


  not
  g303
  (
    n236,
    n97
  );


  buf
  g304
  (
    n154,
    n38
  );


  not
  g305
  (
    n203,
    n39
  );


  buf
  g306
  (
    n321,
    n66
  );


  not
  g307
  (
    n370,
    n59
  );


  not
  g308
  (
    n266,
    n30
  );


  not
  g309
  (
    n261,
    n64
  );


  buf
  g310
  (
    n136,
    n89
  );


  buf
  g311
  (
    n172,
    n27
  );


  not
  g312
  (
    n350,
    n42
  );


  buf
  g313
  (
    n232,
    n42
  );


  not
  g314
  (
    n346,
    n89
  );


  not
  g315
  (
    n323,
    n57
  );


  buf
  g316
  (
    n331,
    n35
  );


  not
  g317
  (
    n335,
    n97
  );


  buf
  g318
  (
    n230,
    n37
  );


  not
  g319
  (
    n105,
    n49
  );


  buf
  g320
  (
    n270,
    n58
  );


  not
  g321
  (
    n395,
    n96
  );


  not
  g322
  (
    n308,
    n74
  );


  not
  g323
  (
    n189,
    n82
  );


  buf
  g324
  (
    n365,
    n77
  );


  buf
  g325
  (
    n284,
    n73
  );


  not
  g326
  (
    n208,
    n50
  );


  not
  g327
  (
    n221,
    n98
  );


  buf
  g328
  (
    n374,
    n76
  );


  not
  g329
  (
    KeyWire_0_19,
    n40
  );


  not
  g330
  (
    n206,
    n47
  );


  not
  g331
  (
    n127,
    n90
  );


  buf
  g332
  (
    n137,
    n72
  );


  buf
  g333
  (
    n174,
    n71
  );


  not
  g334
  (
    n408,
    n95
  );


  buf
  g335
  (
    n138,
    n87
  );


  not
  g336
  (
    n292,
    n51
  );


  not
  g337
  (
    n345,
    n42
  );


  buf
  g338
  (
    n344,
    n56
  );


  not
  g339
  (
    n409,
    n81
  );


  not
  g340
  (
    n333,
    n57
  );


  buf
  g341
  (
    n313,
    n30
  );


  buf
  g342
  (
    n222,
    n50
  );


  buf
  g343
  (
    n135,
    n57
  );


  not
  g344
  (
    n289,
    n74
  );


  buf
  g345
  (
    n283,
    n67
  );


  not
  g346
  (
    n225,
    n63
  );


  buf
  g347
  (
    n325,
    n58
  );


  buf
  g348
  (
    n297,
    n57
  );


  not
  g349
  (
    n320,
    n91
  );


  not
  g350
  (
    n359,
    n88
  );


  buf
  g351
  (
    n294,
    n37
  );


  not
  g352
  (
    n245,
    n92
  );


  not
  g353
  (
    n209,
    n35
  );


  not
  g354
  (
    n406,
    n78
  );


  buf
  g355
  (
    n184,
    n69
  );


  buf
  g356
  (
    n312,
    n47
  );


  not
  g357
  (
    n163,
    n94
  );


  buf
  g358
  (
    n386,
    n27
  );


  not
  g359
  (
    n233,
    n61
  );


  buf
  g360
  (
    n254,
    n68
  );


  not
  g361
  (
    n240,
    n80
  );


  buf
  g362
  (
    n103,
    n24
  );


  not
  g363
  (
    n342,
    n83
  );


  buf
  g364
  (
    n356,
    n80
  );


  not
  g365
  (
    n182,
    n65
  );


  buf
  g366
  (
    KeyWire_0_2,
    n81
  );


  not
  g367
  (
    n210,
    n24
  );


  not
  g368
  (
    n207,
    n65
  );


  buf
  g369
  (
    n201,
    n64
  );


  not
  g370
  (
    n281,
    n27
  );


  buf
  g371
  (
    n378,
    n88
  );


  not
  g372
  (
    n293,
    n79
  );


  buf
  g373
  (
    n299,
    n83
  );


  not
  g374
  (
    n393,
    n36
  );


  buf
  g375
  (
    n115,
    n52
  );


  buf
  g376
  (
    n317,
    n76
  );


  not
  g377
  (
    n259,
    n98
  );


  buf
  g378
  (
    n181,
    n67
  );


  buf
  g379
  (
    n315,
    n98
  );


  buf
  g380
  (
    n170,
    n60
  );


  buf
  g381
  (
    n265,
    n53
  );


  not
  g382
  (
    n177,
    n59
  );


  buf
  g383
  (
    n304,
    n69
  );


  not
  g384
  (
    KeyWire_0_15,
    n31
  );


  not
  g385
  (
    n213,
    n84
  );


  not
  g386
  (
    n301,
    n98
  );


  buf
  g387
  (
    n368,
    n49
  );


  buf
  g388
  (
    n157,
    n36
  );


  not
  g389
  (
    n214,
    n76
  );


  not
  g390
  (
    n169,
    n40
  );


  not
  g391
  (
    n106,
    n70
  );


  buf
  g392
  (
    n130,
    n24
  );


  not
  g393
  (
    n595,
    n344
  );


  buf
  g394
  (
    n755,
    n299
  );


  not
  g395
  (
    n976,
    n137
  );


  not
  g396
  (
    n656,
    n104
  );


  buf
  g397
  (
    n953,
    n240
  );


  not
  g398
  (
    n746,
    n141
  );


  not
  g399
  (
    n795,
    n343
  );


  buf
  g400
  (
    n417,
    n240
  );


  not
  g401
  (
    n599,
    n392
  );


  not
  g402
  (
    n788,
    n147
  );


  buf
  g403
  (
    n843,
    n360
  );


  not
  g404
  (
    n845,
    n414
  );


  buf
  g405
  (
    n929,
    n369
  );


  buf
  g406
  (
    n425,
    n199
  );


  buf
  g407
  (
    n512,
    n195
  );


  buf
  g408
  (
    n711,
    n187
  );


  buf
  g409
  (
    n892,
    n109
  );


  buf
  g410
  (
    n522,
    n355
  );


  buf
  g411
  (
    n846,
    n341
  );


  buf
  g412
  (
    n748,
    n205
  );


  buf
  g413
  (
    n446,
    n109
  );


  not
  g414
  (
    n731,
    n337
  );


  not
  g415
  (
    n634,
    n372
  );


  not
  g416
  (
    n692,
    n394
  );


  not
  g417
  (
    n460,
    n289
  );


  buf
  g418
  (
    n822,
    n151
  );


  buf
  g419
  (
    n850,
    n310
  );


  not
  g420
  (
    n604,
    n246
  );


  not
  g421
  (
    n647,
    n152
  );


  not
  g422
  (
    n616,
    n240
  );


  not
  g423
  (
    n859,
    n204
  );


  not
  g424
  (
    n803,
    n170
  );


  buf
  g425
  (
    n801,
    n128
  );


  not
  g426
  (
    n525,
    n413
  );


  not
  g427
  (
    n776,
    n180
  );


  not
  g428
  (
    n532,
    n311
  );


  not
  g429
  (
    n890,
    n168
  );


  not
  g430
  (
    n907,
    n125
  );


  buf
  g431
  (
    n562,
    n387
  );


  buf
  g432
  (
    n452,
    n225
  );


  not
  g433
  (
    n944,
    n150
  );


  buf
  g434
  (
    n538,
    n188
  );


  not
  g435
  (
    n939,
    n355
  );


  buf
  g436
  (
    n879,
    n272
  );


  buf
  g437
  (
    n772,
    n125
  );


  not
  g438
  (
    n897,
    n395
  );


  buf
  g439
  (
    n483,
    n342
  );


  not
  g440
  (
    n543,
    n188
  );


  not
  g441
  (
    n602,
    n353
  );


  buf
  g442
  (
    KeyWire_0_29,
    n210
  );


  buf
  g443
  (
    n927,
    n323
  );


  not
  g444
  (
    n524,
    n187
  );


  not
  g445
  (
    n913,
    n186
  );


  not
  g446
  (
    n793,
    n255
  );


  buf
  g447
  (
    n967,
    n312
  );


  not
  g448
  (
    n520,
    n224
  );


  not
  g449
  (
    n841,
    n336
  );


  buf
  g450
  (
    n499,
    n167
  );


  not
  g451
  (
    n600,
    n384
  );


  buf
  g452
  (
    n671,
    n406
  );


  not
  g453
  (
    n523,
    n204
  );


  buf
  g454
  (
    n441,
    n117
  );


  buf
  g455
  (
    n884,
    n131
  );


  not
  g456
  (
    n477,
    n288
  );


  not
  g457
  (
    n817,
    n302
  );


  not
  g458
  (
    n982,
    n398
  );


  buf
  g459
  (
    n749,
    n174
  );


  buf
  g460
  (
    n730,
    n129
  );


  buf
  g461
  (
    n804,
    n291
  );


  not
  g462
  (
    n536,
    n319
  );


  buf
  g463
  (
    n871,
    n337
  );


  buf
  g464
  (
    n447,
    n356
  );


  buf
  g465
  (
    n639,
    n265
  );


  not
  g466
  (
    n863,
    n141
  );


  buf
  g467
  (
    n422,
    n181
  );


  not
  g468
  (
    n645,
    n223
  );


  buf
  g469
  (
    KeyWire_0_26,
    n120
  );


  buf
  g470
  (
    n509,
    n380
  );


  not
  g471
  (
    n655,
    n202
  );


  not
  g472
  (
    n474,
    n217
  );


  not
  g473
  (
    n805,
    n224
  );


  buf
  g474
  (
    n491,
    n183
  );


  not
  g475
  (
    n440,
    n316
  );


  buf
  g476
  (
    KeyWire_0_22,
    n335
  );


  not
  g477
  (
    n586,
    n200
  );


  buf
  g478
  (
    n830,
    n313
  );


  not
  g479
  (
    n732,
    n376
  );


  not
  g480
  (
    n878,
    n405
  );


  not
  g481
  (
    n838,
    n174
  );


  buf
  g482
  (
    n462,
    n163
  );


  not
  g483
  (
    n624,
    n383
  );


  buf
  g484
  (
    n559,
    n385
  );


  buf
  g485
  (
    n721,
    n279
  );


  not
  g486
  (
    n739,
    n252
  );


  buf
  g487
  (
    n642,
    n225
  );


  not
  g488
  (
    n426,
    n200
  );


  not
  g489
  (
    n613,
    n275
  );


  buf
  g490
  (
    n966,
    n202
  );


  buf
  g491
  (
    n486,
    n400
  );


  buf
  g492
  (
    n676,
    n249
  );


  not
  g493
  (
    n478,
    n148
  );


  buf
  g494
  (
    n635,
    n287
  );


  buf
  g495
  (
    n651,
    n111
  );


  buf
  g496
  (
    n493,
    n175
  );


  not
  g497
  (
    n661,
    n369
  );


  not
  g498
  (
    n521,
    n332
  );


  buf
  g499
  (
    n787,
    n182
  );


  buf
  g500
  (
    n443,
    n301
  );


  buf
  g501
  (
    n556,
    n138
  );


  not
  g502
  (
    n605,
    n262
  );


  buf
  g503
  (
    n880,
    n227
  );


  buf
  g504
  (
    n872,
    n345
  );


  not
  g505
  (
    KeyWire_0_10,
    n303
  );


  buf
  g506
  (
    n720,
    n288
  );


  buf
  g507
  (
    n771,
    n277
  );


  buf
  g508
  (
    n894,
    n301
  );


  buf
  g509
  (
    n529,
    n374
  );


  buf
  g510
  (
    n958,
    n229
  );


  buf
  g511
  (
    n781,
    n404
  );


  buf
  g512
  (
    n620,
    n192
  );


  buf
  g513
  (
    n456,
    n211
  );


  buf
  g514
  (
    n546,
    n218
  );


  not
  g515
  (
    n714,
    n324
  );


  buf
  g516
  (
    n768,
    n180
  );


  buf
  g517
  (
    n684,
    n172
  );


  not
  g518
  (
    n709,
    n121
  );


  not
  g519
  (
    KeyWire_0_6,
    n297
  );


  not
  g520
  (
    n936,
    n149
  );


  buf
  g521
  (
    n835,
    n145
  );


  buf
  g522
  (
    n530,
    n271
  );


  not
  g523
  (
    n954,
    n267
  );


  buf
  g524
  (
    n856,
    n306
  );


  buf
  g525
  (
    n756,
    n323
  );


  buf
  g526
  (
    n517,
    n290
  );


  buf
  g527
  (
    n681,
    n329
  );


  buf
  g528
  (
    n433,
    n119
  );


  buf
  g529
  (
    n449,
    n175
  );


  not
  g530
  (
    n553,
    n110
  );


  buf
  g531
  (
    n834,
    n217
  );


  buf
  g532
  (
    n912,
    n128
  );


  buf
  g533
  (
    n560,
    n249
  );


  not
  g534
  (
    n459,
    n366
  );


  not
  g535
  (
    n971,
    n309
  );


  not
  g536
  (
    n606,
    n168
  );


  not
  g537
  (
    n563,
    n347
  );


  not
  g538
  (
    n572,
    n156
  );


  not
  g539
  (
    n501,
    n204
  );


  not
  g540
  (
    n866,
    n223
  );


  not
  g541
  (
    n507,
    n289
  );


  buf
  g542
  (
    n535,
    n274
  );


  buf
  g543
  (
    n541,
    n377
  );


  buf
  g544
  (
    n923,
    n250
  );


  buf
  g545
  (
    n796,
    n143
  );


  buf
  g546
  (
    n516,
    n260
  );


  not
  g547
  (
    n854,
    n122
  );


  not
  g548
  (
    n767,
    n144
  );


  buf
  g549
  (
    n965,
    n244
  );


  not
  g550
  (
    n906,
    n365
  );


  not
  g551
  (
    n587,
    n279
  );


  buf
  g552
  (
    n695,
    n176
  );


  buf
  g553
  (
    n947,
    n309
  );


  not
  g554
  (
    n663,
    n348
  );


  not
  g555
  (
    n705,
    n190
  );


  buf
  g556
  (
    n421,
    n108
  );


  not
  g557
  (
    n757,
    n407
  );


  buf
  g558
  (
    n473,
    n351
  );


  buf
  g559
  (
    n636,
    n195
  );


  buf
  g560
  (
    n542,
    n411
  );


  not
  g561
  (
    n598,
    n339
  );


  not
  g562
  (
    n860,
    n161
  );


  not
  g563
  (
    n497,
    n261
  );


  buf
  g564
  (
    n930,
    n192
  );


  not
  g565
  (
    n798,
    n219
  );


  buf
  g566
  (
    n931,
    n243
  );


  not
  g567
  (
    n649,
    n166
  );


  buf
  g568
  (
    n775,
    n359
  );


  not
  g569
  (
    n737,
    n388
  );


  not
  g570
  (
    n814,
    n178
  );


  not
  g571
  (
    n554,
    n385
  );


  buf
  g572
  (
    n873,
    n176
  );


  buf
  g573
  (
    n773,
    n195
  );


  buf
  g574
  (
    n902,
    n215
  );


  buf
  g575
  (
    n573,
    n333
  );


  not
  g576
  (
    n899,
    n400
  );


  not
  g577
  (
    n549,
    n173
  );


  not
  g578
  (
    n677,
    n181
  );


  not
  g579
  (
    n833,
    n168
  );


  buf
  g580
  (
    n943,
    n131
  );


  buf
  g581
  (
    n750,
    n401
  );


  not
  g582
  (
    n961,
    n284
  );


  not
  g583
  (
    n534,
    n144
  );


  not
  g584
  (
    n596,
    n220
  );


  not
  g585
  (
    n733,
    n294
  );


  not
  g586
  (
    n933,
    n144
  );


  not
  g587
  (
    n905,
    n293
  );


  not
  g588
  (
    n765,
    n134
  );


  not
  g589
  (
    n463,
    n164
  );


  not
  g590
  (
    n718,
    n170
  );


  not
  g591
  (
    n875,
    n354
  );


  not
  g592
  (
    n972,
    n152
  );


  not
  g593
  (
    n981,
    n313
  );


  not
  g594
  (
    n815,
    n365
  );


  buf
  g595
  (
    n809,
    n207
  );


  not
  g596
  (
    n802,
    n261
  );


  not
  g597
  (
    n742,
    n265
  );


  not
  g598
  (
    n874,
    n268
  );


  not
  g599
  (
    n650,
    n320
  );


  not
  g600
  (
    n691,
    n216
  );


  buf
  g601
  (
    n423,
    n132
  );


  buf
  g602
  (
    n969,
    n221
  );


  buf
  g603
  (
    KeyWire_0_12,
    n362
  );


  not
  g604
  (
    n480,
    n121
  );


  buf
  g605
  (
    n578,
    n140
  );


  not
  g606
  (
    n886,
    n214
  );


  buf
  g607
  (
    n436,
    n305
  );


  not
  g608
  (
    n794,
    n167
  );


  not
  g609
  (
    n697,
    n289
  );


  buf
  g610
  (
    n494,
    n412
  );


  not
  g611
  (
    n919,
    n332
  );


  buf
  g612
  (
    n607,
    n405
  );


  not
  g613
  (
    n825,
    n186
  );


  buf
  g614
  (
    n581,
    n349
  );


  not
  g615
  (
    n618,
    n190
  );


  buf
  g616
  (
    n580,
    n324
  );


  buf
  g617
  (
    n454,
    n360
  );


  buf
  g618
  (
    n896,
    n300
  );


  not
  g619
  (
    n583,
    n290
  );


  not
  g620
  (
    n481,
    n182
  );


  buf
  g621
  (
    n949,
    n371
  );


  buf
  g622
  (
    n511,
    n402
  );


  not
  g623
  (
    n513,
    n341
  );


  not
  g624
  (
    n461,
    n325
  );


  buf
  g625
  (
    n584,
    n196
  );


  buf
  g626
  (
    n882,
    n208
  );


  buf
  g627
  (
    n544,
    n337
  );


  buf
  g628
  (
    n824,
    n148
  );


  buf
  g629
  (
    n565,
    n379
  );


  buf
  g630
  (
    n675,
    n325
  );


  not
  g631
  (
    n774,
    n240
  );


  buf
  g632
  (
    n485,
    n273
  );


  buf
  g633
  (
    n646,
    n134
  );


  not
  g634
  (
    n503,
    n223
  );


  buf
  g635
  (
    n619,
    n288
  );


  buf
  g636
  (
    n657,
    n320
  );


  not
  g637
  (
    n941,
    n314
  );


  buf
  g638
  (
    n608,
    n194
  );


  buf
  g639
  (
    n434,
    n265
  );


  not
  g640
  (
    n782,
    n176
  );


  not
  g641
  (
    n741,
    n271
  );


  not
  g642
  (
    n910,
    n209
  );


  buf
  g643
  (
    n621,
    n118
  );


  not
  g644
  (
    n617,
    n230
  );


  buf
  g645
  (
    n701,
    n183
  );


  not
  g646
  (
    n960,
    n111
  );


  not
  g647
  (
    n592,
    n154
  );


  not
  g648
  (
    n519,
    n318
  );


  not
  g649
  (
    n561,
    n198
  );


  not
  g650
  (
    n625,
    n368
  );


  not
  g651
  (
    n685,
    n121
  );


  not
  g652
  (
    n492,
    n165
  );


  not
  g653
  (
    n622,
    n135
  );


  not
  g654
  (
    n564,
    n410
  );


  buf
  g655
  (
    n557,
    n222
  );


  buf
  g656
  (
    n807,
    n113
  );


  buf
  g657
  (
    n862,
    n330
  );


  not
  g658
  (
    n855,
    n398
  );


  not
  g659
  (
    n527,
    n204
  );


  buf
  g660
  (
    n864,
    n312
  );


  not
  g661
  (
    n764,
    n378
  );


  not
  g662
  (
    n942,
    n198
  );


  not
  g663
  (
    n895,
    n250
  );


  not
  g664
  (
    n921,
    n336
  );


  not
  g665
  (
    n466,
    n340
  );


  not
  g666
  (
    n652,
    n408
  );


  buf
  g667
  (
    n568,
    n335
  );


  not
  g668
  (
    n799,
    n354
  );


  buf
  g669
  (
    n515,
    n363
  );


  buf
  g670
  (
    n766,
    n192
  );


  buf
  g671
  (
    n870,
    n206
  );


  buf
  g672
  (
    n915,
    n141
  );


  not
  g673
  (
    n448,
    n298
  );


  buf
  g674
  (
    n471,
    n140
  );


  buf
  g675
  (
    n811,
    n213
  );


  not
  g676
  (
    n849,
    n370
  );


  not
  g677
  (
    n745,
    n385
  );


  buf
  g678
  (
    n816,
    n401
  );


  buf
  g679
  (
    n743,
    n314
  );


  not
  g680
  (
    n728,
    n283
  );


  not
  g681
  (
    n648,
    n203
  );


  not
  g682
  (
    n713,
    n262
  );


  not
  g683
  (
    n883,
    n330
  );


  not
  g684
  (
    n783,
    n227
  );


  buf
  g685
  (
    n680,
    n275
  );


  buf
  g686
  (
    n679,
    n358
  );


  buf
  g687
  (
    n903,
    n341
  );


  not
  g688
  (
    KeyWire_0_16,
    n253
  );


  buf
  g689
  (
    n893,
    n216
  );


  not
  g690
  (
    n744,
    n331
  );


  buf
  g691
  (
    n428,
    n130
  );


  not
  g692
  (
    n712,
    n321
  );


  buf
  g693
  (
    n490,
    n364
  );


  not
  g694
  (
    n659,
    n305
  );


  not
  g695
  (
    n689,
    n275
  );


  buf
  g696
  (
    n808,
    n225
  );


  buf
  g697
  (
    n540,
    n237
  );


  not
  g698
  (
    n437,
    n189
  );


  buf
  g699
  (
    n666,
    n332
  );


  not
  g700
  (
    n662,
    n232
  );


  not
  g701
  (
    n740,
    n372
  );


  not
  g702
  (
    n653,
    n278
  );


  not
  g703
  (
    n968,
    n281
  );


  not
  g704
  (
    n752,
    n270
  );


  buf
  g705
  (
    n901,
    n316
  );


  not
  g706
  (
    n665,
    n373
  );


  buf
  g707
  (
    n924,
    n212
  );


  buf
  g708
  (
    n416,
    n338
  );


  buf
  g709
  (
    n612,
    n179
  );


  buf
  g710
  (
    n876,
    n199
  );


  buf
  g711
  (
    n690,
    n374
  );


  not
  g712
  (
    n724,
    n291
  );


  buf
  g713
  (
    n597,
    n198
  );


  buf
  g714
  (
    n827,
    n236
  );


  not
  g715
  (
    n570,
    n188
  );


  buf
  g716
  (
    n738,
    n181
  );


  buf
  g717
  (
    n610,
    n207
  );


  buf
  g718
  (
    n955,
    n216
  );


  buf
  g719
  (
    n442,
    n200
  );


  buf
  g720
  (
    n934,
    n406
  );


  not
  g721
  (
    n547,
    n156
  );


  not
  g722
  (
    n790,
    n224
  );


  buf
  g723
  (
    n696,
    n230
  );


  buf
  g724
  (
    n526,
    n392
  );


  buf
  g725
  (
    n498,
    n411
  );


  buf
  g726
  (
    n614,
    n226
  );


  not
  g727
  (
    n900,
    n203
  );


  buf
  g728
  (
    n703,
    n377
  );


  not
  g729
  (
    n668,
    n302
  );


  buf
  g730
  (
    n674,
    n286
  );


  buf
  g731
  (
    n823,
    n389
  );


  not
  g732
  (
    n725,
    n229
  );


  nor
  g733
  (
    n700,
    n353,
    n141
  );


  nor
  g734
  (
    n593,
    n173,
    n122,
    n326,
    n361
  );


  nor
  g735
  (
    n702,
    n292,
    n154,
    n157,
    n311
  );


  nor
  g736
  (
    n747,
    n403,
    n124,
    n135,
    n409
  );


  xnor
  g737
  (
    n577,
    n129,
    n222,
    n348,
    n376
  );


  xnor
  g738
  (
    n820,
    n193,
    n342,
    n201,
    n269
  );


  and
  g739
  (
    n678,
    n381,
    n254,
    n284,
    n142
  );


  xor
  g740
  (
    n888,
    n331,
    n238,
    n250,
    n375
  );


  or
  g741
  (
    n710,
    n400,
    n143,
    n256,
    n136
  );


  nand
  g742
  (
    n418,
    n146,
    n145,
    n343,
    n409
  );


  nor
  g743
  (
    n539,
    n135,
    n154,
    n112,
    n402
  );


  and
  g744
  (
    n687,
    n186,
    n104,
    n210,
    n135
  );


  xnor
  g745
  (
    n667,
    n410,
    n282,
    n222,
    n369
  );


  nand
  g746
  (
    n751,
    n206,
    n383,
    n169,
    n189
  );


  nand
  g747
  (
    n962,
    n320,
    n345,
    n166,
    n177
  );


  xor
  g748
  (
    n427,
    n348,
    n254,
    n184,
    n160
  );


  or
  g749
  (
    n727,
    n286,
    n167,
    n363,
    n368
  );


  nand
  g750
  (
    n925,
    n111,
    n258,
    n167,
    n152
  );


  and
  g751
  (
    n868,
    n307,
    n351,
    n227,
    n359
  );


  or
  g752
  (
    n977,
    n368,
    n234,
    n280,
    n317
  );


  nand
  g753
  (
    n467,
    n196,
    n217,
    n213,
    n118
  );


  xnor
  g754
  (
    KeyWire_0_0,
    n297,
    n190,
    n164,
    n132
  );


  xnor
  g755
  (
    n819,
    n248,
    n229,
    n363,
    n145
  );


  or
  g756
  (
    n877,
    n137,
    n352,
    n337,
    n138
  );


  nand
  g757
  (
    n506,
    n116,
    n144,
    n105,
    n387
  );


  nor
  g758
  (
    n957,
    n342,
    n233,
    n287,
    n259
  );


  and
  g759
  (
    n851,
    n231,
    n357,
    n235,
    n133
  );


  xnor
  g760
  (
    n660,
    n305,
    n119,
    n165,
    n389
  );


  and
  g761
  (
    n630,
    n262,
    n376,
    n110,
    n311
  );


  nand
  g762
  (
    n837,
    n191,
    n257,
    n205,
    n320
  );


  xor
  g763
  (
    n579,
    n391,
    n331,
    n357,
    n397
  );


  xnor
  g764
  (
    n904,
    n268,
    n110,
    n162,
    n399
  );


  nor
  g765
  (
    n555,
    n184,
    n353,
    n276,
    n269
  );


  xnor
  g766
  (
    KeyWire_0_13,
    n336,
    n206,
    n411,
    n286
  );


  or
  g767
  (
    n495,
    n197,
    n114,
    n112,
    n177
  );


  and
  g768
  (
    n853,
    n272,
    n285,
    n279,
    n277
  );


  nand
  g769
  (
    n891,
    n274,
    n257,
    n242,
    n256
  );


  nor
  g770
  (
    n487,
    n301,
    n300,
    n278,
    n282
  );


  or
  g771
  (
    n754,
    n291,
    n328,
    n276,
    n161
  );


  xnor
  g772
  (
    n469,
    n242,
    n398,
    n406,
    n389
  );


  xor
  g773
  (
    n842,
    n128,
    n126,
    n139,
    n181
  );


  nor
  g774
  (
    n429,
    n244,
    n193,
    n407,
    n202
  );


  nor
  g775
  (
    n909,
    n201,
    n383,
    n352,
    n374
  );


  xnor
  g776
  (
    n956,
    n130,
    n105,
    n210,
    n253
  );


  nand
  g777
  (
    n510,
    n399,
    n249,
    n295,
    n235
  );


  and
  g778
  (
    n980,
    n179,
    n148,
    n346,
    n260
  );


  and
  g779
  (
    n935,
    n155,
    n352,
    n304,
    n313
  );


  xnor
  g780
  (
    n979,
    n283,
    n386,
    n323,
    n184
  );


  xor
  g781
  (
    n928,
    n298,
    n407,
    n160,
    n126
  );


  xor
  g782
  (
    n585,
    n367,
    n160,
    n339,
    n262
  );


  nor
  g783
  (
    n566,
    n292,
    n107,
    n127,
    n218
  );


  nand
  g784
  (
    n881,
    n301,
    n244,
    n214,
    n133
  );


  xnor
  g785
  (
    n780,
    n158,
    n162,
    n255,
    n304
  );


  or
  g786
  (
    n812,
    n130,
    n285,
    n178,
    n345
  );


  nand
  g787
  (
    n719,
    n249,
    n340,
    n176,
    n208
  );


  nand
  g788
  (
    n704,
    n390,
    n321,
    n354,
    n118
  );


  xnor
  g789
  (
    n729,
    n137,
    n330,
    n125,
    n377
  );


  xnor
  g790
  (
    n641,
    n399,
    n148,
    n328,
    n278
  );


  or
  g791
  (
    n505,
    n390,
    n239,
    n382,
    n138
  );


  and
  g792
  (
    n445,
    n299,
    n293,
    n109,
    n133
  );


  nand
  g793
  (
    n688,
    n151,
    n150,
    n119,
    n259
  );


  xnor
  g794
  (
    n920,
    n263,
    n338,
    n304,
    n255
  );


  nand
  g795
  (
    n963,
    n149,
    n308,
    n134,
    n236
  );


  or
  g796
  (
    n569,
    n206,
    n146,
    n414,
    n254
  );


  or
  g797
  (
    n672,
    n334,
    n174,
    n252,
    n299
  );


  nand
  g798
  (
    n785,
    n357,
    n348,
    n107,
    n400
  );


  xnor
  g799
  (
    n762,
    n241,
    n120,
    n365,
    n307
  );


  xor
  g800
  (
    n419,
    n366,
    n129,
    n165,
    n325
  );


  nand
  g801
  (
    n430,
    n413,
    n226,
    n157,
    n230
  );


  nor
  g802
  (
    n465,
    n231,
    n316,
    n162,
    n390
  );


  xor
  g803
  (
    n717,
    n139,
    n258,
    n341,
    n392
  );


  xnor
  g804
  (
    n916,
    n389,
    n395,
    n349,
    n280
  );


  nand
  g805
  (
    n686,
    n187,
    n129,
    n350,
    n356
  );


  xnor
  g806
  (
    n528,
    n327,
    n294,
    n260,
    n194
  );


  xor
  g807
  (
    n974,
    n127,
    n310,
    n333,
    n410
  );


  and
  g808
  (
    n821,
    n385,
    n118,
    n178,
    n295
  );


  or
  g809
  (
    n940,
    n152,
    n276,
    n104,
    n395
  );


  nor
  g810
  (
    n488,
    n219,
    n300,
    n396,
    n270
  );


  nor
  g811
  (
    n500,
    n107,
    n381,
    n159,
    n316
  );


  and
  g812
  (
    n951,
    n153,
    n349,
    n340,
    n280
  );


  nor
  g813
  (
    n615,
    n238,
    n133,
    n251,
    n193
  );


  or
  g814
  (
    KeyWire_0_27,
    n153,
    n189,
    n212,
    n374
  );


  nor
  g815
  (
    n898,
    n178,
    n387,
    n221,
    n122
  );


  or
  g816
  (
    n453,
    n309,
    n319,
    n284,
    n237
  );


  or
  g817
  (
    n777,
    n397,
    n201,
    n168,
    n343
  );


  xor
  g818
  (
    n640,
    n234,
    n117,
    n252,
    n138
  );


  xor
  g819
  (
    n699,
    n371,
    n306,
    n169,
    n171
  );


  nor
  g820
  (
    n887,
    n115,
    n336,
    n215,
    n317
  );


  nand
  g821
  (
    n623,
    n283,
    n158,
    n137,
    n246
  );


  xnor
  g822
  (
    n431,
    n386,
    n269,
    n108,
    n199
  );


  or
  g823
  (
    n826,
    n379,
    n248,
    n308,
    n282
  );


  xnor
  g824
  (
    n844,
    n326,
    n319,
    n179,
    n254
  );


  xnor
  g825
  (
    n847,
    n371,
    n322,
    n123,
    n126
  );


  and
  g826
  (
    n818,
    n279,
    n198,
    n180,
    n388
  );


  xnor
  g827
  (
    n937,
    n212,
    n195,
    n300,
    n211
  );


  and
  g828
  (
    n609,
    n143,
    n245,
    n208,
    n232
  );


  xor
  g829
  (
    n482,
    n282,
    n274,
    n366,
    n368
  );


  or
  g830
  (
    n869,
    n219,
    n147,
    n394
  );


  xor
  g831
  (
    n769,
    n131,
    n157,
    n221,
    n216
  );


  or
  g832
  (
    KeyWire_0_4,
    n294,
    n179,
    n115,
    n142
  );


  xor
  g833
  (
    n643,
    n324,
    n315,
    n270,
    n326
  );


  nor
  g834
  (
    n770,
    n390,
    n360,
    n392,
    n303
  );


  nor
  g835
  (
    n551,
    n218,
    n233,
    n378,
    n373
  );


  nand
  g836
  (
    n435,
    n194,
    n393,
    n292,
    n377
  );


  nand
  g837
  (
    n946,
    n330,
    n402,
    n346,
    n303
  );


  and
  g838
  (
    KeyWire_0_24,
    n386,
    n104,
    n384,
    n313
  );


  xor
  g839
  (
    n574,
    n258,
    n409,
    n285,
    n159
  );


  xnor
  g840
  (
    n632,
    n228,
    n171,
    n373,
    n124
  );


  or
  g841
  (
    n914,
    n397,
    n359,
    n238,
    n271
  );


  xor
  g842
  (
    n633,
    n237,
    n356,
    n246,
    n151
  );


  xnor
  g843
  (
    n537,
    n209,
    n406,
    n267,
    n164
  );


  nand
  g844
  (
    n810,
    n308,
    n403,
    n334,
    n295
  );


  xnor
  g845
  (
    n558,
    n113,
    n384,
    n409,
    n404
  );


  xnor
  g846
  (
    n926,
    n334,
    n272,
    n116,
    n259
  );


  and
  g847
  (
    n734,
    n170,
    n231,
    n318,
    n251
  );


  or
  g848
  (
    n760,
    n413,
    n165,
    n207,
    n105
  );


  nand
  g849
  (
    n644,
    n114,
    n369,
    n205,
    n296
  );


  xor
  g850
  (
    n836,
    n365,
    n372,
    n362,
    n109
  );


  xnor
  g851
  (
    n439,
    n245,
    n146,
    n125,
    n218
  );


  or
  g852
  (
    n832,
    n306,
    n224,
    n295,
    n314
  );


  or
  g853
  (
    n464,
    n367,
    n269,
    n344,
    n403
  );


  nand
  g854
  (
    n784,
    n111,
    n250,
    n302,
    n131
  );


  nor
  g855
  (
    n964,
    n222,
    n139,
    n191,
    n386
  );


  nor
  g856
  (
    n858,
    n247,
    n267,
    n291,
    n396
  );


  nor
  g857
  (
    n758,
    n112,
    n172,
    n263,
    n345
  );


  or
  g858
  (
    n590,
    n350,
    n103,
    n286,
    n268
  );


  and
  g859
  (
    n722,
    n331,
    n258,
    n108,
    n373
  );


  xnor
  g860
  (
    n470,
    n332,
    n172,
    n349,
    n382
  );


  xnor
  g861
  (
    KeyWire_0_8,
    n324,
    n264,
    n191,
    n210
  );


  nor
  g862
  (
    n938,
    n209,
    n197,
    n383,
    n134
  );


  and
  g863
  (
    n852,
    n339,
    n335,
    n401,
    n207
  );


  xnor
  g864
  (
    n857,
    n130,
    n346,
    n395,
    n136
  );


  or
  g865
  (
    n654,
    n404,
    n202,
    n410,
    n215
  );


  nand
  g866
  (
    n716,
    n344,
    n347,
    n175,
    n352
  );


  xnor
  g867
  (
    KeyWire_0_7,
    n156,
    n347,
    n333,
    n106
  );


  xnor
  g868
  (
    n628,
    n289,
    n233,
    n298,
    n328
  );


  or
  g869
  (
    n918,
    n237,
    n293,
    n290,
    n278
  );


  or
  g870
  (
    n627,
    n115,
    n115,
    n318,
    n339
  );


  and
  g871
  (
    n839,
    n311,
    n106,
    n239,
    n230
  );


  nor
  g872
  (
    n786,
    n350,
    n214,
    n326,
    n242
  );


  xnor
  g873
  (
    n806,
    n408,
    n266,
    n264,
    n185
  );


  xor
  g874
  (
    n945,
    n120,
    n112,
    n136,
    n402
  );


  or
  g875
  (
    n550,
    n191,
    n247,
    n183,
    n321
  );


  nor
  g876
  (
    n813,
    n177,
    n358,
    n266,
    n264
  );


  or
  g877
  (
    n683,
    n364,
    n246,
    n227,
    n197
  );


  xnor
  g878
  (
    n950,
    n239,
    n394,
    n166,
    n106
  );


  xor
  g879
  (
    n476,
    n266,
    n317,
    n299,
    n412
  );


  xor
  g880
  (
    n753,
    n317,
    n263,
    n208,
    n335
  );


  nand
  g881
  (
    n450,
    n370,
    n347,
    n401,
    n136
  );


  nand
  g882
  (
    n468,
    n413,
    n381,
    n155,
    n143
  );


  nand
  g883
  (
    KeyWire_0_5,
    n244,
    n362,
    n397,
    n182
  );


  xnor
  g884
  (
    n458,
    n151,
    n173,
    n142
  );


  xnor
  g885
  (
    n514,
    n156,
    n261,
    n242,
    n393
  );


  nand
  g886
  (
    n631,
    n243,
    n163,
    n203,
    n312
  );


  xor
  g887
  (
    KeyWire_0_30,
    n213,
    n297,
    n294,
    n281
  );


  nor
  g888
  (
    n438,
    n403,
    n251,
    n388,
    n343
  );


  or
  g889
  (
    n475,
    n399,
    n362,
    n407,
    n162
  );


  xor
  g890
  (
    n693,
    n213,
    n261,
    n371,
    n103
  );


  or
  g891
  (
    n865,
    n217,
    n375,
    n185,
    n103
  );


  nor
  g892
  (
    n789,
    n114,
    n357,
    n236,
    n370
  );


  xor
  g893
  (
    n970,
    n380,
    n351,
    n226,
    n203
  );


  nand
  g894
  (
    n589,
    n253,
    n338,
    n234,
    n361
  );


  or
  g895
  (
    n736,
    n255,
    n232,
    n379,
    n338
  );


  xnor
  g896
  (
    n707,
    n297,
    n307,
    n106,
    n128
  );


  xnor
  g897
  (
    n848,
    n185,
    n404,
    n225,
    n119
  );


  or
  g898
  (
    n588,
    n376,
    n285,
    n277,
    n361
  );


  and
  g899
  (
    n828,
    n284,
    n280,
    n296,
    n241
  );


  nand
  g900
  (
    n601,
    n355,
    n236,
    n342,
    n124
  );


  and
  g901
  (
    n637,
    n363,
    n140,
    n200,
    n328
  );


  xnor
  g902
  (
    n673,
    n197,
    n196,
    n123,
    n205
  );


  nor
  g903
  (
    n424,
    n161,
    n327,
    n108,
    n247
  );


  xor
  g904
  (
    n444,
    n159,
    n238,
    n199,
    n380
  );


  and
  g905
  (
    n567,
    n155,
    n329,
    n303,
    n149
  );


  or
  g906
  (
    n582,
    n170,
    n310,
    n164
  );


  xor
  g907
  (
    n504,
    n378,
    n209,
    n273,
    n358
  );


  nand
  g908
  (
    n792,
    n211,
    n229,
    n354,
    n149
  );


  and
  g909
  (
    n973,
    n274,
    n271,
    n398,
    n215
  );


  and
  g910
  (
    n451,
    n367,
    n192,
    n378,
    n323
  );


  xor
  g911
  (
    n952,
    n248,
    n160,
    n309,
    n396
  );


  xor
  g912
  (
    n831,
    n127,
    n329,
    n340,
    n233
  );


  or
  g913
  (
    n922,
    n302,
    n296,
    n260,
    n105
  );


  nor
  g914
  (
    n706,
    n161,
    n270,
    n325,
    n123
  );


  xor
  g915
  (
    n533,
    n145,
    n315,
    n290,
    n132
  );


  xor
  g916
  (
    n576,
    n408,
    n277,
    n256,
    n321
  );


  nor
  g917
  (
    n885,
    n150,
    n147,
    n186,
    n235
  );


  and
  g918
  (
    n518,
    n201,
    n393,
    n184,
    n350
  );


  nand
  g919
  (
    n591,
    n226,
    n292,
    n116,
    n117
  );


  nor
  g920
  (
    n479,
    n412,
    n267,
    n281,
    n408
  );


  or
  g921
  (
    n603,
    n116,
    n252,
    n391,
    n360
  );


  nor
  g922
  (
    n670,
    n288,
    n312,
    n219,
    n113
  );


  nor
  g923
  (
    n932,
    n187,
    n265,
    n248,
    n361
  );


  xor
  g924
  (
    n457,
    n220,
    n220,
    n327,
    n188
  );


  xor
  g925
  (
    n638,
    n196,
    n172,
    n123,
    n275
  );


  or
  g926
  (
    n759,
    n124,
    n169,
    n245,
    n387
  );


  xnor
  g927
  (
    n682,
    n245,
    n259,
    n257,
    n190
  );


  xor
  g928
  (
    n735,
    n174,
    n314,
    n322,
    n379
  );


  or
  g929
  (
    n552,
    n266,
    n307,
    n358,
    n268
  );


  and
  g930
  (
    n723,
    n110,
    n189,
    n154,
    n158
  );


  xnor
  g931
  (
    n432,
    n120,
    n346,
    n243,
    n329
  );


  nor
  g932
  (
    n797,
    n155,
    n257,
    n241,
    n163
  );


  xnor
  g933
  (
    n484,
    n381,
    n391,
    n251,
    n366
  );


  nor
  g934
  (
    n911,
    n391,
    n194,
    n272,
    n355
  );


  xor
  g935
  (
    n496,
    n393,
    n122,
    n384,
    n214
  );


  or
  g936
  (
    n715,
    n411,
    n211,
    n298,
    n372
  );


  xnor
  g937
  (
    n626,
    n405,
    n241,
    n234,
    n333
  );


  and
  g938
  (
    n545,
    n287,
    n247,
    n114,
    n405
  );


  nand
  g939
  (
    n420,
    n304,
    n334,
    n243,
    n327
  );


  and
  g940
  (
    n840,
    n153,
    n375,
    n107,
    n228
  );


  or
  g941
  (
    n867,
    n359,
    n281,
    n322,
    n344
  );


  and
  g942
  (
    n472,
    n193,
    n153,
    n113,
    n351
  );


  and
  g943
  (
    n889,
    n296,
    n228,
    n305,
    n171
  );


  nand
  g944
  (
    n611,
    n182,
    n169,
    n177,
    n142
  );


  xnor
  g945
  (
    n975,
    n232,
    n367,
    n364,
    n306
  );


  nand
  g946
  (
    n694,
    n253,
    n231,
    n388,
    n382
  );


  or
  g947
  (
    n959,
    n127,
    n322,
    n171,
    n121
  );


  xor
  g948
  (
    n669,
    n380,
    n132,
    n287,
    n228
  );


  nand
  g949
  (
    n791,
    n157,
    n256,
    n396,
    n223
  );


  xnor
  g950
  (
    n594,
    n220,
    n166,
    n319,
    n103
  );


  and
  g951
  (
    n571,
    n180,
    n140,
    n273,
    n158
  );


  xor
  g952
  (
    n548,
    n315,
    n159,
    n212,
    n221
  );


  xnor
  g953
  (
    n779,
    n139,
    n318,
    n273,
    n382
  );


  nand
  g954
  (
    n708,
    n394,
    n163,
    n263,
    n308
  );


  or
  g955
  (
    n664,
    n264,
    n235,
    n239,
    n293
  );


  or
  g956
  (
    n800,
    n370,
    n276,
    n146,
    n183
  );


  xor
  g957
  (
    n829,
    n315,
    n412,
    n126,
    n283
  );


  or
  g958
  (
    n698,
    n375,
    n175,
    n117,
    n353
  );


  nor
  g959
  (
    KeyWire_0_28,
    n364,
    n356,
    n185,
    n150
  );


  or
  g960
  (
    n1038,
    n955,
    n780,
    n775,
    n824
  );


  nand
  g961
  (
    n1039,
    n575,
    n958,
    n937,
    n969
  );


  nand
  g962
  (
    n1106,
    n435,
    n979,
    n541,
    n779
  );


  xor
  g963
  (
    n1020,
    n430,
    n814,
    n884,
    n933
  );


  nand
  g964
  (
    n1128,
    n549,
    n595,
    n606,
    n728
  );


  xnor
  g965
  (
    n989,
    n950,
    n601,
    n838,
    n694
  );


  nand
  g966
  (
    n986,
    n941,
    n972,
    n464,
    n683
  );


  nand
  g967
  (
    n1091,
    n483,
    n669,
    n661,
    n507
  );


  nand
  g968
  (
    n1016,
    n812,
    n960,
    n791,
    n848
  );


  and
  g969
  (
    n1087,
    n949,
    n782,
    n886,
    n658
  );


  and
  g970
  (
    n1078,
    n654,
    n423,
    n722,
    n681
  );


  and
  g971
  (
    n1133,
    n907,
    n751,
    n913,
    n610
  );


  or
  g972
  (
    n1056,
    n512,
    n932,
    n510,
    n973
  );


  and
  g973
  (
    n1082,
    n684,
    n720,
    n905,
    n816
  );


  nand
  g974
  (
    n1129,
    n740,
    n605,
    n571,
    n518
  );


  xor
  g975
  (
    n1044,
    n826,
    n663,
    n493,
    n880
  );


  nand
  g976
  (
    n1041,
    n650,
    n750,
    n528,
    n965
  );


  nor
  g977
  (
    n1123,
    n578,
    n544,
    n673,
    n719
  );


  xor
  g978
  (
    n1024,
    n540,
    n768,
    n707,
    n440
  );


  nand
  g979
  (
    n1034,
    n645,
    n680,
    n439,
    n966
  );


  nand
  g980
  (
    n1006,
    n754,
    n963,
    n830,
    n504
  );


  nor
  g981
  (
    n1131,
    n685,
    n756,
    n662,
    n781
  );


  and
  g982
  (
    n1124,
    n977,
    n919,
    n726,
    n468
  );


  xnor
  g983
  (
    n1107,
    n490,
    n849,
    n752,
    n948
  );


  nor
  g984
  (
    n1042,
    n427,
    n773,
    n498,
    n534
  );


  xnor
  g985
  (
    n1093,
    n944,
    n557,
    n859,
    n724
  );


  nor
  g986
  (
    n1126,
    n618,
    n603,
    n836,
    n817
  );


  xnor
  g987
  (
    n1003,
    n586,
    n545,
    n898,
    n883
  );


  nor
  g988
  (
    n1119,
    n727,
    n699,
    n833,
    n742
  );


  xnor
  g989
  (
    n1132,
    n964,
    n761,
    n629,
    n585
  );


  nor
  g990
  (
    n1100,
    n776,
    n822,
    n441,
    n567
  );


  xor
  g991
  (
    n994,
    n873,
    n644,
    n521,
    n877
  );


  xnor
  g992
  (
    n1009,
    n729,
    n806,
    n745,
    n978
  );


  nor
  g993
  (
    n1014,
    n636,
    n976,
    n454,
    n743
  );


  and
  g994
  (
    n1004,
    n762,
    n890,
    n596,
    n967
  );


  nor
  g995
  (
    n997,
    n592,
    n482,
    n519,
    n712
  );


  xnor
  g996
  (
    n1115,
    n436,
    n967,
    n637,
    n901
  );


  nor
  g997
  (
    n1049,
    n916,
    n979,
    n965,
    n704
  );


  nand
  g998
  (
    n1089,
    n701,
    n677,
    n546,
    n911
  );


  nor
  g999
  (
    n1057,
    n921,
    n472,
    n691,
    n772
  );


  nand
  g1000
  (
    n1092,
    n656,
    n484,
    n867,
    n450
  );


  nand
  g1001
  (
    n1028,
    n803,
    n463,
    n583,
    n887
  );


  nand
  g1002
  (
    n1063,
    n871,
    n897,
    n591,
    n971
  );


  nor
  g1003
  (
    n1053,
    n974,
    n416,
    n912,
    n469
  );


  nand
  g1004
  (
    n1048,
    n796,
    n640,
    n860,
    n703
  );


  xor
  g1005
  (
    n1122,
    n449,
    n421,
    n809,
    n744
  );


  xnor
  g1006
  (
    n1083,
    n485,
    n931,
    n543,
    n470
  );


  or
  g1007
  (
    KeyWire_0_17,
    n539,
    n844,
    n675,
    n456
  );


  xor
  g1008
  (
    n1075,
    n977,
    n778,
    n965,
    n616
  );


  or
  g1009
  (
    n1137,
    n854,
    n879,
    n893,
    n903
  );


  nor
  g1010
  (
    n1055,
    n581,
    n770,
    n730,
    n520
  );


  nand
  g1011
  (
    n1110,
    n488,
    n710,
    n981,
    n757
  );


  xnor
  g1012
  (
    n1086,
    n457,
    n725,
    n466,
    n551
  );


  and
  g1013
  (
    n996,
    n747,
    n532,
    n598,
    n749
  );


  nand
  g1014
  (
    n1007,
    n785,
    n538,
    n638,
    n715
  );


  xor
  g1015
  (
    n1054,
    n968,
    n914,
    n823,
    n553
  );


  nor
  g1016
  (
    n1138,
    n813,
    n706,
    n758,
    n923
  );


  and
  g1017
  (
    n1022,
    n963,
    n529,
    n835,
    n639
  );


  nor
  g1018
  (
    n1021,
    n633,
    n902,
    n786,
    n980
  );


  nand
  g1019
  (
    n1025,
    n494,
    n582,
    n831,
    n760
  );


  nand
  g1020
  (
    n1103,
    n690,
    n966,
    n574,
    n448
  );


  and
  g1021
  (
    n1035,
    n516,
    n827,
    n547,
    n657
  );


  nor
  g1022
  (
    n1023,
    n878,
    n434,
    n970,
    n925
  );


  or
  g1023
  (
    n983,
    n964,
    n489,
    n579,
    n927
  );


  xor
  g1024
  (
    n1012,
    n899,
    n561,
    n939,
    n965
  );


  xnor
  g1025
  (
    n998,
    n620,
    n954,
    n815,
    n968
  );


  or
  g1026
  (
    n1105,
    n787,
    n508,
    n666,
    n970
  );


  xnor
  g1027
  (
    n1011,
    n973,
    n872,
    n802,
    n731
  );


  and
  g1028
  (
    n1095,
    n794,
    n980,
    n614,
    n531
  );


  xor
  g1029
  (
    n1111,
    n537,
    n788,
    n612,
    n709
  );


  nand
  g1030
  (
    n1037,
    n664,
    n972,
    n597,
    n851
  );


  and
  g1031
  (
    n1008,
    n558,
    n453,
    n444,
    n572
  );


  nor
  g1032
  (
    n1118,
    n665,
    n804,
    n623,
    n888
  );


  and
  g1033
  (
    n1001,
    n594,
    n501,
    n820,
    n962
  );


  xor
  g1034
  (
    n1101,
    n974,
    n853,
    n832,
    n511
  );


  nand
  g1035
  (
    n1060,
    n790,
    n964,
    n692,
    n845
  );


  xor
  g1036
  (
    n1017,
    n801,
    n866,
    n792,
    n678
  );


  xor
  g1037
  (
    n1050,
    n805,
    n562,
    n982,
    n978
  );


  nand
  g1038
  (
    n1032,
    n682,
    n713,
    n542,
    n759
  );


  xor
  g1039
  (
    n1070,
    n930,
    n766,
    n837,
    n865
  );


  xor
  g1040
  (
    n1113,
    n896,
    n478,
    n964,
    n940
  );


  xor
  g1041
  (
    n1033,
    n924,
    n975,
    n968,
    n861
  );


  and
  g1042
  (
    n1015,
    n467,
    n789,
    n739,
    n548
  );


  nand
  g1043
  (
    n993,
    n475,
    n563,
    n746,
    n972
  );


  or
  g1044
  (
    n1045,
    n447,
    n573,
    n956,
    n615
  );


  xor
  g1045
  (
    n1108,
    n635,
    n981,
    n741,
    n971
  );


  xnor
  g1046
  (
    n1031,
    n431,
    n695,
    n882,
    n630
  );


  xnor
  g1047
  (
    n1002,
    n868,
    n885,
    n723,
    n978
  );


  nand
  g1048
  (
    n1139,
    n753,
    n696,
    n850,
    n609
  );


  nor
  g1049
  (
    n1084,
    n425,
    n676,
    n588,
    n499
  );


  or
  g1050
  (
    n1030,
    n735,
    n818,
    n980,
    n648
  );


  nor
  g1051
  (
    n1026,
    n671,
    n611,
    n895,
    n975
  );


  or
  g1052
  (
    n1067,
    n840,
    n556,
    n641,
    n651
  );


  or
  g1053
  (
    n1099,
    n559,
    n733,
    n569,
    n771
  );


  xor
  g1054
  (
    n1068,
    n589,
    n855,
    n777,
    n798
  );


  xnor
  g1055
  (
    n1005,
    n973,
    n767,
    n908,
    n474
  );


  nor
  g1056
  (
    n1069,
    n881,
    n917,
    n875,
    n976
  );


  and
  g1057
  (
    n1013,
    n975,
    n736,
    n819,
    n473
  );


  xnor
  g1058
  (
    n1134,
    n433,
    n522,
    n506,
    n961
  );


  xnor
  g1059
  (
    n1097,
    n672,
    n446,
    n535,
    n580
  );


  nand
  g1060
  (
    n1010,
    n689,
    n846,
    n647,
    n734
  );


  and
  g1061
  (
    n1094,
    n763,
    n442,
    n769,
    n705
  );


  xnor
  g1062
  (
    n985,
    n962,
    n934,
    n870,
    n688
  );


  nor
  g1063
  (
    n1018,
    n622,
    n513,
    n967,
    n462
  );


  xnor
  g1064
  (
    n1114,
    n514,
    n617,
    n492,
    n619
  );


  nand
  g1065
  (
    n1058,
    n653,
    n634,
    n936,
    n452
  );


  or
  g1066
  (
    n1000,
    n797,
    n564,
    n968,
    n977
  );


  nor
  g1067
  (
    n1130,
    n418,
    n910,
    n714,
    n643
  );


  xnor
  g1068
  (
    n1079,
    n503,
    n975,
    n477,
    n969
  );


  and
  g1069
  (
    n992,
    n500,
    n811,
    n737,
    n976
  );


  nand
  g1070
  (
    n1098,
    n807,
    n497,
    n970,
    n821
  );


  and
  g1071
  (
    n1073,
    n828,
    n947,
    n981,
    n738
  );


  xor
  g1072
  (
    n1102,
    n560,
    n938,
    n847,
    n668
  );


  xnor
  g1073
  (
    n999,
    n892,
    n979,
    n566,
    n445
  );


  xor
  g1074
  (
    n1047,
    n957,
    n697,
    n889,
    n834
  );


  or
  g1075
  (
    n991,
    n945,
    n667,
    n509,
    n718
  );


  or
  g1076
  (
    n1109,
    n642,
    n825,
    n981,
    n795
  );


  and
  g1077
  (
    n1027,
    n602,
    n891,
    n920,
    n783
  );


  xor
  g1078
  (
    n1046,
    n732,
    n977,
    n550,
    n979
  );


  xnor
  g1079
  (
    n1085,
    n967,
    n460,
    n496,
    n451
  );


  xnor
  g1080
  (
    n1076,
    n533,
    n784,
    n852,
    n829
  );


  xnor
  g1081
  (
    n1062,
    n962,
    n842,
    n590,
    n570
  );


  xnor
  g1082
  (
    n1125,
    n922,
    n659,
    n443,
    n686
  );


  xnor
  g1083
  (
    n1061,
    n963,
    n869,
    n523,
    n461
  );


  xnor
  g1084
  (
    n1127,
    n915,
    n765,
    n874,
    n693
  );


  xnor
  g1085
  (
    n1120,
    n437,
    n621,
    n943,
    n465
  );


  nor
  g1086
  (
    n1036,
    n717,
    n978,
    n679,
    n942
  );


  or
  g1087
  (
    n1065,
    n670,
    n593,
    n970,
    n702
  );


  nor
  g1088
  (
    n1052,
    n458,
    n455,
    n929,
    n505
  );


  nor
  g1089
  (
    n1090,
    n774,
    n980,
    n649,
    n959
  );


  nor
  g1090
  (
    n1104,
    n565,
    n530,
    n969,
    n608
  );


  nand
  g1091
  (
    n1040,
    n721,
    n841,
    n480,
    n487
  );


  and
  g1092
  (
    n1136,
    n515,
    n971,
    n536,
    n417
  );


  nand
  g1093
  (
    n1112,
    n904,
    n962,
    n843,
    n502
  );


  nor
  g1094
  (
    n1117,
    n876,
    n525,
    n491,
    n517
  );


  or
  g1095
  (
    n1077,
    n632,
    n864,
    n576,
    n972
  );


  and
  g1096
  (
    n984,
    n625,
    n856,
    n613,
    n607
  );


  or
  g1097
  (
    n1116,
    n428,
    n974,
    n476,
    n963
  );


  nand
  g1098
  (
    n987,
    n422,
    n584,
    n863,
    n587
  );


  or
  g1099
  (
    n1135,
    n894,
    n900,
    n966,
    n793
  );


  and
  g1100
  (
    n1081,
    n626,
    n527,
    n858,
    n432
  );


  nor
  g1101
  (
    n1096,
    n600,
    n652,
    n526,
    n935
  );


  or
  g1102
  (
    n1071,
    n909,
    n624,
    n687,
    n486
  );


  xor
  g1103
  (
    n1121,
    n926,
    n764,
    n808,
    n946
  );


  xnor
  g1104
  (
    n1064,
    n426,
    n604,
    n552,
    n599
  );


  and
  g1105
  (
    n1080,
    n700,
    n471,
    n424,
    n438
  );


  or
  g1106
  (
    n1072,
    n631,
    n419,
    n479,
    n524
  );


  nor
  g1107
  (
    n1029,
    n660,
    n973,
    n906,
    n971
  );


  and
  g1108
  (
    n1066,
    n568,
    n674,
    n862,
    n716
  );


  and
  g1109
  (
    n995,
    n800,
    n708,
    n918,
    n755
  );


  nand
  g1110
  (
    n1043,
    n420,
    n495,
    n982,
    n969
  );


  xnor
  g1111
  (
    n1074,
    n974,
    n839,
    n655,
    n698
  );


  or
  g1112
  (
    n1051,
    n966,
    n481,
    n810,
    n627
  );


  nor
  g1113
  (
    n1059,
    n748,
    n646,
    n953,
    n429
  );


  and
  g1114
  (
    n1019,
    n799,
    n952,
    n857,
    n577
  );


  nor
  g1115
  (
    n988,
    n628,
    n459,
    n951,
    n711
  );


  or
  g1116
  (
    n990,
    n554,
    n976,
    n928,
    n555
  );


  not
  g1117
  (
    n1170,
    n1001
  );


  buf
  g1118
  (
    n1162,
    n1124
  );


  not
  g1119
  (
    n1173,
    n1026
  );


  not
  g1120
  (
    n1159,
    n1076
  );


  buf
  g1121
  (
    n1231,
    n1115
  );


  buf
  g1122
  (
    n1148,
    n1134
  );


  not
  g1123
  (
    n1230,
    n1009
  );


  not
  g1124
  (
    n1186,
    n1052
  );


  buf
  g1125
  (
    n1169,
    n1128
  );


  not
  g1126
  (
    n1259,
    n990
  );


  buf
  g1127
  (
    n1166,
    n1124
  );


  buf
  g1128
  (
    n1226,
    n1120
  );


  buf
  g1129
  (
    n1165,
    n1043
  );


  buf
  g1130
  (
    n1156,
    n1090
  );


  not
  g1131
  (
    n1207,
    n1088
  );


  not
  g1132
  (
    n1176,
    n1116
  );


  buf
  g1133
  (
    n1233,
    n1103
  );


  buf
  g1134
  (
    n1228,
    n1111
  );


  buf
  g1135
  (
    n1179,
    n1080
  );


  not
  g1136
  (
    n1189,
    n1065
  );


  not
  g1137
  (
    n1172,
    n1123
  );


  not
  g1138
  (
    n1155,
    n1133
  );


  not
  g1139
  (
    n1224,
    n1081
  );


  not
  g1140
  (
    n1193,
    n1024
  );


  not
  g1141
  (
    n1229,
    n1139
  );


  not
  g1142
  (
    n1145,
    n1115
  );


  not
  g1143
  (
    n1249,
    n1036
  );


  buf
  g1144
  (
    n1171,
    n1012
  );


  buf
  g1145
  (
    n1214,
    n1015
  );


  not
  g1146
  (
    n1158,
    n1122
  );


  not
  g1147
  (
    n1164,
    n1028
  );


  not
  g1148
  (
    n1185,
    n1132
  );


  not
  g1149
  (
    n1160,
    n1098
  );


  buf
  g1150
  (
    n1178,
    n984
  );


  buf
  g1151
  (
    n1199,
    n1058
  );


  buf
  g1152
  (
    n1246,
    n983
  );


  not
  g1153
  (
    n1237,
    n1048
  );


  not
  g1154
  (
    n1146,
    n1027
  );


  not
  g1155
  (
    n1152,
    n1139
  );


  buf
  g1156
  (
    n1167,
    n1137
  );


  buf
  g1157
  (
    n1206,
    n1018
  );


  not
  g1158
  (
    n1168,
    n1046
  );


  not
  g1159
  (
    n1143,
    n1135
  );


  buf
  g1160
  (
    n1250,
    n989
  );


  not
  g1161
  (
    n1217,
    n1072
  );


  buf
  g1162
  (
    n1157,
    n1138
  );


  not
  g1163
  (
    n1212,
    n1111
  );


  not
  g1164
  (
    n1204,
    n1086
  );


  buf
  g1165
  (
    n1208,
    n1135
  );


  not
  g1166
  (
    n1256,
    n1134
  );


  buf
  g1167
  (
    n1209,
    n1040
  );


  not
  g1168
  (
    n1253,
    n1084
  );


  buf
  g1169
  (
    n1175,
    n1112
  );


  not
  g1170
  (
    n1195,
    n1139
  );


  not
  g1171
  (
    n1177,
    n1127
  );


  buf
  g1172
  (
    n1235,
    n1078
  );


  not
  g1173
  (
    n1234,
    n1131
  );


  not
  g1174
  (
    n1187,
    n1126
  );


  not
  g1175
  (
    n1221,
    n1124
  );


  not
  g1176
  (
    n1254,
    n1074
  );


  not
  g1177
  (
    n1190,
    n1091
  );


  not
  g1178
  (
    n1241,
    n1070
  );


  not
  g1179
  (
    n1184,
    n1032
  );


  not
  g1180
  (
    n1258,
    n1095
  );


  buf
  g1181
  (
    n1205,
    n1130
  );


  buf
  g1182
  (
    n1174,
    n1119
  );


  not
  g1183
  (
    n1257,
    n1123
  );


  buf
  g1184
  (
    n1180,
    n1139
  );


  buf
  g1185
  (
    n1201,
    n1118
  );


  buf
  g1186
  (
    n1192,
    n1115
  );


  buf
  g1187
  (
    n1202,
    n1016
  );


  buf
  g1188
  (
    n1163,
    n1128
  );


  buf
  g1189
  (
    n1151,
    n1117
  );


  buf
  g1190
  (
    n1218,
    n998
  );


  not
  g1191
  (
    n1194,
    n1121
  );


  buf
  g1192
  (
    n1222,
    n1017
  );


  not
  g1193
  (
    n1227,
    n1075
  );


  not
  g1194
  (
    n1239,
    n1120
  );


  not
  g1195
  (
    n1188,
    n1000
  );


  not
  g1196
  (
    n1255,
    n1059
  );


  nor
  g1197
  (
    n1150,
    n1093,
    n1127,
    n1117,
    n1096
  );


  xor
  g1198
  (
    n1248,
    n1044,
    n1113,
    n1083,
    n1051
  );


  nand
  g1199
  (
    n1240,
    n1137,
    n997,
    n1131,
    n1006
  );


  xnor
  g1200
  (
    n1238,
    n1069,
    n1113,
    n1066,
    n1132
  );


  nand
  g1201
  (
    n1183,
    n1124,
    n1094,
    n1039,
    n1112
  );


  xor
  g1202
  (
    n1191,
    n1119,
    n1008,
    n1138,
    n1041
  );


  or
  g1203
  (
    n1232,
    n1120,
    n1061,
    n1129,
    n1114
  );


  and
  g1204
  (
    n1225,
    n1104,
    n1120,
    n1056,
    n1129
  );


  xor
  g1205
  (
    n1245,
    n1136,
    n1109,
    n1053,
    n1073
  );


  xnor
  g1206
  (
    n1210,
    n1025,
    n1127,
    n1121,
    n1114
  );


  xnor
  g1207
  (
    KeyWire_0_23,
    n1116,
    n1047,
    n991,
    n1107
  );


  and
  g1208
  (
    n1252,
    n1005,
    n995,
    n1100,
    n1019
  );


  nand
  g1209
  (
    n1182,
    n1127,
    n1108,
    n1020,
    n1099
  );


  nand
  g1210
  (
    n1236,
    n1119,
    n1014,
    n1125,
    n1114
  );


  nand
  g1211
  (
    n1144,
    n1087,
    n1133,
    n1138,
    n1063
  );


  nor
  g1212
  (
    n1215,
    n1038,
    n1117,
    n1057,
    n1004
  );


  and
  g1213
  (
    n1200,
    n1064,
    n1034,
    n1030,
    n1102
  );


  nor
  g1214
  (
    n1220,
    n1126,
    n1060,
    n1055,
    n1092
  );


  xor
  g1215
  (
    n1223,
    n1136,
    n1054,
    n1116,
    n1118
  );


  nand
  g1216
  (
    n1149,
    n1089,
    n1129,
    n993,
    n985
  );


  and
  g1217
  (
    n1244,
    n1113,
    n986,
    n1133,
    n1125
  );


  nor
  g1218
  (
    n1251,
    n1114,
    n1132,
    n1126
  );


  xor
  g1219
  (
    n1161,
    n1128,
    n1101,
    n1077,
    n1116
  );


  and
  g1220
  (
    n1154,
    n1122,
    n1136,
    n1013,
    n1045
  );


  nand
  g1221
  (
    n1142,
    n1135,
    n1130,
    n1022,
    n1021
  );


  nand
  g1222
  (
    n1243,
    n1105,
    n1130,
    n1033,
    n1125
  );


  xor
  g1223
  (
    n1219,
    n1126,
    n1085,
    n1106,
    n1135
  );


  xor
  g1224
  (
    n1198,
    n1023,
    n1118,
    n1079,
    n1037
  );


  nor
  g1225
  (
    n1147,
    n1123,
    n1067,
    n1134,
    n1118
  );


  or
  g1226
  (
    n1196,
    n1131,
    n1136,
    n1003,
    n1113
  );


  and
  g1227
  (
    n1213,
    n992,
    n1082,
    n1121,
    n1122
  );


  xor
  g1228
  (
    n1216,
    n1133,
    n1002,
    n1119,
    n988
  );


  nand
  g1229
  (
    n1153,
    n1138,
    n1117,
    n994,
    n1031
  );


  nor
  g1230
  (
    n1141,
    n1129,
    n1115,
    n1137,
    n996
  );


  xnor
  g1231
  (
    n1242,
    n1121,
    n1137,
    n1128,
    n1007
  );


  xnor
  g1232
  (
    n1181,
    n1049,
    n1123,
    n1071,
    n1042
  );


  nor
  g1233
  (
    n1197,
    n1122,
    n1134,
    n1050,
    n1125
  );


  or
  g1234
  (
    n1203,
    n1131,
    n987,
    n1011,
    n1062
  );


  nand
  g1235
  (
    n1211,
    n1010,
    n999,
    n1029,
    n1068
  );


  nor
  g1236
  (
    n1247,
    n1130,
    n1097,
    n1110,
    n1035
  );


  and
  g1237
  (
    n1271,
    n1188,
    n1161
  );


  nand
  g1238
  (
    n1270,
    n1190,
    n1222,
    n1164,
    n1180
  );


  nand
  g1239
  (
    n1272,
    n1143,
    n1165,
    n1212,
    n1226
  );


  xnor
  g1240
  (
    n1269,
    n1229,
    n1241,
    n1202,
    n1249
  );


  or
  g1241
  (
    n1265,
    n1174,
    n1197,
    n1173,
    n1178
  );


  xnor
  g1242
  (
    n1263,
    n1232,
    n1237,
    n1230,
    n1218
  );


  xor
  g1243
  (
    n1276,
    n1169,
    n1141,
    n1170,
    n1167
  );


  or
  g1244
  (
    n1291,
    n1244,
    n1228,
    n1242,
    n1231
  );


  and
  g1245
  (
    n1274,
    n1181,
    n1171,
    n1149,
    n1177
  );


  xnor
  g1246
  (
    n1288,
    n1193,
    n1259,
    n1223,
    n1203
  );


  nand
  g1247
  (
    n1268,
    n1146,
    n1240,
    n1205,
    n1182
  );


  xor
  g1248
  (
    n1266,
    n1186,
    n1259,
    n1215,
    n1191
  );


  xnor
  g1249
  (
    n1280,
    n1211,
    n1142,
    n1199,
    n1243
  );


  and
  g1250
  (
    n1264,
    n1185,
    n1145,
    n1227,
    n1162
  );


  and
  g1251
  (
    n1287,
    n1158,
    n1201,
    n1166,
    n1250
  );


  and
  g1252
  (
    n1281,
    n1156,
    n1152,
    n1213,
    n1256
  );


  and
  g1253
  (
    n1289,
    n1183,
    n1209,
    n1224,
    n1208
  );


  xor
  g1254
  (
    n1286,
    n101,
    n1238,
    n1163,
    n1258
  );


  nand
  g1255
  (
    n1275,
    n1159,
    n1168,
    n1154,
    n1259
  );


  xor
  g1256
  (
    n1283,
    n1247,
    n1179,
    n1189,
    n1140
  );


  xor
  g1257
  (
    n1261,
    n1216,
    n1210,
    n1148,
    n1239
  );


  or
  g1258
  (
    n1279,
    n1144,
    n101,
    n1245,
    n1151
  );


  xnor
  g1259
  (
    n1284,
    n1204,
    n1225,
    n1253,
    n1257
  );


  xor
  g1260
  (
    n1285,
    n1220,
    n1252,
    n1175,
    n1206
  );


  and
  g1261
  (
    n1277,
    n1236,
    n1219,
    n1217,
    n1176
  );


  nor
  g1262
  (
    n1262,
    n1194,
    n1195,
    n1172,
    n1150
  );


  nand
  g1263
  (
    n1273,
    n1214,
    n1192,
    n1155,
    n1248
  );


  nand
  g1264
  (
    n1278,
    n1184,
    n1196,
    n1255,
    n1147
  );


  nand
  g1265
  (
    n1290,
    n1187,
    n1254,
    n1198,
    n1234
  );


  xnor
  g1266
  (
    n1282,
    n1200,
    n1207,
    n1160,
    n1235
  );


  nand
  g1267
  (
    n1260,
    n1251,
    n1221,
    n1246,
    n1157
  );


  and
  g1268
  (
    n1267,
    n1233,
    n1153,
    n1259,
    n101
  );


  buf
  g1269
  (
    n1297,
    n1282
  );


  not
  g1270
  (
    n1300,
    n1286
  );


  not
  g1271
  (
    n1293,
    n1283
  );


  not
  g1272
  (
    n1294,
    n1285
  );


  buf
  g1273
  (
    n1292,
    n1284
  );


  not
  g1274
  (
    n1298,
    n1288
  );


  buf
  g1275
  (
    n1301,
    n1287
  );


  buf
  g1276
  (
    n1299,
    n1289
  );


  not
  g1277
  (
    n1295,
    n1291
  );


  not
  g1278
  (
    n1296,
    n1290
  );


  not
  g1279
  (
    n1315,
    n1293
  );


  not
  g1280
  (
    n1310,
    n1297
  );


  not
  g1281
  (
    n1307,
    n1297
  );


  buf
  g1282
  (
    n1311,
    n1298
  );


  not
  g1283
  (
    n1306,
    n1297
  );


  not
  g1284
  (
    n1313,
    n1296
  );


  not
  g1285
  (
    n1314,
    n1294
  );


  buf
  g1286
  (
    n1309,
    n1296
  );


  buf
  g1287
  (
    n1312,
    n1292
  );


  not
  g1288
  (
    n1302,
    n1298
  );


  buf
  g1289
  (
    n1304,
    n1298
  );


  buf
  g1290
  (
    n1308,
    n1297
  );


  buf
  g1291
  (
    n1305,
    n1299
  );


  buf
  g1292
  (
    n1316,
    n1295
  );


  not
  g1293
  (
    n1303,
    n1299
  );


  buf
  g1294
  (
    n1317,
    n1298
  );


  buf
  g1295
  (
    n1319,
    n1302
  );


  buf
  g1296
  (
    n1320,
    n1305
  );


  not
  g1297
  (
    n1323,
    n1305
  );


  not
  g1298
  (
    n1321,
    n1305
  );


  buf
  g1299
  (
    n1322,
    n1303
  );


  buf
  g1300
  (
    n1318,
    n1304
  );


  not
  g1301
  (
    n1335,
    n1322
  );


  buf
  g1302
  (
    n1325,
    n1307
  );


  not
  g1303
  (
    KeyWire_0_20,
    n1306
  );


  not
  g1304
  (
    n1340,
    n1307
  );


  not
  g1305
  (
    n1339,
    n1308
  );


  buf
  g1306
  (
    n1328,
    n1322
  );


  buf
  g1307
  (
    n1332,
    n1318
  );


  buf
  g1308
  (
    n1324,
    n1320
  );


  and
  g1309
  (
    n1330,
    n415,
    n1309,
    n414,
    n1308
  );


  nor
  g1310
  (
    n1331,
    n1300,
    n1306,
    n1323,
    n1322
  );


  and
  g1311
  (
    n1326,
    n415,
    n21,
    n1321,
    n1306
  );


  nor
  g1312
  (
    n1334,
    n1318,
    n1319,
    n1300,
    n1321
  );


  xor
  g1313
  (
    n1337,
    n1320,
    n415,
    n1321
  );


  xnor
  g1314
  (
    n1329,
    n1319,
    n1321,
    n1323,
    n1318
  );


  nand
  g1315
  (
    n1338,
    n1308,
    n1320,
    n1306,
    n1319
  );


  xor
  g1316
  (
    n1333,
    n1299,
    n1323,
    n1318
  );


  nand
  g1317
  (
    n1327,
    n1307,
    n414,
    n1322,
    n1309
  );


  nor
  g1318
  (
    n1342,
    n1320,
    n21,
    n1308,
    n1307
  );


  xor
  g1319
  (
    n1336,
    n1299,
    n1305,
    n1319,
    n21
  );


  xor
  g1320
  (
    n1360,
    n1334,
    n1331,
    n1328
  );


  nand
  g1321
  (
    n1350,
    n1326,
    n1328,
    n1337,
    n1327
  );


  xor
  g1322
  (
    n1359,
    n1309,
    n1326,
    n1325,
    n1336
  );


  nor
  g1323
  (
    n1352,
    n1342,
    n1333,
    n1310,
    n1326
  );


  xnor
  g1324
  (
    n1347,
    n1342,
    n1329,
    n1333,
    n1331
  );


  nor
  g1325
  (
    n1362,
    n1336,
    n1339,
    n1328,
    n1334
  );


  nand
  g1326
  (
    n1344,
    n1332,
    n1337,
    n1328,
    n1340
  );


  nand
  g1327
  (
    n1353,
    n1340,
    n1310,
    n1341,
    n1339
  );


  xnor
  g1328
  (
    n1343,
    n1311,
    n1341,
    n1310,
    n1339
  );


  xor
  g1329
  (
    n1351,
    n1335,
    n1311,
    n1334,
    n1327
  );


  and
  g1330
  (
    n1354,
    n1309,
    n1337,
    n1329,
    n1335
  );


  nand
  g1331
  (
    n1349,
    n1333,
    n1330,
    n1327,
    n1332
  );


  xnor
  g1332
  (
    n1357,
    n1336,
    n1330,
    n1342,
    n1338
  );


  nor
  g1333
  (
    n1346,
    n1336,
    n1338,
    n1327,
    n1329
  );


  or
  g1334
  (
    n1345,
    n1335,
    n1340,
    n1334,
    n1339
  );


  nor
  g1335
  (
    n1356,
    n1337,
    n1331,
    n1341,
    n1310
  );


  and
  g1336
  (
    n1355,
    n1329,
    n1330,
    n1332,
    n1341
  );


  xnor
  g1337
  (
    KeyWire_0_18,
    n1326,
    n1324,
    n1311,
    n1335
  );


  or
  g1338
  (
    n1361,
    n1330,
    n1332,
    n1338
  );


  xnor
  g1339
  (
    n1348,
    n1311,
    n1340,
    n1333,
    n1342
  );


  buf
  g1340
  (
    n1366,
    n1350
  );


  buf
  g1341
  (
    n1363,
    n1343
  );


  not
  g1342
  (
    n1372,
    n1345
  );


  not
  g1343
  (
    n1365,
    n1351
  );


  buf
  g1344
  (
    n1364,
    n1347
  );


  buf
  g1345
  (
    n1369,
    n1348
  );


  buf
  g1346
  (
    n1367,
    n1354
  );


  not
  g1347
  (
    n1368,
    n1346
  );


  and
  g1348
  (
    n1370,
    n1344,
    n1353
  );


  nand
  g1349
  (
    n1371,
    n1352,
    n1349
  );


  xnor
  g1350
  (
    n1373,
    n1365,
    n1367,
    n1364,
    n1366
  );


  nor
  g1351
  (
    n1374,
    n1366,
    n1366,
    n1365,
    n1367
  );


  or
  g1352
  (
    n1376,
    n1363,
    n1365,
    n1364
  );


  xor
  g1353
  (
    n1375,
    n1364,
    n1364,
    n1366,
    n1367
  );


  nand
  g1354
  (
    n1379,
    n1376,
    n1355
  );


  or
  g1355
  (
    n1385,
    n22,
    n982,
    n1313
  );


  xor
  g1356
  (
    n1384,
    n22,
    n1313
  );


  xor
  g1357
  (
    n1382,
    n1375,
    n1312,
    n1376
  );


  xnor
  g1358
  (
    n1377,
    n1373,
    n1374,
    n1314
  );


  and
  g1359
  (
    n1383,
    n22,
    n1313,
    n982
  );


  xnor
  g1360
  (
    n1381,
    n1355,
    n1312,
    n21
  );


  and
  g1361
  (
    n1378,
    n22,
    n1314,
    n1376,
    n1375
  );


  xor
  g1362
  (
    n1380,
    n1355,
    n1312,
    n1374,
    n1376
  );


  nand
  g1363
  (
    n1395,
    n1368,
    n1356,
    n1315,
    n1371
  );


  or
  g1364
  (
    n1407,
    n1300,
    n1377,
    n102,
    n1357
  );


  nand
  g1365
  (
    n1399,
    n1359,
    n1301,
    n1370,
    n1385
  );


  nor
  g1366
  (
    n1398,
    n1383,
    n102,
    n1384,
    n1380
  );


  nand
  g1367
  (
    n1401,
    n1371,
    n1315,
    n1381,
    n1385
  );


  nand
  g1368
  (
    n1406,
    n1368,
    n1357,
    n1378,
    n1371
  );


  xor
  g1369
  (
    n1402,
    n1384,
    n1385,
    n1378,
    n1357
  );


  nor
  g1370
  (
    n1397,
    n1358,
    n1357,
    n1316,
    n1377
  );


  xor
  g1371
  (
    n1391,
    n1380,
    n1371,
    n1370,
    n1359
  );


  xnor
  g1372
  (
    n1408,
    n1383,
    n1381,
    n1300,
    n1369
  );


  nand
  g1373
  (
    n1392,
    n1316,
    n1383,
    n1369,
    n1370
  );


  nor
  g1374
  (
    n1394,
    n1368,
    n1301,
    n1372,
    n1358
  );


  or
  g1375
  (
    n1387,
    n1368,
    n1379,
    n1384,
    n102
  );


  or
  g1376
  (
    n1388,
    n1382,
    n1356,
    n1369
  );


  and
  g1377
  (
    n1389,
    n1358,
    n1316,
    n1378
  );


  and
  g1378
  (
    n1400,
    n1381,
    n1301,
    n1378
  );


  and
  g1379
  (
    n1390,
    n1385,
    n1380,
    n1382,
    n1315
  );


  and
  g1380
  (
    n1393,
    n1367,
    n1315,
    n1356,
    n1314
  );


  xnor
  g1381
  (
    n1386,
    n1380,
    n1379,
    n1372,
    n102
  );


  xor
  g1382
  (
    n1396,
    n1370,
    n1379,
    n1372,
    n1382
  );


  nor
  g1383
  (
    n1404,
    n1314,
    n1369,
    n1372,
    n1358
  );


  or
  g1384
  (
    KeyWire_0_9,
    n1379,
    n1359,
    n1384,
    n1383
  );


  nor
  g1385
  (
    n1405,
    n1377,
    n1377,
    n1381,
    n1382
  );


  xnor
  g1386
  (
    n1418,
    n1407,
    n1317,
    n1359,
    n1395
  );


  or
  g1387
  (
    n1417,
    n1317,
    n1391,
    n1401,
    n1386
  );


  xor
  g1388
  (
    n1416,
    n1399,
    n1362,
    n1390,
    n1398
  );


  xnor
  g1389
  (
    n1412,
    n1361,
    n1360,
    n1362
  );


  or
  g1390
  (
    n1415,
    n1362,
    n1396,
    n1408,
    n1317
  );


  xor
  g1391
  (
    n1413,
    n1397,
    n1406,
    n1362,
    n1388
  );


  xor
  g1392
  (
    n1414,
    n1392,
    n1402,
    n1361
  );


  or
  g1393
  (
    n1411,
    n1389,
    n1403,
    n1360
  );


  or
  g1394
  (
    n1409,
    n1400,
    n1393,
    n1361,
    n1405
  );


  and
  g1395
  (
    n1410,
    n1394,
    n1387,
    n1404,
    n1317
  );


  xor
  KeyGate_0_0
  (
    n575,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n122,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n196,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n256,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n726,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n948,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n778,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n629,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n761,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1403,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n978,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n328,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n658,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n861,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n45,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n357,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n917,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1088,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1358,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n318,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1341,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n116,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n502,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n1140,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n489,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n227,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n455,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n531,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n908,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n508,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n763,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n70,
    KeyNOTWire_0_31
  );


endmodule

