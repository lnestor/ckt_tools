// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_153 written by SynthGen on 2021/04/05 11:08:34
module Stat_1000_153( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1004, n991, n988, n990, n992, n995, n1005, n1010,
 n987, n1009, n996, n1014, n994, n1012, n989, n1008,
 n1001, n1015, n1013, n1017, n998, n1019, n1007, n993,
 n1011, n1018, n1020, n1022, n1024, n1025, n1032, n1031);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1004, n991, n988, n990, n992, n995, n1005, n1010,
 n987, n1009, n996, n1014, n994, n1012, n989, n1008,
 n1001, n1015, n1013, n1017, n998, n1019, n1007, n993,
 n1011, n1018, n1020, n1022, n1024, n1025, n1032, n1031;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n997, n999, n1000, n1002, n1003, n1006,
 n1016, n1021, n1023, n1026, n1027, n1028, n1029, n1030;

buf  g0 (n108, n17);
buf  g1 (n40, n23);
buf  g2 (n139, n11);
buf  g3 (n36, n9);
not  g4 (n126, n14);
buf  g5 (n54, n20);
buf  g6 (n85, n3);
not  g7 (n98, n20);
buf  g8 (n34, n4);
not  g9 (n128, n7);
not  g10 (n41, n5);
buf  g11 (n71, n26);
buf  g12 (n148, n10);
buf  g13 (n152, n29);
buf  g14 (n47, n25);
buf  g15 (n63, n24);
buf  g16 (n94, n23);
not  g17 (n107, n30);
not  g18 (n33, n13);
buf  g19 (n127, n14);
not  g20 (n142, n5);
not  g21 (n84, n21);
not  g22 (n109, n21);
buf  g23 (n104, n6);
not  g24 (n42, n21);
buf  g25 (n61, n15);
not  g26 (n100, n9);
not  g27 (n120, n20);
not  g28 (n66, n15);
buf  g29 (n86, n6);
buf  g30 (n87, n12);
not  g31 (n133, n3);
not  g32 (n93, n25);
not  g33 (n44, n19);
buf  g34 (n48, n14);
not  g35 (n143, n16);
buf  g36 (n39, n1);
not  g37 (n82, n19);
buf  g38 (n130, n7);
buf  g39 (n81, n17);
not  g40 (n96, n31);
buf  g41 (n146, n9);
buf  g42 (n149, n16);
buf  g43 (n125, n14);
not  g44 (n45, n9);
not  g45 (n80, n16);
buf  g46 (n118, n5);
not  g47 (n60, n7);
buf  g48 (n52, n2);
not  g49 (n132, n16);
not  g50 (n70, n15);
buf  g51 (n90, n10);
buf  g52 (n105, n29);
not  g53 (n151, n27);
buf  g54 (n123, n31);
buf  g55 (n131, n22);
buf  g56 (n53, n1);
buf  g57 (n67, n19);
buf  g58 (n88, n17);
not  g59 (n141, n29);
not  g60 (n113, n11);
not  g61 (n116, n13);
not  g62 (n137, n24);
buf  g63 (n62, n26);
buf  g64 (n49, n19);
buf  g65 (n124, n30);
not  g66 (n57, n22);
buf  g67 (n144, n23);
buf  g68 (n35, n30);
not  g69 (n46, n4);
buf  g70 (n112, n8);
buf  g71 (n77, n12);
not  g72 (n64, n28);
not  g73 (n83, n18);
not  g74 (n135, n8);
buf  g75 (n145, n13);
buf  g76 (n99, n18);
not  g77 (n37, n4);
not  g78 (n69, n20);
buf  g79 (n68, n31);
buf  g80 (n122, n22);
buf  g81 (n89, n7);
buf  g82 (n138, n6);
buf  g83 (n72, n8);
buf  g84 (n121, n30);
not  g85 (n91, n4);
not  g86 (n140, n21);
not  g87 (n101, n26);
not  g88 (n103, n3);
not  g89 (n58, n1);
buf  g90 (n43, n18);
buf  g91 (n136, n25);
buf  g92 (n97, n11);
buf  g93 (n129, n12);
buf  g94 (n117, n26);
buf  g95 (n55, n11);
not  g96 (n38, n8);
not  g97 (n119, n2);
buf  g98 (n92, n5);
buf  g99 (n65, n23);
not  g100 (n147, n24);
not  g101 (n111, n6);
buf  g102 (n56, n10);
not  g103 (n74, n15);
buf  g104 (n51, n28);
not  g105 (n114, n27);
not  g106 (n106, n18);
buf  g107 (n102, n10);
not  g108 (n110, n28);
buf  g109 (n73, n29);
buf  g110 (n79, n12);
buf  g111 (n150, n17);
buf  g112 (n59, n28);
not  g113 (n134, n27);
not  g114 (n115, n24);
not  g115 (n75, n13);
not  g116 (n95, n22);
buf  g117 (n76, n25);
buf  g118 (n78, n27);
not  g119 (n50, n2);
not  g120 (n291, n56);
not  g121 (n327, n33);
buf  g122 (n233, n40);
buf  g123 (n303, n34);
buf  g124 (n219, n63);
buf  g125 (n260, n37);
buf  g126 (n302, n56);
buf  g127 (n316, n46);
not  g128 (n189, n35);
buf  g129 (n325, n52);
buf  g130 (n211, n73);
not  g131 (n156, n73);
buf  g132 (n162, n46);
not  g133 (n193, n62);
buf  g134 (n235, n38);
buf  g135 (n241, n70);
not  g136 (n209, n47);
buf  g137 (n246, n56);
not  g138 (n312, n40);
buf  g139 (n252, n56);
not  g140 (n282, n69);
not  g141 (n185, n76);
buf  g142 (n247, n54);
not  g143 (n216, n42);
buf  g144 (n323, n64);
not  g145 (n250, n50);
not  g146 (n321, n65);
not  g147 (n191, n45);
not  g148 (n256, n50);
buf  g149 (n217, n71);
not  g150 (n164, n47);
not  g151 (n244, n51);
buf  g152 (n227, n53);
not  g153 (n163, n57);
not  g154 (n290, n75);
not  g155 (n236, n59);
not  g156 (n218, n72);
not  g157 (n175, n51);
not  g158 (n172, n37);
not  g159 (n157, n68);
buf  g160 (n258, n67);
buf  g161 (n155, n36);
buf  g162 (n311, n50);
buf  g163 (n269, n53);
buf  g164 (n285, n48);
buf  g165 (n314, n52);
buf  g166 (n309, n68);
not  g167 (n170, n62);
buf  g168 (n226, n48);
buf  g169 (n153, n37);
not  g170 (n243, n49);
not  g171 (n300, n35);
not  g172 (n166, n63);
buf  g173 (n293, n55);
buf  g174 (n232, n41);
buf  g175 (n313, n76);
not  g176 (n305, n38);
not  g177 (n186, n73);
not  g178 (n284, n36);
buf  g179 (n304, n68);
buf  g180 (n322, n75);
buf  g181 (n263, n74);
buf  g182 (n173, n52);
not  g183 (n165, n49);
not  g184 (n265, n53);
not  g185 (n274, n61);
not  g186 (n308, n48);
not  g187 (n229, n58);
buf  g188 (n295, n66);
not  g189 (n206, n74);
buf  g190 (n286, n51);
not  g191 (n188, n35);
not  g192 (n329, n63);
buf  g193 (n196, n63);
buf  g194 (n179, n45);
buf  g195 (n177, n33);
buf  g196 (n223, n41);
not  g197 (n181, n46);
buf  g198 (n264, n75);
buf  g199 (n254, n36);
buf  g200 (n310, n35);
buf  g201 (n301, n70);
buf  g202 (n326, n55);
not  g203 (n272, n62);
not  g204 (n294, n57);
not  g205 (n180, n61);
buf  g206 (n242, n61);
buf  g207 (n195, n37);
not  g208 (n281, n34);
not  g209 (n324, n36);
not  g210 (n200, n44);
not  g211 (n187, n42);
buf  g212 (n296, n38);
not  g213 (n237, n38);
buf  g214 (n292, n54);
buf  g215 (n255, n76);
not  g216 (n280, n66);
buf  g217 (n205, n45);
not  g218 (n299, n43);
buf  g219 (n184, n57);
not  g220 (n202, n71);
buf  g221 (n198, n48);
buf  g222 (n262, n65);
not  g223 (n270, n44);
not  g224 (n306, n46);
buf  g225 (n214, n70);
not  g226 (n231, n72);
not  g227 (n251, n39);
buf  g228 (n288, n42);
buf  g229 (n176, n77);
buf  g230 (n277, n53);
buf  g231 (n230, n62);
not  g232 (n275, n64);
buf  g233 (n317, n33);
not  g234 (n192, n59);
not  g235 (n276, n58);
buf  g236 (n319, n42);
not  g237 (n183, n45);
not  g238 (n215, n68);
buf  g239 (n154, n73);
buf  g240 (n210, n41);
buf  g241 (n182, n52);
buf  g242 (n289, n41);
not  g243 (n208, n71);
not  g244 (n160, n69);
buf  g245 (n174, n44);
not  g246 (n261, n71);
buf  g247 (n167, n43);
not  g248 (n224, n47);
not  g249 (n178, n49);
buf  g250 (n245, n47);
buf  g251 (n161, n39);
not  g252 (n328, n65);
buf  g253 (n213, n61);
not  g254 (n225, n39);
buf  g255 (n234, n39);
buf  g256 (n283, n74);
buf  g257 (n253, n34);
not  g258 (n279, n72);
buf  g259 (n320, n51);
buf  g260 (n257, n57);
buf  g261 (n239, n34);
buf  g262 (n228, n65);
buf  g263 (n220, n59);
buf  g264 (n287, n43);
not  g265 (n197, n58);
not  g266 (n240, n70);
buf  g267 (n297, n60);
not  g268 (n271, n66);
buf  g269 (n199, n64);
buf  g270 (n273, n49);
not  g271 (n158, n50);
buf  g272 (n318, n66);
buf  g273 (n278, n69);
buf  g274 (n204, n76);
buf  g275 (n203, n58);
not  g276 (n159, n75);
buf  g277 (n267, n55);
buf  g278 (n268, n72);
buf  g279 (n307, n69);
not  g280 (n201, n59);
not  g281 (n207, n55);
not  g282 (n222, n74);
not  g283 (n315, n40);
buf  g284 (n194, n33);
buf  g285 (n190, n60);
buf  g286 (n238, n67);
buf  g287 (n248, n60);
not  g288 (n249, n54);
not  g289 (n259, n67);
buf  g290 (n221, n67);
not  g291 (n212, n43);
buf  g292 (n298, n40);
buf  g293 (n168, n60);
buf  g294 (n266, n54);
buf  g295 (n171, n64);
buf  g296 (n169, n44);
not  g297 (n519, n220);
buf  g298 (n476, n322);
not  g299 (n345, n227);
not  g300 (n516, n189);
buf  g301 (n405, n290);
buf  g302 (n397, n307);
not  g303 (n420, n303);
not  g304 (n391, n265);
buf  g305 (n571, n262);
not  g306 (n555, n266);
buf  g307 (n562, n279);
buf  g308 (n483, n274);
buf  g309 (n374, n183);
buf  g310 (n347, n160);
not  g311 (n379, n254);
buf  g312 (n518, n286);
buf  g313 (n498, n164);
buf  g314 (n487, n191);
not  g315 (n552, n203);
buf  g316 (n439, n82);
buf  g317 (n400, n313);
not  g318 (n526, n235);
buf  g319 (n393, n313);
buf  g320 (n425, n168);
not  g321 (n448, n288);
not  g322 (n422, n274);
buf  g323 (n511, n199);
not  g324 (n560, n169);
buf  g325 (n394, n252);
buf  g326 (n433, n292);
buf  g327 (n482, n247);
buf  g328 (n428, n200);
not  g329 (n427, n154);
not  g330 (n356, n234);
not  g331 (n340, n218);
not  g332 (n419, n318);
buf  g333 (n387, n266);
buf  g334 (n543, n325);
buf  g335 (n554, n79);
not  g336 (n401, n306);
buf  g337 (n495, n296);
not  g338 (n556, n300);
buf  g339 (n354, n222);
not  g340 (n375, n261);
buf  g341 (n463, n294);
not  g342 (n440, n154);
buf  g343 (n453, n301);
not  g344 (n462, n189);
buf  g345 (n536, n291);
not  g346 (n538, n267);
not  g347 (n565, n168);
buf  g348 (n456, n232);
not  g349 (n540, n82);
not  g350 (n435, n298);
not  g351 (n352, n295);
buf  g352 (n344, n277);
buf  g353 (n521, n276);
buf  g354 (n541, n304);
not  g355 (n572, n223);
buf  g356 (n468, n320);
not  g357 (n331, n299);
not  g358 (n548, n260);
not  g359 (n492, n264);
not  g360 (n535, n239);
not  g361 (n349, n296);
not  g362 (n359, n218);
not  g363 (n389, n210);
not  g364 (n549, n188);
buf  g365 (n564, n317);
not  g366 (n402, n246);
not  g367 (n355, n77);
buf  g368 (n348, n214);
not  g369 (n525, n294);
buf  g370 (n574, n204);
buf  g371 (n496, n282);
buf  g372 (n413, n316);
not  g373 (n534, n299);
buf  g374 (n503, n296);
not  g375 (n467, n239);
not  g376 (n418, n209);
buf  g377 (n371, n166);
buf  g378 (n406, n288);
buf  g379 (n442, n177);
not  g380 (n411, n267);
not  g381 (n542, n302);
not  g382 (n522, n272);
buf  g383 (n444, n271);
buf  g384 (n415, n303);
not  g385 (n514, n324);
not  g386 (n508, n277);
not  g387 (n458, n255);
not  g388 (n491, n292);
buf  g389 (n424, n228);
not  g390 (n373, n187);
not  g391 (n333, n195);
not  g392 (n421, n273);
buf  g393 (n545, n325);
buf  g394 (n550, n309);
buf  g395 (n377, n300);
buf  g396 (n409, n78);
buf  g397 (n489, n246);
not  g398 (n475, n207);
not  g399 (n523, n259);
not  g400 (n396, n315);
not  g401 (n416, n298);
not  g402 (n384, n236);
not  g403 (n392, n322);
buf  g404 (n423, n309);
not  g405 (n484, n291);
not  g406 (n513, n221);
buf  g407 (n461, n219);
not  g408 (n412, n193);
buf  g409 (n343, n271);
not  g410 (n459, n165);
not  g411 (n460, n305);
buf  g412 (n517, n170);
not  g413 (n330, n157);
not  g414 (n366, n264);
not  g415 (n553, n268);
not  g416 (n529, n318);
not  g417 (n378, n323);
not  g418 (n507, n81);
not  g419 (n465, n187);
buf  g420 (n395, n160);
buf  g421 (n334, n259);
buf  g422 (n474, n257);
not  g423 (n557, n246);
not  g424 (n342, n269);
buf  g425 (n382, n224);
not  g426 (n490, n194);
buf  g427 (n341, n170);
buf  g428 (n486, n190);
not  g429 (n500, n78);
not  g430 (n504, n242);
buf  g431 (n501, n202);
buf  g432 (n417, n242);
buf  g433 (n469, n310);
not  g434 (n568, n299);
buf  g435 (n376, n198);
not  g436 (n351, n223);
buf  g437 (n505, n240);
not  g438 (n558, n248);
not  g439 (n403, n196);
not  g440 (n383, n311);
not  g441 (n559, n317);
buf  g442 (n499, n272);
not  g443 (n451, n270);
buf  g444 (n528, n286);
xor  g445 (n436, n295, n282);
and  g446 (n502, n290, n263, n302, n307);
nand g447 (n365, n181, n153, n278, n155);
nor  g448 (n477, n83, n245, n215, n180);
and  g449 (n539, n297, n283, n313, n236);
nor  g450 (n357, n277, n202, n249, n78);
nor  g451 (n480, n316, n305, n297, n269);
or   g452 (n446, n208, n214, n273, n321);
or   g453 (n399, n323, n285, n312, n294);
xor  g454 (n338, n283, n295, n176, n196);
nor  g455 (n404, n269, n226, n186, n212);
or   g456 (n488, n288, n296, n317, n251);
or   g457 (n443, n216, n324, n182, n79);
nor  g458 (n367, n321, n173, n279, n250);
xnor g459 (n429, n260, n285, n175, n259);
or   g460 (n370, n306, n181, n158, n263);
and  g461 (n431, n258, n291, n203, n235);
nand g462 (n390, n311, n219, n251, n276);
nand g463 (n533, n247, n184, n193, n228);
or   g464 (n547, n294, n284, n314, n216);
or   g465 (n524, n254, n307, n268, n303);
xor  g466 (n455, n276, n178, n255, n308);
and  g467 (n509, n258, n210, n261, n243);
or   g468 (n479, n270, n81, n293, n302);
and  g469 (n454, n318, n317, n319, n284);
and  g470 (n407, n275, n211, n174, n213);
xnor g471 (n364, n234, n322, n199, n251);
xor  g472 (n358, n310, n323, n250, n185);
nand g473 (n532, n229, n278, n287, n163);
nand g474 (n493, n311, n265, n263, n171);
xnor g475 (n449, n319, n320, n162, n293);
nor  g476 (n481, n293, n309, n180, n253);
or   g477 (n437, n325, n245, n237, n82);
nor  g478 (n438, n271, n287, n300, n265);
xor  g479 (n464, n278, n253, n262, n306);
and  g480 (n512, n191, n291, n255, n252);
nand g481 (n339, n184, n221, n268, n204);
and  g482 (n473, n194, n78, n289, n224);
nand g483 (n527, n307, n249, n217, n175);
nor  g484 (n494, n232, n246, n308, n230);
xor  g485 (n472, n258, n325, n312, n226);
or   g486 (n398, n179, n249, n188, n222);
nor  g487 (n369, n82, n273, n304, n233);
nor  g488 (n537, n192, n164, n79, n283);
nor  g489 (n381, n310, n304, n270, n79);
or   g490 (n506, n281, n297, n306, n282);
or   g491 (n388, n314, n285, n161, n230);
nor  g492 (n368, n295, n81, n257, n270);
xor  g493 (n569, n272, n323, n250, n286);
or   g494 (n441, n261, n83, n256, n299);
and  g495 (n361, n266, n280, n319, n315);
or   g496 (n497, n269, n243, n183, n309);
and  g497 (n567, n217, n192, n279, n247);
and  g498 (n386, n312, n254, n206, n205);
xnor g499 (n573, n162, n205, n267, n238);
or   g500 (n466, n318, n182, n215, n167);
xor  g501 (n337, n247, n157, n301, n195);
nor  g502 (n563, n253, n271, n206, n283);
nand g503 (n531, n281, n256, n166, n304);
or   g504 (n510, n158, n301, n163, n197);
or   g505 (n372, n240, n264, n248, n281);
xor  g506 (n434, n263, n171, n290, n314);
xnor g507 (n350, n298, n80, n177, n268);
or   g508 (n362, n256, n179, n305, n253);
xor  g509 (n546, n77, n297, n290, n316);
and  g510 (n457, n282, n261, n185, n280);
nand g511 (n426, n190, n287, n314, n264);
or   g512 (n385, n213, n267, n159, n81);
and  g513 (n478, n178, n275, n249, n197);
nor  g514 (n551, n244, n324, n308, n156);
xnor g515 (n408, n227, n259, n319, n153);
and  g516 (n335, n172, n159, n280, n208);
nor  g517 (n353, n167, n200, n315, n322);
xor  g518 (n515, n279, n275, n265, n284);
or   g519 (n450, n320, n252, n241, n251);
and  g520 (n380, n315, n165, n161, n237);
and  g521 (n430, n198, n155, n241, n245);
or   g522 (n544, n281, n209, n248, n257);
nor  g523 (n447, n320, n258, n186, n248);
nand g524 (n346, n276, n274, n289, n312);
or   g525 (n410, n176, n316, n284, n254);
nand g526 (n470, n308, n300, n288, n231);
xor  g527 (n414, n262, n156, n321, n225);
and  g528 (n432, n313, n238, n273, n174);
and  g529 (n520, n292, n278, n262, n287);
xnor g530 (n452, n289, n274, n303, n201);
nor  g531 (n530, n77, n266, n301, n260);
xor  g532 (n336, n244, n83, n321, n277);
or   g533 (n360, n293, n220, n280, n286);
and  g534 (n471, n311, n80, n298, n229);
xnor g535 (n445, n289, n256, n207, n250);
or   g536 (n561, n275, n272, n305, n245);
nand g537 (n485, n173, n302, n255, n80);
nor  g538 (n566, n324, n201, n260, n80);
nand g539 (n570, n169, n225, n285, n257);
or   g540 (n332, n233, n252, n172, n231);
nor  g541 (n363, n212, n211, n310, n292);
buf  g542 (n635, n360);
buf  g543 (n584, n384);
buf  g544 (n620, n380);
not  g545 (n631, n389);
buf  g546 (n597, n346);
buf  g547 (n610, n377);
not  g548 (n578, n393);
not  g549 (n608, n333);
buf  g550 (n590, n368);
not  g551 (n607, n334);
not  g552 (n602, n379);
buf  g553 (n595, n330);
not  g554 (n592, n371);
buf  g555 (n589, n349);
not  g556 (n626, n359);
not  g557 (n624, n372);
buf  g558 (n616, n373);
not  g559 (n579, n352);
not  g560 (n600, n358);
buf  g561 (n614, n344);
buf  g562 (n606, n388);
not  g563 (n588, n347);
not  g564 (n605, n362);
buf  g565 (n632, n331);
not  g566 (n638, n361);
not  g567 (n599, n375);
buf  g568 (n612, n381);
not  g569 (n630, n338);
not  g570 (n634, n351);
buf  g571 (n586, n365);
not  g572 (n625, n386);
not  g573 (n576, n363);
buf  g574 (n598, n383);
not  g575 (n617, n336);
buf  g576 (n596, n376);
buf  g577 (n637, n355);
buf  g578 (n583, n335);
not  g579 (n636, n369);
not  g580 (n581, n392);
not  g581 (n613, n366);
buf  g582 (n619, n354);
not  g583 (n627, n345);
buf  g584 (n615, n337);
buf  g585 (n580, n356);
buf  g586 (n601, n350);
buf  g587 (n633, n348);
not  g588 (n594, n364);
buf  g589 (n593, n339);
buf  g590 (n621, n341);
not  g591 (n587, n374);
not  g592 (n628, n343);
buf  g593 (n577, n370);
buf  g594 (n591, n357);
buf  g595 (n604, n387);
not  g596 (n575, n340);
buf  g597 (n618, n353);
buf  g598 (n609, n378);
buf  g599 (n603, n391);
buf  g600 (n611, n390);
buf  g601 (n582, n382);
not  g602 (n585, n342);
buf  g603 (n622, n367);
not  g604 (n629, n385);
buf  g605 (n623, n332);
or   g606 (n643, n469, n584);
and  g607 (n662, n467, n406, n499, n416);
xor  g608 (n677, n577, n585, n578, n441);
xor  g609 (n651, n517, n408, n581, n491);
or   g610 (n676, n493, n395, n494, n409);
xor  g611 (n639, n421, n453, n470, n579);
nand g612 (n647, n457, n412, n446, n497);
and  g613 (n640, n584, n437, n580, n521);
xnor g614 (n660, n503, n581, n508, n468);
xor  g615 (n671, n501, n496, n460, n576);
and  g616 (n667, n450, n403, n415, n397);
and  g617 (n670, n523, n433, n476, n413);
nor  g618 (n658, n514, n522, n473, n455);
xor  g619 (n650, n502, n480, n579, n581);
or   g620 (n661, n575, n513, n492, n444);
or   g621 (n656, n472, n509, n580, n479);
nand g622 (n675, n424, n405, n442, n581);
nor  g623 (n668, n586, n434, n454, n578);
and  g624 (n665, n448, n486, n582, n427);
xnor g625 (n646, n440, n422, n520, n585);
xor  g626 (n681, n498, n584, n426, n474);
xor  g627 (n652, n483, n585, n582, n402);
nand g628 (n655, n583, n425, n580, n459);
nand g629 (n679, n414, n515, n394, n429);
xnor g630 (n644, n586, n464, n435, n452);
nor  g631 (n678, n505, n458, n439, n478);
nand g632 (n663, n461, n506, n485, n579);
nor  g633 (n674, n420, n451, n575, n510);
or   g634 (n664, n576, n511, n518, n577);
xnor g635 (n645, n585, n430, n436, n431);
xnor g636 (n654, n418, n404, n399, n456);
nand g637 (n682, n417, n583, n481, n423);
and  g638 (n669, n471, n487, n443, n578);
xnor g639 (n672, n577, n512, n576, n438);
or   g640 (n680, n407, n462, n584, n477);
nand g641 (n659, n504, n400, n580, n583);
nor  g642 (n653, n495, n582, n445, n432);
or   g643 (n649, n419, n447, n582, n583);
nand g644 (n642, n484, n475, n579, n428);
and  g645 (n666, n488, n578, n482, n489);
nor  g646 (n648, n396, n500, n516, n465);
nand g647 (n657, n519, n449, n401, n411);
xor  g648 (n673, n463, n466, n507, n490);
xnor g649 (n641, n575, n410, n398, n577);
xnor g650 (n693, n629, n621, n627, n607);
xnor g651 (n690, n88, n588, n631, n93);
nor  g652 (n725, n587, n603, n681, n628);
xor  g653 (n685, n657, n624, n609, n663);
nor  g654 (n747, n670, n587, n88, n86);
or   g655 (n717, n596, n613, n622, n611);
and  g656 (n754, n525, n617, n603, n622);
and  g657 (n759, n605, n637, n675, n594);
xor  g658 (n756, n604, n96, n631, n635);
or   g659 (n692, n604, n593, n587, n616);
xnor g660 (n694, n592, n594, n85);
nand g661 (n689, n606, n679, n603, n93);
and  g662 (n684, n644, n653, n595, n651);
nand g663 (n738, n598, n93, n607, n591);
or   g664 (n696, n606, n591, n94, n587);
nand g665 (n723, n592, n643, n636, n590);
xnor g666 (n757, n619, n615, n654, n86);
xnor g667 (n760, n660, n590, n602, n623);
or   g668 (n710, n593, n629, n661, n588);
nor  g669 (n709, n93, n91, n597);
nor  g670 (n708, n679, n92, n88, n610);
and  g671 (n722, n660, n634, n90, n627);
and  g672 (n711, n599, n624, n597, n623);
or   g673 (n700, n662, n597, n97, n589);
nor  g674 (n719, n671, n681, n632, n611);
xnor g675 (n765, n674, n640, n614, n88);
nand g676 (n727, n649, n601, n592, n607);
xor  g677 (n745, n594, n618, n605);
and  g678 (n713, n608, n600, n603, n590);
nor  g679 (n712, n608, n621, n596, n84);
xnor g680 (n720, n592, n90, n658, n87);
nand g681 (n763, n616, n624, n595, n610);
xnor g682 (n751, n677, n90, n675, n602);
or   g683 (n715, n682, n84, n646, n680);
nor  g684 (n691, n613, n666, n655, n625);
or   g685 (n770, n640, n662, n86, n621);
and  g686 (n766, n89, n614, n672, n616);
xnor g687 (n737, n664, n87, n639, n629);
and  g688 (n698, n665, n615, n668, n651);
nor  g689 (n743, n586, n635, n598, n605);
xnor g690 (n721, n666, n682, n627, n626);
and  g691 (n686, n669, n671, n524, n599);
or   g692 (n697, n604, n596, n622, n94);
nand g693 (n705, n602, n673, n664, n649);
or   g694 (n687, n613, n634, n657, n648);
and  g695 (n731, n620, n627, n631, n594);
xnor g696 (n706, n614, n623, n631, n630);
xnor g697 (n724, n605, n680, n616, n619);
xor  g698 (n702, n85, n95, n87, n633);
nor  g699 (n740, n635, n91, n673, n90);
xor  g700 (n703, n621, n644, n628, n611);
nand g701 (n750, n632, n614, n647, n600);
nand g702 (n729, n95, n628, n647, n615);
or   g703 (n758, n637, n593, n591, n588);
nand g704 (n714, n643, n609, n650, n639);
nand g705 (n716, n630, n674, n611, n89);
xor  g706 (n739, n648, n658, n94, n625);
xnor g707 (n707, n628, n676, n608, n597);
and  g708 (n768, n615, n610, n677, n618);
nand g709 (n683, n642, n91, n676, n89);
and  g710 (n762, n604, n656, n601, n620);
nor  g711 (n755, n590, n617, n596, n645);
xor  g712 (n733, n595, n625, n600, n652);
and  g713 (n732, n618, n667, n665, n642);
xor  g714 (n726, n85, n96, n669, n617);
xor  g715 (n704, n613, n632, n593, n620);
or   g716 (n753, n622, n624, n84, n87);
nand g717 (n748, n600, n650, n92, n653);
nor  g718 (n695, n89, n645, n670, n598);
or   g719 (n761, n608, n678, n652, n667);
and  g720 (n746, n94, n96, n609, n655);
and  g721 (n764, n599, n626, n659, n617);
nand g722 (n742, n610, n663, n620, n601);
and  g723 (n718, n634, n635, n612, n591);
xor  g724 (n688, n606, n661, n612, n630);
nand g725 (n730, n659, n589, n92, n602);
nor  g726 (n734, n95, n84, n619, n641);
or   g727 (n741, n633, n601, n632, n612);
nand g728 (n767, n625, n656, n86, n646);
xnor g729 (n744, n678, n641, n607, n634);
xor  g730 (n728, n629, n619, n96, n83);
or   g731 (n769, n95, n92, n588, n595);
xor  g732 (n699, n626, n589, n668, n609);
or   g733 (n736, n636, n598, n599, n672);
xnor g734 (n752, n589, n633, n637);
or   g735 (n749, n606, n626, n97, n612);
xnor g736 (n701, n636, n586, n633, n630);
xnor g737 (n735, n623, n97, n654, n636);
and  g738 (n849, n720, n735, n756, n721);
xnor g739 (n773, n124, n739, n106, n756);
and  g740 (n861, n733, n108, n140, n750);
nand g741 (n800, n138, n754, n740, n103);
xnor g742 (n822, n707, n730, n755, n749);
xnor g743 (n825, n121, n140, n128, n722);
nor  g744 (n821, n692, n105, n757, n117);
xnor g745 (n791, n101, n709, n737, n722);
xor  g746 (n854, n715, n98, n104, n118);
or   g747 (n788, n683, n107, n726, n757);
and  g748 (n840, n120, n693, n140, n133);
xor  g749 (n864, n704, n749, n119, n103);
or   g750 (n806, n705, n121, n130, n748);
xor  g751 (n789, n103, n106, n132, n700);
and  g752 (n792, n704, n145, n111, n703);
nor  g753 (n834, n119, n735, n716, n743);
and  g754 (n809, n123, n762, n711, n769);
xnor g755 (n829, n752, n762, n694, n120);
and  g756 (n855, n110, n738, n142, n766);
xor  g757 (n823, n114, n683, n142, n689);
nor  g758 (n814, n133, n746, n144, n103);
xor  g759 (n799, n131, n709, n729, n759);
and  g760 (n803, n730, n765, n713, n685);
or   g761 (n815, n134, n133, n110, n144);
xor  g762 (n862, n747, n723, n99, n126);
xor  g763 (n782, n723, n718, n748, n125);
and  g764 (n816, n100, n135, n766, n687);
xor  g765 (n836, n131, n144, n696, n684);
and  g766 (n824, n695, n143, n741);
xor  g767 (n796, n770, n761, n727, n714);
xor  g768 (n798, n684, n768, n132, n114);
xor  g769 (n801, n108, n726, n146, n757);
xor  g770 (n843, n690, n736, n105, n145);
xnor g771 (n784, n689, n692, n98, n115);
and  g772 (n802, n764, n99, n751, n118);
nor  g773 (n812, n135, n128, n143, n132);
or   g774 (n851, n715, n751, n97, n755);
nor  g775 (n804, n729, n113, n765, n731);
xor  g776 (n847, n740, n117, n697, n758);
or   g777 (n790, n123, n731, n145, n702);
or   g778 (n805, n104, n750, n130, n121);
or   g779 (n837, n767, n121, n763);
nand g780 (n839, n697, n770, n129, n139);
nor  g781 (n841, n714, n125, n713, n129);
or   g782 (n863, n701, n768, n116, n98);
and  g783 (n771, n109, n753, n754, n744);
nor  g784 (n781, n100, n105, n762, n131);
xor  g785 (n830, n759, n760, n104, n758);
nor  g786 (n795, n142, n686, n102, n756);
nand g787 (n844, n702, n769, n742, n112);
or   g788 (n860, n101, n712, n741, n761);
or   g789 (n820, n122, n701, n111, n127);
or   g790 (n777, n750, n109, n703, n717);
xnor g791 (n867, n752, n136, n127, n690);
nor  g792 (n794, n101, n767, n128, n122);
xor  g793 (n865, n119, n124, n753, n734);
xor  g794 (n858, n685, n122, n746, n753);
nor  g795 (n783, n707, n698, n114, n691);
nand g796 (n866, n137, n136, n724, n130);
and  g797 (n852, n134, n124, n705, n107);
or   g798 (n832, n108, n770, n110, n112);
xor  g799 (n828, n126, n135, n109, n100);
nor  g800 (n817, n719, n141, n105, n694);
nor  g801 (n835, n126, n687, n717, n99);
and  g802 (n780, n113, n139, n131, n695);
xnor g803 (n786, n123, n732, n725, n126);
nand g804 (n811, n127, n768, n102, n112);
nor  g805 (n859, n754, n696, n738, n708);
or   g806 (n838, n130, n111, n109);
nor  g807 (n797, n767, n120, n133, n747);
xnor g808 (n857, n129, n108, n132, n102);
and  g809 (n776, n765, n710, n693, n739);
xnor g810 (n833, n728, n724, n118, n113);
nor  g811 (n842, n137, n107, n706, n699);
nor  g812 (n810, n769, n140, n137, n764);
and  g813 (n819, n708, n110, n101, n760);
nor  g814 (n779, n755, n141, n142, n734);
nor  g815 (n807, n124, n115, n135, n112);
nor  g816 (n827, n706, n116, n691, n136);
or   g817 (n785, n733, n764, n727, n106);
and  g818 (n774, n99, n766, n123, n719);
xor  g819 (n787, n710, n125, n744, n698);
xnor g820 (n775, n146, n138, n117, n120);
or   g821 (n831, n114, n116, n134, n145);
nand g822 (n818, n721, n115, n116, n104);
or   g823 (n772, n737, n712, n763, n761);
or   g824 (n868, n751, n138, n127, n102);
or   g825 (n850, n143, n128, n745, n139);
nand g826 (n845, n758, n736, n106, n699);
nor  g827 (n808, n141, n688, n686, n752);
and  g828 (n793, n98, n136, n100, n759);
nor  g829 (n846, n745, n134, n688, n760);
xnor g830 (n856, n138, n139, n725, n144);
and  g831 (n778, n742, n129, n118, n107);
xor  g832 (n853, n117, n720, n728, n732);
xnor g833 (n848, n716, n125, n113, n137);
xor  g834 (n826, n115, n141, n122, n743);
nor  g835 (n813, n718, n711, n700, n119);
buf  g836 (n878, n816);
buf  g837 (n887, n821);
not  g838 (n884, n781);
not  g839 (n879, n771);
buf  g840 (n896, n812);
not  g841 (n882, n845);
nand g842 (n892, n789, n834);
and  g843 (n886, n798, n783, n785);
nor  g844 (n885, n833, n807, n830);
nand g845 (n895, n844, n815, n786);
and  g846 (n899, n776, n843, n838);
and  g847 (n893, n823, n809, n795);
xor  g848 (n874, n841, n832, n819);
or   g849 (n880, n835, n784, n808);
or   g850 (n877, n849, n790, n846);
or   g851 (n870, n824, n774, n836);
nand g852 (n890, n829, n817, n788);
nor  g853 (n871, n782, n794, n837);
xor  g854 (n875, n803, n806, n822);
and  g855 (n891, n802, n792, n825);
xnor g856 (n883, n775, n791, n813);
nand g857 (n888, n811, n820, n800);
or   g858 (n869, n810, n827, n840);
xnor g859 (n881, n772, n826, n793);
or   g860 (n898, n778, n796, n805);
nand g861 (n876, n799, n847, n839);
or   g862 (n894, n801, n842, n797);
nand g863 (n889, n831, n787, n804);
or   g864 (n872, n773, n818, n828);
nand g865 (n897, n850, n814, n780);
or   g866 (n873, n779, n777, n848);
not  g867 (n926, n534);
not  g868 (n916, n563);
buf  g869 (n919, n537);
buf  g870 (n924, n874);
or   g871 (n901, n875, n874);
nand g872 (n911, n558, n549, n876);
xor  g873 (n928, n556, n540, n560, n527);
xnor g874 (n922, n552, n535, n871);
nor  g875 (n909, n872, n562, n877, n873);
xnor g876 (n927, n876, n528, n547, n533);
nor  g877 (n920, n872, n872, n551, n545);
nand g878 (n915, n877, n877, n557, n560);
xor  g879 (n929, n878, n536, n877, n561);
nand g880 (n900, n547, n564, n542, n875);
or   g881 (n910, n536, n878, n546, n540);
and  g882 (n925, n550, n875, n873, n871);
xnor g883 (n921, n870, n869, n533, n553);
nand g884 (n914, n874, n556, n550, n554);
xor  g885 (n907, n544, n538, n548, n534);
and  g886 (n903, n554, n555, n875, n537);
nor  g887 (n904, n553, n543, n546, n530);
nand g888 (n906, n543, n538, n870);
nand g889 (n902, n545, n869, n871, n559);
nand g890 (n913, n562, n539, n549);
xnor g891 (n908, n872, n558, n557, n559);
xor  g892 (n912, n870, n873, n561, n876);
nor  g893 (n905, n542, n548, n544, n529);
xnor g894 (n923, n532, n552, n871, n551);
and  g895 (n917, n541, n555, n563, n526);
nor  g896 (n918, n873, n531, n874, n541);
and  g897 (n937, n896, n892, n908);
or   g898 (n946, n882, n893, n884);
xor  g899 (n931, n895, n919, n906, n917);
nand g900 (n935, n881, n897, n879);
nor  g901 (n955, n883, n925, n886, n920);
or   g902 (n934, n891, n915, n884, n898);
nor  g903 (n939, n912, n896, n905);
xor  g904 (n938, n894, n897, n890);
xor  g905 (n930, n889, n893, n926, n887);
nand g906 (n945, n888, n911, n887, n890);
xnor g907 (n957, n898, n891, n893, n887);
xor  g908 (n952, n904, n903, n881, n922);
and  g909 (n949, n880, n890, n900, n894);
xor  g910 (n951, n882, n879, n902, n884);
xnor g911 (n942, n878, n885, n881, n910);
and  g912 (n940, n909, n884, n888, n881);
and  g913 (n941, n880, n898, n887, n899);
nand g914 (n953, n886, n878, n899, n885);
nand g915 (n936, n892, n927, n897, n889);
nand g916 (n947, n895, n883, n898, n888);
and  g917 (n950, n901, n883, n907, n914);
nand g918 (n948, n880, n894, n921, n886);
xor  g919 (n933, n879, n883, n889, n888);
xnor g920 (n944, n924, n880, n923, n885);
nand g921 (n956, n894, n916, n882, n886);
xor  g922 (n932, n891, n913, n896, n889);
nor  g923 (n954, n885, n895, n918);
xor  g924 (n943, n892, n891, n882, n890);
buf  g925 (n978, n32);
buf  g926 (n958, n328);
not  g927 (n967, n929);
buf  g928 (n969, n148);
buf  g929 (n964, n942);
buf  g930 (n972, n933);
buf  g931 (n979, n329);
buf  g932 (n984, n329);
buf  g933 (n966, n566);
buf  g934 (n973, n936);
buf  g935 (n975, n326);
not  g936 (n959, n928);
nand g937 (n976, n32, n147, n940, n567);
xnor g938 (n981, n944, n954, n949, n568);
or   g939 (n971, n327, n570, n569, n957);
or   g940 (n983, n326, n932, n328, n568);
or   g941 (n962, n148, n931, n947, n570);
nand g942 (n980, n572, n950, n957, n945);
and  g943 (n982, n930, n326, n147);
nor  g944 (n965, n327, n328, n571, n565);
xor  g945 (n970, n569, n327, n934, n938);
xnor g946 (n977, n943, n147, n939, n927);
or   g947 (n985, n929, n146, n564);
nand g948 (n963, n948, n956, n327, n851);
nor  g949 (n986, n937, n329, n566, n953);
or   g950 (n974, n565, n571, n32, n328);
nand g951 (n968, n946, n32, n951, n928);
and  g952 (n960, n147, n567, n935, n952);
xnor g953 (n961, n329, n955, n941, n31);
xnor g954 (n993, n149, n974, n982, n980);
xnor g955 (n995, n150, n150, n972, n966);
and  g956 (n1011, n976, n976, n979, n983);
or   g957 (n1003, n970, n151, n961, n959);
xnor g958 (n1018, n985, n960, n979, n965);
xor  g959 (n1006, n984, n148, n968, n151);
and  g960 (n1005, n983, n971, n977, n980);
or   g961 (n1004, n964, n978, n573, n965);
xnor g962 (n1010, n958, n981, n971, n974);
nor  g963 (n999, n972, n971, n961, n964);
xnor g964 (n997, n978, n982, n974, n852);
and  g965 (n1016, n973, n985, n983, n969);
xnor g966 (n1008, n973, n981, n977, n980);
and  g967 (n992, n965, n958, n969, n964);
and  g968 (n991, n974, n149, n975, n960);
xnor g969 (n1020, n964, n959, n152, n961);
nor  g970 (n1013, n572, n573, n971, n960);
nand g971 (n990, n968, n958, n970, n980);
and  g972 (n1012, n970, n961, n149, n152);
xor  g973 (n994, n976, n982, n963);
nor  g974 (n1014, n981, n977, n976, n966);
xnor g975 (n989, n959, n985, n969);
nand g976 (n1000, n962, n978, n152, n975);
nor  g977 (n1017, n966, n977, n149, n968);
xnor g978 (n1009, n981, n150, n984, n962);
nand g979 (n1007, n963, n968, n967, n972);
nand g980 (n1015, n962, n967, n152, n969);
xnor g981 (n1019, n975, n962, n963, n979);
xnor g982 (n1001, n150, n983, n973, n574);
nor  g983 (n998, n986, n967, n970, n973);
or   g984 (n1002, n984, n967, n151, n965);
or   g985 (n987, n984, n151, n972, n978);
xnor g986 (n996, n958, n975, n959, n960);
xor  g987 (n988, n982, n966, n148, n979);
xnor g988 (n1027, n854, n1018, n986, n1019);
xor  g989 (n1026, n861, n1016, n856, n860);
nand g990 (n1022, n1014, n867, n868, n857);
nor  g991 (n1025, n864, n899, n866, n859);
and  g992 (n1023, n1015, n858, n863, n862);
xor  g993 (n1021, n853, n1020, n865, n855);
nand g994 (n1024, n1017, n986, n899);
buf  g995 (n1030, n574);
not  g996 (n1028, n1025);
nand g997 (n1029, n1024, n1026);
and  g998 (n1032, n1027, n1028, n638);
xnor g999 (n1031, n1029, n638, n1030);
endmodule
