

module Stat_1057_14_11
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n771,
  n1065,
  n1076,
  n1074,
  n1071,
  n1070,
  n1067,
  n1069,
  n1075,
  n1073,
  n1061,
  n1057,
  n1064,
  n1068,
  n1072,
  n1058,
  n1066,
  n1055,
  n1056,
  n1063,
  n1062,
  n1059,
  n1060,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n771;
  output n1065;
  output n1076;
  output n1074;
  output n1071;
  output n1070;
  output n1067;
  output n1069;
  output n1075;
  output n1073;
  output n1061;
  output n1057;
  output n1064;
  output n1068;
  output n1072;
  output n1058;
  output n1066;
  output n1055;
  output n1056;
  output n1063;
  output n1062;
  output n1059;
  output n1060;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n90,
    n11
  );


  not
  g1
  (
    n93,
    n8
  );


  not
  g2
  (
    n79,
    n4
  );


  not
  g3
  (
    n53,
    n13
  );


  buf
  g4
  (
    n49,
    n10
  );


  not
  g5
  (
    n77,
    n18
  );


  buf
  g6
  (
    n70,
    n15
  );


  not
  g7
  (
    n33,
    n12
  );


  buf
  g8
  (
    n60,
    n9
  );


  not
  g9
  (
    n34,
    n5
  );


  buf
  g10
  (
    n78,
    n14
  );


  buf
  g11
  (
    n65,
    n19
  );


  buf
  g12
  (
    n21,
    n16
  );


  not
  g13
  (
    n61,
    n19
  );


  not
  g14
  (
    n75,
    n19
  );


  buf
  g15
  (
    n26,
    n14
  );


  buf
  g16
  (
    n32,
    n4
  );


  buf
  g17
  (
    KeyWire_0_20,
    n5
  );


  not
  g18
  (
    n76,
    n8
  );


  not
  g19
  (
    n43,
    n1
  );


  buf
  g20
  (
    n48,
    n13
  );


  not
  g21
  (
    n30,
    n14
  );


  not
  g22
  (
    n41,
    n15
  );


  buf
  g23
  (
    n91,
    n3
  );


  not
  g24
  (
    KeyWire_0_34,
    n15
  );


  buf
  g25
  (
    n51,
    n7
  );


  not
  g26
  (
    n67,
    n12
  );


  not
  g27
  (
    n58,
    n1
  );


  buf
  g28
  (
    n69,
    n2
  );


  not
  g29
  (
    n22,
    n13
  );


  not
  g30
  (
    n94,
    n7
  );


  buf
  g31
  (
    n52,
    n7
  );


  not
  g32
  (
    n27,
    n18
  );


  not
  g33
  (
    n42,
    n4
  );


  buf
  g34
  (
    n59,
    n3
  );


  buf
  g35
  (
    n84,
    n4
  );


  not
  g36
  (
    n71,
    n8
  );


  not
  g37
  (
    n56,
    n6
  );


  buf
  g38
  (
    n82,
    n12
  );


  not
  g39
  (
    n20,
    n11
  );


  buf
  g40
  (
    n39,
    n8
  );


  not
  g41
  (
    n57,
    n6
  );


  buf
  g42
  (
    n92,
    n2
  );


  buf
  g43
  (
    n38,
    n17
  );


  buf
  g44
  (
    n73,
    n9
  );


  not
  g45
  (
    n68,
    n7
  );


  not
  g46
  (
    n87,
    n17
  );


  buf
  g47
  (
    KeyWire_0_54,
    n1
  );


  buf
  g48
  (
    n95,
    n19
  );


  buf
  g49
  (
    n64,
    n2
  );


  not
  g50
  (
    n72,
    n6
  );


  not
  g51
  (
    n83,
    n15
  );


  not
  g52
  (
    n31,
    n14
  );


  not
  g53
  (
    n88,
    n6
  );


  not
  g54
  (
    n40,
    n16
  );


  buf
  g55
  (
    n74,
    n1
  );


  buf
  g56
  (
    n89,
    n9
  );


  not
  g57
  (
    n36,
    n3
  );


  buf
  g58
  (
    n37,
    n17
  );


  buf
  g59
  (
    n25,
    n5
  );


  buf
  g60
  (
    n47,
    n16
  );


  buf
  g61
  (
    n62,
    n17
  );


  not
  g62
  (
    n44,
    n10
  );


  buf
  g63
  (
    n24,
    n18
  );


  not
  g64
  (
    n63,
    n5
  );


  buf
  g65
  (
    n45,
    n18
  );


  not
  g66
  (
    n29,
    n10
  );


  not
  g67
  (
    n23,
    n16
  );


  buf
  g68
  (
    n35,
    n12
  );


  not
  g69
  (
    n46,
    n11
  );


  not
  g70
  (
    n28,
    n2
  );


  buf
  g71
  (
    n66,
    n10
  );


  buf
  g72
  (
    n81,
    n13
  );


  buf
  g73
  (
    KeyWire_0_46,
    n9
  );


  not
  g74
  (
    n85,
    n11
  );


  not
  g75
  (
    n80,
    n3
  );


  buf
  g76
  (
    n322,
    n56
  );


  not
  g77
  (
    n366,
    n91
  );


  buf
  g78
  (
    n265,
    n23
  );


  not
  g79
  (
    KeyWire_0_38,
    n41
  );


  not
  g80
  (
    n237,
    n22
  );


  buf
  g81
  (
    n104,
    n47
  );


  buf
  g82
  (
    n157,
    n33
  );


  not
  g83
  (
    n128,
    n68
  );


  not
  g84
  (
    n107,
    n57
  );


  buf
  g85
  (
    n148,
    n93
  );


  buf
  g86
  (
    n315,
    n89
  );


  not
  g87
  (
    n217,
    n50
  );


  not
  g88
  (
    n290,
    n53
  );


  not
  g89
  (
    n206,
    n57
  );


  not
  g90
  (
    n369,
    n80
  );


  buf
  g91
  (
    n150,
    n46
  );


  not
  g92
  (
    n133,
    n42
  );


  not
  g93
  (
    n121,
    n32
  );


  not
  g94
  (
    n342,
    n94
  );


  not
  g95
  (
    n240,
    n28
  );


  buf
  g96
  (
    n296,
    n90
  );


  not
  g97
  (
    n362,
    n56
  );


  buf
  g98
  (
    n295,
    n49
  );


  not
  g99
  (
    n102,
    n22
  );


  buf
  g100
  (
    n360,
    n20
  );


  buf
  g101
  (
    n142,
    n72
  );


  not
  g102
  (
    n226,
    n30
  );


  buf
  g103
  (
    n147,
    n59
  );


  not
  g104
  (
    n208,
    n24
  );


  not
  g105
  (
    n381,
    n89
  );


  not
  g106
  (
    n307,
    n56
  );


  buf
  g107
  (
    n215,
    n77
  );


  buf
  g108
  (
    n389,
    n32
  );


  buf
  g109
  (
    n123,
    n83
  );


  not
  g110
  (
    n251,
    n21
  );


  not
  g111
  (
    n122,
    n73
  );


  not
  g112
  (
    n168,
    n47
  );


  not
  g113
  (
    n309,
    n48
  );


  not
  g114
  (
    n340,
    n82
  );


  buf
  g115
  (
    n98,
    n73
  );


  not
  g116
  (
    n328,
    n75
  );


  buf
  g117
  (
    n184,
    n28
  );


  not
  g118
  (
    n269,
    n80
  );


  not
  g119
  (
    n278,
    n34
  );


  buf
  g120
  (
    n117,
    n85
  );


  not
  g121
  (
    n187,
    n83
  );


  buf
  g122
  (
    n285,
    n27
  );


  not
  g123
  (
    n384,
    n36
  );


  not
  g124
  (
    n140,
    n39
  );


  not
  g125
  (
    n195,
    n44
  );


  not
  g126
  (
    n186,
    n63
  );


  buf
  g127
  (
    n247,
    n52
  );


  not
  g128
  (
    n266,
    n64
  );


  not
  g129
  (
    n308,
    n51
  );


  buf
  g130
  (
    KeyWire_0_22,
    n84
  );


  not
  g131
  (
    n116,
    n90
  );


  buf
  g132
  (
    n234,
    n44
  );


  buf
  g133
  (
    n352,
    n89
  );


  not
  g134
  (
    n270,
    n26
  );


  not
  g135
  (
    n317,
    n55
  );


  not
  g136
  (
    n106,
    n88
  );


  buf
  g137
  (
    n244,
    n40
  );


  buf
  g138
  (
    n219,
    n91
  );


  buf
  g139
  (
    n159,
    n60
  );


  buf
  g140
  (
    KeyWire_0_53,
    n41
  );


  not
  g141
  (
    n292,
    n36
  );


  not
  g142
  (
    n203,
    n69
  );


  not
  g143
  (
    n262,
    n75
  );


  buf
  g144
  (
    n174,
    n33
  );


  not
  g145
  (
    n141,
    n30
  );


  not
  g146
  (
    n127,
    n45
  );


  not
  g147
  (
    n232,
    n48
  );


  not
  g148
  (
    n139,
    n93
  );


  buf
  g149
  (
    KeyWire_0_35,
    n39
  );


  not
  g150
  (
    n109,
    n58
  );


  not
  g151
  (
    n151,
    n63
  );


  buf
  g152
  (
    n349,
    n74
  );


  buf
  g153
  (
    KeyWire_0_15,
    n38
  );


  buf
  g154
  (
    n257,
    n61
  );


  buf
  g155
  (
    n129,
    n94
  );


  not
  g156
  (
    n275,
    n47
  );


  buf
  g157
  (
    n385,
    n63
  );


  buf
  g158
  (
    n331,
    n62
  );


  not
  g159
  (
    n394,
    n57
  );


  buf
  g160
  (
    n119,
    n49
  );


  buf
  g161
  (
    KeyWire_0_12,
    n80
  );


  not
  g162
  (
    KeyWire_0_13,
    n62
  );


  buf
  g163
  (
    n303,
    n77
  );


  not
  g164
  (
    n231,
    n25
  );


  buf
  g165
  (
    n306,
    n45
  );


  not
  g166
  (
    n281,
    n71
  );


  not
  g167
  (
    n143,
    n23
  );


  not
  g168
  (
    KeyWire_0_19,
    n92
  );


  not
  g169
  (
    n361,
    n54
  );


  not
  g170
  (
    n101,
    n31
  );


  not
  g171
  (
    n166,
    n71
  );


  buf
  g172
  (
    n372,
    n34
  );


  buf
  g173
  (
    n393,
    n61
  );


  buf
  g174
  (
    n209,
    n42
  );


  not
  g175
  (
    n132,
    n70
  );


  buf
  g176
  (
    n334,
    n92
  );


  not
  g177
  (
    n387,
    n58
  );


  buf
  g178
  (
    n204,
    n84
  );


  not
  g179
  (
    n347,
    n29
  );


  not
  g180
  (
    n351,
    n52
  );


  buf
  g181
  (
    n239,
    n54
  );


  buf
  g182
  (
    n355,
    n79
  );


  not
  g183
  (
    n200,
    n58
  );


  not
  g184
  (
    n326,
    n25
  );


  not
  g185
  (
    KeyWire_0_1,
    n38
  );


  not
  g186
  (
    n249,
    n52
  );


  buf
  g187
  (
    n344,
    n55
  );


  not
  g188
  (
    n310,
    n73
  );


  not
  g189
  (
    n259,
    n45
  );


  not
  g190
  (
    n210,
    n90
  );


  buf
  g191
  (
    n377,
    n70
  );


  buf
  g192
  (
    n304,
    n83
  );


  not
  g193
  (
    n131,
    n42
  );


  not
  g194
  (
    n300,
    n71
  );


  buf
  g195
  (
    n325,
    n35
  );


  buf
  g196
  (
    n96,
    n54
  );


  buf
  g197
  (
    n291,
    n87
  );


  buf
  g198
  (
    n346,
    n66
  );


  buf
  g199
  (
    n162,
    n43
  );


  buf
  g200
  (
    n341,
    n93
  );


  not
  g201
  (
    n316,
    n64
  );


  buf
  g202
  (
    n323,
    n82
  );


  buf
  g203
  (
    n177,
    n46
  );


  not
  g204
  (
    n164,
    n53
  );


  not
  g205
  (
    n336,
    n88
  );


  not
  g206
  (
    n379,
    n35
  );


  not
  g207
  (
    n190,
    n29
  );


  not
  g208
  (
    KeyWire_0_58,
    n74
  );


  buf
  g209
  (
    n179,
    n30
  );


  buf
  g210
  (
    n343,
    n94
  );


  not
  g211
  (
    n213,
    n61
  );


  not
  g212
  (
    n156,
    n67
  );


  buf
  g213
  (
    n192,
    n69
  );


  not
  g214
  (
    n223,
    n42
  );


  not
  g215
  (
    KeyWire_0_28,
    n20
  );


  not
  g216
  (
    KeyWire_0_25,
    n38
  );


  buf
  g217
  (
    n264,
    n46
  );


  buf
  g218
  (
    n335,
    n84
  );


  buf
  g219
  (
    n197,
    n67
  );


  buf
  g220
  (
    n145,
    n86
  );


  not
  g221
  (
    n297,
    n81
  );


  buf
  g222
  (
    n161,
    n91
  );


  buf
  g223
  (
    n294,
    n23
  );


  not
  g224
  (
    n312,
    n55
  );


  not
  g225
  (
    n155,
    n66
  );


  not
  g226
  (
    n365,
    n34
  );


  buf
  g227
  (
    n238,
    n81
  );


  buf
  g228
  (
    n110,
    n70
  );


  buf
  g229
  (
    n392,
    n21
  );


  not
  g230
  (
    n178,
    n31
  );


  not
  g231
  (
    n152,
    n50
  );


  not
  g232
  (
    n271,
    n80
  );


  not
  g233
  (
    n327,
    n55
  );


  buf
  g234
  (
    n284,
    n34
  );


  buf
  g235
  (
    n373,
    n35
  );


  buf
  g236
  (
    n207,
    n47
  );


  not
  g237
  (
    n134,
    n86
  );


  not
  g238
  (
    n380,
    n60
  );


  buf
  g239
  (
    n391,
    n37
  );


  not
  g240
  (
    n277,
    n29
  );


  not
  g241
  (
    n293,
    n95
  );


  buf
  g242
  (
    n205,
    n51
  );


  buf
  g243
  (
    n321,
    n72
  );


  buf
  g244
  (
    n286,
    n78
  );


  buf
  g245
  (
    n170,
    n60
  );


  buf
  g246
  (
    n337,
    n85
  );


  not
  g247
  (
    n339,
    n86
  );


  not
  g248
  (
    n202,
    n58
  );


  not
  g249
  (
    n144,
    n85
  );


  buf
  g250
  (
    n256,
    n25
  );


  not
  g251
  (
    n149,
    n71
  );


  not
  g252
  (
    n263,
    n78
  );


  buf
  g253
  (
    n158,
    n33
  );


  buf
  g254
  (
    n198,
    n88
  );


  not
  g255
  (
    n287,
    n75
  );


  not
  g256
  (
    n242,
    n76
  );


  buf
  g257
  (
    n398,
    n65
  );


  buf
  g258
  (
    n279,
    n95
  );


  buf
  g259
  (
    n189,
    n72
  );


  not
  g260
  (
    KeyWire_0_45,
    n43
  );


  not
  g261
  (
    n105,
    n24
  );


  not
  g262
  (
    n350,
    n84
  );


  buf
  g263
  (
    KeyWire_0_10,
    n29
  );


  buf
  g264
  (
    KeyWire_0_33,
    n62
  );


  not
  g265
  (
    n274,
    n41
  );


  buf
  g266
  (
    n248,
    n92
  );


  not
  g267
  (
    n114,
    n76
  );


  buf
  g268
  (
    n193,
    n40
  );


  buf
  g269
  (
    n333,
    n93
  );


  not
  g270
  (
    n224,
    n36
  );


  buf
  g271
  (
    n188,
    n37
  );


  not
  g272
  (
    n367,
    n50
  );


  not
  g273
  (
    n358,
    n75
  );


  buf
  g274
  (
    n97,
    n59
  );


  buf
  g275
  (
    n301,
    n57
  );


  buf
  g276
  (
    n314,
    n59
  );


  buf
  g277
  (
    KeyWire_0_55,
    n65
  );


  buf
  g278
  (
    KeyWire_0_17,
    n78
  );


  buf
  g279
  (
    n163,
    n61
  );


  not
  g280
  (
    n115,
    n67
  );


  buf
  g281
  (
    n108,
    n28
  );


  buf
  g282
  (
    n368,
    n33
  );


  buf
  g283
  (
    KeyWire_0_41,
    n30
  );


  buf
  g284
  (
    n216,
    n21
  );


  not
  g285
  (
    n130,
    n50
  );


  not
  g286
  (
    n330,
    n24
  );


  not
  g287
  (
    n260,
    n73
  );


  not
  g288
  (
    n126,
    n54
  );


  buf
  g289
  (
    n99,
    n65
  );


  buf
  g290
  (
    n235,
    n82
  );


  buf
  g291
  (
    n222,
    n69
  );


  buf
  g292
  (
    n250,
    n68
  );


  not
  g293
  (
    n298,
    n83
  );


  not
  g294
  (
    KeyWire_0_2,
    n40
  );


  not
  g295
  (
    n374,
    n22
  );


  buf
  g296
  (
    n230,
    n79
  );


  buf
  g297
  (
    n169,
    n81
  );


  not
  g298
  (
    n338,
    n78
  );


  not
  g299
  (
    n364,
    n68
  );


  buf
  g300
  (
    n112,
    n74
  );


  not
  g301
  (
    n243,
    n43
  );


  not
  g302
  (
    n218,
    n67
  );


  buf
  g303
  (
    n345,
    n25
  );


  not
  g304
  (
    n329,
    n32
  );


  not
  g305
  (
    n245,
    n26
  );


  not
  g306
  (
    n182,
    n36
  );


  not
  g307
  (
    n252,
    n76
  );


  not
  g308
  (
    n241,
    n51
  );


  buf
  g309
  (
    n185,
    n45
  );


  buf
  g310
  (
    n227,
    n90
  );


  buf
  g311
  (
    n319,
    n81
  );


  buf
  g312
  (
    n288,
    n31
  );


  not
  g313
  (
    n376,
    n53
  );


  buf
  g314
  (
    KeyWire_0_5,
    n87
  );


  buf
  g315
  (
    n214,
    n38
  );


  buf
  g316
  (
    n370,
    n27
  );


  buf
  g317
  (
    n354,
    n27
  );


  buf
  g318
  (
    n153,
    n74
  );


  buf
  g319
  (
    n280,
    n79
  );


  not
  g320
  (
    n258,
    n92
  );


  not
  g321
  (
    n318,
    n77
  );


  not
  g322
  (
    n302,
    n49
  );


  buf
  g323
  (
    n118,
    n64
  );


  not
  g324
  (
    n255,
    n39
  );


  buf
  g325
  (
    n113,
    n64
  );


  buf
  g326
  (
    n103,
    n56
  );


  buf
  g327
  (
    n220,
    n39
  );


  not
  g328
  (
    n324,
    n89
  );


  buf
  g329
  (
    KeyWire_0_44,
    n20
  );


  buf
  g330
  (
    n383,
    n35
  );


  not
  g331
  (
    n160,
    n77
  );


  buf
  g332
  (
    n313,
    n52
  );


  not
  g333
  (
    n191,
    n66
  );


  buf
  g334
  (
    n283,
    n70
  );


  buf
  g335
  (
    n356,
    n59
  );


  not
  g336
  (
    n136,
    n79
  );


  buf
  g337
  (
    n268,
    n63
  );


  not
  g338
  (
    n261,
    n23
  );


  buf
  g339
  (
    n276,
    n37
  );


  not
  g340
  (
    n311,
    n46
  );


  not
  g341
  (
    n375,
    n49
  );


  buf
  g342
  (
    n289,
    n21
  );


  buf
  g343
  (
    n173,
    n48
  );


  buf
  g344
  (
    n175,
    n69
  );


  not
  g345
  (
    n194,
    n82
  );


  buf
  g346
  (
    n267,
    n87
  );


  not
  g347
  (
    n183,
    n60
  );


  not
  g348
  (
    n236,
    n62
  );


  buf
  g349
  (
    n167,
    n22
  );


  buf
  g350
  (
    n390,
    n26
  );


  not
  g351
  (
    KeyWire_0_32,
    n40
  );


  not
  g352
  (
    n353,
    n88
  );


  not
  g353
  (
    n212,
    n72
  );


  buf
  g354
  (
    n154,
    n24
  );


  buf
  g355
  (
    n357,
    n43
  );


  buf
  g356
  (
    n371,
    n65
  );


  not
  g357
  (
    n135,
    n20
  );


  buf
  g358
  (
    n172,
    n27
  );


  not
  g359
  (
    n171,
    n41
  );


  not
  g360
  (
    n273,
    n76
  );


  buf
  g361
  (
    n397,
    n86
  );


  not
  g362
  (
    n348,
    n95
  );


  not
  g363
  (
    KeyWire_0_51,
    n28
  );


  buf
  g364
  (
    n146,
    n44
  );


  buf
  g365
  (
    KeyWire_0_57,
    n94
  );


  not
  g366
  (
    n138,
    n44
  );


  buf
  g367
  (
    n395,
    n37
  );


  buf
  g368
  (
    n386,
    n87
  );


  buf
  g369
  (
    n137,
    n53
  );


  buf
  g370
  (
    n120,
    n31
  );


  not
  g371
  (
    n229,
    n85
  );


  buf
  g372
  (
    n359,
    n66
  );


  not
  g373
  (
    n221,
    n32
  );


  not
  g374
  (
    n272,
    n48
  );


  not
  g375
  (
    n196,
    n68
  );


  buf
  g376
  (
    n165,
    n26
  );


  buf
  g377
  (
    n228,
    n51
  );


  buf
  g378
  (
    n201,
    n91
  );


  buf
  g379
  (
    n624,
    n299
  );


  not
  g380
  (
    n580,
    n357
  );


  not
  g381
  (
    KeyWire_0_52,
    n391
  );


  buf
  g382
  (
    n412,
    n333
  );


  not
  g383
  (
    n546,
    n376
  );


  buf
  g384
  (
    n420,
    n313
  );


  buf
  g385
  (
    n692,
    n215
  );


  buf
  g386
  (
    n621,
    n191
  );


  not
  g387
  (
    n493,
    n97
  );


  not
  g388
  (
    n726,
    n380
  );


  not
  g389
  (
    n471,
    n358
  );


  not
  g390
  (
    n419,
    n369
  );


  not
  g391
  (
    n442,
    n370
  );


  not
  g392
  (
    n399,
    n390
  );


  buf
  g393
  (
    n633,
    n221
  );


  buf
  g394
  (
    n522,
    n253
  );


  not
  g395
  (
    n504,
    n106
  );


  not
  g396
  (
    n694,
    n201
  );


  not
  g397
  (
    n429,
    n380
  );


  not
  g398
  (
    n541,
    n133
  );


  buf
  g399
  (
    n464,
    n199
  );


  not
  g400
  (
    n590,
    n305
  );


  buf
  g401
  (
    n611,
    n236
  );


  buf
  g402
  (
    n698,
    n331
  );


  buf
  g403
  (
    n720,
    n352
  );


  not
  g404
  (
    n618,
    n359
  );


  buf
  g405
  (
    n413,
    n357
  );


  not
  g406
  (
    n647,
    n352
  );


  not
  g407
  (
    n655,
    n372
  );


  buf
  g408
  (
    KeyWire_0_29,
    n185
  );


  buf
  g409
  (
    n542,
    n183
  );


  buf
  g410
  (
    n450,
    n225
  );


  not
  g411
  (
    n607,
    n143
  );


  not
  g412
  (
    n482,
    n208
  );


  buf
  g413
  (
    n461,
    n390
  );


  buf
  g414
  (
    n718,
    n272
  );


  buf
  g415
  (
    n729,
    n322
  );


  not
  g416
  (
    n747,
    n373
  );


  buf
  g417
  (
    n595,
    n279
  );


  not
  g418
  (
    n717,
    n368
  );


  buf
  g419
  (
    n731,
    n114
  );


  buf
  g420
  (
    n660,
    n344
  );


  not
  g421
  (
    n734,
    n351
  );


  not
  g422
  (
    n416,
    n149
  );


  buf
  g423
  (
    n564,
    n275
  );


  not
  g424
  (
    n439,
    n101
  );


  not
  g425
  (
    n634,
    n388
  );


  buf
  g426
  (
    KeyWire_0_60,
    n323
  );


  buf
  g427
  (
    n437,
    n381
  );


  buf
  g428
  (
    n689,
    n379
  );


  not
  g429
  (
    KeyWire_0_27,
    n285
  );


  not
  g430
  (
    n481,
    n338
  );


  not
  g431
  (
    n579,
    n281
  );


  not
  g432
  (
    n536,
    n301
  );


  buf
  g433
  (
    n631,
    n232
  );


  not
  g434
  (
    n679,
    n391
  );


  buf
  g435
  (
    n555,
    n138
  );


  not
  g436
  (
    n661,
    n386
  );


  buf
  g437
  (
    n581,
    n240
  );


  not
  g438
  (
    KeyWire_0_18,
    n246
  );


  not
  g439
  (
    n530,
    n242
  );


  not
  g440
  (
    KeyWire_0_47,
    n354
  );


  buf
  g441
  (
    n709,
    n342
  );


  buf
  g442
  (
    n714,
    n359
  );


  not
  g443
  (
    n430,
    n227
  );


  buf
  g444
  (
    n737,
    n355
  );


  not
  g445
  (
    n742,
    n361
  );


  buf
  g446
  (
    n405,
    n375
  );


  buf
  g447
  (
    n623,
    n388
  );


  not
  g448
  (
    n514,
    n283
  );


  buf
  g449
  (
    n699,
    n269
  );


  buf
  g450
  (
    n575,
    n344
  );


  not
  g451
  (
    n697,
    n117
  );


  not
  g452
  (
    n646,
    n142
  );


  not
  g453
  (
    n553,
    n200
  );


  buf
  g454
  (
    n677,
    n147
  );


  buf
  g455
  (
    n500,
    n145
  );


  not
  g456
  (
    n417,
    n366
  );


  buf
  g457
  (
    n423,
    n336
  );


  buf
  g458
  (
    n670,
    n156
  );


  buf
  g459
  (
    n507,
    n315
  );


  buf
  g460
  (
    n441,
    n312
  );


  not
  g461
  (
    n418,
    n166
  );


  not
  g462
  (
    n715,
    n367
  );


  not
  g463
  (
    n627,
    n186
  );


  buf
  g464
  (
    n604,
    n198
  );


  buf
  g465
  (
    n733,
    n338
  );


  not
  g466
  (
    n577,
    n298
  );


  not
  g467
  (
    n512,
    n123
  );


  not
  g468
  (
    n434,
    n377
  );


  not
  g469
  (
    n616,
    n254
  );


  buf
  g470
  (
    n691,
    n274
  );


  buf
  g471
  (
    n465,
    n357
  );


  not
  g472
  (
    n613,
    n118
  );


  buf
  g473
  (
    n445,
    n293
  );


  buf
  g474
  (
    n549,
    n360
  );


  buf
  g475
  (
    KeyWire_0_4,
    n165
  );


  not
  g476
  (
    n738,
    n104
  );


  buf
  g477
  (
    n444,
    n126
  );


  not
  g478
  (
    n603,
    n245
  );


  buf
  g479
  (
    n723,
    n169
  );


  buf
  g480
  (
    n470,
    n328
  );


  not
  g481
  (
    n548,
    n243
  );


  buf
  g482
  (
    n711,
    n390
  );


  buf
  g483
  (
    n705,
    n140
  );


  not
  g484
  (
    n727,
    n187
  );


  not
  g485
  (
    n440,
    n181
  );


  buf
  g486
  (
    KeyWire_0_16,
    n152
  );


  buf
  g487
  (
    n523,
    n360
  );


  buf
  g488
  (
    n732,
    n369
  );


  buf
  g489
  (
    n710,
    n192
  );


  buf
  g490
  (
    n740,
    n116
  );


  not
  g491
  (
    n642,
    n334
  );


  buf
  g492
  (
    n659,
    n353
  );


  buf
  g493
  (
    n678,
    n220
  );


  not
  g494
  (
    n400,
    n105
  );


  not
  g495
  (
    n456,
    n378
  );


  buf
  g496
  (
    n645,
    n373
  );


  buf
  g497
  (
    n712,
    n290
  );


  not
  g498
  (
    n650,
    n150
  );


  buf
  g499
  (
    n432,
    n125
  );


  not
  g500
  (
    n612,
    n174
  );


  not
  g501
  (
    n680,
    n99
  );


  not
  g502
  (
    n508,
    n136
  );


  buf
  g503
  (
    n449,
    n258
  );


  buf
  g504
  (
    n630,
    n334
  );


  buf
  g505
  (
    n510,
    n311
  );


  buf
  g506
  (
    n498,
    n259
  );


  buf
  g507
  (
    n495,
    n160
  );


  buf
  g508
  (
    n436,
    n226
  );


  buf
  g509
  (
    n672,
    n154
  );


  buf
  g510
  (
    n540,
    n383
  );


  buf
  g511
  (
    n640,
    n379
  );


  not
  g512
  (
    n473,
    n110
  );


  not
  g513
  (
    n695,
    n155
  );


  not
  g514
  (
    n704,
    n261
  );


  not
  g515
  (
    n414,
    n196
  );


  buf
  g516
  (
    n489,
    n251
  );


  buf
  g517
  (
    n597,
    n282
  );


  not
  g518
  (
    n629,
    n324
  );


  not
  g519
  (
    KeyWire_0_61,
    n341
  );


  buf
  g520
  (
    n518,
    n300
  );


  buf
  g521
  (
    n739,
    n354
  );


  not
  g522
  (
    n703,
    n108
  );


  buf
  g523
  (
    n681,
    n264
  );


  not
  g524
  (
    n584,
    n382
  );


  buf
  g525
  (
    KeyWire_0_7,
    n375
  );


  not
  g526
  (
    n422,
    n205
  );


  buf
  g527
  (
    n520,
    n332
  );


  buf
  g528
  (
    n525,
    n129
  );


  not
  g529
  (
    n455,
    n249
  );


  buf
  g530
  (
    n503,
    n379
  );


  buf
  g531
  (
    n639,
    n276
  );


  not
  g532
  (
    n543,
    n350
  );


  buf
  g533
  (
    n499,
    n361
  );


  not
  g534
  (
    n620,
    n308
  );


  buf
  g535
  (
    n665,
    n364
  );


  buf
  g536
  (
    n528,
    n347
  );


  not
  g537
  (
    n632,
    n332
  );


  not
  g538
  (
    KeyWire_0_50,
    n351
  );


  buf
  g539
  (
    n466,
    n389
  );


  buf
  g540
  (
    n459,
    n137
  );


  not
  g541
  (
    n669,
    n378
  );


  buf
  g542
  (
    n708,
    n189
  );


  buf
  g543
  (
    n526,
    n350
  );


  not
  g544
  (
    n609,
    n153
  );


  not
  g545
  (
    n447,
    n250
  );


  buf
  g546
  (
    n568,
    n273
  );


  not
  g547
  (
    n566,
    n384
  );


  buf
  g548
  (
    n599,
    n223
  );


  not
  g549
  (
    n651,
    n139
  );


  not
  g550
  (
    n683,
    n386
  );


  not
  g551
  (
    n668,
    n376
  );


  not
  g552
  (
    n676,
    n372
  );


  not
  g553
  (
    n690,
    n134
  );


  buf
  g554
  (
    n460,
    n381
  );


  buf
  g555
  (
    n454,
    n387
  );


  buf
  g556
  (
    KeyWire_0_49,
    n361
  );


  buf
  g557
  (
    n602,
    n268
  );


  buf
  g558
  (
    n664,
    n260
  );


  not
  g559
  (
    n467,
    n348
  );


  not
  g560
  (
    n476,
    n288
  );


  buf
  g561
  (
    n598,
    n96
  );


  not
  g562
  (
    n558,
    n204
  );


  not
  g563
  (
    n741,
    n121
  );


  buf
  g564
  (
    n527,
    n190
  );


  buf
  g565
  (
    n744,
    n325
  );


  not
  g566
  (
    n538,
    n148
  );


  not
  g567
  (
    n474,
    n157
  );


  not
  g568
  (
    KeyWire_0_42,
    n228
  );


  buf
  g569
  (
    n673,
    n381
  );


  buf
  g570
  (
    n657,
    n337
  );


  buf
  g571
  (
    n516,
    n385
  );


  buf
  g572
  (
    n517,
    n144
  );


  buf
  g573
  (
    n625,
    n321
  );


  buf
  g574
  (
    n614,
    n314
  );


  not
  g575
  (
    n636,
    n202
  );


  not
  g576
  (
    n529,
    n341
  );


  not
  g577
  (
    n656,
    n267
  );


  not
  g578
  (
    n666,
    n329
  );


  not
  g579
  (
    n452,
    n365
  );


  buf
  g580
  (
    KeyWire_0_48,
    n368
  );


  not
  g581
  (
    n728,
    n241
  );


  not
  g582
  (
    n572,
    n318
  );


  buf
  g583
  (
    n571,
    n359
  );


  buf
  g584
  (
    n674,
    n257
  );


  buf
  g585
  (
    n589,
    n178
  );


  buf
  g586
  (
    n648,
    n280
  );


  buf
  g587
  (
    n426,
    n353
  );


  not
  g588
  (
    n610,
    n319
  );


  buf
  g589
  (
    n537,
    n384
  );


  buf
  g590
  (
    n750,
    n320
  );


  not
  g591
  (
    n688,
    n331
  );


  buf
  g592
  (
    n685,
    n349
  );


  not
  g593
  (
    n539,
    n327
  );


  not
  g594
  (
    KeyWire_0_26,
    n211
  );


  buf
  g595
  (
    n684,
    n231
  );


  not
  g596
  (
    n488,
    n238
  );


  not
  g597
  (
    n535,
    n107
  );


  not
  g598
  (
    n743,
    n307
  );


  buf
  g599
  (
    n506,
    n385
  );


  buf
  g600
  (
    n573,
    n214
  );


  buf
  g601
  (
    n494,
    n162
  );


  not
  g602
  (
    KeyWire_0_59,
    n366
  );


  buf
  g603
  (
    n588,
    n369
  );


  buf
  g604
  (
    n578,
    n224
  );


  not
  g605
  (
    n463,
    n376
  );


  not
  g606
  (
    n401,
    n353
  );


  not
  g607
  (
    n706,
    n367
  );


  buf
  g608
  (
    n561,
    n203
  );


  not
  g609
  (
    n424,
    n374
  );


  not
  g610
  (
    n600,
    n336
  );


  buf
  g611
  (
    n722,
    n248
  );


  buf
  g612
  (
    n713,
    n366
  );


  buf
  g613
  (
    n736,
    n335
  );


  buf
  g614
  (
    n428,
    n349
  );


  not
  g615
  (
    n560,
    n339
  );


  buf
  g616
  (
    n457,
    n387
  );


  not
  g617
  (
    KeyWire_0_8,
    n306
  );


  not
  g618
  (
    n567,
    n286
  );


  buf
  g619
  (
    KeyWire_0_43,
    n291
  );


  not
  g620
  (
    n485,
    n345
  );


  not
  g621
  (
    n586,
    n380
  );


  not
  g622
  (
    n487,
    n345
  );


  not
  g623
  (
    n591,
    n363
  );


  not
  g624
  (
    n408,
    n364
  );


  buf
  g625
  (
    n702,
    n218
  );


  not
  g626
  (
    n596,
    n180
  );


  buf
  g627
  (
    n663,
    n158
  );


  not
  g628
  (
    n582,
    n230
  );


  buf
  g629
  (
    n626,
    n141
  );


  not
  g630
  (
    n545,
    n330
  );


  buf
  g631
  (
    n643,
    n164
  );


  not
  g632
  (
    n745,
    n216
  );


  not
  g633
  (
    n667,
    n115
  );


  buf
  g634
  (
    n622,
    n333
  );


  not
  g635
  (
    n484,
    n170
  );


  not
  g636
  (
    n653,
    n98
  );


  not
  g637
  (
    n721,
    n206
  );


  not
  g638
  (
    n480,
    n175
  );


  buf
  g639
  (
    n521,
    n302
  );


  not
  g640
  (
    n477,
    n168
  );


  buf
  g641
  (
    n403,
    n335
  );


  buf
  g642
  (
    n707,
    n340
  );


  not
  g643
  (
    n451,
    n365
  );


  not
  g644
  (
    n701,
    n256
  );


  buf
  g645
  (
    n601,
    n356
  );


  not
  g646
  (
    KeyWire_0_40,
    n365
  );


  not
  g647
  (
    n511,
    n348
  );


  buf
  g648
  (
    n411,
    n102
  );


  buf
  g649
  (
    n402,
    n383
  );


  buf
  g650
  (
    n443,
    n356
  );


  not
  g651
  (
    n431,
    n292
  );


  not
  g652
  (
    KeyWire_0_56,
    n316
  );


  buf
  g653
  (
    n565,
    n362
  );


  buf
  g654
  (
    n554,
    n284
  );


  not
  g655
  (
    n483,
    n351
  );


  not
  g656
  (
    n658,
    n130
  );


  not
  g657
  (
    n746,
    n378
  );


  buf
  g658
  (
    n519,
    n161
  );


  not
  g659
  (
    n749,
    n239
  );


  not
  g660
  (
    n559,
    n119
  );


  buf
  g661
  (
    n587,
    n207
  );


  not
  g662
  (
    n700,
    n382
  );


  not
  g663
  (
    n409,
    n159
  );


  not
  g664
  (
    n682,
    n194
  );


  buf
  g665
  (
    n433,
    n271
  );


  buf
  g666
  (
    n592,
    n358
  );


  not
  g667
  (
    n628,
    n343
  );


  not
  g668
  (
    n421,
    n128
  );


  not
  g669
  (
    n675,
    n382
  );


  buf
  g670
  (
    n593,
    n263
  );


  buf
  g671
  (
    n513,
    n339
  );


  not
  g672
  (
    n550,
    n362
  );


  not
  g673
  (
    n492,
    n103
  );


  not
  g674
  (
    n583,
    n184
  );


  not
  g675
  (
    n515,
    n247
  );


  buf
  g676
  (
    n427,
    n213
  );


  not
  g677
  (
    n478,
    n372
  );


  not
  g678
  (
    KeyWire_0_23,
    n296
  );


  not
  g679
  (
    n615,
    n167
  );


  buf
  g680
  (
    n608,
    n289
  );


  not
  g681
  (
    n425,
    n352
  );


  not
  g682
  (
    n435,
    n370
  );


  not
  g683
  (
    n562,
    n131
  );


  buf
  g684
  (
    n491,
    n265
  );


  not
  g685
  (
    n662,
    n360
  );


  buf
  g686
  (
    n570,
    n368
  );


  not
  g687
  (
    n547,
    n132
  );


  buf
  g688
  (
    n475,
    n337
  );


  not
  g689
  (
    n533,
    n217
  );


  not
  g690
  (
    KeyWire_0_30,
    n355
  );


  buf
  g691
  (
    n637,
    n244
  );


  buf
  g692
  (
    n563,
    n347
  );


  not
  g693
  (
    n644,
    n277
  );


  buf
  g694
  (
    n641,
    n358
  );


  buf
  g695
  (
    n649,
    n188
  );


  not
  g696
  (
    n605,
    n342
  );


  not
  g697
  (
    n531,
    n356
  );


  not
  g698
  (
    n407,
    n177
  );


  not
  g699
  (
    n719,
    n210
  );


  not
  g700
  (
    n585,
    n252
  );


  not
  g701
  (
    n509,
    n171
  );


  buf
  g702
  (
    n410,
    n349
  );


  not
  g703
  (
    n524,
    n287
  );


  buf
  g704
  (
    n490,
    n255
  );


  not
  g705
  (
    n652,
    n163
  );


  buf
  g706
  (
    n635,
    n383
  );


  not
  g707
  (
    n735,
    n363
  );


  not
  g708
  (
    n619,
    n303
  );


  buf
  g709
  (
    n557,
    n377
  );


  not
  g710
  (
    n406,
    n384
  );


  buf
  g711
  (
    n671,
    n135
  );


  buf
  g712
  (
    n486,
    n309
  );


  not
  g713
  (
    n472,
    n237
  );


  buf
  g714
  (
    n654,
    n374
  );


  or
  g715
  (
    n462,
    n389,
    n295,
    n355,
    n127
  );


  nand
  g716
  (
    n438,
    n151,
    n362,
    n179,
    n233
  );


  xnor
  g717
  (
    n468,
    n120,
    n367,
    n386,
    n310
  );


  and
  g718
  (
    n446,
    n219,
    n350,
    n370,
    n304
  );


  and
  g719
  (
    n693,
    n377,
    n374,
    n270,
    n266
  );


  and
  g720
  (
    n687,
    n262,
    n375,
    n193,
    n173
  );


  nor
  g721
  (
    n552,
    n278,
    n209,
    n124,
    n195
  );


  or
  g722
  (
    n569,
    n387,
    n234,
    n172,
    n389
  );


  nand
  g723
  (
    n404,
    n112,
    n176,
    n348,
    n297
  );


  xnor
  g724
  (
    n725,
    n222,
    n182,
    n326,
    n294
  );


  xnor
  g725
  (
    n617,
    n122,
    n100,
    n146,
    n235
  );


  nand
  g726
  (
    n696,
    n113,
    n197,
    n346,
    n317
  );


  xnor
  g727
  (
    n716,
    n373,
    n371,
    n111,
    n346
  );


  nand
  g728
  (
    n576,
    n371,
    n385,
    n212,
    n363
  );


  nand
  g729
  (
    n724,
    n229,
    n109,
    n388,
    n340
  );


  nand
  g730
  (
    n551,
    n364,
    n343,
    n354,
    n371
  );


  xnor
  g731
  (
    n754,
    n433,
    n480,
    n439,
    n502
  );


  and
  g732
  (
    n760,
    n469,
    n495,
    n478,
    n421
  );


  and
  g733
  (
    n767,
    n509,
    n526,
    n504,
    n527
  );


  nor
  g734
  (
    n777,
    n416,
    n473,
    n459,
    n520
  );


  nand
  g735
  (
    n753,
    n529,
    n420,
    n506,
    n419
  );


  nor
  g736
  (
    n765,
    n496,
    n524,
    n413,
    n431
  );


  nand
  g737
  (
    n758,
    n513,
    n514,
    n485,
    n501
  );


  or
  g738
  (
    n771,
    n487,
    n425,
    n445,
    n522
  );


  and
  g739
  (
    n768,
    n517,
    n458,
    n424,
    n508
  );


  xnor
  g740
  (
    n751,
    n484,
    n400,
    n523,
    n452
  );


  and
  g741
  (
    n757,
    n482,
    n438,
    n455,
    n410
  );


  and
  g742
  (
    n772,
    n449,
    n494,
    n491,
    n462
  );


  xnor
  g743
  (
    n755,
    n446,
    n476,
    n401,
    n479
  );


  xnor
  g744
  (
    n759,
    n407,
    n515,
    n481,
    n429
  );


  and
  g745
  (
    n761,
    n486,
    n456,
    n464,
    n411
  );


  or
  g746
  (
    n781,
    n519,
    n525,
    n500,
    n426
  );


  xor
  g747
  (
    n778,
    n471,
    n403,
    n448,
    n460
  );


  xor
  g748
  (
    n773,
    n530,
    n470,
    n477,
    n443
  );


  nor
  g749
  (
    n775,
    n488,
    n434,
    n518,
    n512
  );


  nand
  g750
  (
    n756,
    n427,
    n467,
    n493,
    n475
  );


  nor
  g751
  (
    n769,
    n447,
    n503,
    n505,
    n441
  );


  and
  g752
  (
    n776,
    n414,
    n440,
    n406,
    n490
  );


  xor
  g753
  (
    n766,
    n450,
    n428,
    n474,
    n528
  );


  nor
  g754
  (
    n752,
    n489,
    n498,
    n417,
    n451
  );


  nand
  g755
  (
    n770,
    n453,
    n466,
    n454,
    n497
  );


  nand
  g756
  (
    n779,
    n408,
    n405,
    n442,
    n510
  );


  nor
  g757
  (
    n782,
    n444,
    n507,
    n492,
    n465
  );


  xor
  g758
  (
    n774,
    n472,
    n511,
    n432,
    n483
  );


  or
  g759
  (
    n783,
    n516,
    n415,
    n521,
    n499
  );


  nor
  g760
  (
    n763,
    n436,
    n461,
    n422,
    n457
  );


  nand
  g761
  (
    n762,
    n463,
    n430,
    n399,
    n412
  );


  and
  g762
  (
    n764,
    n423,
    n468,
    n402,
    n418
  );


  and
  g763
  (
    n780,
    n409,
    n435,
    n437,
    n404
  );


  or
  g764
  (
    n812,
    n553,
    n545,
    n591,
    n574
  );


  xor
  g765
  (
    n796,
    n609,
    n758,
    n778,
    n589
  );


  nand
  g766
  (
    n802,
    n606,
    n623,
    n780,
    n611
  );


  or
  g767
  (
    n787,
    n766,
    n603,
    n575,
    n626
  );


  and
  g768
  (
    n785,
    n586,
    n578,
    n579,
    n563
  );


  xnor
  g769
  (
    n795,
    n543,
    n617,
    n776,
    n584
  );


  and
  g770
  (
    n814,
    n752,
    n595,
    n567,
    n583
  );


  xor
  g771
  (
    n804,
    n544,
    n767,
    n756,
    n592
  );


  and
  g772
  (
    n811,
    n775,
    n624,
    n546,
    n548
  );


  or
  g773
  (
    n792,
    n618,
    n601,
    n533,
    n572
  );


  nand
  g774
  (
    n808,
    n566,
    n772,
    n612,
    n588
  );


  xnor
  g775
  (
    n789,
    n620,
    n764,
    n607,
    n569
  );


  xnor
  g776
  (
    n784,
    n759,
    n549,
    n762,
    n757
  );


  or
  g777
  (
    n810,
    n550,
    n782,
    n777,
    n753
  );


  xnor
  g778
  (
    n809,
    n577,
    n593,
    n604,
    n568
  );


  or
  g779
  (
    n800,
    n608,
    n561,
    n783,
    n538
  );


  and
  g780
  (
    n801,
    n769,
    n770,
    n570,
    n536
  );


  xor
  g781
  (
    n807,
    n754,
    n555,
    n779,
    n773
  );


  xnor
  g782
  (
    n815,
    n594,
    n587,
    n547,
    n534
  );


  xnor
  g783
  (
    n793,
    n613,
    n616,
    n560,
    n576
  );


  nand
  g784
  (
    KeyWire_0_36,
    n597,
    n622,
    n571,
    n581
  );


  xor
  g785
  (
    n794,
    n539,
    n556,
    n541,
    n559
  );


  xor
  g786
  (
    n788,
    n552,
    n771,
    n573,
    n535
  );


  nand
  g787
  (
    n803,
    n781,
    n557,
    n760,
    n619
  );


  and
  g788
  (
    n805,
    n598,
    n554,
    n537,
    n602
  );


  nand
  g789
  (
    n786,
    n605,
    n551,
    n614,
    n585
  );


  and
  g790
  (
    n799,
    n540,
    n564,
    n558,
    n582
  );


  nand
  g791
  (
    n790,
    n768,
    n755,
    n531,
    n625
  );


  and
  g792
  (
    n791,
    n600,
    n532,
    n580,
    n763
  );


  and
  g793
  (
    n797,
    n774,
    n621,
    n761,
    n610
  );


  or
  g794
  (
    n806,
    n565,
    n562,
    n615,
    n599
  );


  or
  g795
  (
    n798,
    n542,
    n765,
    n596,
    n590
  );


  buf
  g796
  (
    n843,
    n805
  );


  buf
  g797
  (
    n830,
    n798
  );


  buf
  g798
  (
    n838,
    n788
  );


  buf
  g799
  (
    n850,
    n800
  );


  not
  g800
  (
    n840,
    n801
  );


  buf
  g801
  (
    n837,
    n804
  );


  not
  g802
  (
    n819,
    n796
  );


  not
  g803
  (
    n845,
    n802
  );


  buf
  g804
  (
    n853,
    n789
  );


  not
  g805
  (
    n820,
    n802
  );


  buf
  g806
  (
    n832,
    n786
  );


  buf
  g807
  (
    n839,
    n800
  );


  buf
  g808
  (
    n821,
    n794
  );


  not
  g809
  (
    n855,
    n808
  );


  buf
  g810
  (
    n828,
    n805
  );


  not
  g811
  (
    n856,
    n790
  );


  buf
  g812
  (
    n834,
    n801
  );


  buf
  g813
  (
    n844,
    n795
  );


  not
  g814
  (
    n859,
    n797
  );


  not
  g815
  (
    n842,
    n806
  );


  not
  g816
  (
    n816,
    n796
  );


  buf
  g817
  (
    n846,
    n810
  );


  buf
  g818
  (
    n848,
    n786
  );


  not
  g819
  (
    n825,
    n804
  );


  xor
  g820
  (
    n818,
    n795,
    n793,
    n785,
    n807
  );


  nor
  g821
  (
    n857,
    n798,
    n786,
    n791,
    n803
  );


  xor
  g822
  (
    n824,
    n791,
    n788,
    n809
  );


  xor
  g823
  (
    KeyWire_0_62,
    n809,
    n787,
    n784,
    n803
  );


  or
  g824
  (
    n858,
    n794,
    n794,
    n801,
    n807
  );


  and
  g825
  (
    n831,
    n785,
    n806,
    n791,
    n810
  );


  nor
  g826
  (
    n827,
    n802,
    n806,
    n795,
    n797
  );


  xor
  g827
  (
    n860,
    n790,
    n788,
    n784,
    n792
  );


  or
  g828
  (
    n836,
    n808,
    n799,
    n798,
    n793
  );


  nand
  g829
  (
    n823,
    n806,
    n785,
    n810,
    n790
  );


  xnor
  g830
  (
    n849,
    n785,
    n796,
    n789,
    n791
  );


  nor
  g831
  (
    n841,
    n804,
    n809,
    n801,
    n786
  );


  or
  g832
  (
    n822,
    n803,
    n799,
    n794,
    n792
  );


  xnor
  g833
  (
    KeyWire_0_21,
    n792,
    n784,
    n807
  );


  xnor
  g834
  (
    n852,
    n800,
    n799,
    n808,
    n789
  );


  and
  g835
  (
    n833,
    n793,
    n803,
    n799,
    n804
  );


  or
  g836
  (
    n835,
    n807,
    n805,
    n810,
    n797
  );


  xnor
  g837
  (
    n847,
    n805,
    n798,
    n787,
    n808
  );


  or
  g838
  (
    n817,
    n797,
    n790,
    n787,
    n792
  );


  xnor
  g839
  (
    n826,
    n802,
    n809,
    n796,
    n793
  );


  nor
  g840
  (
    n851,
    n787,
    n789,
    n800,
    n795
  );


  not
  g841
  (
    n864,
    n832
  );


  buf
  g842
  (
    n867,
    n824
  );


  not
  g843
  (
    n874,
    n823
  );


  buf
  g844
  (
    n876,
    n825
  );


  buf
  g845
  (
    n879,
    n826
  );


  not
  g846
  (
    n877,
    n828
  );


  not
  g847
  (
    n875,
    n817
  );


  buf
  g848
  (
    n863,
    n822
  );


  not
  g849
  (
    n861,
    n835
  );


  not
  g850
  (
    n873,
    n819
  );


  not
  g851
  (
    n880,
    n818
  );


  not
  g852
  (
    n868,
    n827
  );


  buf
  g853
  (
    n870,
    n820
  );


  not
  g854
  (
    n865,
    n829
  );


  buf
  g855
  (
    n878,
    n830
  );


  buf
  g856
  (
    n866,
    n834
  );


  buf
  g857
  (
    n871,
    n831
  );


  not
  g858
  (
    n872,
    n816
  );


  not
  g859
  (
    n862,
    n833
  );


  buf
  g860
  (
    n869,
    n821
  );


  not
  g861
  (
    n882,
    n868
  );


  buf
  g862
  (
    n886,
    n874
  );


  buf
  g863
  (
    n895,
    n866
  );


  not
  g864
  (
    n893,
    n863
  );


  buf
  g865
  (
    n897,
    n870
  );


  buf
  g866
  (
    n898,
    n864
  );


  buf
  g867
  (
    KeyWire_0_6,
    n873
  );


  buf
  g868
  (
    n885,
    n873
  );


  not
  g869
  (
    n892,
    n861
  );


  not
  g870
  (
    n894,
    n870
  );


  not
  g871
  (
    n896,
    n869
  );


  buf
  g872
  (
    n884,
    n867
  );


  not
  g873
  (
    n881,
    n862
  );


  not
  g874
  (
    n888,
    n872
  );


  not
  g875
  (
    n887,
    n872
  );


  not
  g876
  (
    KeyWire_0_0,
    n871
  );


  not
  g877
  (
    KeyWire_0_39,
    n865
  );


  not
  g878
  (
    n889,
    n871
  );


  not
  g879
  (
    n938,
    n896
  );


  buf
  g880
  (
    n950,
    n889
  );


  not
  g881
  (
    n932,
    n875
  );


  not
  g882
  (
    n934,
    n883
  );


  not
  g883
  (
    n918,
    n885
  );


  not
  g884
  (
    n926,
    n889
  );


  buf
  g885
  (
    n953,
    n892
  );


  buf
  g886
  (
    KeyWire_0_31,
    n893
  );


  buf
  g887
  (
    n946,
    n890
  );


  not
  g888
  (
    n903,
    n887
  );


  buf
  g889
  (
    n941,
    n886
  );


  not
  g890
  (
    n900,
    n886
  );


  buf
  g891
  (
    n925,
    n883
  );


  buf
  g892
  (
    n930,
    n887
  );


  buf
  g893
  (
    n921,
    n893
  );


  not
  g894
  (
    n949,
    n897
  );


  not
  g895
  (
    n937,
    n891
  );


  not
  g896
  (
    n924,
    n898
  );


  not
  g897
  (
    n913,
    n888
  );


  buf
  g898
  (
    n951,
    n882
  );


  buf
  g899
  (
    n919,
    n882
  );


  buf
  g900
  (
    KeyWire_0_9,
    n888
  );


  not
  g901
  (
    n948,
    n881
  );


  not
  g902
  (
    n911,
    n893
  );


  buf
  g903
  (
    n909,
    n881
  );


  buf
  g904
  (
    n929,
    n874
  );


  buf
  g905
  (
    n905,
    n886
  );


  buf
  g906
  (
    n935,
    n895
  );


  not
  g907
  (
    n923,
    n885
  );


  not
  g908
  (
    n943,
    n897
  );


  not
  g909
  (
    n942,
    n890
  );


  not
  g910
  (
    n917,
    n876
  );


  buf
  g911
  (
    n899,
    n889
  );


  not
  g912
  (
    n933,
    n892
  );


  buf
  g913
  (
    n939,
    n884
  );


  not
  g914
  (
    n904,
    n896
  );


  buf
  g915
  (
    n947,
    n875
  );


  not
  g916
  (
    n902,
    n898
  );


  buf
  g917
  (
    n944,
    n876
  );


  not
  g918
  (
    n914,
    n891
  );


  not
  g919
  (
    n927,
    n898
  );


  buf
  g920
  (
    n922,
    n887
  );


  not
  g921
  (
    n931,
    n895
  );


  buf
  g922
  (
    n952,
    n894
  );


  buf
  g923
  (
    n912,
    n882
  );


  not
  g924
  (
    n915,
    n888
  );


  not
  g925
  (
    n910,
    n894
  );


  buf
  g926
  (
    n936,
    n892
  );


  buf
  g927
  (
    n906,
    n884
  );


  not
  g928
  (
    n901,
    n896
  );


  buf
  g929
  (
    n908,
    n895
  );


  buf
  g930
  (
    n916,
    n885
  );


  not
  g931
  (
    n945,
    n894
  );


  nand
  g932
  (
    n940,
    n890,
    n891,
    n881
  );


  xor
  g933
  (
    n920,
    n897,
    n884,
    n898,
    n883
  );


  nand
  g934
  (
    n967,
    n926,
    n919,
    n904,
    n910
  );


  and
  g935
  (
    n964,
    n928,
    n918,
    n906,
    n923
  );


  and
  g936
  (
    n957,
    n916,
    n917,
    n926,
    n902
  );


  xor
  g937
  (
    n954,
    n911,
    n907,
    n913,
    n899
  );


  and
  g938
  (
    KeyWire_0_37,
    n914,
    n927,
    n916,
    n929
  );


  xor
  g939
  (
    n956,
    n904,
    n900,
    n905,
    n920
  );


  xor
  g940
  (
    n965,
    n899,
    n925,
    n908,
    n906
  );


  or
  g941
  (
    n966,
    n907,
    n925,
    n914,
    n931
  );


  and
  g942
  (
    n955,
    n932,
    n902,
    n912,
    n901
  );


  xor
  g943
  (
    n970,
    n910,
    n920,
    n931,
    n919
  );


  and
  g944
  (
    KeyWire_0_63,
    n915,
    n913,
    n927,
    n912
  );


  nand
  g945
  (
    n968,
    n930,
    n930,
    n909,
    n911
  );


  nor
  g946
  (
    n962,
    n900,
    n903,
    n915,
    n917
  );


  nand
  g947
  (
    n958,
    n932,
    n901,
    n928,
    n929
  );


  xnor
  g948
  (
    n961,
    n905,
    n918,
    n903,
    n921
  );


  nand
  g949
  (
    n969,
    n909,
    n921,
    n923,
    n922
  );


  or
  g950
  (
    n959,
    n908,
    n924,
    n922
  );


  buf
  g951
  (
    n971,
    n957
  );


  buf
  g952
  (
    n974,
    n954
  );


  not
  g953
  (
    n972,
    n955
  );


  not
  g954
  (
    n973,
    n956
  );


  xnor
  g955
  (
    n975,
    n971,
    n971,
    n967,
    n974
  );


  xnor
  g956
  (
    n985,
    n391,
    n966,
    n396,
    n965
  );


  and
  g957
  (
    n983,
    n973,
    n974,
    n971,
    n878
  );


  xor
  g958
  (
    n981,
    n974,
    n960,
    n392
  );


  xor
  g959
  (
    n990,
    n973,
    n974,
    n395,
    n971
  );


  xnor
  g960
  (
    n988,
    n393,
    n972,
    n395
  );


  nand
  g961
  (
    n984,
    n812,
    n392,
    n972,
    n393
  );


  xor
  g962
  (
    n980,
    n393,
    n878,
    n812,
    n811
  );


  xor
  g963
  (
    n978,
    n972,
    n630,
    n629,
    n811
  );


  and
  g964
  (
    n987,
    n812,
    n877,
    n811,
    n933
  );


  xnor
  g965
  (
    n989,
    n962,
    n396,
    n973,
    n395
  );


  nand
  g966
  (
    n982,
    n877,
    n961,
    n964,
    n969
  );


  nand
  g967
  (
    n977,
    n631,
    n879,
    n394,
    n811
  );


  or
  g968
  (
    n986,
    n394,
    n973,
    n963,
    n397
  );


  xor
  g969
  (
    n976,
    n959,
    n968,
    n396,
    n958
  );


  xor
  g970
  (
    n979,
    n970,
    n628,
    n394,
    n627
  );


  or
  g971
  (
    n1050,
    n648,
    n989,
    n710,
    n979
  );


  xnor
  g972
  (
    n1022,
    n977,
    n983,
    n666,
    n684
  );


  or
  g973
  (
    n1026,
    n698,
    n688,
    n879,
    n686
  );


  xor
  g974
  (
    KeyWire_0_14,
    n661,
    n851,
    n986,
    n978
  );


  and
  g975
  (
    n998,
    n669,
    n697,
    n683,
    n646
  );


  and
  g976
  (
    n1008,
    n939,
    n986,
    n95,
    n815
  );


  nor
  g977
  (
    n1023,
    n691,
    n938,
    n981,
    n934
  );


  and
  g978
  (
    n1018,
    n744,
    n815,
    n681,
    n814
  );


  xnor
  g979
  (
    n1054,
    n651,
    n977,
    n838,
    n983
  );


  or
  g980
  (
    n1005,
    n741,
    n937,
    n846,
    n702
  );


  nor
  g981
  (
    KeyWire_0_3,
    n813,
    n990,
    n842,
    n978
  );


  or
  g982
  (
    n992,
    n935,
    n654,
    n855,
    n976
  );


  and
  g983
  (
    n1035,
    n397,
    n985,
    n662,
    n841
  );


  and
  g984
  (
    n1028,
    n655,
    n987,
    n849,
    n978
  );


  nor
  g985
  (
    n1048,
    n658,
    n656,
    n732,
    n843
  );


  nand
  g986
  (
    n1027,
    n986,
    n815,
    n975,
    n671
  );


  and
  g987
  (
    n1000,
    n712,
    n984,
    n728,
    n689
  );


  nand
  g988
  (
    n1030,
    n736,
    n980,
    n636,
    n988
  );


  or
  g989
  (
    n1047,
    n659,
    n660,
    n981,
    n976
  );


  xnor
  g990
  (
    n1036,
    n982,
    n944,
    n813,
    n977
  );


  nand
  g991
  (
    n1031,
    n679,
    n813,
    n853,
    n990
  );


  xnor
  g992
  (
    n1024,
    n943,
    n632,
    n694,
    n980
  );


  xnor
  g993
  (
    n994,
    n937,
    n717,
    n680,
    n747
  );


  nand
  g994
  (
    n999,
    n750,
    n701,
    n734,
    n722
  );


  or
  g995
  (
    n1034,
    n715,
    n976,
    n941,
    n668
  );


  xor
  g996
  (
    n1044,
    n936,
    n988,
    n721,
    n985
  );


  nor
  g997
  (
    KeyWire_0_11,
    n638,
    n735,
    n719,
    n738
  );


  nand
  g998
  (
    n1051,
    n985,
    n707,
    n645,
    n814
  );


  and
  g999
  (
    n1012,
    n988,
    n685,
    n979,
    n672
  );


  xor
  g1000
  (
    n1052,
    n975,
    n398,
    n649
  );


  nand
  g1001
  (
    n1014,
    n637,
    n983,
    n844,
    n988
  );


  nand
  g1002
  (
    n995,
    n980,
    n731,
    n982,
    n700
  );


  xor
  g1003
  (
    n1025,
    n814,
    n852,
    n644,
    n714
  );


  or
  g1004
  (
    n1032,
    n989,
    n639,
    n837,
    n749
  );


  nor
  g1005
  (
    n1010,
    n979,
    n980,
    n984,
    n812
  );


  nand
  g1006
  (
    n1017,
    n858,
    n946,
    n641,
    n720
  );


  or
  g1007
  (
    n1019,
    n941,
    n942,
    n705,
    n981
  );


  and
  g1008
  (
    n1045,
    n938,
    n746,
    n989,
    n990
  );


  or
  g1009
  (
    n1021,
    n984,
    n836,
    n982,
    n675
  );


  nor
  g1010
  (
    n1049,
    n987,
    n860,
    n989,
    n737
  );


  and
  g1011
  (
    n1002,
    n730,
    n667,
    n983,
    n703
  );


  xnor
  g1012
  (
    n997,
    n665,
    n944,
    n742,
    n642
  );


  and
  g1013
  (
    n1038,
    n945,
    n985,
    n723,
    n740
  );


  xor
  g1014
  (
    n993,
    n936,
    n946,
    n633,
    n945
  );


  or
  g1015
  (
    n1029,
    n690,
    n942,
    n978,
    n848
  );


  nor
  g1016
  (
    n1037,
    n673,
    n854,
    n724,
    n981
  );


  nand
  g1017
  (
    n1003,
    n711,
    n934,
    n856,
    n634
  );


  xnor
  g1018
  (
    n1013,
    n696,
    n726,
    n814,
    n713
  );


  or
  g1019
  (
    KeyWire_0_24,
    n975,
    n682,
    n397,
    n987
  );


  xnor
  g1020
  (
    n1041,
    n725,
    n743,
    n990,
    n933
  );


  xor
  g1021
  (
    n1040,
    n940,
    n745,
    n739,
    n706
  );


  or
  g1022
  (
    n996,
    n678,
    n815,
    n845,
    n733
  );


  nor
  g1023
  (
    n1020,
    n704,
    n687,
    n670,
    n748
  );


  and
  g1024
  (
    n1016,
    n813,
    n664,
    n943,
    n709
  );


  xor
  g1025
  (
    n1009,
    n699,
    n940,
    n986,
    n663
  );


  xnor
  g1026
  (
    n1053,
    n946,
    n643,
    n987,
    n653
  );


  xor
  g1027
  (
    n1046,
    n939,
    n647,
    n859,
    n979
  );


  and
  g1028
  (
    n1007,
    n635,
    n976,
    n984,
    n982
  );


  nand
  g1029
  (
    n991,
    n657,
    n716,
    n729,
    n727
  );


  or
  g1030
  (
    n1043,
    n708,
    n650,
    n695,
    n975
  );


  nor
  g1031
  (
    n1015,
    n718,
    n839,
    n935,
    n847
  );


  xor
  g1032
  (
    n1004,
    n677,
    n676,
    n693,
    n850
  );


  xor
  g1033
  (
    n1001,
    n857,
    n674,
    n652,
    n692
  );


  and
  g1034
  (
    n1042,
    n840,
    n640,
    n977,
    n945
  );


  xor
  g1035
  (
    n1058,
    n1023,
    n948,
    n1008,
    n1028
  );


  nor
  g1036
  (
    n1060,
    n1038,
    n1053,
    n999,
    n1045
  );


  nor
  g1037
  (
    n1057,
    n1009,
    n947,
    n1043,
    n1046
  );


  and
  g1038
  (
    n1070,
    n992,
    n1037,
    n951,
    n952
  );


  and
  g1039
  (
    n1073,
    n1001,
    n1027,
    n1050,
    n1051
  );


  nor
  g1040
  (
    n1066,
    n1035,
    n947,
    n998,
    n948
  );


  xnor
  g1041
  (
    n1076,
    n1014,
    n1021,
    n1026,
    n1025
  );


  xor
  g1042
  (
    n1065,
    n1042,
    n949,
    n1017,
    n1034
  );


  xor
  g1043
  (
    n1072,
    n948,
    n950,
    n1012
  );


  nor
  g1044
  (
    n1067,
    n1039,
    n398,
    n952,
    n1004
  );


  or
  g1045
  (
    n1055,
    n1054,
    n949,
    n1030,
    n996
  );


  nand
  g1046
  (
    n1064,
    n952,
    n949,
    n953,
    n1011
  );


  xor
  g1047
  (
    n1063,
    n880,
    n1016,
    n1013,
    n1019
  );


  xnor
  g1048
  (
    n1075,
    n1036,
    n1010,
    n1040,
    n947
  );


  nor
  g1049
  (
    n1061,
    n1031,
    n1033,
    n1006,
    n1000
  );


  or
  g1050
  (
    n1059,
    n953,
    n880,
    n994,
    n1015
  );


  or
  g1051
  (
    n1068,
    n1022,
    n1032,
    n1020,
    n995
  );


  or
  g1052
  (
    n1074,
    n1049,
    n1005,
    n1041,
    n1024
  );


  nand
  g1053
  (
    n1071,
    n1029,
    n1048,
    n953,
    n1018
  );


  and
  g1054
  (
    n1069,
    n1047,
    n993,
    n1044,
    n1002
  );


  xor
  g1055
  (
    n1062,
    n950,
    n951,
    n997
  );


  nand
  g1056
  (
    n1056,
    n1003,
    n1052,
    n1007,
    n991
  );


  xnor
  KeyGate_0_0
  (
    n890,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n254,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n305,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1011,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n448,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n181,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n883,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n469,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n730,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n907,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n111,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1039,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n396,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n332,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1006,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n199,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n532,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n125,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n497,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n388,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n86,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n829,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n363,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n534,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n1033,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n233,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n496,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n638,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n176,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n502,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n453,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n928,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n100,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n320,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n50,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n282,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n813,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n960,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n299,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n891,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n415,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n180,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n594,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n505,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n378,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n246,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n55,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n748,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n574,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n458,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n606,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n211,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n556,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n382,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n54,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n253,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n686,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n225,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n124,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n479,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n544,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n501,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n854,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n963,
    KeyNOTWire_0_63
  );


endmodule

