// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_46 written by SynthGen on 2021/04/05 11:08:37
module Stat_100_46( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n70, n69, n120, n102, n121, n106, n108, n112,
 n114, n109, n85, n83, n94, n111, n99, n115,
 n92, n116, n89, n86, n110, n119, n125, n123,
 n127, n131, n128, n126, n124, n132, n130, n129);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n70, n69, n120, n102, n121, n106, n108, n112,
 n114, n109, n85, n83, n94, n111, n99, n115,
 n92, n116, n89, n86, n110, n119, n125, n123,
 n127, n131, n128, n126, n124, n132, n130, n129;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n84, n87, n88, n90, n91, n93, n95, n96,
 n97, n98, n100, n101, n103, n104, n105, n107,
 n113, n117, n118, n122;

buf  g0 (n42, n3);
not  g1 (n35, n1);
not  g2 (n43, n10);
not  g3 (n36, n5);
buf  g4 (n37, n4);
buf  g5 (n40, n9);
buf  g6 (n33, n7);
not  g7 (n41, n6);
buf  g8 (n39, n2);
not  g9 (n34, n11);
not  g10 (n38, n8);
not  g11 (n48, n36);
buf  g12 (n55, n35);
buf  g13 (n56, n37);
not  g14 (n63, n36);
buf  g15 (n71, n43);
buf  g16 (n62, n41);
buf  g17 (n70, n41);
not  g18 (n57, n34);
not  g19 (n68, n42);
buf  g20 (n64, n38);
not  g21 (n59, n35);
buf  g22 (n75, n38);
not  g23 (n47, n41);
buf  g24 (n74, n39);
buf  g25 (n45, n43);
buf  g26 (n73, n39);
not  g27 (n44, n36);
not  g28 (n81, n40);
buf  g29 (n78, n37);
buf  g30 (n79, n43);
buf  g31 (n69, n42);
not  g32 (n61, n35);
buf  g33 (n49, n35);
not  g34 (n51, n38);
buf  g35 (n76, n37);
not  g36 (n60, n34);
not  g37 (n80, n38);
buf  g38 (n65, n34);
not  g39 (n50, n42);
buf  g40 (n46, n41);
buf  g41 (n82, n36);
buf  g42 (n66, n39);
buf  g43 (n72, n39);
buf  g44 (n54, n43);
buf  g45 (n77, n34);
buf  g46 (n58, n37);
not  g47 (n67, n40);
buf  g48 (n52, n42);
buf  g49 (n53, n40);
not  g50 (n110, n70);
buf  g51 (n91, n56);
xor  g52 (n95, n55, n72, n71);
nor  g53 (n108, n77, n82, n69, n65);
nor  g54 (n109, n46, n63, n60, n77);
xor  g55 (n84, n46, n66, n58, n71);
xnor g56 (n86, n78, n77, n50);
or   g57 (n83, n61, n47, n62, n68);
or   g58 (n98, n79, n78, n55, n50);
or   g59 (n104, n57, n81, n68);
nor  g60 (n93, n78, n76, n79, n61);
nor  g61 (n101, n62, n73, n55, n57);
xnor g62 (n119, n70, n56, n49, n48);
xor  g63 (n85, n59, n56, n80, n58);
and  g64 (n105, n67, n64, n81, n62);
xnor g65 (n120, n75, n70, n60, n63);
or   g66 (n100, n79, n81, n51, n54);
or   g67 (n117, n64, n59, n74, n82);
or   g68 (n122, n64, n76, n75, n73);
xnor g69 (n99, n55, n75, n59, n64);
nand g70 (n112, n48, n79, n71, n69);
xor  g71 (n121, n57, n45, n49, n73);
or   g72 (n116, n72, n80, n62, n74);
xnor g73 (n118, n75, n60, n45, n69);
or   g74 (n113, n49, n51, n53);
xor  g75 (n92, n65, n47, n51, n66);
nor  g76 (n89, n54, n54, n82, n50);
and  g77 (n90, n80, n66, n57);
xor  g78 (n106, n53, n50, n47, n12);
xnor g79 (n114, n72, n82, n61, n63);
xor  g80 (n111, n65, n49, n76, n60);
nand g81 (n96, n45, n71, n48, n47);
or   g82 (n97, n58, n67, n53, n61);
or   g83 (n107, n67, n46, n69, n45);
or   g84 (n88, n76, n52, n73);
nor  g85 (n115, n78, n56, n58, n68);
nand g86 (n102, n59, n74, n80, n54);
xnor g87 (n87, n74, n65, n52, n70);
xnor g88 (n94, n48, n68, n53, n67);
nand g89 (n103, n52, n72, n46, n63);
xnor g90 (n126, n13, n105, n108, n110);
nor  g91 (n129, n115, n24, n119, n19);
nand g92 (n124, n30, n113, n104, n28);
nor  g93 (n123, n114, n25, n111, n109);
or   g94 (n130, n122, n117, n29, n15);
nand g95 (n131, n120, n14, n103, n16);
or   g96 (n128, n112, n17, n26, n121);
xor  g97 (n127, n31, n20, n21, n23);
or   g98 (n132, n107, n116, n106, n118);
and  g99 (n125, n27, n22, n32, n18);
endmodule
