

module Stat_913_268
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n681,
  n686,
  n684,
  n682,
  n690,
  n693,
  n696,
  n692,
  n691,
  n699,
  n695,
  n698,
  n865,
  n943,
  n938,
  n945,
  n941,
  n940,
  n937,
  n942,
  n935,
  n936,
  n939,
  n944
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n681;output n686;output n684;output n682;output n690;output n693;output n696;output n692;output n691;output n699;output n695;output n698;output n865;output n943;output n938;output n945;output n941;output n940;output n937;output n942;output n935;output n936;output n939;output n944;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n683;wire n685;wire n687;wire n688;wire n689;wire n694;wire n697;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;

  buf
  g0
  (
    n157,
    n10
  );


  not
  g1
  (
    n94,
    n26
  );


  buf
  g2
  (
    n121,
    n1
  );


  not
  g3
  (
    n125,
    n21
  );


  buf
  g4
  (
    n47,
    n27
  );


  buf
  g5
  (
    n151,
    n15
  );


  not
  g6
  (
    n37,
    n29
  );


  buf
  g7
  (
    n111,
    n25
  );


  buf
  g8
  (
    n80,
    n18
  );


  not
  g9
  (
    KeyWire_0_1,
    n31
  );


  not
  g10
  (
    n128,
    n28
  );


  not
  g11
  (
    n103,
    n30
  );


  not
  g12
  (
    n150,
    n14
  );


  not
  g13
  (
    n38,
    n5
  );


  not
  g14
  (
    n105,
    n23
  );


  not
  g15
  (
    n132,
    n15
  );


  buf
  g16
  (
    KeyWire_0_10,
    n6
  );


  not
  g17
  (
    n137,
    n26
  );


  not
  g18
  (
    n41,
    n24
  );


  not
  g19
  (
    n81,
    n12
  );


  not
  g20
  (
    n99,
    n4
  );


  not
  g21
  (
    n88,
    n23
  );


  not
  g22
  (
    n71,
    n32
  );


  not
  g23
  (
    n139,
    n15
  );


  not
  g24
  (
    n146,
    n6
  );


  buf
  g25
  (
    n98,
    n28
  );


  buf
  g26
  (
    n122,
    n3
  );


  buf
  g27
  (
    n54,
    n29
  );


  buf
  g28
  (
    n113,
    n21
  );


  not
  g29
  (
    n66,
    n11
  );


  buf
  g30
  (
    n119,
    n25
  );


  not
  g31
  (
    n69,
    n16
  );


  buf
  g32
  (
    n110,
    n7
  );


  not
  g33
  (
    n72,
    n14
  );


  buf
  g34
  (
    n44,
    n10
  );


  buf
  g35
  (
    n90,
    n28
  );


  buf
  g36
  (
    n148,
    n19
  );


  not
  g37
  (
    n63,
    n22
  );


  buf
  g38
  (
    n67,
    n28
  );


  buf
  g39
  (
    n89,
    n12
  );


  not
  g40
  (
    n97,
    n31
  );


  not
  g41
  (
    n65,
    n31
  );


  not
  g42
  (
    n142,
    n10
  );


  not
  g43
  (
    n33,
    n18
  );


  buf
  g44
  (
    n159,
    n9
  );


  buf
  g45
  (
    n73,
    n1
  );


  not
  g46
  (
    n87,
    n9
  );


  not
  g47
  (
    n149,
    n5
  );


  buf
  g48
  (
    n102,
    n14
  );


  not
  g49
  (
    n61,
    n24
  );


  not
  g50
  (
    n147,
    n13
  );


  buf
  g51
  (
    n108,
    n7
  );


  buf
  g52
  (
    n124,
    n13
  );


  buf
  g53
  (
    n93,
    n5
  );


  not
  g54
  (
    n43,
    n25
  );


  not
  g55
  (
    n153,
    n29
  );


  not
  g56
  (
    n145,
    n21
  );


  not
  g57
  (
    n130,
    n11
  );


  buf
  g58
  (
    n135,
    n32
  );


  buf
  g59
  (
    n158,
    n14
  );


  not
  g60
  (
    n64,
    n8
  );


  not
  g61
  (
    n106,
    n27
  );


  buf
  g62
  (
    n136,
    n8
  );


  buf
  g63
  (
    n129,
    n3
  );


  not
  g64
  (
    n50,
    n30
  );


  not
  g65
  (
    n49,
    n15
  );


  not
  g66
  (
    n144,
    n20
  );


  buf
  g67
  (
    n74,
    n27
  );


  not
  g68
  (
    n82,
    n18
  );


  not
  g69
  (
    n95,
    n24
  );


  buf
  g70
  (
    n115,
    n4
  );


  not
  g71
  (
    n116,
    n32
  );


  not
  g72
  (
    n83,
    n7
  );


  not
  g73
  (
    n48,
    n18
  );


  not
  g74
  (
    n91,
    n8
  );


  not
  g75
  (
    n101,
    n26
  );


  buf
  g76
  (
    n117,
    n27
  );


  not
  g77
  (
    n59,
    n31
  );


  not
  g78
  (
    n127,
    n17
  );


  buf
  g79
  (
    n52,
    n23
  );


  buf
  g80
  (
    n155,
    n16
  );


  not
  g81
  (
    n160,
    n22
  );


  not
  g82
  (
    n36,
    n26
  );


  not
  g83
  (
    n78,
    n32
  );


  not
  g84
  (
    n70,
    n2
  );


  buf
  g85
  (
    n141,
    n9
  );


  buf
  g86
  (
    n34,
    n1
  );


  not
  g87
  (
    n143,
    n25
  );


  buf
  g88
  (
    n56,
    n30
  );


  buf
  g89
  (
    n68,
    n13
  );


  not
  g90
  (
    n60,
    n16
  );


  buf
  g91
  (
    n120,
    n2
  );


  buf
  g92
  (
    n77,
    n12
  );


  buf
  g93
  (
    n112,
    n19
  );


  not
  g94
  (
    n86,
    n3
  );


  buf
  g95
  (
    n51,
    n4
  );


  not
  g96
  (
    n55,
    n20
  );


  buf
  g97
  (
    n109,
    n1
  );


  not
  g98
  (
    n75,
    n23
  );


  not
  g99
  (
    n42,
    n17
  );


  buf
  g100
  (
    n46,
    n11
  );


  buf
  g101
  (
    n85,
    n4
  );


  not
  g102
  (
    n126,
    n29
  );


  buf
  g103
  (
    n39,
    n22
  );


  not
  g104
  (
    n62,
    n20
  );


  not
  g105
  (
    n76,
    n12
  );


  buf
  g106
  (
    n57,
    n17
  );


  not
  g107
  (
    n92,
    n10
  );


  buf
  g108
  (
    n45,
    n3
  );


  not
  g109
  (
    n134,
    n30
  );


  buf
  g110
  (
    n138,
    n21
  );


  not
  g111
  (
    n114,
    n22
  );


  not
  g112
  (
    n58,
    n19
  );


  not
  g113
  (
    n53,
    n2
  );


  not
  g114
  (
    n100,
    n9
  );


  buf
  g115
  (
    n154,
    n6
  );


  buf
  g116
  (
    n140,
    n7
  );


  not
  g117
  (
    n131,
    n16
  );


  not
  g118
  (
    n107,
    n24
  );


  not
  g119
  (
    n133,
    n13
  );


  buf
  g120
  (
    n79,
    n17
  );


  not
  g121
  (
    n123,
    n19
  );


  buf
  g122
  (
    n40,
    n8
  );


  not
  g123
  (
    n156,
    n11
  );


  buf
  g124
  (
    n35,
    n20
  );


  not
  g125
  (
    n96,
    n6
  );


  not
  g126
  (
    n104,
    n5
  );


  not
  g127
  (
    n118,
    n2
  );


  not
  g128
  (
    n392,
    n33
  );


  buf
  g129
  (
    n213,
    n142
  );


  not
  g130
  (
    n306,
    n75
  );


  not
  g131
  (
    n202,
    n51
  );


  buf
  g132
  (
    n182,
    n67
  );


  buf
  g133
  (
    n429,
    n45
  );


  not
  g134
  (
    n442,
    n61
  );


  buf
  g135
  (
    n178,
    n117
  );


  buf
  g136
  (
    n322,
    n56
  );


  buf
  g137
  (
    n342,
    n144
  );


  not
  g138
  (
    n169,
    n148
  );


  buf
  g139
  (
    n179,
    n136
  );


  not
  g140
  (
    n247,
    n128
  );


  buf
  g141
  (
    n210,
    n74
  );


  not
  g142
  (
    n272,
    n137
  );


  not
  g143
  (
    n197,
    n99
  );


  buf
  g144
  (
    n358,
    n136
  );


  not
  g145
  (
    n257,
    n35
  );


  buf
  g146
  (
    n294,
    n46
  );


  buf
  g147
  (
    n302,
    n50
  );


  not
  g148
  (
    n451,
    n145
  );


  not
  g149
  (
    n377,
    n47
  );


  buf
  g150
  (
    n224,
    n147
  );


  buf
  g151
  (
    n414,
    n122
  );


  not
  g152
  (
    n276,
    n126
  );


  not
  g153
  (
    n323,
    n107
  );


  not
  g154
  (
    n352,
    n84
  );


  buf
  g155
  (
    n223,
    n68
  );


  buf
  g156
  (
    n399,
    n53
  );


  not
  g157
  (
    n436,
    n37
  );


  not
  g158
  (
    n419,
    n91
  );


  buf
  g159
  (
    n263,
    n113
  );


  not
  g160
  (
    n389,
    n56
  );


  buf
  g161
  (
    n232,
    n76
  );


  not
  g162
  (
    n295,
    n91
  );


  not
  g163
  (
    n362,
    n42
  );


  not
  g164
  (
    n338,
    n91
  );


  not
  g165
  (
    n382,
    n108
  );


  buf
  g166
  (
    n349,
    n90
  );


  buf
  g167
  (
    n471,
    n72
  );


  buf
  g168
  (
    n261,
    n146
  );


  buf
  g169
  (
    n446,
    n140
  );


  not
  g170
  (
    n353,
    n113
  );


  not
  g171
  (
    n395,
    n94
  );


  not
  g172
  (
    n415,
    n88
  );


  buf
  g173
  (
    n273,
    n147
  );


  not
  g174
  (
    n423,
    n82
  );


  buf
  g175
  (
    n312,
    n91
  );


  not
  g176
  (
    n246,
    n147
  );


  not
  g177
  (
    n435,
    n81
  );


  not
  g178
  (
    n360,
    n132
  );


  not
  g179
  (
    n409,
    n142
  );


  not
  g180
  (
    n385,
    n65
  );


  not
  g181
  (
    n404,
    n145
  );


  buf
  g182
  (
    n443,
    n129
  );


  buf
  g183
  (
    n198,
    n86
  );


  buf
  g184
  (
    n420,
    n120
  );


  not
  g185
  (
    n229,
    n142
  );


  buf
  g186
  (
    n316,
    n118
  );


  buf
  g187
  (
    n344,
    n96
  );


  buf
  g188
  (
    n403,
    n37
  );


  not
  g189
  (
    n278,
    n34
  );


  buf
  g190
  (
    n464,
    n126
  );


  buf
  g191
  (
    n196,
    n38
  );


  buf
  g192
  (
    n245,
    n48
  );


  buf
  g193
  (
    n175,
    n97
  );


  not
  g194
  (
    n287,
    n49
  );


  not
  g195
  (
    n288,
    n39
  );


  not
  g196
  (
    n274,
    n116
  );


  not
  g197
  (
    n383,
    n72
  );


  buf
  g198
  (
    n172,
    n150
  );


  not
  g199
  (
    n215,
    n122
  );


  not
  g200
  (
    n356,
    n124
  );


  buf
  g201
  (
    n239,
    n88
  );


  not
  g202
  (
    n265,
    n106
  );


  not
  g203
  (
    n454,
    n115
  );


  buf
  g204
  (
    n388,
    n138
  );


  not
  g205
  (
    n386,
    n135
  );


  not
  g206
  (
    n290,
    n84
  );


  buf
  g207
  (
    n235,
    n69
  );


  not
  g208
  (
    n381,
    n95
  );


  not
  g209
  (
    n199,
    n124
  );


  not
  g210
  (
    n244,
    n107
  );


  buf
  g211
  (
    n359,
    n81
  );


  not
  g212
  (
    n298,
    n47
  );


  buf
  g213
  (
    n397,
    n43
  );


  not
  g214
  (
    n343,
    n123
  );


  not
  g215
  (
    n328,
    n128
  );


  buf
  g216
  (
    n194,
    n126
  );


  buf
  g217
  (
    n432,
    n109
  );


  buf
  g218
  (
    n363,
    n34
  );


  not
  g219
  (
    n333,
    n117
  );


  not
  g220
  (
    n228,
    n71
  );


  not
  g221
  (
    n309,
    n92
  );


  buf
  g222
  (
    n268,
    n49
  );


  not
  g223
  (
    n410,
    n88
  );


  buf
  g224
  (
    n264,
    n154
  );


  not
  g225
  (
    n424,
    n34
  );


  not
  g226
  (
    n472,
    n89
  );


  buf
  g227
  (
    n440,
    n66
  );


  buf
  g228
  (
    n171,
    n102
  );


  not
  g229
  (
    n254,
    n127
  );


  not
  g230
  (
    n369,
    n40
  );


  not
  g231
  (
    n260,
    n67
  );


  buf
  g232
  (
    n332,
    n114
  );


  buf
  g233
  (
    KeyWire_0_8,
    n37
  );


  buf
  g234
  (
    n370,
    n148
  );


  buf
  g235
  (
    n315,
    n103
  );


  buf
  g236
  (
    n378,
    n45
  );


  buf
  g237
  (
    n475,
    n66
  );


  not
  g238
  (
    KeyWire_0_7,
    n151
  );


  buf
  g239
  (
    n325,
    n60
  );


  buf
  g240
  (
    n321,
    n79
  );


  buf
  g241
  (
    n307,
    n46
  );


  buf
  g242
  (
    n331,
    n77
  );


  buf
  g243
  (
    n310,
    n96
  );


  not
  g244
  (
    n296,
    n36
  );


  buf
  g245
  (
    n350,
    n120
  );


  buf
  g246
  (
    n188,
    n74
  );


  not
  g247
  (
    n367,
    n92
  );


  not
  g248
  (
    n402,
    n111
  );


  not
  g249
  (
    n262,
    n83
  );


  buf
  g250
  (
    n324,
    n69
  );


  not
  g251
  (
    n366,
    n65
  );


  not
  g252
  (
    n418,
    n79
  );


  buf
  g253
  (
    n167,
    n69
  );


  buf
  g254
  (
    n201,
    n124
  );


  not
  g255
  (
    n177,
    n127
  );


  not
  g256
  (
    n444,
    n55
  );


  buf
  g257
  (
    n200,
    n125
  );


  not
  g258
  (
    n463,
    n122
  );


  buf
  g259
  (
    n212,
    n152
  );


  buf
  g260
  (
    n161,
    n41
  );


  not
  g261
  (
    n162,
    n106
  );


  not
  g262
  (
    n303,
    n47
  );


  not
  g263
  (
    n330,
    n76
  );


  not
  g264
  (
    n434,
    n83
  );


  not
  g265
  (
    n391,
    n38
  );


  buf
  g266
  (
    n291,
    n131
  );


  buf
  g267
  (
    n227,
    n41
  );


  not
  g268
  (
    n318,
    n36
  );


  buf
  g269
  (
    n368,
    n43
  );


  not
  g270
  (
    n271,
    n115
  );


  not
  g271
  (
    n340,
    n78
  );


  buf
  g272
  (
    n433,
    n150
  );


  not
  g273
  (
    n181,
    n84
  );


  not
  g274
  (
    n209,
    n136
  );


  buf
  g275
  (
    n412,
    n40
  );


  not
  g276
  (
    n237,
    n94
  );


  not
  g277
  (
    n173,
    n148
  );


  buf
  g278
  (
    n455,
    n44
  );


  buf
  g279
  (
    n190,
    n104
  );


  buf
  g280
  (
    n374,
    n131
  );


  not
  g281
  (
    n259,
    n53
  );


  buf
  g282
  (
    n365,
    n105
  );


  buf
  g283
  (
    n417,
    n67
  );


  not
  g284
  (
    n279,
    n107
  );


  not
  g285
  (
    n217,
    n85
  );


  not
  g286
  (
    n241,
    n151
  );


  buf
  g287
  (
    KeyWire_0_4,
    n134
  );


  buf
  g288
  (
    n207,
    n95
  );


  not
  g289
  (
    n387,
    n102
  );


  not
  g290
  (
    n300,
    n152
  );


  not
  g291
  (
    n460,
    n103
  );


  not
  g292
  (
    n336,
    n68
  );


  buf
  g293
  (
    n269,
    n63
  );


  not
  g294
  (
    KeyWire_0_15,
    n59
  );


  buf
  g295
  (
    n408,
    n59
  );


  buf
  g296
  (
    n345,
    n141
  );


  buf
  g297
  (
    n170,
    n114
  );


  not
  g298
  (
    n165,
    n143
  );


  buf
  g299
  (
    n219,
    n129
  );


  buf
  g300
  (
    n281,
    n35
  );


  not
  g301
  (
    n384,
    n100
  );


  buf
  g302
  (
    n208,
    n100
  );


  buf
  g303
  (
    n448,
    n98
  );


  not
  g304
  (
    n411,
    n44
  );


  not
  g305
  (
    n441,
    n38
  );


  buf
  g306
  (
    n252,
    n52
  );


  not
  g307
  (
    n299,
    n40
  );


  not
  g308
  (
    n308,
    n121
  );


  not
  g309
  (
    n248,
    n87
  );


  not
  g310
  (
    n311,
    n109
  );


  not
  g311
  (
    n327,
    n89
  );


  buf
  g312
  (
    n275,
    n134
  );


  buf
  g313
  (
    n166,
    n110
  );


  buf
  g314
  (
    n314,
    n76
  );


  buf
  g315
  (
    n192,
    n108
  );


  not
  g316
  (
    n204,
    n75
  );


  not
  g317
  (
    n430,
    n80
  );


  buf
  g318
  (
    n355,
    n65
  );


  not
  g319
  (
    KeyWire_0_12,
    n127
  );


  not
  g320
  (
    n280,
    n119
  );


  not
  g321
  (
    n428,
    n90
  );


  buf
  g322
  (
    n230,
    n98
  );


  not
  g323
  (
    n465,
    n80
  );


  buf
  g324
  (
    n238,
    n134
  );


  buf
  g325
  (
    n211,
    n62
  );


  buf
  g326
  (
    n317,
    n56
  );


  buf
  g327
  (
    n461,
    n133
  );


  not
  g328
  (
    n250,
    n101
  );


  not
  g329
  (
    n220,
    n50
  );


  buf
  g330
  (
    n176,
    n105
  );


  not
  g331
  (
    n185,
    n109
  );


  buf
  g332
  (
    n351,
    n139
  );


  not
  g333
  (
    n187,
    n149
  );


  not
  g334
  (
    n427,
    n102
  );


  buf
  g335
  (
    n186,
    n122
  );


  buf
  g336
  (
    n270,
    n56
  );


  not
  g337
  (
    n469,
    n82
  );


  not
  g338
  (
    n406,
    n124
  );


  not
  g339
  (
    n214,
    n71
  );


  buf
  g340
  (
    n329,
    n76
  );


  buf
  g341
  (
    n297,
    n84
  );


  not
  g342
  (
    n462,
    n140
  );


  not
  g343
  (
    n304,
    n139
  );


  buf
  g344
  (
    n163,
    n78
  );


  not
  g345
  (
    n354,
    n55
  );


  not
  g346
  (
    n305,
    n86
  );


  buf
  g347
  (
    n242,
    n73
  );


  buf
  g348
  (
    n277,
    n68
  );


  not
  g349
  (
    n174,
    n52
  );


  not
  g350
  (
    n326,
    n89
  );


  not
  g351
  (
    n470,
    n152
  );


  not
  g352
  (
    n438,
    n107
  );


  buf
  g353
  (
    n337,
    n146
  );


  not
  g354
  (
    n361,
    n120
  );


  not
  g355
  (
    n218,
    n139
  );


  buf
  g356
  (
    n205,
    n82
  );


  not
  g357
  (
    n400,
    n60
  );


  buf
  g358
  (
    n286,
    n64
  );


  buf
  g359
  (
    n236,
    n80
  );


  buf
  g360
  (
    n258,
    n94
  );


  not
  g361
  (
    n206,
    n78
  );


  not
  g362
  (
    n347,
    n146
  );


  buf
  g363
  (
    n289,
    n114
  );


  not
  g364
  (
    n180,
    n61
  );


  not
  g365
  (
    n203,
    n121
  );


  buf
  g366
  (
    n293,
    n132
  );


  not
  g367
  (
    n393,
    n63
  );


  not
  g368
  (
    n221,
    n136
  );


  buf
  g369
  (
    n466,
    n120
  );


  buf
  g370
  (
    n346,
    n70
  );


  not
  g371
  (
    n447,
    n55
  );


  not
  g372
  (
    n253,
    n106
  );


  buf
  g373
  (
    n425,
    n135
  );


  not
  g374
  (
    n422,
    n60
  );


  buf
  g375
  (
    n401,
    n111
  );


  buf
  g376
  (
    n183,
    n109
  );


  buf
  g377
  (
    n283,
    n39
  );


  buf
  g378
  (
    n474,
    n47
  );


  buf
  g379
  (
    n292,
    n73
  );


  not
  g380
  (
    n375,
    n113
  );


  not
  g381
  (
    n320,
    n51
  );


  not
  g382
  (
    n473,
    n73
  );


  not
  g383
  (
    n467,
    n64
  );


  buf
  g384
  (
    n371,
    n125
  );


  not
  g385
  (
    n284,
    n42
  );


  nor
  g386
  (
    n357,
    n62,
    n137,
    n59
  );


  xor
  g387
  (
    n439,
    n51,
    n39,
    n42,
    n103
  );


  or
  g388
  (
    n431,
    n110,
    n39,
    n137,
    n64
  );


  and
  g389
  (
    n376,
    n118,
    n45,
    n44,
    n104
  );


  xor
  g390
  (
    n233,
    n70,
    n133,
    n75,
    n130
  );


  nand
  g391
  (
    n421,
    n137,
    n74,
    n115,
    n57
  );


  xnor
  g392
  (
    n164,
    n58,
    n99,
    n121,
    n110
  );


  xor
  g393
  (
    n226,
    n87,
    n61,
    n96,
    n101
  );


  xnor
  g394
  (
    n319,
    n135,
    n141,
    n112,
    n134
  );


  nand
  g395
  (
    n450,
    n112,
    n57,
    n104,
    n138
  );


  xor
  g396
  (
    n168,
    n104,
    n121,
    n48,
    n41
  );


  and
  g397
  (
    n243,
    n149,
    n85,
    n111,
    n130
  );


  and
  g398
  (
    n416,
    n132,
    n85,
    n118,
    n130
  );


  or
  g399
  (
    n453,
    n38,
    n49,
    n98,
    n130
  );


  xor
  g400
  (
    n407,
    n149,
    n138,
    n147,
    n69
  );


  xnor
  g401
  (
    n234,
    n149,
    n75,
    n60,
    n140
  );


  nand
  g402
  (
    n458,
    n116,
    n145,
    n153,
    n72
  );


  and
  g403
  (
    n437,
    n92,
    n95,
    n67,
    n62
  );


  xnor
  g404
  (
    n282,
    n81,
    n52,
    n79,
    n53
  );


  and
  g405
  (
    n189,
    n112,
    n119,
    n64,
    n68
  );


  or
  g406
  (
    n255,
    n62,
    n113,
    n105,
    n36
  );


  nand
  g407
  (
    n364,
    n123,
    n117,
    n111,
    n131
  );


  xnor
  g408
  (
    n348,
    n96,
    n94,
    n140,
    n63
  );


  nor
  g409
  (
    n452,
    n135,
    n33,
    n119,
    n143
  );


  or
  g410
  (
    n313,
    n141,
    n70,
    n34,
    n108
  );


  xor
  g411
  (
    n426,
    n78,
    n44,
    n98,
    n77
  );


  xor
  g412
  (
    n339,
    n101,
    n43,
    n99,
    n61
  );


  nor
  g413
  (
    n240,
    n37,
    n86,
    n41,
    n152
  );


  nand
  g414
  (
    n222,
    n114,
    n93,
    n106,
    n82
  );


  nor
  g415
  (
    n398,
    n89,
    n46,
    n97,
    n73
  );


  nor
  g416
  (
    n468,
    n151,
    n87,
    n116,
    n153
  );


  nor
  g417
  (
    n301,
    n123,
    n139,
    n50,
    n142
  );


  or
  g418
  (
    n193,
    n129,
    n51,
    n133,
    n59
  );


  xor
  g419
  (
    n372,
    n48,
    n48,
    n54,
    n63
  );


  nand
  g420
  (
    n459,
    n126,
    n112,
    n93,
    n153
  );


  or
  g421
  (
    n445,
    n43,
    n97,
    n74,
    n110
  );


  or
  g422
  (
    n390,
    n144,
    n58,
    n80,
    n33
  );


  xor
  g423
  (
    n231,
    n58,
    n151,
    n93,
    n70
  );


  and
  g424
  (
    n256,
    n35,
    n128,
    n85,
    n86
  );


  and
  g425
  (
    n449,
    n58,
    n148,
    n146,
    n55
  );


  xnor
  g426
  (
    n373,
    n77,
    n100,
    n145,
    n57
  );


  and
  g427
  (
    n285,
    n52,
    n35,
    n88,
    n99
  );


  nor
  g428
  (
    n379,
    n54,
    n66,
    n138,
    n117
  );


  xor
  g429
  (
    n380,
    n131,
    n118,
    n81,
    n144
  );


  and
  g430
  (
    n266,
    n132,
    n79,
    n54,
    n108
  );


  xor
  g431
  (
    KeyWire_0_3,
    n93,
    n153,
    n115,
    n150
  );


  xor
  g432
  (
    n216,
    n123,
    n66,
    n87,
    n105
  );


  and
  g433
  (
    n341,
    n72,
    n71,
    n102,
    n83
  );


  xor
  g434
  (
    n225,
    n133,
    n144,
    n129,
    n97
  );


  nor
  g435
  (
    n335,
    n45,
    n150,
    n116,
    n71
  );


  xor
  g436
  (
    n249,
    n57,
    n119,
    n125,
    n143
  );


  xnor
  g437
  (
    n191,
    n83,
    n128,
    n65,
    n92
  );


  or
  g438
  (
    n413,
    n127,
    n77,
    n33,
    n90
  );


  and
  g439
  (
    n457,
    n143,
    n49,
    n125,
    n50
  );


  nand
  g440
  (
    n251,
    n53,
    n103,
    n100,
    n101
  );


  nand
  g441
  (
    n394,
    n90,
    n36,
    n40,
    n141
  );


  nand
  g442
  (
    n396,
    n95,
    n42,
    n46,
    n54
  );


  nand
  g443
  (
    n491,
    n178,
    n181,
    n220,
    n222
  );


  or
  g444
  (
    n490,
    n162,
    n170,
    n217,
    n200
  );


  nand
  g445
  (
    n484,
    n212,
    n186,
    n184,
    n227
  );


  nor
  g446
  (
    n492,
    n183,
    n205,
    n175,
    n190
  );


  xor
  g447
  (
    n478,
    n214,
    n196,
    n163,
    n216
  );


  or
  g448
  (
    n476,
    n179,
    n191,
    n206,
    n164
  );


  xnor
  g449
  (
    n488,
    n177,
    n172,
    n182,
    n161
  );


  nor
  g450
  (
    n493,
    n180,
    n202,
    n174,
    n219
  );


  xor
  g451
  (
    n479,
    n204,
    n228,
    n171,
    n207
  );


  xor
  g452
  (
    n483,
    n213,
    n209,
    n169,
    n166
  );


  nor
  g453
  (
    n477,
    n185,
    n195,
    n199,
    n229
  );


  xnor
  g454
  (
    n481,
    n197,
    n173,
    n225,
    n232
  );


  nand
  g455
  (
    n489,
    n176,
    n230,
    n189,
    n211
  );


  xnor
  g456
  (
    n485,
    n165,
    n223,
    n188,
    n194
  );


  xor
  g457
  (
    n486,
    n208,
    n167,
    n201,
    n224
  );


  xor
  g458
  (
    n482,
    n226,
    n192,
    n210,
    n218
  );


  xor
  g459
  (
    n487,
    n168,
    n193,
    n198,
    n203
  );


  xnor
  g460
  (
    KeyWire_0_13,
    n231,
    n187,
    n215,
    n221
  );


  not
  g461
  (
    KeyWire_0_0,
    n155
  );


  buf
  g462
  (
    n501,
    n156
  );


  buf
  g463
  (
    n502,
    n154
  );


  buf
  g464
  (
    n495,
    n481
  );


  not
  g465
  (
    n505,
    n485
  );


  buf
  g466
  (
    n497,
    n479
  );


  or
  g467
  (
    n496,
    n487,
    n157
  );


  or
  g468
  (
    n498,
    n484,
    n478,
    n155,
    n156
  );


  xnor
  g469
  (
    n500,
    n480,
    n158,
    n482,
    n157
  );


  or
  g470
  (
    n499,
    n486,
    n155,
    n156
  );


  or
  g471
  (
    n504,
    n157,
    n155,
    n154
  );


  nand
  g472
  (
    n503,
    n477,
    n476,
    n483,
    n157
  );


  not
  g473
  (
    n507,
    n495
  );


  buf
  g474
  (
    n515,
    n495
  );


  buf
  g475
  (
    n509,
    n494
  );


  not
  g476
  (
    n508,
    n496
  );


  buf
  g477
  (
    n511,
    n494
  );


  buf
  g478
  (
    n513,
    n496
  );


  buf
  g479
  (
    n512,
    n496
  );


  buf
  g480
  (
    n506,
    n495
  );


  buf
  g481
  (
    n516,
    n495
  );


  buf
  g482
  (
    n514,
    n494
  );


  not
  g483
  (
    n510,
    n494
  );


  buf
  g484
  (
    n531,
    n508
  );


  not
  g485
  (
    n532,
    n489
  );


  buf
  g486
  (
    n521,
    n507
  );


  buf
  g487
  (
    n527,
    n508
  );


  not
  g488
  (
    n523,
    n506
  );


  not
  g489
  (
    n526,
    n506
  );


  buf
  g490
  (
    n517,
    n509
  );


  not
  g491
  (
    n518,
    n509
  );


  buf
  g492
  (
    n530,
    n507
  );


  not
  g493
  (
    n522,
    n509
  );


  buf
  g494
  (
    KeyWire_0_9,
    n509
  );


  buf
  g495
  (
    n525,
    n507
  );


  not
  g496
  (
    n519,
    n507
  );


  not
  g497
  (
    n529,
    n506
  );


  not
  g498
  (
    n524,
    n508
  );


  or
  g499
  (
    KeyWire_0_11,
    n506,
    n488,
    n508,
    n490
  );


  not
  g500
  (
    n536,
    n497
  );


  not
  g501
  (
    n537,
    n519
  );


  not
  g502
  (
    n539,
    n518
  );


  buf
  g503
  (
    n541,
    n500
  );


  nor
  g504
  (
    n533,
    n499,
    n497
  );


  nand
  g505
  (
    n538,
    n491,
    n518,
    n500
  );


  or
  g506
  (
    n534,
    n501,
    n498,
    n518
  );


  or
  g507
  (
    n540,
    n499,
    n497,
    n498,
    n518
  );


  xnor
  g508
  (
    n535,
    n499,
    n497,
    n517
  );


  nor
  g509
  (
    n543,
    n498,
    n519,
    n517
  );


  and
  g510
  (
    n542,
    n500,
    n519,
    n499,
    n496
  );


  not
  g511
  (
    n546,
    n503
  );


  buf
  g512
  (
    n566,
    n543
  );


  not
  g513
  (
    n564,
    n542
  );


  buf
  g514
  (
    n548,
    n540
  );


  not
  g515
  (
    n568,
    n543
  );


  buf
  g516
  (
    n559,
    n504
  );


  buf
  g517
  (
    n565,
    n537
  );


  not
  g518
  (
    n553,
    n510
  );


  not
  g519
  (
    n561,
    n503
  );


  buf
  g520
  (
    n558,
    n503
  );


  buf
  g521
  (
    n551,
    n505
  );


  buf
  g522
  (
    n545,
    n535
  );


  buf
  g523
  (
    n544,
    n541
  );


  buf
  g524
  (
    n569,
    n510
  );


  buf
  g525
  (
    n560,
    n539
  );


  not
  g526
  (
    n555,
    n511
  );


  nand
  g527
  (
    n557,
    n542,
    n501,
    n543
  );


  xor
  g528
  (
    n552,
    n504,
    n539,
    n501,
    n505
  );


  xnor
  g529
  (
    n567,
    n511,
    n234,
    n502,
    n235
  );


  xnor
  g530
  (
    n547,
    n533,
    n502,
    n501,
    n504
  );


  or
  g531
  (
    n562,
    n541,
    n504,
    n502,
    n511
  );


  nor
  g532
  (
    n549,
    n540,
    n503,
    n542,
    n233
  );


  xnor
  g533
  (
    n563,
    n502,
    n541,
    n539,
    n534
  );


  and
  g534
  (
    n550,
    n505,
    n536,
    n538,
    n511
  );


  nand
  g535
  (
    n554,
    n540,
    n510
  );


  and
  g536
  (
    n556,
    n541,
    n542,
    n539,
    n505
  );


  not
  g537
  (
    n575,
    n547
  );


  buf
  g538
  (
    n585,
    n545
  );


  buf
  g539
  (
    n589,
    n520
  );


  buf
  g540
  (
    n572,
    n548
  );


  not
  g541
  (
    n588,
    n520
  );


  buf
  g542
  (
    n571,
    n521
  );


  buf
  g543
  (
    n578,
    n547
  );


  buf
  g544
  (
    n590,
    n546
  );


  not
  g545
  (
    n576,
    n545
  );


  not
  g546
  (
    n574,
    n520
  );


  buf
  g547
  (
    n570,
    n549
  );


  buf
  g548
  (
    n573,
    n548
  );


  buf
  g549
  (
    n587,
    n548
  );


  not
  g550
  (
    n580,
    n544
  );


  buf
  g551
  (
    n584,
    n546
  );


  buf
  g552
  (
    n581,
    n544
  );


  not
  g553
  (
    n577,
    n548
  );


  not
  g554
  (
    n579,
    n521
  );


  or
  g555
  (
    n582,
    n544,
    n519
  );


  or
  g556
  (
    n586,
    n522,
    n544,
    n545
  );


  xnor
  g557
  (
    n591,
    n547,
    n521,
    n520
  );


  or
  g558
  (
    n583,
    n547,
    n546,
    n549
  );


  buf
  g559
  (
    n613,
    n572
  );


  buf
  g560
  (
    n596,
    n572
  );


  not
  g561
  (
    n611,
    n570
  );


  buf
  g562
  (
    n603,
    n573
  );


  buf
  g563
  (
    n593,
    n574
  );


  not
  g564
  (
    n595,
    n528
  );


  not
  g565
  (
    n601,
    n527
  );


  not
  g566
  (
    n614,
    n528
  );


  not
  g567
  (
    n592,
    n528
  );


  not
  g568
  (
    n597,
    n570
  );


  not
  g569
  (
    n604,
    n526
  );


  not
  g570
  (
    n608,
    n574
  );


  not
  g571
  (
    n609,
    n523
  );


  and
  g572
  (
    n612,
    n573,
    n525
  );


  and
  g573
  (
    n602,
    n529,
    n570,
    n522,
    n524
  );


  nand
  g574
  (
    n598,
    n523,
    n571,
    n574,
    n573
  );


  nand
  g575
  (
    n607,
    n528,
    n573,
    n574,
    n572
  );


  nor
  g576
  (
    n606,
    n525,
    n570,
    n575,
    n571
  );


  nand
  g577
  (
    n605,
    n571,
    n572,
    n575,
    n524
  );


  nor
  g578
  (
    n615,
    n524,
    n529,
    n571,
    n527
  );


  nand
  g579
  (
    n610,
    n523,
    n529,
    n522,
    n526
  );


  and
  g580
  (
    n594,
    n530,
    n524,
    n526
  );


  or
  g581
  (
    n599,
    n525,
    n527,
    n529,
    n575
  );


  nor
  g582
  (
    n600,
    n523,
    n522,
    n527,
    n575
  );


  or
  g583
  (
    n629,
    n594,
    n236,
    n558,
    n593
  );


  nor
  g584
  (
    n628,
    n597,
    n595,
    n554,
    n549
  );


  xor
  g585
  (
    n637,
    n558,
    n564,
    n563,
    n592
  );


  xor
  g586
  (
    n643,
    n594,
    n515,
    n557
  );


  and
  g587
  (
    n618,
    n514,
    n595,
    n554
  );


  xor
  g588
  (
    n630,
    n599,
    n564,
    n596,
    n600
  );


  xnor
  g589
  (
    n639,
    n562,
    n565,
    n239,
    n563
  );


  xor
  g590
  (
    n640,
    n515,
    n562,
    n595,
    n592
  );


  nor
  g591
  (
    n634,
    n563,
    n513,
    n554
  );


  xnor
  g592
  (
    n616,
    n551,
    n598,
    n600,
    n564
  );


  xor
  g593
  (
    n649,
    n561,
    n557,
    n562,
    n237
  );


  nor
  g594
  (
    n624,
    n514,
    n569,
    n592,
    n566
  );


  nor
  g595
  (
    n617,
    n559,
    n564,
    n599
  );


  nor
  g596
  (
    n632,
    n550,
    n552,
    n599,
    n566
  );


  xnor
  g597
  (
    n642,
    n556,
    n555,
    n563,
    n242
  );


  or
  g598
  (
    n625,
    n566,
    n562,
    n550,
    n560
  );


  nor
  g599
  (
    n648,
    n559,
    n550,
    n567,
    n568
  );


  and
  g600
  (
    n644,
    n596,
    n561,
    n559,
    n594
  );


  xnor
  g601
  (
    n635,
    n555,
    n569,
    n596,
    n592
  );


  nor
  g602
  (
    n631,
    n553,
    n569,
    n551,
    n243
  );


  xnor
  g603
  (
    n623,
    n552,
    n559,
    n240,
    n514
  );


  xnor
  g604
  (
    n645,
    n558,
    n568,
    n551,
    n512
  );


  nor
  g605
  (
    n650,
    n569,
    n513,
    n593,
    n556
  );


  xnor
  g606
  (
    n641,
    n597,
    n568,
    n560
  );


  and
  g607
  (
    n646,
    n555,
    n565,
    n552,
    n566
  );


  and
  g608
  (
    n619,
    n512,
    n551,
    n600,
    n560
  );


  or
  g609
  (
    n626,
    n561,
    n241,
    n554,
    n512
  );


  and
  g610
  (
    KeyWire_0_5,
    n244,
    n553,
    n598,
    n512
  );


  xnor
  g611
  (
    n621,
    n594,
    n552,
    n567,
    n513
  );


  nor
  g612
  (
    n647,
    n514,
    n598,
    n567,
    n565
  );


  xor
  g613
  (
    n622,
    n567,
    n597,
    n556,
    n555
  );


  nor
  g614
  (
    n620,
    n553,
    n593,
    n565,
    n556
  );


  nor
  g615
  (
    n638,
    n561,
    n557,
    n550,
    n598
  );


  nand
  g616
  (
    n627,
    n596,
    n553,
    n558,
    n560
  );


  xor
  g617
  (
    n636,
    n549,
    n593,
    n597,
    n238
  );


  xnor
  g618
  (
    n652,
    n581,
    n581,
    n578,
    n623
  );


  xnor
  g619
  (
    n656,
    n618,
    n582,
    n577,
    n621
  );


  and
  g620
  (
    n655,
    n622,
    n579,
    n576
  );


  xnor
  g621
  (
    n657,
    n580,
    n577,
    n581
  );


  xor
  g622
  (
    n659,
    n582,
    n578,
    n580
  );


  nor
  g623
  (
    n658,
    n624,
    n582,
    n580,
    n577
  );


  xor
  g624
  (
    n651,
    n581,
    n576,
    n578
  );


  xor
  g625
  (
    n654,
    n619,
    n576,
    n620,
    n616
  );


  xor
  g626
  (
    n653,
    n617,
    n580,
    n579
  );


  not
  g627
  (
    n669,
    n654
  );


  buf
  g628
  (
    n667,
    n653
  );


  buf
  g629
  (
    n665,
    n652
  );


  not
  g630
  (
    n668,
    n653
  );


  not
  g631
  (
    n679,
    n651
  );


  not
  g632
  (
    n660,
    n654
  );


  not
  g633
  (
    n672,
    n652
  );


  buf
  g634
  (
    n671,
    n600
  );


  buf
  g635
  (
    n675,
    n651
  );


  buf
  g636
  (
    n673,
    n652
  );


  buf
  g637
  (
    n677,
    n653
  );


  not
  g638
  (
    n674,
    n601
  );


  buf
  g639
  (
    n666,
    n601
  );


  not
  g640
  (
    n661,
    n601
  );


  buf
  g641
  (
    n662,
    n651
  );


  buf
  g642
  (
    n663,
    n653
  );


  not
  g643
  (
    n664,
    n602
  );


  buf
  g644
  (
    n676,
    n654
  );


  nor
  g645
  (
    n678,
    n651,
    n655
  );


  xor
  g646
  (
    n670,
    n652,
    n601,
    n655,
    n654
  );


  nor
  g647
  (
    n686,
    n625,
    n603,
    n660
  );


  xnor
  g648
  (
    n685,
    n605,
    n604,
    n603,
    n661
  );


  xnor
  g649
  (
    n682,
    n660,
    n604,
    n602,
    n606
  );


  and
  g650
  (
    n680,
    n602,
    n605,
    n604,
    n661
  );


  nand
  g651
  (
    n684,
    n604,
    n606,
    n603,
    n605
  );


  xor
  g652
  (
    n681,
    n627,
    n605,
    n603,
    n660
  );


  xor
  g653
  (
    n683,
    n661,
    n626,
    n606,
    n602
  );


  nand
  g654
  (
    n689,
    n631,
    n632,
    n684,
    n630
  );


  and
  g655
  (
    n688,
    n629,
    n635,
    n628,
    n636
  );


  xor
  g656
  (
    n687,
    n633,
    n634,
    n685,
    n686
  );


  xnor
  g657
  (
    n701,
    n669,
    n689,
    n665,
    n662
  );


  or
  g658
  (
    n691,
    n663,
    n669,
    n687
  );


  or
  g659
  (
    n697,
    n670,
    n668,
    n666,
    n664
  );


  or
  g660
  (
    n693,
    n668,
    n688,
    n665,
    n662
  );


  xor
  g661
  (
    n698,
    n662,
    n689,
    n670,
    n666
  );


  nor
  g662
  (
    n692,
    n667,
    n666,
    n687
  );


  nor
  g663
  (
    n694,
    n670,
    n664,
    n667,
    n665
  );


  and
  g664
  (
    n699,
    n662,
    n666,
    n689,
    n663
  );


  xor
  g665
  (
    n690,
    n661,
    n688,
    n664,
    n669
  );


  and
  g666
  (
    n696,
    n669,
    n688,
    n664,
    n665
  );


  or
  g667
  (
    n700,
    n663,
    n689,
    n668
  );


  nor
  g668
  (
    n695,
    n663,
    n688,
    n667
  );


  nand
  g669
  (
    n705,
    n671,
    n672,
    n673
  );


  nand
  g670
  (
    n703,
    n701,
    n672,
    n670
  );


  xnor
  g671
  (
    n704,
    n671,
    n673,
    n699
  );


  nand
  g672
  (
    n702,
    n671,
    n671,
    n698,
    n700
  );


  nor
  g673
  (
    n707,
    n704,
    n656,
    n609,
    n608
  );


  nand
  g674
  (
    n714,
    n609,
    n585,
    n640,
    n644
  );


  or
  g675
  (
    n719,
    n608,
    n608,
    n515,
    n584
  );


  xor
  g676
  (
    n718,
    n607,
    n702,
    n583,
    n639
  );


  and
  g677
  (
    n715,
    n705,
    n638,
    n703,
    n704
  );


  nor
  g678
  (
    n712,
    n656,
    n606,
    n637,
    n607
  );


  nand
  g679
  (
    n711,
    n610,
    n583,
    n656,
    n643
  );


  nor
  g680
  (
    n716,
    n656,
    n642,
    n612,
    n702
  );


  xnor
  g681
  (
    n717,
    n583,
    n705,
    n607,
    n611
  );


  nor
  g682
  (
    n706,
    n609,
    n582,
    n611,
    n607
  );


  xnor
  g683
  (
    n721,
    n611,
    n608,
    n703,
    n609
  );


  xnor
  g684
  (
    n710,
    n516,
    n515,
    n703,
    n610
  );


  nor
  g685
  (
    n709,
    n704,
    n702,
    n584
  );


  xnor
  g686
  (
    n720,
    n611,
    n610,
    n705,
    n702
  );


  xnor
  g687
  (
    n708,
    n704,
    n641,
    n703,
    n705
  );


  or
  g688
  (
    n713,
    n584,
    n610,
    n612,
    n583
  );


  not
  g689
  (
    n742,
    n710
  );


  buf
  g690
  (
    n734,
    n706
  );


  not
  g691
  (
    n745,
    n706
  );


  not
  g692
  (
    n726,
    n708
  );


  not
  g693
  (
    n747,
    n708
  );


  not
  g694
  (
    n744,
    n711
  );


  buf
  g695
  (
    n746,
    n707
  );


  not
  g696
  (
    n727,
    n709
  );


  not
  g697
  (
    n739,
    n707
  );


  buf
  g698
  (
    n724,
    n710
  );


  not
  g699
  (
    n735,
    n712
  );


  not
  g700
  (
    n725,
    n706
  );


  not
  g701
  (
    n738,
    n706
  );


  not
  g702
  (
    n731,
    n709
  );


  not
  g703
  (
    n736,
    n707
  );


  not
  g704
  (
    n737,
    n711
  );


  not
  g705
  (
    n740,
    n710
  );


  buf
  g706
  (
    n730,
    n711
  );


  not
  g707
  (
    n723,
    n712
  );


  not
  g708
  (
    n729,
    n708
  );


  buf
  g709
  (
    n741,
    n708
  );


  buf
  g710
  (
    n733,
    n710
  );


  buf
  g711
  (
    n728,
    n707
  );


  not
  g712
  (
    n743,
    n711
  );


  buf
  g713
  (
    n722,
    n709
  );


  not
  g714
  (
    n732,
    n709
  );


  xor
  g715
  (
    n780,
    n726,
    n741,
    n673
  );


  xnor
  g716
  (
    n766,
    n727,
    n461,
    n159,
    n349
  );


  nor
  g717
  (
    n797,
    n736,
    n727,
    n399,
    n739
  );


  xnor
  g718
  (
    n807,
    n730,
    n614,
    n740,
    n376
  );


  xnor
  g719
  (
    n816,
    n587,
    n467,
    n746,
    n423
  );


  xnor
  g720
  (
    n764,
    n739,
    n585,
    n471,
    n492
  );


  or
  g721
  (
    n753,
    n379,
    n472,
    n160,
    n587
  );


  or
  g722
  (
    n817,
    n733,
    n417,
    n732,
    n470
  );


  xnor
  g723
  (
    KeyWire_0_2,
    n462,
    n329,
    n269,
    n734
  );


  or
  g724
  (
    n782,
    n158,
    n442,
    n273,
    n675
  );


  and
  g725
  (
    n837,
    n254,
    n263,
    n590,
    n431
  );


  nand
  g726
  (
    n819,
    n308,
    n374,
    n403,
    n460
  );


  xor
  g727
  (
    n841,
    n428,
    n742,
    n588,
    n586
  );


  xnor
  g728
  (
    n788,
    n388,
    n474,
    n355,
    n331
  );


  and
  g729
  (
    n781,
    n313,
    n725,
    n372,
    n456
  );


  xnor
  g730
  (
    n755,
    n474,
    n464,
    n415,
    n412
  );


  and
  g731
  (
    n750,
    n418,
    n457,
    n675,
    n470
  );


  or
  g732
  (
    n846,
    n741,
    n731,
    n251,
    n726
  );


  xnor
  g733
  (
    n825,
    n395,
    n435,
    n304,
    n358
  );


  and
  g734
  (
    n751,
    n317,
    n336,
    n407,
    n436
  );


  xnor
  g735
  (
    n834,
    n587,
    n275,
    n531,
    n590
  );


  nor
  g736
  (
    n770,
    n250,
    n339,
    n409,
    n327
  );


  nor
  g737
  (
    n773,
    n742,
    n290,
    n466,
    n738
  );


  nand
  g738
  (
    n802,
    n745,
    n475,
    n253
  );


  xnor
  g739
  (
    n769,
    n341,
    n159,
    n274,
    n326
  );


  nor
  g740
  (
    n848,
    n258,
    n448,
    n724,
    n314
  );


  or
  g741
  (
    n811,
    n402,
    n398,
    n743,
    n255
  );


  and
  g742
  (
    n795,
    n366,
    n383,
    n247,
    n282
  );


  nand
  g743
  (
    n784,
    n674,
    n345,
    n588,
    n731
  );


  nor
  g744
  (
    n789,
    n324,
    n724,
    n293,
    n734
  );


  or
  g745
  (
    n844,
    n265,
    n350,
    n472,
    n449
  );


  xor
  g746
  (
    n815,
    n472,
    n722,
    n411,
    n249
  );


  xor
  g747
  (
    n809,
    n260,
    n318,
    n424,
    n724
  );


  xnor
  g748
  (
    n783,
    n733,
    n419,
    n737,
    n248
  );


  nor
  g749
  (
    n775,
    n335,
    n433,
    n322,
    n589
  );


  nor
  g750
  (
    n771,
    n320,
    n421,
    n730,
    n347
  );


  and
  g751
  (
    n785,
    n729,
    n158,
    n441,
    n740
  );


  xor
  g752
  (
    n831,
    n729,
    n590,
    n589,
    n312
  );


  xor
  g753
  (
    n828,
    n444,
    n286,
    n256,
    n453
  );


  nor
  g754
  (
    n799,
    n408,
    n585,
    n613,
    n473
  );


  and
  g755
  (
    n761,
    n612,
    n728,
    n735,
    n473
  );


  and
  g756
  (
    n787,
    n300,
    n723,
    n385,
    n724
  );


  nand
  g757
  (
    n804,
    n741,
    n261,
    n160,
    n739
  );


  and
  g758
  (
    n835,
    n471,
    n343,
    n532,
    n591
  );


  xor
  g759
  (
    n774,
    n746,
    n381,
    n736,
    n323
  );


  xor
  g760
  (
    n845,
    n726,
    n295,
    n737,
    n272
  );


  xor
  g761
  (
    n779,
    n392,
    n373,
    n731,
    n727
  );


  xor
  g762
  (
    n801,
    n420,
    n612,
    n732,
    n585
  );


  xnor
  g763
  (
    n850,
    n746,
    n405,
    n438,
    n397
  );


  or
  g764
  (
    n810,
    n369,
    n287,
    n736,
    n303
  );


  nor
  g765
  (
    n759,
    n382,
    n736,
    n340,
    n354
  );


  or
  g766
  (
    n752,
    n674,
    n396,
    n586,
    n365
  );


  nor
  g767
  (
    n760,
    n443,
    n613,
    n380,
    n262
  );


  xnor
  g768
  (
    n793,
    n288,
    n743,
    n451,
    n298
  );


  xnor
  g769
  (
    n765,
    n532,
    n257,
    n353,
    n375
  );


  xor
  g770
  (
    n851,
    n384,
    n416,
    n732,
    n531
  );


  nor
  g771
  (
    n824,
    n296,
    n377,
    n734,
    n268
  );


  nor
  g772
  (
    n756,
    n747,
    n352,
    n738,
    n252
  );


  xor
  g773
  (
    n826,
    n281,
    n731,
    n342,
    n474
  );


  and
  g774
  (
    n822,
    n276,
    n446,
    n725,
    n469
  );


  nor
  g775
  (
    n832,
    n746,
    n356,
    n306,
    n271
  );


  or
  g776
  (
    n827,
    n390,
    n738,
    n472,
    n413
  );


  nor
  g777
  (
    n758,
    n739,
    n733,
    n246,
    n292
  );


  nand
  g778
  (
    n805,
    n159,
    n589,
    n289,
    n735
  );


  nand
  g779
  (
    n767,
    n532,
    n730,
    n747,
    n325
  );


  and
  g780
  (
    n838,
    n470,
    n674,
    n530,
    n744
  );


  xnor
  g781
  (
    n768,
    n725,
    n294,
    n676,
    n359
  );


  nor
  g782
  (
    n763,
    n722,
    n455,
    n264,
    n747
  );


  xnor
  g783
  (
    n791,
    n410,
    n588,
    n330,
    n307
  );


  or
  g784
  (
    n833,
    n590,
    n742,
    n722,
    n591
  );


  and
  g785
  (
    n820,
    n302,
    n465,
    n471,
    n735
  );


  xnor
  g786
  (
    n748,
    n473,
    n531,
    n351,
    n160
  );


  xor
  g787
  (
    n849,
    n645,
    n309,
    n328,
    n371
  );


  or
  g788
  (
    n840,
    n743,
    n440,
    n474,
    n277
  );


  or
  g789
  (
    n754,
    n463,
    n744,
    n266,
    n613
  );


  xor
  g790
  (
    n772,
    n728,
    n725,
    n473,
    n425
  );


  nor
  g791
  (
    n806,
    n723,
    n338,
    n445,
    n422
  );


  nor
  g792
  (
    n762,
    n297,
    n737,
    n728,
    n259
  );


  xnor
  g793
  (
    n808,
    n439,
    n387,
    n319,
    n613
  );


  and
  g794
  (
    n839,
    n738,
    n735,
    n159,
    n301
  );


  xor
  g795
  (
    n792,
    n344,
    n400,
    n391,
    n311
  );


  or
  g796
  (
    n794,
    n740,
    n727,
    n316,
    n279
  );


  nor
  g797
  (
    n778,
    n468,
    n426,
    n434,
    n406
  );


  or
  g798
  (
    n796,
    n429,
    n722,
    n675,
    n432
  );


  nor
  g799
  (
    n818,
    n733,
    n437,
    n321,
    n742
  );


  and
  g800
  (
    n803,
    n732,
    n357,
    n530,
    n283
  );


  and
  g801
  (
    n800,
    n745,
    n346,
    n530,
    n452
  );


  nand
  g802
  (
    n798,
    n404,
    n299,
    n378,
    n160
  );


  and
  g803
  (
    n776,
    n734,
    n587,
    n245,
    n723
  );


  or
  g804
  (
    n823,
    n348,
    n740,
    n459,
    n393
  );


  or
  g805
  (
    n786,
    n744,
    n267,
    n728,
    n729
  );


  xnor
  g806
  (
    n821,
    n367,
    n532,
    n729,
    n414
  );


  xnor
  g807
  (
    n749,
    n386,
    n447,
    n270,
    n744
  );


  and
  g808
  (
    n842,
    n285,
    n360,
    n743,
    n745
  );


  and
  g809
  (
    KeyWire_0_14,
    n747,
    n370,
    n586,
    n458
  );


  and
  g810
  (
    n812,
    n401,
    n280,
    n361,
    n589
  );


  and
  g811
  (
    n814,
    n531,
    n368,
    n586,
    n475
  );


  xnor
  g812
  (
    n843,
    n394,
    n745,
    n315,
    n450
  );


  nor
  g813
  (
    n777,
    n334,
    n332,
    n364,
    n284
  );


  nor
  g814
  (
    n813,
    n427,
    n737,
    n291,
    n675
  );


  xor
  g815
  (
    n847,
    n730,
    n278,
    n362,
    n310
  );


  xor
  g816
  (
    n830,
    n389,
    n363,
    n726,
    n454
  );


  nand
  g817
  (
    n836,
    n333,
    n158,
    n337,
    n430
  );


  and
  g818
  (
    n757,
    n674,
    n588,
    n305,
    n723
  );


  and
  g819
  (
    n854,
    n713,
    n754
  );


  xor
  g820
  (
    n852,
    n714,
    n716,
    n713,
    n750
  );


  xnor
  g821
  (
    n855,
    n753,
    n749,
    n715,
    n712
  );


  and
  g822
  (
    n858,
    n717,
    n716,
    n714,
    n713
  );


  xor
  g823
  (
    n857,
    n716,
    n715,
    n717
  );


  xnor
  g824
  (
    n853,
    n715,
    n748,
    n714,
    n716
  );


  xor
  g825
  (
    n859,
    n755,
    n752,
    n717
  );


  nor
  g826
  (
    n856,
    n714,
    n751,
    n713,
    n712
  );


  xor
  g827
  (
    n863,
    n718,
    n719,
    n591,
    n721
  );


  xor
  g828
  (
    n864,
    n591,
    n721,
    n855
  );


  nor
  g829
  (
    n860,
    n855,
    n719
  );


  nor
  g830
  (
    n861,
    n718,
    n720,
    n853,
    n855
  );


  xnor
  g831
  (
    n865,
    n854,
    n720,
    n721
  );


  xnor
  g832
  (
    n862,
    n852,
    n718,
    n720
  );


  or
  g833
  (
    n866,
    n757,
    n759,
    n766,
    n762
  );


  xnor
  g834
  (
    n867,
    n863,
    n862,
    n768,
    n770
  );


  xnor
  g835
  (
    n870,
    n758,
    n769,
    n865,
    n861
  );


  or
  g836
  (
    n869,
    n767,
    n760,
    n764,
    n763
  );


  nor
  g837
  (
    n868,
    n765,
    n756,
    n761,
    n864
  );


  and
  g838
  (
    n876,
    n789,
    n867,
    n779,
    n787
  );


  and
  g839
  (
    n890,
    n797,
    n783,
    n784,
    n788
  );


  and
  g840
  (
    n882,
    n870,
    n830,
    n866,
    n828
  );


  nor
  g841
  (
    n883,
    n870,
    n804,
    n829,
    n816
  );


  nand
  g842
  (
    n874,
    n802,
    n867,
    n866
  );


  xor
  g843
  (
    n871,
    n818,
    n793,
    n819,
    n782
  );


  or
  g844
  (
    n887,
    n869,
    n866,
    n868,
    n780
  );


  xor
  g845
  (
    n879,
    n800,
    n795,
    n796,
    n869
  );


  nand
  g846
  (
    n886,
    n791,
    n812,
    n823,
    n870
  );


  and
  g847
  (
    n885,
    n867,
    n868,
    n821
  );


  xnor
  g848
  (
    n878,
    n799,
    n810,
    n808,
    n794
  );


  or
  g849
  (
    n881,
    n775,
    n869,
    n820,
    n814
  );


  xor
  g850
  (
    n880,
    n869,
    n807,
    n822,
    n785
  );


  xnor
  g851
  (
    n875,
    n773,
    n798,
    n781,
    n774
  );


  nor
  g852
  (
    n884,
    n824,
    n790,
    n866,
    n803
  );


  nand
  g853
  (
    n877,
    n815,
    n827,
    n771,
    n811
  );


  xnor
  g854
  (
    n872,
    n813,
    n778,
    n801,
    n868
  );


  nand
  g855
  (
    n889,
    n817,
    n825,
    n809,
    n772
  );


  xnor
  g856
  (
    n888,
    n792,
    n805,
    n777,
    n776
  );


  or
  g857
  (
    n873,
    n786,
    n826,
    n806,
    n870
  );


  nand
  g858
  (
    n907,
    n837,
    n850,
    n856,
    n843
  );


  xnor
  g859
  (
    n903,
    n678,
    n887,
    n832,
    n657
  );


  xor
  g860
  (
    n928,
    n840,
    n834,
    n657,
    n516
  );


  nand
  g861
  (
    n902,
    n659,
    n848,
    n858,
    n658
  );


  and
  g862
  (
    n892,
    n658,
    n887,
    n882,
    n614
  );


  or
  g863
  (
    KeyWire_0_6,
    n835,
    n851,
    n882,
    n847
  );


  nand
  g864
  (
    n904,
    n843,
    n849,
    n887,
    n879
  );


  or
  g865
  (
    n906,
    n881,
    n844,
    n883,
    n677
  );


  and
  g866
  (
    n909,
    n856,
    n659,
    n615,
    n475
  );


  nand
  g867
  (
    n893,
    n657,
    n886,
    n648,
    n888
  );


  xor
  g868
  (
    n921,
    n840,
    n840,
    n659,
    n646
  );


  nor
  g869
  (
    n923,
    n841,
    n885,
    n872,
    n850
  );


  or
  g870
  (
    n918,
    n833,
    n881,
    n851,
    n859
  );


  or
  g871
  (
    n898,
    n845,
    n878,
    n676,
    n842
  );


  nand
  g872
  (
    n894,
    n880,
    n859,
    n849,
    n841
  );


  xnor
  g873
  (
    n934,
    n846,
    n844,
    n881,
    n885
  );


  and
  g874
  (
    n891,
    n846,
    n848,
    n856,
    n658
  );


  xnor
  g875
  (
    n905,
    n886,
    n846,
    n890,
    n883
  );


  or
  g876
  (
    n930,
    n880,
    n881,
    n839,
    n858
  );


  nand
  g877
  (
    n915,
    n615,
    n838,
    n845,
    n884
  );


  nand
  g878
  (
    n927,
    n848,
    n851,
    n884
  );


  xor
  g879
  (
    n908,
    n879,
    n845,
    n871,
    n840
  );


  nand
  g880
  (
    n901,
    n882,
    n858,
    n873
  );


  nand
  g881
  (
    n931,
    n888,
    n890,
    n847,
    n883
  );


  nand
  g882
  (
    n929,
    n676,
    n831,
    n847,
    n845
  );


  and
  g883
  (
    n911,
    n676,
    n659,
    n857,
    n877
  );


  nand
  g884
  (
    n920,
    n883,
    n882,
    n890,
    n842
  );


  nand
  g885
  (
    n895,
    n844,
    n842,
    n857,
    n884
  );


  or
  g886
  (
    n913,
    n677,
    n649,
    n859,
    n847
  );


  xnor
  g887
  (
    n912,
    n851,
    n677,
    n678,
    n679
  );


  nand
  g888
  (
    n925,
    n887,
    n876,
    n890,
    n889
  );


  or
  g889
  (
    n924,
    n889,
    n647,
    n839,
    n855
  );


  nor
  g890
  (
    n916,
    n842,
    n850,
    n886,
    n889
  );


  xnor
  g891
  (
    n914,
    n493,
    n885,
    n857,
    n657
  );


  xnor
  g892
  (
    n900,
    n857,
    n849,
    n516,
    n678
  );


  xor
  g893
  (
    n897,
    n856,
    n874,
    n516,
    n614
  );


  nor
  g894
  (
    n919,
    n886,
    n679,
    n880,
    n615
  );


  or
  g895
  (
    n933,
    n879,
    n614,
    n885,
    n679
  );


  xor
  g896
  (
    n896,
    n839,
    n888,
    n849,
    n880
  );


  and
  g897
  (
    n910,
    n679,
    n888,
    n848,
    n650
  );


  xnor
  g898
  (
    n922,
    n843,
    n875,
    n841,
    n836
  );


  nand
  g899
  (
    n932,
    n859,
    n841,
    n844,
    n846
  );


  nand
  g900
  (
    n917,
    n678,
    n658,
    n889,
    n850
  );


  nor
  g901
  (
    n899,
    n677,
    n615,
    n839,
    n843
  );


  nand
  g902
  (
    n939,
    n931,
    n891,
    n933,
    n929
  );


  nand
  g903
  (
    n937,
    n906,
    n927,
    n896,
    n893
  );


  xnor
  g904
  (
    n935,
    n923,
    n932,
    n897,
    n904
  );


  xnor
  g905
  (
    n940,
    n912,
    n902,
    n921,
    n908
  );


  or
  g906
  (
    n942,
    n913,
    n895,
    n918,
    n920
  );


  and
  g907
  (
    n943,
    n930,
    n911,
    n907,
    n901
  );


  xor
  g908
  (
    n936,
    n892,
    n925,
    n915,
    n934
  );


  nor
  g909
  (
    n941,
    n924,
    n894,
    n899,
    n898
  );


  xor
  g910
  (
    n944,
    n903,
    n916,
    n905,
    n909
  );


  nor
  g911
  (
    n945,
    n900,
    n914,
    n917,
    n928
  );


  nor
  g912
  (
    n938,
    n910,
    n922,
    n919,
    n926
  );


  xor
  KeyGate_0_0
  (
    n494,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n84,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n790,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n184,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n195,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n633,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n926,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n405,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n334,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n520,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n152,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n528,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n267,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n480,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n829,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n456,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


