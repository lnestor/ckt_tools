

module Stat_100_510
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n86,
  n96,
  n117,
  n111,
  n81,
  n80,
  n108,
  n97,
  n92,
  n85,
  n94,
  n93,
  n106,
  n114,
  n107,
  n104,
  n95,
  n113,
  n102,
  n110,
  n90,
  n84,
  n82,
  n91,
  n88,
  n83,
  n118,
  n101,
  n105,
  n100,
  n132,
  n131
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n86;output n96;output n117;output n111;output n81;output n80;output n108;output n97;output n92;output n85;output n94;output n93;output n106;output n114;output n107;output n104;output n95;output n113;output n102;output n110;output n90;output n84;output n82;output n91;output n88;output n83;output n118;output n101;output n105;output n100;output n132;output n131;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n87;wire n89;wire n98;wire n99;wire n103;wire n109;wire n112;wire n115;wire n116;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    n38,
    n13
  );


  not
  g1
  (
    n48,
    n13
  );


  buf
  g2
  (
    KeyWire_0_9,
    n25
  );


  not
  g3
  (
    KeyWire_0_61,
    n27
  );


  not
  g4
  (
    n71,
    n25
  );


  buf
  g5
  (
    KeyWire_0_63,
    n14
  );


  buf
  g6
  (
    n50,
    n8
  );


  buf
  g7
  (
    KeyWire_0_37,
    n14
  );


  buf
  g8
  (
    KeyWire_0_47,
    n20
  );


  buf
  g9
  (
    n65,
    n1
  );


  not
  g10
  (
    KeyWire_0_8,
    n10
  );


  buf
  g11
  (
    KeyWire_0_20,
    n17
  );


  not
  g12
  (
    KeyWire_0_38,
    n19
  );


  not
  g13
  (
    n53,
    n30
  );


  not
  g14
  (
    KeyWire_0_4,
    n25
  );


  not
  g15
  (
    KeyWire_0_58,
    n18
  );


  buf
  g16
  (
    n76,
    n30
  );


  buf
  g17
  (
    KeyWire_0_59,
    n31
  );


  not
  g18
  (
    KeyWire_0_1,
    n10
  );


  buf
  g19
  (
    n77,
    n4
  );


  buf
  g20
  (
    n46,
    n16
  );


  or
  g21
  (
    n59,
    n10,
    n3,
    n23
  );


  and
  g22
  (
    KeyWire_0_35,
    n23,
    n1,
    n20,
    n30
  );


  and
  g23
  (
    n66,
    n29,
    n26,
    n14,
    n13
  );


  xor
  g24
  (
    KeyWire_0_60,
    n17,
    n2,
    n23,
    n24
  );


  and
  g25
  (
    KeyWire_0_28,
    n19,
    n31,
    n28,
    n7
  );


  xor
  g26
  (
    n79,
    n17,
    n26,
    n31,
    n3
  );


  and
  g27
  (
    n62,
    n9,
    n11,
    n22,
    n3
  );


  xnor
  g28
  (
    KeyWire_0_13,
    n6,
    n15,
    n28,
    n16
  );


  nor
  g29
  (
    n45,
    n6,
    n19,
    n18,
    n1
  );


  xor
  g30
  (
    KeyWire_0_14,
    n10,
    n4,
    n8,
    n16
  );


  xnor
  g31
  (
    KeyWire_0_62,
    n18,
    n9,
    n22,
    n14
  );


  nand
  g32
  (
    KeyWire_0_23,
    n24,
    n12,
    n23,
    n29
  );


  xor
  g33
  (
    n33,
    n11,
    n5,
    n25
  );


  xor
  g34
  (
    KeyWire_0_15,
    n24,
    n11,
    n12,
    n5
  );


  and
  g35
  (
    KeyWire_0_51,
    n21,
    n29,
    n18,
    n7
  );


  nand
  g36
  (
    KeyWire_0_45,
    n9,
    n6
  );


  and
  g37
  (
    KeyWire_0_5,
    n12,
    n21,
    n19
  );


  nand
  g38
  (
    KeyWire_0_24,
    n5,
    n20,
    n17,
    n1
  );


  nand
  g39
  (
    KeyWire_0_2,
    n22,
    n2,
    n16,
    n24
  );


  and
  g40
  (
    n73,
    n27,
    n28,
    n11,
    n13
  );


  nand
  g41
  (
    KeyWire_0_32,
    n29,
    n3,
    n8
  );


  nand
  g42
  (
    n39,
    n15,
    n22,
    n7,
    n27
  );


  nand
  g43
  (
    n58,
    n4,
    n30,
    n28,
    n31
  );


  nor
  g44
  (
    KeyWire_0_10,
    n12,
    n20,
    n15
  );


  nand
  g45
  (
    KeyWire_0_6,
    n4,
    n2,
    n27,
    n21
  );


  nand
  g46
  (
    KeyWire_0_34,
    n2,
    n26,
    n7
  );


  nor
  g47
  (
    n94,
    n53,
    n58,
    n51,
    n52
  );


  or
  g48
  (
    KeyWire_0_42,
    n50,
    n67,
    n45,
    n59
  );


  nor
  g49
  (
    KeyWire_0_12,
    n63,
    n53,
    n59,
    n70
  );


  nand
  g50
  (
    n114,
    n41,
    n64,
    n38,
    n74
  );


  nor
  g51
  (
    KeyWire_0_36,
    n69,
    n68,
    n66,
    n48
  );


  or
  g52
  (
    KeyWire_0_0,
    n46,
    n58,
    n52,
    n65
  );


  or
  g53
  (
    n116,
    n39,
    n36,
    n75,
    n43
  );


  xnor
  g54
  (
    n104,
    n73,
    n52,
    n57,
    n60
  );


  xnor
  g55
  (
    KeyWire_0_55,
    n71,
    n65,
    n60,
    n77
  );


  or
  g56
  (
    KeyWire_0_39,
    n78,
    n54,
    n43,
    n53
  );


  or
  g57
  (
    KeyWire_0_30,
    n48,
    n78,
    n47,
    n67
  );


  xnor
  g58
  (
    KeyWire_0_11,
    n48,
    n56,
    n50,
    n78
  );


  xnor
  g59
  (
    KeyWire_0_53,
    n55,
    n47,
    n70,
    n74
  );


  xor
  g60
  (
    KeyWire_0_7,
    n54,
    n77,
    n62,
    n47
  );


  nand
  g61
  (
    KeyWire_0_57,
    n62,
    n67,
    n76,
    n42
  );


  nor
  g62
  (
    KeyWire_0_19,
    n61,
    n75,
    n76,
    n34
  );


  xor
  g63
  (
    n100,
    n38,
    n56,
    n55,
    n68
  );


  and
  g64
  (
    KeyWire_0_26,
    n41,
    n76,
    n64,
    n75
  );


  or
  g65
  (
    n88,
    n61,
    n66,
    n37,
    n73
  );


  xnor
  g66
  (
    KeyWire_0_54,
    n45,
    n46,
    n56,
    n77
  );


  nor
  g67
  (
    n92,
    n58,
    n73,
    n51
  );


  or
  g68
  (
    KeyWire_0_3,
    n79,
    n60,
    n66,
    n40
  );


  nor
  g69
  (
    KeyWire_0_22,
    n57,
    n50,
    n73,
    n48
  );


  xor
  g70
  (
    n106,
    n64,
    n59,
    n39,
    n57
  );


  xnor
  g71
  (
    n103,
    n60,
    n63,
    n55,
    n36
  );


  nand
  g72
  (
    KeyWire_0_48,
    n51,
    n69,
    n74,
    n59
  );


  xnor
  g73
  (
    KeyWire_0_40,
    n68,
    n37,
    n54,
    n50
  );


  or
  g74
  (
    n95,
    n49,
    n74,
    n79,
    n75
  );


  nand
  g75
  (
    KeyWire_0_31,
    n78,
    n64,
    n61,
    n70
  );


  nor
  g76
  (
    KeyWire_0_43,
    n35,
    n72,
    n79,
    n52
  );


  or
  g77
  (
    KeyWire_0_29,
    n57,
    n35,
    n49,
    n71
  );


  nand
  g78
  (
    KeyWire_0_50,
    n58,
    n33,
    n44,
    n62
  );


  nand
  g79
  (
    KeyWire_0_33,
    n44,
    n61,
    n33,
    n65
  );


  xnor
  g80
  (
    KeyWire_0_56,
    n66,
    n67,
    n53,
    n49
  );


  nand
  g81
  (
    KeyWire_0_16,
    n69,
    n55,
    n72,
    n70
  );


  nand
  g82
  (
    KeyWire_0_25,
    n77,
    n68,
    n40,
    n65
  );


  and
  g83
  (
    KeyWire_0_44,
    n62,
    n71,
    n34,
    n49
  );


  nor
  g84
  (
    KeyWire_0_18,
    n47,
    n79,
    n69,
    n71
  );


  nor
  g85
  (
    KeyWire_0_21,
    n72,
    n63,
    n76,
    n54
  );


  and
  g86
  (
    n98,
    n56,
    n72,
    n42,
    n63
  );


  buf
  g87
  (
    KeyWire_0_46,
    n111
  );


  not
  g88
  (
    n121,
    n114
  );


  buf
  g89
  (
    n124,
    n113
  );


  not
  g90
  (
    n123,
    n112
  );


  not
  g91
  (
    n120,
    n110
  );


  nor
  g92
  (
    n129,
    n121,
    n123,
    n117
  );


  or
  g93
  (
    n130,
    n124,
    n32,
    n122,
    n115
  );


  xnor
  g94
  (
    KeyWire_0_41,
    n121,
    n119,
    n32,
    n120
  );


  or
  g95
  (
    KeyWire_0_27,
    n124,
    n32
  );


  xor
  g96
  (
    KeyWire_0_52,
    n121,
    n120,
    n124,
    n118
  );


  and
  g97
  (
    KeyWire_0_49,
    n116,
    n123,
    n122
  );


  xor
  g98
  (
    n132,
    n128,
    n130,
    n129,
    n126
  );


  xnor
  g99
  (
    KeyWire_0_17,
    n127,
    n130,
    n129,
    n125
  );


  xnor
  KeyGate_0_0
  (
    n117,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n61,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n44,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n87,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n75,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n72,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n47,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n111,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n69,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n37,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n78,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n102,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n97,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n63,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n35,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n41,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n82,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n131,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n99,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n118,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n74,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n112,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n90,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n67,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n70,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n105,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n101,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n128,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n57,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n91,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n109,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n84,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n60,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n115,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n49,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n36,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n81,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n55,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n40,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n86,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n89,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n127,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n80,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n119,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n96,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n51,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n122,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n56,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n85,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n125,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n108,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n64,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n126,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n83,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n113,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n110,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n93,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n107,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n68,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n42,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n34,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n52,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n43,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n54,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


