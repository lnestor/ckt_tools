// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_229 written by SynthGen on 2021/04/05 11:23:27
module Stat_2000_229( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n442, n418, n445, n423, n400, n395, n437, n443,
 n450, n430, n454, n1451, n2013, n2014, n1996, n2026,
 n2020, n2024, n2028, n2023, n2027, n2032, n2029, n2021,
 n2031, n2030, n2019, n2017, n2022, n2025, n2016, n2018);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n442, n418, n445, n423, n400, n395, n437, n443,
 n450, n430, n454, n1451, n2013, n2014, n1996, n2026,
 n2020, n2024, n2028, n2023, n2027, n2032, n2029, n2021,
 n2031, n2030, n2019, n2017, n2022, n2025, n2016, n2018;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n396, n397, n398, n399, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n419,
 n420, n421, n422, n424, n425, n426, n427, n428,
 n429, n431, n432, n433, n434, n435, n436, n438,
 n439, n440, n441, n444, n446, n447, n448, n449,
 n451, n452, n453, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n634, n635,
 n636, n637, n638, n639, n640, n641, n642, n643,
 n644, n645, n646, n647, n648, n649, n650, n651,
 n652, n653, n654, n655, n656, n657, n658, n659,
 n660, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685, n686, n687, n688, n689, n690, n691,
 n692, n693, n694, n695, n696, n697, n698, n699,
 n700, n701, n702, n703, n704, n705, n706, n707,
 n708, n709, n710, n711, n712, n713, n714, n715,
 n716, n717, n718, n719, n720, n721, n722, n723,
 n724, n725, n726, n727, n728, n729, n730, n731,
 n732, n733, n734, n735, n736, n737, n738, n739,
 n740, n741, n742, n743, n744, n745, n746, n747,
 n748, n749, n750, n751, n752, n753, n754, n755,
 n756, n757, n758, n759, n760, n761, n762, n763,
 n764, n765, n766, n767, n768, n769, n770, n771,
 n772, n773, n774, n775, n776, n777, n778, n779,
 n780, n781, n782, n783, n784, n785, n786, n787,
 n788, n789, n790, n791, n792, n793, n794, n795,
 n796, n797, n798, n799, n800, n801, n802, n803,
 n804, n805, n806, n807, n808, n809, n810, n811,
 n812, n813, n814, n815, n816, n817, n818, n819,
 n820, n821, n822, n823, n824, n825, n826, n827,
 n828, n829, n830, n831, n832, n833, n834, n835,
 n836, n837, n838, n839, n840, n841, n842, n843,
 n844, n845, n846, n847, n848, n849, n850, n851,
 n852, n853, n854, n855, n856, n857, n858, n859,
 n860, n861, n862, n863, n864, n865, n866, n867,
 n868, n869, n870, n871, n872, n873, n874, n875,
 n876, n877, n878, n879, n880, n881, n882, n883,
 n884, n885, n886, n887, n888, n889, n890, n891,
 n892, n893, n894, n895, n896, n897, n898, n899,
 n900, n901, n902, n903, n904, n905, n906, n907,
 n908, n909, n910, n911, n912, n913, n914, n915,
 n916, n917, n918, n919, n920, n921, n922, n923,
 n924, n925, n926, n927, n928, n929, n930, n931,
 n932, n933, n934, n935, n936, n937, n938, n939,
 n940, n941, n942, n943, n944, n945, n946, n947,
 n948, n949, n950, n951, n952, n953, n954, n955,
 n956, n957, n958, n959, n960, n961, n962, n963,
 n964, n965, n966, n967, n968, n969, n970, n971,
 n972, n973, n974, n975, n976, n977, n978, n979,
 n980, n981, n982, n983, n984, n985, n986, n987,
 n988, n989, n990, n991, n992, n993, n994, n995,
 n996, n997, n998, n999, n1000, n1001, n1002, n1003,
 n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
 n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
 n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
 n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
 n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
 n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
 n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
 n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
 n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
 n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
 n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
 n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
 n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
 n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
 n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
 n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
 n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
 n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
 n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
 n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
 n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
 n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
 n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
 n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
 n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
 n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
 n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
 n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
 n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
 n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
 n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
 n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
 n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
 n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
 n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
 n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
 n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
 n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
 n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
 n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
 n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
 n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
 n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
 n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
 n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
 n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
 n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
 n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
 n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
 n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
 n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
 n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
 n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
 n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
 n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
 n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1452,
 n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
 n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
 n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
 n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
 n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
 n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
 n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
 n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
 n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
 n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
 n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
 n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
 n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
 n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
 n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
 n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
 n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
 n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
 n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
 n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
 n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
 n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
 n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
 n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
 n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
 n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
 n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
 n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
 n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
 n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
 n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
 n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
 n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
 n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
 n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
 n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
 n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
 n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
 n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
 n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
 n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
 n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
 n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
 n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
 n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
 n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
 n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
 n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
 n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
 n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
 n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
 n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
 n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
 n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
 n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
 n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
 n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
 n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
 n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
 n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
 n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
 n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
 n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
 n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
 n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
 n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
 n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
 n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1997,
 n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
 n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2015;

buf  g0 (n44, n1);
buf  g1 (n41, n3);
buf  g2 (n39, n3);
buf  g3 (n40, n2);
buf  g4 (n42, n1);
buf  g5 (n34, n3);
not  g6 (n35, n2);
buf  g7 (n38, n4);
not  g8 (n36, n1);
buf  g9 (n43, n2);
buf  g10 (n46, n3);
buf  g11 (n33, n2);
buf  g12 (n37, n1);
not  g13 (n45, n4);
not  g14 (n53, n41);
buf  g15 (n55, n34);
not  g16 (n87, n35);
buf  g17 (n63, n40);
buf  g18 (n86, n36);
buf  g19 (n85, n36);
buf  g20 (n48, n38);
buf  g21 (n67, n35);
buf  g22 (n62, n35);
not  g23 (n71, n44);
not  g24 (n57, n35);
not  g25 (n60, n42);
not  g26 (n59, n43);
buf  g27 (n79, n44);
not  g28 (n76, n42);
buf  g29 (n74, n42);
buf  g30 (n89, n43);
buf  g31 (n64, n38);
buf  g32 (n61, n39);
not  g33 (n95, n34);
buf  g34 (n75, n44);
not  g35 (n58, n41);
not  g36 (n77, n43);
not  g37 (n92, n37);
not  g38 (n51, n40);
not  g39 (n65, n34);
buf  g40 (n70, n40);
buf  g41 (n50, n40);
not  g42 (n68, n37);
not  g43 (n78, n39);
not  g44 (n91, n36);
buf  g45 (n83, n45);
buf  g46 (n84, n37);
not  g47 (n66, n43);
not  g48 (n93, n41);
buf  g49 (n81, n44);
not  g50 (n90, n38);
not  g51 (n49, n33);
buf  g52 (n54, n42);
buf  g53 (n52, n33);
buf  g54 (n73, n38);
buf  g55 (n80, n34);
buf  g56 (n47, n39);
buf  g57 (n72, n37);
not  g58 (n56, n33);
not  g59 (n94, n39);
not  g60 (n69, n33);
not  g61 (n88, n36);
buf  g62 (n82, n41);
xor  g63 (n97, n51, n55);
xor  g64 (n96, n55, n56, n53, n50);
xor  g65 (n112, n64, n49, n65, n60);
and  g66 (n106, n49, n52, n54, n53);
nand g67 (n102, n65, n56, n61, n60);
xor  g68 (n109, n56, n63, n58, n52);
nor  g69 (n108, n57, n57, n49, n54);
nor  g70 (n105, n50, n59, n54, n64);
xor  g71 (n99, n63, n55, n61, n56);
xor  g72 (n114, n50, n48, n60);
xnor g73 (n100, n48, n57, n47, n50);
nand g74 (n111, n53, n59, n52, n64);
and  g75 (n110, n49, n59, n54, n61);
nand g76 (n113, n63, n62, n58, n64);
xor  g77 (n107, n63, n47, n62);
xnor g78 (n101, n62, n57, n58, n59);
nand g79 (n103, n48, n62, n52, n61);
xnor g80 (n104, n58, n51);
and  g81 (n98, n48, n55, n47, n53);
not  g82 (n123, n101);
buf  g83 (n118, n109);
not  g84 (n116, n113);
not  g85 (n125, n103);
buf  g86 (n120, n100);
nor  g87 (n122, n111, n112, n107);
and  g88 (n119, n98, n112, n113);
xnor g89 (n121, n113, n113, n106, n108);
or   g90 (n115, n111, n111, n110, n112);
xor  g91 (n117, n97, n104, n99, n96);
xnor g92 (n124, n105, n111, n102, n110);
buf  g93 (n135, n116);
not  g94 (n149, n122);
not  g95 (n152, n66);
buf  g96 (n148, n121);
buf  g97 (n128, n67);
not  g98 (n137, n65);
not  g99 (n140, n117);
buf  g100 (n129, n65);
not  g101 (n139, n67);
not  g102 (n131, n119);
buf  g103 (n147, n117);
not  g104 (n154, n124);
buf  g105 (n146, n122);
not  g106 (n155, n120);
not  g107 (n151, n116);
not  g108 (n153, n118);
not  g109 (n143, n120);
not  g110 (n127, n124);
not  g111 (n158, n115);
not  g112 (n134, n117);
not  g113 (n130, n118);
not  g114 (n142, n123);
buf  g115 (n159, n66);
buf  g116 (n156, n66);
not  g117 (n144, n120);
buf  g118 (n145, n68);
not  g119 (n141, n117);
not  g120 (n150, n121);
not  g121 (n157, n67);
or   g122 (n138, n118, n124, n121);
nor  g123 (n126, n66, n68, n119, n123);
nor  g124 (n133, n119, n67, n68, n121);
nor  g125 (n132, n119, n122, n118, n68);
nor  g126 (n136, n120, n122, n123);
buf  g127 (n200, n142);
buf  g128 (n198, n133);
buf  g129 (n187, n130);
not  g130 (n211, n133);
not  g131 (n167, n127);
buf  g132 (n212, n127);
buf  g133 (n221, n128);
buf  g134 (n227, n134);
buf  g135 (n170, n129);
not  g136 (n225, n134);
buf  g137 (n199, n128);
buf  g138 (n219, n143);
not  g139 (n226, n130);
buf  g140 (n223, n129);
not  g141 (n179, n143);
not  g142 (n178, n130);
buf  g143 (n162, n128);
not  g144 (n180, n136);
buf  g145 (n197, n138);
not  g146 (n160, n144);
buf  g147 (n204, n128);
buf  g148 (n171, n145);
buf  g149 (n216, n138);
not  g150 (n190, n144);
buf  g151 (n175, n132);
buf  g152 (n169, n144);
not  g153 (n214, n129);
not  g154 (n208, n132);
not  g155 (n176, n139);
not  g156 (n164, n139);
buf  g157 (n184, n135);
buf  g158 (n163, n133);
not  g159 (n189, n135);
not  g160 (n205, n126);
not  g161 (n215, n126);
buf  g162 (n168, n140);
not  g163 (n177, n141);
not  g164 (n210, n126);
buf  g165 (n166, n131);
not  g166 (n217, n134);
not  g167 (n191, n143);
not  g168 (n202, n137);
buf  g169 (n218, n132);
buf  g170 (n172, n143);
buf  g171 (n196, n132);
not  g172 (n192, n139);
not  g173 (n195, n140);
buf  g174 (n224, n141);
not  g175 (n174, n136);
buf  g176 (n188, n140);
buf  g177 (n165, n137);
buf  g178 (n194, n142);
buf  g179 (n201, n131);
not  g180 (n213, n134);
buf  g181 (n203, n127);
buf  g182 (n193, n141);
not  g183 (n207, n126);
not  g184 (n220, n137);
not  g185 (n209, n135);
not  g186 (n228, n136);
buf  g187 (n222, n144);
buf  g188 (n182, n135);
buf  g189 (n186, n138);
buf  g190 (n185, n131);
buf  g191 (n173, n129);
not  g192 (n161, n142);
nor  g193 (n206, n133, n127, n142, n145);
or   g194 (n183, n140, n137, n130, n131);
and  g195 (n181, n136, n139, n138, n141);
buf  g196 (n252, n165);
not  g197 (n248, n169);
not  g198 (n238, n173);
buf  g199 (n244, n169);
buf  g200 (n237, n171);
not  g201 (n233, n166);
not  g202 (n229, n165);
buf  g203 (n241, n168);
not  g204 (n239, n166);
buf  g205 (n235, n174);
not  g206 (n254, n166);
buf  g207 (n250, n164);
buf  g208 (n236, n172);
buf  g209 (n251, n174);
buf  g210 (n246, n168);
buf  g211 (n245, n167);
buf  g212 (n234, n173);
buf  g213 (n231, n170);
or   g214 (n249, n168, n166);
nand g215 (n243, n163, n160);
or   g216 (n253, n171, n161, n165, n172);
and  g217 (n232, n171, n169, n173, n172);
and  g218 (n230, n174, n165, n162, n167);
xor  g219 (n242, n169, n168, n171, n170);
xnor g220 (n240, n167, n170, n174, n172);
and  g221 (n247, n167, n175, n173, n170);
buf  g222 (n267, n232);
buf  g223 (n268, n232);
buf  g224 (n258, n233);
not  g225 (n272, n234);
not  g226 (n261, n233);
not  g227 (n259, n231);
buf  g228 (n264, n234);
buf  g229 (n260, n231);
buf  g230 (n263, n232);
buf  g231 (n262, n231);
buf  g232 (n265, n231);
not  g233 (n256, n234);
not  g234 (n271, n230);
buf  g235 (n257, n232);
not  g236 (n270, n234);
buf  g237 (n266, n233);
not  g238 (n255, n233);
buf  g239 (n269, n229);
nand g240 (n273, n187, n267, n193);
xor  g241 (n319, n218, n261, n178, n210);
nor  g242 (n298, n255, n204, n207, n219);
nor  g243 (n274, n213, n197, n267, n270);
or   g244 (n275, n188, n208, n198, n192);
nand g245 (n284, n262, n206, n197, n257);
nor  g246 (n297, n210, n263, n217, n177);
or   g247 (n321, n214, n191, n189, n263);
and  g248 (n325, n220, n205, n189, n216);
and  g249 (n289, n199, n260, n264, n192);
or   g250 (n283, n191, n185, n206, n175);
or   g251 (n334, n212, n256, n269, n177);
and  g252 (n277, n208, n182, n177, n211);
or   g253 (n278, n203, n199, n180, n258);
and  g254 (n302, n220, n221, n269, n265);
nand g255 (n292, n259, n210, n266, n186);
or   g256 (n287, n266, n202, n262, n218);
xor  g257 (n282, n221, n184, n206, n215);
or   g258 (n331, n176, n259, n205, n220);
nand g259 (n330, n185, n258, n270, n198);
nor  g260 (n291, n183, n178, n218, n201);
xnor g261 (n301, n207, n222, n184, n175);
xor  g262 (n333, n191, n195, n268, n267);
or   g263 (n310, n216, n260, n175, n187);
xnor g264 (n322, n186, n205, n257, n187);
xnor g265 (n303, n189, n219, n195, n266);
or   g266 (n311, n215, n270, n176, n214);
or   g267 (n314, n192, n262, n199, n220);
and  g268 (n305, n212, n188, n208, n269);
and  g269 (n312, n182, n198, n184, n206);
or   g270 (n323, n211, n193, n203);
xnor g271 (n295, n196, n219, n199, n257);
and  g272 (n324, n177, n213, n189, n190);
nand g273 (n328, n183, n214, n207, n193);
xor  g274 (n332, n258, n255, n262, n182);
nor  g275 (n315, n256, n260, n270, n215);
and  g276 (n317, n202, n256, n210, n258);
xnor g277 (n313, n223, n261, n265, n186);
and  g278 (n307, n181, n200, n183, n211);
xor  g279 (n279, n255, n192, n179, n196);
nand g280 (n288, n257, n266, n259, n200);
nor  g281 (n281, n200, n179, n190, n191);
or   g282 (n327, n201, n209, n204, n188);
or   g283 (n335, n200, n211, n204, n218);
or   g284 (n320, n213, n185, n195, n265);
nand g285 (n326, n222, n194, n217, n221);
nor  g286 (n294, n263, n264, n194, n216);
and  g287 (n304, n197, n195, n181);
or   g288 (n309, n269, n180, n181, n190);
nor  g289 (n285, n194, n205, n221, n209);
xor  g290 (n306, n179, n180, n264, n209);
nand g291 (n296, n214, n203, n212, n183);
xnor g292 (n318, n222, n263, n255, n212);
nor  g293 (n286, n187, n261, n197, n268);
nor  g294 (n299, n256, n185, n213, n259);
nor  g295 (n316, n182, n202, n194, n201);
nand g296 (n336, n265, n204, n178, n208);
nand g297 (n293, n268, n268, n178, n180);
or   g298 (n290, n176, n179, n219, n188);
xor  g299 (n308, n198, n215, n201, n190);
nand g300 (n300, n196, n264, n261, n207);
xor  g301 (n276, n184, n217, n209, n222);
nand g302 (n280, n260, n267, n186, n202);
xnor g303 (n329, n176, n196, n217, n216);
or   g304 (n354, n154, n151, n244, n147);
or   g305 (n353, n147, n148, n236);
nand g306 (n350, n237, n145, n150, n240);
xor  g307 (n351, n153, n147, n154, n275);
nor  g308 (n360, n273, n276, n243, n236);
nand g309 (n346, n146, n235, n243);
and  g310 (n337, n150, n276, n146, n279);
xnor g311 (n352, n150, n274, n243, n151);
nor  g312 (n355, n145, n148, n153, n239);
or   g313 (n347, n235, n151, n239, n154);
and  g314 (n357, n236, n239, n277, n274);
xor  g315 (n342, n242, n279, n152, n241);
nor  g316 (n341, n150, n149, n242, n277);
and  g317 (n348, n149, n146, n278, n241);
nand g318 (n345, n153, n147, n239, n148);
or   g319 (n359, n154, n242, n241, n277);
nand g320 (n340, n243, n273, n237);
nor  g321 (n362, n237, n278, n238, n244);
and  g322 (n339, n152, n276, n241, n238);
or   g323 (n338, n240, n278, n275);
or   g324 (n358, n240, n238, n149, n153);
nor  g325 (n361, n277, n278, n242, n237);
nor  g326 (n343, n149, n151, n244, n275);
xor  g327 (n349, n152, n238, n276, n146);
and  g328 (n344, n152, n273, n244, n236);
nor  g329 (n356, n235, n240, n274);
not  g330 (n375, n343);
buf  g331 (n366, n340);
buf  g332 (n380, n341);
not  g333 (n365, n343);
buf  g334 (n382, n340);
not  g335 (n381, n341);
buf  g336 (n363, n340);
not  g337 (n371, n340);
not  g338 (n369, n342);
buf  g339 (n368, n342);
buf  g340 (n367, n343);
buf  g341 (n370, n339);
not  g342 (n364, n343);
not  g343 (n384, n344);
not  g344 (n383, n342);
not  g345 (n373, n338);
not  g346 (n372, n344);
not  g347 (n374, n344);
buf  g348 (n378, n341);
not  g349 (n377, n342);
not  g350 (n376, n341);
buf  g351 (n379, n344);
nor  g352 (n463, n303, n346, n320, n334);
nand g353 (n393, n297, n384, n289, n299);
xnor g354 (n451, n297, n299, n248, n287);
xor  g355 (n413, n374, n318, n287, n284);
and  g356 (n386, n318, n287, n371, n293);
nor  g357 (n443, n248, n247, n291, n328);
nor  g358 (n388, n332, n375, n316, n369);
xnor g359 (n390, n347, n333, n224, n286);
xor  g360 (n432, n307, n283, n282, n327);
and  g361 (n406, n291, n312, n310, n329);
xor  g362 (n452, n285, n331, n246, n286);
nor  g363 (n408, n379, n314, n324);
or   g364 (n419, n309, n297, n282, n333);
nor  g365 (n392, n380, n292, n249, n321);
and  g366 (n445, n247, n308, n297, n293);
xor  g367 (n421, n371, n315, n312, n280);
nor  g368 (n398, n294, n300, n369, n373);
xor  g369 (n423, n372, n376, n381, n306);
nand g370 (n409, n327, n246, n329, n363);
nor  g371 (n444, n308, n379, n301, n292);
nor  g372 (n449, n316, n223, n298, n326);
nand g373 (n457, n303, n315, n333, n373);
xor  g374 (n431, n324, n333, n245, n377);
xnor g375 (n453, n293, n366, n245, n250);
xor  g376 (n426, n289, n325, n291, n331);
nand g377 (n469, n246, n332, n345, n310);
or   g378 (n425, n367, n364, n249, n370);
or   g379 (n415, n294, n290, n328, n317);
nand g380 (n420, n346, n309, n282, n325);
nor  g381 (n417, n308, n377, n288, n279);
xor  g382 (n436, n332, n346, n323, n368);
xnor g383 (n471, n301, n305, n383, n378);
or   g384 (n395, n322, n313, n328, n321);
xor  g385 (n434, n320, n290, n306, n345);
nor  g386 (n428, n365, n384, n373, n370);
nand g387 (n411, n304, n304, n288, n322);
xor  g388 (n412, n323, n365, n374, n306);
or   g389 (n472, n371, n281, n329, n327);
and  g390 (n407, n334, n283, n330, n368);
and  g391 (n416, n295, n281, n382, n305);
nand g392 (n446, n298, n310, n302, n285);
nor  g393 (n470, n299, n365, n324, n368);
nor  g394 (n418, n317, n285, n346, n323);
xor  g395 (n462, n245, n223, n284, n325);
or   g396 (n399, n316, n319, n309, n279);
and  g397 (n433, n289, n284, n326, n320);
and  g398 (n402, n296, n249, n245, n375);
and  g399 (n430, n312, n307, n223, n364);
nand g400 (n385, n302, n317, n322, n326);
or   g401 (n429, n303, n292, n314, n369);
nand g402 (n466, n246, n325, n334, n300);
nand g403 (n459, n380, n364, n372, n376);
xnor g404 (n404, n224, n301, n311, n287);
or   g405 (n410, n313, n384, n315, n379);
or   g406 (n439, n281, n293, n288, n317);
or   g407 (n467, n321, n281, n308, n290);
xnor g408 (n403, n298, n306, n319, n377);
nand g409 (n391, n383, n373, n315, n370);
nor  g410 (n396, n310, n250, n305, n312);
xor  g411 (n447, n280, n324, n304, n382);
and  g412 (n405, n313, n331, n295, n296);
or   g413 (n401, n382, n378, n291, n311);
xor  g414 (n435, n319, n366, n247, n372);
xor  g415 (n397, n374, n307, n314, n248);
or   g416 (n465, n305, n383, n294, n345);
xor  g417 (n387, n247, n329, n374, n367);
xor  g418 (n448, n376, n384, n371, n282);
xnor g419 (n389, n330, n365, n311, n322);
or   g420 (n441, n378, n318, n295, n364);
nand g421 (n464, n369, n347, n303, n224);
and  g422 (n437, n334, n248, n326, n225);
xor  g423 (n414, n311, n283, n327, n375);
xnor g424 (n456, n286, n302, n380, n330);
xnor g425 (n461, n332, n321, n294, n292);
nand g426 (n460, n381, n331, n304, n289);
and  g427 (n427, n367, n345, n335, n316);
and  g428 (n454, n313, n377, n283, n368);
xor  g429 (n440, n318, n363, n370, n323);
and  g430 (n422, n376, n285, n288, n330);
xor  g431 (n455, n366, n319, n299, n363);
nor  g432 (n450, n363, n366, n290, n302);
xor  g433 (n400, n379, n284, n375, n296);
or   g434 (n438, n300, n249, n301, n382);
xor  g435 (n424, n300, n309, n320, n347);
or   g436 (n458, n380, n296, n298, n367);
and  g437 (n442, n295, n307, n280, n224);
nor  g438 (n394, n280, n381, n372);
xor  g439 (n468, n328, n383, n378, n286);
not  g440 (n511, n354);
buf  g441 (n510, n349);
buf  g442 (n530, n348);
buf  g443 (n490, n354);
not  g444 (n523, n357);
buf  g445 (n526, n455);
not  g446 (n486, n439);
not  g447 (n494, n415);
buf  g448 (n541, n404);
not  g449 (n542, n447);
buf  g450 (n518, n440);
buf  g451 (n528, n399);
buf  g452 (n517, n355);
not  g453 (n491, n349);
buf  g454 (n529, n400);
buf  g455 (n540, n428);
buf  g456 (n475, n355);
buf  g457 (n543, n457);
not  g458 (n536, n398);
buf  g459 (n545, n466);
not  g460 (n502, n435);
buf  g461 (n506, n401);
not  g462 (n527, n357);
buf  g463 (n479, n411);
buf  g464 (n505, n353);
not  g465 (n495, n358);
not  g466 (n499, n353);
not  g467 (n489, n470);
not  g468 (n476, n354);
not  g469 (n493, n420);
not  g470 (n509, n452);
not  g471 (n483, n416);
not  g472 (n513, n405);
not  g473 (n482, n430);
buf  g474 (n537, n412);
buf  g475 (n539, n352);
buf  g476 (n474, n463);
buf  g477 (n531, n352);
not  g478 (n544, n443);
buf  g479 (n535, n421);
not  g480 (n520, n418);
buf  g481 (n512, n438);
not  g482 (n522, n355);
not  g483 (n496, n468);
buf  g484 (n521, n458);
buf  g485 (n549, n358);
not  g486 (n538, n347);
not  g487 (n533, n357);
not  g488 (n484, n422);
not  g489 (n508, n351);
buf  g490 (n546, n349);
buf  g491 (n478, n414);
buf  g492 (n514, n353);
not  g493 (n500, n413);
buf  g494 (n515, n351);
buf  g495 (n485, n437);
not  g496 (n497, n449);
buf  g497 (n488, n432);
buf  g498 (n524, n453);
buf  g499 (n548, n434);
buf  g500 (n487, n355);
buf  g501 (n498, n441);
and  g502 (n503, n424, n350, n349, n357);
xor  g503 (n501, n356, n348, n448, n465);
nand g504 (n525, n352, n445, n469, n451);
nor  g505 (n480, n442, n467, n417, n350);
nand g506 (n547, n356, n425, n444, n471);
nand g507 (n492, n351, n403, n450, n409);
nand g508 (n519, n433, n464, n436, n348);
xnor g509 (n481, n456, n460, n354, n429);
and  g510 (n516, n356, n350, n459);
xor  g511 (n477, n472, n446, n462, n353);
xor  g512 (n532, n407, n358, n410, n426);
and  g513 (n507, n358, n431, n406, n348);
xor  g514 (n473, n397, n356, n461, n454);
nor  g515 (n504, n423, n419, n408, n351);
or   g516 (n534, n402, n396, n352, n427);
not  g517 (n603, n498);
not  g518 (n731, n17);
buf  g519 (n628, n31);
not  g520 (n649, n533);
buf  g521 (n689, n524);
not  g522 (n687, n500);
buf  g523 (n688, n538);
not  g524 (n698, n8);
not  g525 (n680, n336);
buf  g526 (n661, n251);
buf  g527 (n604, n478);
buf  g528 (n735, n509);
buf  g529 (n660, n493);
buf  g530 (n624, n516);
buf  g531 (n684, n14);
not  g532 (n627, n544);
buf  g533 (n676, n22);
buf  g534 (n612, n15);
buf  g535 (n703, n536);
buf  g536 (n618, n507);
buf  g537 (n717, n24);
not  g538 (n577, n359);
buf  g539 (n711, n530);
not  g540 (n696, n523);
buf  g541 (n576, n250);
not  g542 (n588, n482);
buf  g543 (n583, n538);
not  g544 (n555, n530);
buf  g545 (n646, n23);
not  g546 (n574, n504);
buf  g547 (n682, n501);
not  g548 (n550, n548);
not  g549 (n742, n519);
not  g550 (n672, n520);
buf  g551 (n600, n336);
not  g552 (n747, n527);
not  g553 (n563, n11);
buf  g554 (n651, n490);
not  g555 (n573, n519);
buf  g556 (n630, n227);
buf  g557 (n585, n487);
not  g558 (n738, n499);
not  g559 (n566, n499);
buf  g560 (n611, n31);
not  g561 (n652, n253);
not  g562 (n732, n29);
not  g563 (n657, n155);
not  g564 (n751, n537);
not  g565 (n675, n501);
buf  g566 (n620, n536);
buf  g567 (n667, n487);
buf  g568 (n659, n474);
not  g569 (n599, n503);
not  g570 (n720, n492);
not  g571 (n638, n478);
not  g572 (n671, n530);
not  g573 (n610, n156);
not  g574 (n565, n30);
not  g575 (n743, n515);
not  g576 (n551, n496);
buf  g577 (n592, n535);
buf  g578 (n699, n477);
not  g579 (n741, n516);
buf  g580 (n626, n484);
not  g581 (n633, n542);
not  g582 (n558, n519);
buf  g583 (n737, n24);
buf  g584 (n733, n16);
buf  g585 (n632, n485);
not  g586 (n724, n19);
not  g587 (n595, n480);
not  g588 (n679, n520);
buf  g589 (n674, n503);
not  g590 (n669, n533);
buf  g591 (n613, n545);
buf  g592 (n727, n531);
not  g593 (n704, n539);
buf  g594 (n719, n17);
buf  g595 (n609, n498);
not  g596 (n665, n525);
buf  g597 (n695, n521);
not  g598 (n601, n22);
buf  g599 (n647, n535);
not  g600 (n634, n543);
not  g601 (n560, n19);
not  g602 (n643, n517);
buf  g603 (n656, n546);
buf  g604 (n581, n480);
not  g605 (n608, n544);
not  g606 (n655, n360);
buf  g607 (n635, n17);
buf  g608 (n640, n477);
buf  g609 (n637, n492);
not  g610 (n567, n32);
not  g611 (n716, n475);
not  g612 (n553, n529);
not  g613 (n714, n251);
buf  g614 (n664, n541);
not  g615 (n697, n517);
buf  g616 (n622, n5);
not  g617 (n561, n518);
buf  g618 (n653, n527);
not  g619 (n584, n227);
not  g620 (n605, n20);
xnor g621 (n616, n13, n251, n4);
nor  g622 (n700, n225, n503, n25);
xnor g623 (n562, n17, n490, n511, n18);
nand g624 (n739, n362, n524, n513, n31);
xnor g625 (n606, n27, n46, n7, n502);
nor  g626 (n663, n525, n543, n541, n513);
nand g627 (n648, n546, n508, n496, n492);
or   g628 (n598, n9, n16, n481, n250);
or   g629 (n752, n8, n18, n485);
or   g630 (n715, n46, n5, n271, n30);
xor  g631 (n692, n501, n45, n24, n541);
xnor g632 (n569, n534, n272, n492, n500);
nand g633 (n587, n545, n539, n505, n27);
xnor g634 (n590, n11, n510, n523, n155);
and  g635 (n572, n543, n359, n272, n528);
xor  g636 (n641, n30, n499, n15, n253);
and  g637 (n694, n46, n227, n253, n498);
nand g638 (n708, n6, n549, n506, n226);
xnor g639 (n631, n23, n504, n497, n26);
xor  g640 (n644, n542, n507, n6, n547);
nor  g641 (n570, n28, n514, n362, n513);
and  g642 (n668, n359, n503, n486, n539);
and  g643 (n701, n520, n488, n497, n518);
nor  g644 (n691, n489, n529, n8, n496);
nor  g645 (n615, n11, n12, n361, n480);
nand g646 (n639, n487, n272, n510, n491);
nand g647 (n725, n524, n28, n22, n69);
xor  g648 (n706, n477, n497, n14, n28);
nand g649 (n591, n498, n8, n540, n514);
nor  g650 (n580, n497, n522, n533, n495);
and  g651 (n625, n483, n252, n506, n529);
or   g652 (n681, n479, n514, n526, n532);
nand g653 (n607, n524, n251, n335, n483);
nand g654 (n619, n481, n254, n228, n252);
nand g655 (n740, n20, n474, n488, n483);
and  g656 (n753, n547, n489, n490, n496);
xor  g657 (n666, n502, n517, n254, n473);
xnor g658 (n670, n31, n528, n544, n535);
and  g659 (n746, n69, n495, n493, n482);
xnor g660 (n723, n514, n518, n360, n13);
xnor g661 (n557, n474, n26, n21, n482);
xor  g662 (n683, n509, n226, n479, n114);
or   g663 (n552, n529, n21, n535, n537);
xor  g664 (n678, n21, n522, n501, n549);
or   g665 (n589, n491, n486, n533, n484);
xnor g666 (n712, n482, n45, n540, n483);
xor  g667 (n710, n548, n4, n481, n479);
xor  g668 (n594, n225, n537, n359, n546);
or   g669 (n709, n271, n16, n508, n25);
xor  g670 (n586, n7, n23, n502, n32);
nor  g671 (n730, n15, n515, n523, n475);
nand g672 (n554, n534, n536, n494);
xor  g673 (n636, n46, n516, n10, n512);
or   g674 (n748, n537, n362, n14, n542);
or   g675 (n685, n28, n9, n10, n543);
or   g676 (n617, n532, n360, n6, n507);
nor  g677 (n745, n547, n252, n542, n13);
nand g678 (n690, n508, n525, n528, n549);
xnor g679 (n729, n526, n522, n495, n271);
or   g680 (n702, n494, n491, n476, n525);
nor  g681 (n559, n511, n521, n480, n488);
and  g682 (n596, n486, n361, n511);
nand g683 (n658, n475, n19, n545, n512);
nor  g684 (n707, n547, n517, n540, n493);
and  g685 (n571, n45, n253, n538, n476);
xor  g686 (n749, n489, n494, n531);
nand g687 (n654, n272, n519, n531, n29);
or   g688 (n722, n155, n13, n26, n25);
and  g689 (n614, n549, n486, n5, n506);
nor  g690 (n602, n11, n476, n474, n512);
xnor g691 (n734, n507, n493, n532, n479);
or   g692 (n728, n544, n500, n26, n22);
nand g693 (n718, n540, n30, n484, n520);
nand g694 (n593, n271, n505, n6, n29);
xnor g695 (n642, n548, n9, n522, n227);
nand g696 (n623, n509, n155, n15, n12);
xnor g697 (n736, n114, n29, n516, n510);
xnor g698 (n686, n27, n504, n528, n484);
xor  g699 (n578, n491, n548, n521, n12);
xor  g700 (n645, n504, n509, n473, n539);
xnor g701 (n597, n114, n25, n10, n27);
or   g702 (n662, n505, n476, n473, n485);
nor  g703 (n564, n20, n18, n226, n495);
nor  g704 (n575, n490, n521, n487, n475);
or   g705 (n621, n505, n510, n360, n23);
nand g706 (n556, n32, n526, n534, n499);
nand g707 (n705, n538, n7, n513, n478);
nor  g708 (n582, n19, n335, n500, n546);
or   g709 (n744, n477, n512, n254, n545);
xnor g710 (n673, n336, n228, n10, n511);
nor  g711 (n713, n531, n530, n489, n527);
xnor g712 (n568, n114, n534, n481, n523);
nand g713 (n579, n506, n515, n527, n7);
or   g714 (n693, n225, n32, n21, n515);
xor  g715 (n721, n485, n502, n14, n254);
nor  g716 (n629, n478, n518, n5, n488);
xnor g717 (n650, n336, n226, n16, n20);
xnor g718 (n677, n252, n541, n9, n361);
xor  g719 (n750, n508, n473, n12, n24);
and  g720 (n726, n532, n362, n335, n526);
xor  g721 (n817, n744, n729, n740, n684);
and  g722 (n946, n643, n667, n732, n702);
xnor g723 (n900, n673, n564, n646, n633);
xnor g724 (n834, n696, n741, n722, n610);
nor  g725 (n947, n651, n656, n717, n718);
nand g726 (n790, n573, n599, n676, n690);
xnor g727 (n943, n662, n662, n637, n701);
nand g728 (n853, n574, n737, n685, n591);
nor  g729 (n833, n614, n604, n557, n593);
xnor g730 (n801, n709, n604, n725, n552);
or   g731 (n887, n724, n592, n615, n554);
xnor g732 (n886, n681, n586, n625, n617);
nor  g733 (n821, n738, n589, n595, n722);
xnor g734 (n938, n653, n700, n745, n660);
or   g735 (n941, n634, n698, n598, n719);
and  g736 (n806, n690, n615, n725, n650);
or   g737 (n936, n572, n701, n680, n661);
xor  g738 (n885, n734, n606, n634, n731);
xor  g739 (n772, n697, n695, n707, n653);
or   g740 (n765, n578, n720, n638, n572);
and  g741 (n917, n711, n636, n716, n715);
or   g742 (n892, n641, n645, n732, n573);
and  g743 (n774, n737, n666, n659, n681);
xor  g744 (n896, n613, n693, n638, n660);
or   g745 (n915, n734, n620, n623);
nand g746 (n763, n651, n668, n714, n615);
xor  g747 (n762, n659, n724, n645, n562);
xor  g748 (n828, n729, n628, n705, n706);
or   g749 (n795, n631, n609, n603, n710);
xnor g750 (n856, n647, n704, n743, n700);
xnor g751 (n913, n702, n666, n601, n664);
xnor g752 (n756, n604, n576, n710, n654);
xor  g753 (n788, n645, n594, n660, n564);
nor  g754 (n781, n596, n639, n633, n643);
or   g755 (n820, n678, n715, n658);
xor  g756 (n819, n555, n686, n570, n729);
xor  g757 (n842, n626, n730, n643, n632);
nor  g758 (n912, n607, n734, n568, n710);
and  g759 (n793, n677, n733, n575, n687);
nor  g760 (n816, n591, n651, n650, n728);
and  g761 (n901, n629, n602, n581, n746);
nand g762 (n870, n686, n625, n616, n637);
and  g763 (n868, n727, n662, n624, n742);
nand g764 (n893, n739, n741, n726, n666);
and  g765 (n875, n683, n682, n627, n689);
xnor g766 (n832, n580, n711, n694);
xnor g767 (n823, n706, n579, n657, n711);
nand g768 (n903, n685, n623, n682, n617);
nor  g769 (n789, n691, n660, n635, n671);
xor  g770 (n888, n738, n669, n562, n559);
nor  g771 (n775, n608, n680, n576, n574);
nand g772 (n771, n616, n621, n695, n678);
nor  g773 (n931, n665, n645, n554, n628);
nor  g774 (n845, n550, n705, n558, n634);
and  g775 (n773, n579, n670, n576, n693);
and  g776 (n792, n712, n640, n656, n718);
or   g777 (n862, n665, n621, n694, n554);
and  g778 (n778, n656, n650, n596, n608);
nor  g779 (n928, n727, n675, n746, n717);
xnor g780 (n920, n591, n667, n603, n628);
xnor g781 (n841, n649, n692, n565, n558);
xor  g782 (n935, n681, n703, n556, n678);
nor  g783 (n785, n570, n626, n607, n585);
nor  g784 (n805, n653, n613, n576, n583);
or   g785 (n837, n730, n657, n653, n593);
and  g786 (n881, n725, n627, n567, n640);
nand g787 (n754, n667, n586, n661, n655);
xnor g788 (n876, n558, n569, n643, n577);
or   g789 (n867, n721, n628, n613, n633);
and  g790 (n949, n713, n639, n590, n609);
xor  g791 (n871, n707, n734, n672, n635);
xor  g792 (n826, n649, n708, n673, n641);
xnor g793 (n923, n738, n611, n590, n722);
nor  g794 (n940, n710, n599, n608, n638);
xor  g795 (n846, n617, n691, n658, n604);
or   g796 (n797, n744, n741, n667, n706);
xor  g797 (n909, n605, n714, n718, n732);
xor  g798 (n770, n584, n663, n672, n568);
nand g799 (n847, n678, n730, n703, n652);
nand g800 (n861, n620, n601, n685, n579);
and  g801 (n878, n614, n641, n708, n624);
xnor g802 (n844, n636, n618, n624, n575);
xor  g803 (n898, n566, n583, n683, n601);
and  g804 (n884, n691, n612, n702, n597);
or   g805 (n944, n625, n597, n590, n716);
or   g806 (n905, n735, n614, n685, n740);
nand g807 (n916, n570, n606, n571, n669);
nand g808 (n919, n562, n629, n666, n716);
nand g809 (n840, n559, n738, n578, n720);
nand g810 (n836, n563, n686, n568, n698);
xor  g811 (n776, n674, n627, n584, n670);
and  g812 (n796, n609, n574, n599, n572);
and  g813 (n812, n584, n654, n629, n565);
xor  g814 (n921, n578, n618, n726, n602);
or   g815 (n902, n739, n632, n617, n593);
or   g816 (n942, n625, n567, n727, n595);
xor  g817 (n780, n675, n661, n707, n571);
nand g818 (n798, n697, n658, n600, n664);
nand g819 (n835, n587, n562, n572, n646);
or   g820 (n922, n644, n632, n647, n621);
xor  g821 (n910, n742, n669, n557, n688);
nor  g822 (n760, n743, n654, n695, n726);
and  g823 (n894, n591, n745, n641, n671);
or   g824 (n764, n599, n691, n730, n596);
nor  g825 (n877, n690, n728, n632, n619);
nand g826 (n777, n610, n677, n589, n657);
nor  g827 (n880, n631, n642, n671, n652);
xor  g828 (n859, n684, n593, n647, n665);
and  g829 (n945, n575, n704, n651, n569);
nand g830 (n883, n578, n672, n620, n588);
or   g831 (n874, n740, n614, n670, n693);
xor  g832 (n794, n638, n582, n580, n655);
nand g833 (n873, n713, n716, n586, n564);
nand g834 (n767, n639, n648, n550, n717);
and  g835 (n891, n634, n704, n665, n649);
xnor g836 (n889, n598, n595, n557, n693);
nand g837 (n934, n630, n606, n689, n605);
nor  g838 (n786, n726, n676, n592, n699);
nand g839 (n851, n664, n563, n635, n640);
nor  g840 (n897, n687, n622, n696, n736);
nor  g841 (n911, n675, n597, n690, n587);
xnor g842 (n825, n631, n602, n573);
or   g843 (n854, n560, n605, n656, n742);
nand g844 (n830, n668, n717, n612, n619);
xnor g845 (n924, n594, n636, n680, n575);
nor  g846 (n803, n571, n679, n731, n705);
and  g847 (n855, n559, n689, n673, n610);
and  g848 (n899, n649, n565, n580, n637);
or   g849 (n918, n555, n592, n673, n736);
nand g850 (n782, n630, n733, n692, n598);
nand g851 (n864, n611, n664, n630, n581);
nor  g852 (n869, n657, n705, n655, n580);
xor  g853 (n814, n619, n719, n743, n703);
nor  g854 (n758, n636, n642, n723, n676);
xnor g855 (n926, n713, n719, n626, n712);
nor  g856 (n848, n627, n567, n621, n733);
xor  g857 (n895, n719, n619, n596, n559);
and  g858 (n827, n686, n588, n680, n709);
nand g859 (n800, n583, n721, n571, n679);
and  g860 (n779, n644, n683, n682, n611);
xor  g861 (n759, n583, n631, n681, n612);
nand g862 (n810, n737, n739, n552, n736);
and  g863 (n809, n677, n674, n551, n732);
nor  g864 (n824, n588, n577, n553, n708);
and  g865 (n890, n581, n682, n724, n556);
or   g866 (n860, n745, n652, n568, n699);
and  g867 (n925, n647, n560, n715, n742);
xnor g868 (n808, n700, n701, n737, n646);
nand g869 (n849, n695, n676, n736, n696);
and  g870 (n783, n607, n561, n699, n721);
nand g871 (n757, n741, n689, n677, n585);
xnor g872 (n937, n563, n701, n603, n553);
nor  g873 (n839, n563, n607, n702, n744);
nand g874 (n852, n708, n587, n697, n616);
nand g875 (n791, n698, n609, n605, n706);
and  g876 (n950, n569, n699, n671, n561);
xnor g877 (n929, n692, n644, n557, n570);
xnor g878 (n939, n746, n640, n744, n556);
or   g879 (n815, n692, n574, n622, n735);
or   g880 (n914, n594, n560, n561, n720);
xor  g881 (n818, n674, n700, n551, n615);
nor  g882 (n755, n694, n633, n731, n740);
nand g883 (n882, n551, n644, n600, n564);
or   g884 (n838, n648, n637, n561, n552);
xnor g885 (n766, n608, n713, n674, n712);
nor  g886 (n768, n590, n623, n723, n577);
or   g887 (n787, n612, n554, n735, n715);
or   g888 (n904, n581, n553, n698, n556);
or   g889 (n811, n724, n582, n626);
and  g890 (n829, n565, n594, n723, n603);
and  g891 (n863, n600, n642, n727, n566);
xnor g892 (n930, n683, n723, n551, n670);
nand g893 (n879, n550, n655, n577, n582);
or   g894 (n807, n661, n725, n567, n648);
and  g895 (n799, n585, n550, n659, n668);
nand g896 (n933, n624, n712, n579, n663);
nor  g897 (n872, n659, n592, n587, n586);
nor  g898 (n908, n718, n662, n669, n642);
or   g899 (n784, n684, n618, n622, n687);
xor  g900 (n906, n668, n630, n721, n553);
nand g901 (n857, n696, n687, n733, n731);
nor  g902 (n850, n639, n672, n589, n654);
xnor g903 (n907, n735, n635, n618, n688);
nor  g904 (n761, n555, n566, n558, n739);
and  g905 (n858, n613, n560, n652, n709);
xnor g906 (n769, n714, n595, n688, n555);
xor  g907 (n948, n585, n711, n722, n679);
and  g908 (n831, n610, n675, n606, n697);
xor  g909 (n927, n611, n569, n745, n650);
xnor g910 (n843, n743, n597, n663, n707);
nor  g911 (n866, n703, n552, n663, n598);
nand g912 (n932, n729, n728, n646, n622);
nor  g913 (n804, n688, n616, n679, n704);
and  g914 (n865, n709, n566, n600, n588);
nand g915 (n802, n629, n648, n746, n728);
and  g916 (n813, n601, n602, n589, n684);
nand g917 (n822, n584, n623, n714, n720);
not  g918 (n1031, n936);
not  g919 (n1053, n788);
not  g920 (n1130, n881);
not  g921 (n1080, n810);
buf  g922 (n981, n785);
buf  g923 (n1034, n73);
not  g924 (n1051, n926);
buf  g925 (n972, n82);
buf  g926 (n975, n917);
not  g927 (n1063, n83);
buf  g928 (n1146, n773);
buf  g929 (n1056, n944);
buf  g930 (n1043, n859);
not  g931 (n1082, n857);
buf  g932 (n970, n890);
buf  g933 (n1040, n891);
not  g934 (n1083, n875);
not  g935 (n957, n796);
buf  g936 (n1020, n795);
not  g937 (n1089, n943);
buf  g938 (n1116, n885);
buf  g939 (n1052, n790);
not  g940 (n1047, n820);
buf  g941 (n1109, n887);
buf  g942 (n1045, n764);
not  g943 (n1137, n892);
buf  g944 (n1131, n82);
not  g945 (n1028, n812);
buf  g946 (n1114, n77);
not  g947 (n1105, n830);
not  g948 (n1097, n770);
not  g949 (n1081, n873);
not  g950 (n1029, n69);
buf  g951 (n977, n841);
buf  g952 (n964, n80);
buf  g953 (n1099, n828);
not  g954 (n1087, n907);
not  g955 (n1016, n901);
buf  g956 (n1027, n851);
buf  g957 (n979, n77);
not  g958 (n1094, n902);
buf  g959 (n1098, n900);
not  g960 (n1007, n72);
not  g961 (n1019, n755);
not  g962 (n1122, n769);
not  g963 (n1125, n78);
buf  g964 (n1133, n79);
not  g965 (n1003, n777);
not  g966 (n1011, n883);
not  g967 (n1004, n789);
buf  g968 (n1023, n80);
not  g969 (n961, n776);
not  g970 (n1127, n767);
not  g971 (n1103, n914);
buf  g972 (n1135, n836);
not  g973 (n1120, n805);
not  g974 (n1074, n807);
buf  g975 (n1046, n74);
buf  g976 (n1073, n782);
buf  g977 (n1128, n861);
buf  g978 (n1041, n825);
not  g979 (n953, n70);
buf  g980 (n1036, n79);
not  g981 (n1093, n950);
not  g982 (n1044, n922);
buf  g983 (n1060, n77);
buf  g984 (n1129, n945);
not  g985 (n983, n910);
not  g986 (n1124, n870);
not  g987 (n973, n813);
buf  g988 (n1049, n821);
not  g989 (n1091, n838);
not  g990 (n1070, n85);
not  g991 (n1111, n905);
not  g992 (n1033, n792);
buf  g993 (n1014, n806);
not  g994 (n1005, n76);
buf  g995 (n1104, n74);
buf  g996 (n1144, n886);
buf  g997 (n985, n768);
not  g998 (n1138, n787);
buf  g999 (n989, n837);
not  g1000 (n1022, n935);
not  g1001 (n1030, n804);
not  g1002 (n1054, n920);
not  g1003 (n1143, n81);
buf  g1004 (n1096, n82);
not  g1005 (n1134, n876);
not  g1006 (n1050, n889);
buf  g1007 (n966, n758);
buf  g1008 (n990, n898);
buf  g1009 (n1084, n933);
buf  g1010 (n1078, n754);
buf  g1011 (n991, n784);
not  g1012 (n1008, n940);
buf  g1013 (n1048, n853);
buf  g1014 (n1072, n893);
buf  g1015 (n952, n930);
buf  g1016 (n1059, n868);
not  g1017 (n994, n903);
buf  g1018 (n1075, n948);
not  g1019 (n1092, n867);
not  g1020 (n980, n75);
buf  g1021 (n1119, n896);
buf  g1022 (n1140, n763);
not  g1023 (n1058, n929);
not  g1024 (n1001, n835);
not  g1025 (n971, n947);
buf  g1026 (n1062, n84);
buf  g1027 (n967, n878);
buf  g1028 (n1035, n76);
buf  g1029 (n1141, n874);
not  g1030 (n1101, n84);
not  g1031 (n1018, n882);
not  g1032 (n993, n80);
not  g1033 (n992, n80);
not  g1034 (n1064, n83);
buf  g1035 (n1112, n832);
not  g1036 (n1017, n70);
not  g1037 (n987, n82);
buf  g1038 (n1024, n879);
buf  g1039 (n997, n923);
buf  g1040 (n984, n75);
not  g1041 (n1021, n924);
buf  g1042 (n995, n760);
buf  g1043 (n1117, n778);
buf  g1044 (n968, n843);
not  g1045 (n1113, n70);
not  g1046 (n1085, n872);
not  g1047 (n1013, n85);
buf  g1048 (n1106, n781);
buf  g1049 (n976, n942);
buf  g1050 (n1002, n783);
not  g1051 (n1095, n817);
buf  g1052 (n1123, n844);
not  g1053 (n1012, n800);
buf  g1054 (n1067, n762);
buf  g1055 (n1032, n794);
buf  g1056 (n1042, n76);
buf  g1057 (n1107, n79);
buf  g1058 (n1057, n73);
not  g1059 (n1102, n81);
buf  g1060 (n1115, n84);
buf  g1061 (n1025, n74);
buf  g1062 (n982, n765);
buf  g1063 (n1039, n869);
not  g1064 (n1026, n927);
not  g1065 (n1009, n72);
buf  g1066 (n958, n864);
not  g1067 (n954, n818);
not  g1068 (n1077, n809);
buf  g1069 (n1139, n848);
not  g1070 (n1055, n76);
buf  g1071 (n1121, n849);
not  g1072 (n999, n909);
not  g1073 (n1066, n831);
not  g1074 (n956, n949);
buf  g1075 (n951, n79);
buf  g1076 (n988, n906);
not  g1077 (n959, n888);
buf  g1078 (n1038, n756);
not  g1079 (n1006, n803);
not  g1080 (n1100, n855);
not  g1081 (n1108, n827);
buf  g1082 (n1132, n815);
not  g1083 (n1068, n941);
buf  g1084 (n1000, n829);
not  g1085 (n1069, n774);
not  g1086 (n1076, n78);
buf  g1087 (n965, n83);
not  g1088 (n1086, n75);
buf  g1089 (n1088, n816);
not  g1090 (n1142, n834);
not  g1091 (n974, n852);
xor  g1092 (n978, n801, n799, n850, n69);
nor  g1093 (n955, n802, n932, n921, n822);
or   g1094 (n1126, n72, n819, n793, n71);
xor  g1095 (n998, n797, n761, n808, n928);
xnor g1096 (n996, n84, n775, n71, n880);
nor  g1097 (n1079, n919, n871, n911, n81);
nand g1098 (n1010, n854, n70, n858, n824);
nand g1099 (n962, n860, n894, n842, n938);
and  g1100 (n1118, n83, n73, n863, n77);
nor  g1101 (n1071, n826, n913, n759, n912);
xnor g1102 (n1061, n884, n78, n72, n71);
or   g1103 (n960, n846, n772, n771, n823);
or   g1104 (n1037, n897, n865, n798, n78);
xor  g1105 (n1090, n845, n934, n939, n757);
xor  g1106 (n1145, n908, n895, n833, n946);
xor  g1107 (n1015, n918, n899, n85, n814);
and  g1108 (n963, n916, n780, n779, n81);
xnor g1109 (n1065, n766, n877, n811, n73);
nor  g1110 (n1110, n866, n847, n931, n925);
or   g1111 (n1136, n937, n840, n75, n915);
xnor g1112 (n986, n791, n786, n71, n862);
xor  g1113 (n969, n74, n856, n839, n904);
not  g1114 (n1311, n1025);
buf  g1115 (n1286, n1000);
not  g1116 (n1280, n753);
buf  g1117 (n1276, n993);
not  g1118 (n1282, n972);
buf  g1119 (n1237, n993);
not  g1120 (n1297, n1008);
buf  g1121 (n1313, n1040);
buf  g1122 (n1373, n982);
buf  g1123 (n1227, n968);
not  g1124 (n1290, n957);
buf  g1125 (n1193, n962);
not  g1126 (n1263, n1007);
not  g1127 (n1339, n1038);
buf  g1128 (n1296, n996);
buf  g1129 (n1180, n1010);
buf  g1130 (n1255, n974);
buf  g1131 (n1405, n752);
buf  g1132 (n1302, n969);
buf  g1133 (n1248, n982);
buf  g1134 (n1314, n1030);
not  g1135 (n1316, n1038);
not  g1136 (n1184, n967);
not  g1137 (n1164, n994);
not  g1138 (n1204, n957);
not  g1139 (n1249, n1018);
buf  g1140 (n1269, n995);
buf  g1141 (n1403, n973);
buf  g1142 (n1327, n983);
not  g1143 (n1163, n1027);
not  g1144 (n1289, n964);
buf  g1145 (n1258, n970);
not  g1146 (n1247, n975);
not  g1147 (n1400, n955);
not  g1148 (n1185, n1031);
buf  g1149 (n1354, n1032);
buf  g1150 (n1241, n1040);
not  g1151 (n1391, n998);
not  g1152 (n1179, n953);
buf  g1153 (n1293, n1027);
not  g1154 (n1157, n1015);
buf  g1155 (n1343, n1024);
not  g1156 (n1190, n1026);
not  g1157 (n1226, n1041);
not  g1158 (n1332, n991);
buf  g1159 (n1234, n979);
buf  g1160 (n1315, n1009);
not  g1161 (n1394, n975);
not  g1162 (n1261, n978);
buf  g1163 (n1246, n981);
not  g1164 (n1397, n1013);
not  g1165 (n1324, n994);
buf  g1166 (n1162, n953);
not  g1167 (n1168, n957);
not  g1168 (n1380, n1027);
buf  g1169 (n1377, n965);
not  g1170 (n1155, n1017);
buf  g1171 (n1298, n1005);
buf  g1172 (n1338, n972);
not  g1173 (n1195, n1026);
not  g1174 (n1360, n1002);
buf  g1175 (n1275, n974);
buf  g1176 (n1328, n954);
buf  g1177 (n1250, n1018);
not  g1178 (n1378, n1013);
buf  g1179 (n1148, n1023);
buf  g1180 (n1156, n993);
buf  g1181 (n1172, n1023);
not  g1182 (n1294, n1028);
not  g1183 (n1173, n974);
not  g1184 (n1308, n984);
not  g1185 (n1174, n1017);
buf  g1186 (n1270, n959);
buf  g1187 (n1187, n750);
buf  g1188 (n1346, n997);
not  g1189 (n1287, n977);
buf  g1190 (n1228, n1019);
not  g1191 (n1166, n1004);
buf  g1192 (n1303, n1028);
not  g1193 (n1205, n1019);
not  g1194 (n1387, n1037);
not  g1195 (n1375, n967);
not  g1196 (n1238, n980);
buf  g1197 (n1370, n961);
buf  g1198 (n1331, n750);
buf  g1199 (n1178, n990);
buf  g1200 (n1356, n973);
buf  g1201 (n1323, n1005);
not  g1202 (n1344, n1042);
not  g1203 (n1288, n1005);
not  g1204 (n1169, n956);
not  g1205 (n1197, n1040);
not  g1206 (n1279, n962);
buf  g1207 (n1398, n961);
buf  g1208 (n1264, n974);
not  g1209 (n1257, n1019);
buf  g1210 (n1242, n958);
not  g1211 (n1244, n970);
not  g1212 (n1272, n998);
not  g1213 (n1212, n1003);
not  g1214 (n1167, n1030);
buf  g1215 (n1299, n1000);
buf  g1216 (n1215, n971);
buf  g1217 (n1367, n971);
buf  g1218 (n1229, n1034);
not  g1219 (n1231, n954);
not  g1220 (n1158, n1038);
not  g1221 (n1194, n984);
not  g1222 (n1199, n1037);
not  g1223 (n1353, n966);
buf  g1224 (n1281, n991);
not  g1225 (n1235, n1032);
buf  g1226 (n1364, n960);
not  g1227 (n1189, n964);
buf  g1228 (n1236, n996);
not  g1229 (n1183, n1006);
buf  g1230 (n1191, n1003);
buf  g1231 (n1301, n976);
not  g1232 (n1218, n1026);
not  g1233 (n1347, n963);
not  g1234 (n1350, n988);
buf  g1235 (n1390, n981);
buf  g1236 (n1222, n988);
not  g1237 (n1351, n1016);
not  g1238 (n1192, n999);
buf  g1239 (n1319, n1029);
not  g1240 (n1355, n753);
buf  g1241 (n1225, n993);
not  g1242 (n1150, n1014);
buf  g1243 (n1152, n1039);
not  g1244 (n1216, n977);
buf  g1245 (n1147, n976);
buf  g1246 (n1243, n1000);
not  g1247 (n1240, n959);
buf  g1248 (n1340, n1017);
buf  g1249 (n1278, n752);
buf  g1250 (n1304, n1024);
not  g1251 (n1366, n995);
not  g1252 (n1300, n976);
not  g1253 (n1233, n987);
buf  g1254 (n1345, n975);
not  g1255 (n1379, n961);
buf  g1256 (n1392, n989);
buf  g1257 (n1160, n967);
buf  g1258 (n1369, n1022);
buf  g1259 (n1200, n989);
buf  g1260 (n1371, n979);
not  g1261 (n1395, n1041);
not  g1262 (n1309, n1009);
not  g1263 (n1386, n979);
not  g1264 (n1165, n977);
buf  g1265 (n1196, n1015);
buf  g1266 (n1224, n1007);
not  g1267 (n1352, n1035);
buf  g1268 (n1306, n967);
not  g1269 (n1161, n749);
not  g1270 (n1388, n1004);
not  g1271 (n1251, n985);
not  g1272 (n1273, n1012);
not  g1273 (n1383, n1002);
not  g1274 (n1341, n1005);
buf  g1275 (n1358, n1001);
not  g1276 (n1334, n1007);
buf  g1277 (n1262, n983);
buf  g1278 (n1385, n970);
buf  g1279 (n1349, n963);
not  g1280 (n1271, n749);
buf  g1281 (n1203, n1013);
buf  g1282 (n1359, n1009);
buf  g1283 (n1329, n1036);
not  g1284 (n1317, n1006);
buf  g1285 (n1362, n747);
not  g1286 (n1266, n747);
buf  g1287 (n1188, n1035);
not  g1288 (n1210, n1037);
not  g1289 (n1333, n964);
buf  g1290 (n1211, n1016);
buf  g1291 (n1177, n968);
not  g1292 (n1335, n990);
buf  g1293 (n1245, n969);
buf  g1294 (n1342, n1032);
not  g1295 (n1292, n980);
buf  g1296 (n1223, n989);
not  g1297 (n1322, n997);
buf  g1298 (n1206, n1009);
not  g1299 (n1283, n977);
buf  g1300 (n1337, n751);
buf  g1301 (n1406, n1024);
buf  g1302 (n1284, n1013);
not  g1303 (n1368, n1022);
buf  g1304 (n1348, n1024);
not  g1305 (n1259, n981);
buf  g1306 (n1176, n1028);
buf  g1307 (n1267, n1038);
not  g1308 (n1381, n1008);
buf  g1309 (n1357, n1040);
not  g1310 (n1363, n1030);
not  g1311 (n1149, n1000);
not  g1312 (n1399, n999);
not  g1313 (n1365, n1021);
not  g1314 (n1312, n969);
buf  g1315 (n1201, n1017);
buf  g1316 (n1171, n1021);
not  g1317 (n1326, n1042);
buf  g1318 (n1291, n1004);
not  g1319 (n1252, n1006);
not  g1320 (n1401, n1001);
not  g1321 (n1151, n1003);
not  g1322 (n1208, n985);
not  g1323 (n1159, n982);
buf  g1324 (n1310, n751);
not  g1325 (n1374, n962);
buf  g1326 (n1361, n1033);
not  g1327 (n1295, n975);
buf  g1328 (n1320, n1041);
not  g1329 (n1170, n984);
buf  g1330 (n1407, n1003);
xor  g1331 (n1376, n1033, n1034);
xnor g1332 (n1372, n965, n1032, n992, n751);
xnor g1333 (n1256, n751, n1031, n1039, n997);
nand g1334 (n1209, n1026, n992, n986, n750);
xnor g1335 (n1325, n995, n973, n1011, n987);
or   g1336 (n1207, n1030, n973, n1029, n966);
xnor g1337 (n1285, n1010, n1006, n1035, n957);
xnor g1338 (n1404, n972, n952, n1012, n750);
xnor g1339 (n1274, n986, n978, n968, n1011);
xor  g1340 (n1254, n1020, n951, n976, n1023);
nor  g1341 (n1214, n998, n1042, n956, n966);
xor  g1342 (n1305, n1015, n1008, n1037, n753);
nand g1343 (n1219, n1011, n1039, n958, n954);
xor  g1344 (n1307, n964, n1014, n1001, n1039);
and  g1345 (n1198, n1012, n992, n748, n959);
nand g1346 (n1384, n1029, n983, n990, n994);
nor  g1347 (n1253, n1012, n991, n1020, n1029);
xor  g1348 (n1213, n997, n989, n753, n959);
xor  g1349 (n1396, n1022, n1033, n995, n752);
xor  g1350 (n1220, n972, n978, n1036, n963);
nor  g1351 (n1202, n747, n1018, n979, n1020);
nor  g1352 (n1230, n965, n1036, n982, n962);
nor  g1353 (n1221, n980, n1041, n988, n1021);
xnor g1354 (n1330, n954, n960, n749, n1025);
nand g1355 (n1336, n1034, n1034, n958, n978);
nor  g1356 (n1182, n987, n1020, n955, n1023);
or   g1357 (n1217, n963, n958, n955, n1031);
or   g1358 (n1382, n980, n996, n1001, n956);
xnor g1359 (n1181, n990, n1025, n1027);
or   g1360 (n1393, n1016, n1011, n749, n992);
or   g1361 (n1186, n1010, n1042, n1004, n986);
or   g1362 (n1389, n1002, n999, n1014, n1016);
xor  g1363 (n1239, n998, n985, n969, n1036);
nor  g1364 (n1318, n1043, n981, n1019, n971);
xnor g1365 (n1402, n970, n1028, n968, n984);
or   g1366 (n1277, n955, n994, n999, n971);
xnor g1367 (n1153, n752, n747, n1010, n1007);
and  g1368 (n1268, n966, n987, n1002, n985);
nand g1369 (n1175, n1015, n960, n983, n1031);
xnor g1370 (n1265, n991, n996, n1033, n961);
and  g1371 (n1154, n1018, n748, n988, n960);
xor  g1372 (n1232, n1021, n986, n953);
xor  g1373 (n1260, n1035, n1008, n748, n1014);
xnor g1374 (n1321, n748, n956, n1022, n965);
not  g1375 (n1516, n1295);
buf  g1376 (n1534, n1325);
not  g1377 (n1484, n1272);
buf  g1378 (n1515, n1365);
buf  g1379 (n1589, n1296);
not  g1380 (n1554, n1253);
not  g1381 (n1597, n1292);
not  g1382 (n1560, n1329);
not  g1383 (n1549, n1260);
not  g1384 (n1457, n1326);
not  g1385 (n1466, n1246);
not  g1386 (n1533, n1255);
not  g1387 (n1531, n1209);
not  g1388 (n1444, n1223);
not  g1389 (n1604, n1342);
xnor g1390 (n1553, n1188, n1383, n1155, n1378);
and  g1391 (n1591, n1393, n1376, n1257, n1389);
nor  g1392 (n1525, n1330, n1287, n1358, n1318);
xnor g1393 (n1426, n1298, n1296, n1371, n1378);
nand g1394 (n1448, n1364, n1374, n1402, n1396);
nor  g1395 (n1432, n1150, n1296, n1357, n1339);
xnor g1396 (n1417, n1379, n1352, n1320, n1267);
xor  g1397 (n1546, n1346, n1349, n1336, n1319);
nor  g1398 (n1571, n1372, n1210, n1322, n1313);
xor  g1399 (n1409, n1242, n1394, n1315, n1294);
or   g1400 (n1419, n1264, n1251, n1278, n1252);
and  g1401 (n1411, n1342, n1343, n1386);
and  g1402 (n1593, n1338, n1270, n1395, n1388);
or   g1403 (n1539, n1367, n1391, n1393, n1381);
and  g1404 (n1514, n1365, n1286, n1267, n1256);
xor  g1405 (n1465, n1328, n1304, n1339, n1265);
xnor g1406 (n1559, n1382, n1167, n1293, n1183);
xnor g1407 (n1480, n1399, n1313, n1252, n1287);
and  g1408 (n1552, n1307, n1375, n1372, n1186);
and  g1409 (n1522, n1233, n1392, n1400, n1376);
xnor g1410 (n1478, n1283, n1219, n1318, n1310);
xnor g1411 (n1583, n1198, n1371, n1380, n1215);
and  g1412 (n1418, n1353, n1251, n1290, n1311);
and  g1413 (n1575, n1363, n1290, n1204, n1259);
xor  g1414 (n1600, n1394, n1339, n1348, n1396);
xor  g1415 (n1471, n1312, n1369, n1320, n1268);
and  g1416 (n1595, n1403, n1312, n1151, n1282);
xnor g1417 (n1430, n1269, n1282, n1358, n1352);
xnor g1418 (n1468, n1281, n1291, n1341, n1349);
nor  g1419 (n1492, n1354, n1384, n1256, n1270);
xor  g1420 (n1558, n1152, n1200, n1403, n1239);
and  g1421 (n1524, n1229, n1374, n1336, n1333);
nor  g1422 (n1474, n1376, n1304, n1299, n1251);
nand g1423 (n1528, n1358, n1371, n1269, n1391);
xnor g1424 (n1453, n1402, n1262, n1386, n1363);
and  g1425 (n1491, n1361, n1319, n1308, n1347);
nand g1426 (n1450, n1331, n1322, n1302, n1349);
nor  g1427 (n1503, n1272, n1370, n1175, n1298);
xnor g1428 (n1562, n1281, n1171, n1221, n1182);
xnor g1429 (n1423, n1399, n1354, n1343, n1191);
and  g1430 (n1573, n1316, n1300, n1266, n1311);
nand g1431 (n1537, n1257, n1348, n1261, n1360);
xnor g1432 (n1499, n1336, n1306, n1401, n1383);
nand g1433 (n1523, n1263, n1289, n1346, n1302);
nand g1434 (n1508, n1280, n1199, n1333, n1406);
xor  g1435 (n1526, n1395, n1332, n1214, n1389);
xnor g1436 (n1479, n1291, n1161, n1327, n1254);
or   g1437 (n1420, n1366, n1165, n1332, n1269);
or   g1438 (n1487, n1313, n1398, n1322, n1260);
xnor g1439 (n1585, n1330, n1254, n1377, n1392);
xnor g1440 (n1544, n1294, n1362, n1335, n1301);
nor  g1441 (n1603, n1197, n1383, n1225, n1367);
xor  g1442 (n1550, n1323, n1231, n1379, n1149);
xnor g1443 (n1572, n1216, n1370, n1380, n1361);
xor  g1444 (n1581, n1385, n1387, n1355, n125);
xnor g1445 (n1477, n1227, n1299, n1240, n1258);
and  g1446 (n1455, n1342, n1286, n1327, n1377);
nor  g1447 (n1433, n1360, n1345, n1319, n1397);
nor  g1448 (n1565, n1332, n1380, n1283, n1327);
and  g1449 (n1441, n1399, n1345, n1190, n1338);
and  g1450 (n1601, n1218, n1334, n1222, n1405);
xor  g1451 (n1584, n1329, n1235, n1398, n1181);
xor  g1452 (n1529, n1275, n1268, n1159, n1307);
or   g1453 (n1472, n1311, n1350, n1317, n1304);
xnor g1454 (n1551, n1264, n1271, n1236, n1317);
nor  g1455 (n1509, n1253, n1373, n1291, n1319);
and  g1456 (n1429, n1351, n1364, n1270, n1292);
xor  g1457 (n1594, n1327, n1237, n1400, n1404);
xnor g1458 (n1570, n1324, n1196, n1278, n1245);
xor  g1459 (n1592, n1251, n1259, n1340, n1344);
xor  g1460 (n1540, n1271, n1368, n1305, n1324);
nand g1461 (n1431, n1262, n1368, n1379, n1340);
or   g1462 (n1460, n1288, n1192, n1201, n1337);
xnor g1463 (n1434, n1275, n1257, n1346, n1301);
or   g1464 (n1462, n1348, n1266, n1250, n1290);
or   g1465 (n1543, n1313, n1407, n1234, n1187);
or   g1466 (n1599, n1244, n1367, n1212, n1368);
and  g1467 (n1556, n1250, n1232, n1407, n1335);
or   g1468 (n1451, n1355, n1312, n1160, n1406);
and  g1469 (n1459, n1243, n1357, n1312, n1203);
or   g1470 (n1510, n1309, n1179, n1303, n1178);
or   g1471 (n1415, n1355, n1352, n1373, n1297);
or   g1472 (n1446, n1390, n1405, n1287, n1334);
or   g1473 (n1440, n1250, n1305, n125, n1277);
xnor g1474 (n1596, n1375, n1396, n1406, n1255);
xnor g1475 (n1435, n1169, n1277, n124, n1359);
and  g1476 (n1475, n1369, n1259, n1256, n1329);
nor  g1477 (n1467, n1337, n1289, n1284, n1363);
xnor g1478 (n1502, n1308, n1156, n1314, n1265);
or   g1479 (n1458, n1241, n1311, n1392, n1372);
xor  g1480 (n1413, n1307, n1282, n1324, n1295);
nor  g1481 (n1447, n1302, n1374, n1364, n1370);
nor  g1482 (n1507, n1353, n1335, n1226, n1339);
or   g1483 (n1427, n1360, n1257, n1180, n1255);
or   g1484 (n1513, n1366, n1341, n1394, n1276);
or   g1485 (n1587, n1390, n1362, n1353, n1220);
nand g1486 (n1437, n1286, n1334, n1388, n1389);
nor  g1487 (n1456, n1207, n1359, n1249, n1263);
nand g1488 (n1410, n1389, n1318, n1306, n1345);
and  g1489 (n1489, n1276, n1260, n1297, n1264);
nand g1490 (n1494, n1276, n1266, n1382, n1340);
and  g1491 (n1481, n1324, n1351, n1332, n1275);
xnor g1492 (n1485, n1367, n1362, n1347, n1344);
xor  g1493 (n1443, n1279, n1306, n1315, n1309);
nor  g1494 (n1439, n1371, n1405, n1318, n1249);
nand g1495 (n1495, n1377, n1300, n1351, n1381);
nor  g1496 (n1517, n1293, n1357, n1315, n1387);
or   g1497 (n1476, n1407, n1393, n1390, n1279);
xor  g1498 (n1445, n1325, n1285, n1164, n1310);
xor  g1499 (n1530, n1285, n1258, n1353, n1287);
xnor g1500 (n1582, n1252, n1293, n1331, n1291);
nor  g1501 (n1412, n1280, n1337, n1230, n1297);
and  g1502 (n1473, n1396, n1383, n1351, n1259);
and  g1503 (n1545, n1157, n1323, n1399, n1299);
or   g1504 (n1557, n1286, n1387, n1345, n1158);
xor  g1505 (n1578, n1261, n1195, n1272, n1267);
xor  g1506 (n1535, n1315, n1385, n1395, n1282);
nand g1507 (n1577, n1398, n1281, n1288, n1331);
xnor g1508 (n1470, n1397, n1350, n1249, n1185);
xnor g1509 (n1496, n1350, n1265, n1172, n1323);
nor  g1510 (n1438, n1302, n1328, n1323, n1290);
xor  g1511 (n1486, n1379, n1354, n1295, n1333);
nor  g1512 (n1576, n1303, n1301, n1208, n1382);
or   g1513 (n1461, n1273, n1348, n1316, n1279);
xor  g1514 (n1511, n1363, n1381, n1372, n1391);
nor  g1515 (n1536, n1365, n1362, n1384, n1273);
xor  g1516 (n1602, n1276, n1403, n1289, n1385);
or   g1517 (n1580, n1274, n1385, n1250, n1392);
or   g1518 (n1463, n1253, n1299, n1340, n1310);
xnor g1519 (n1501, n1262, n1361, n1316, n1253);
nand g1520 (n1422, n1238, n1341, n1213, n1306);
xnor g1521 (n1421, n1405, n1292, n1344, n1329);
nor  g1522 (n1414, n1269, n1272, n1321, n1263);
nand g1523 (n1416, n1330, n1337, n1394, n1301);
nor  g1524 (n1598, n1305, n1252, n1382, n1356);
xnor g1525 (n1547, n1369, n1261, n1378, n1400);
nor  g1526 (n1505, n1364, n1289, n1281, n1277);
nand g1527 (n1521, n1254, n1278, n1356, n1403);
nand g1528 (n1454, n1260, n1268, n1397, n1407);
nor  g1529 (n1520, n1262, n1369, n1298, n1320);
xnor g1530 (n1493, n1366, n1202, n1248, n1294);
xnor g1531 (n1532, n1266, n1336, n1387, n1193);
nor  g1532 (n1436, n1258, n1314, n1247, n1401);
nor  g1533 (n1488, n1325, n1346, n1211, n1321);
xnor g1534 (n1518, n1406, n1402, n1359, n1366);
xor  g1535 (n1555, n1330, n1303, n1395, n1374);
or   g1536 (n1500, n1373, n1217, n1184, n1314);
or   g1537 (n1541, n1354, n1267, n1397, n1168);
or   g1538 (n1498, n1404, n1365, n1376, n1170);
xor  g1539 (n1497, n1352, n1249, n1273, n1271);
xnor g1540 (n1563, n1373, n1309, n1386, n1333);
xor  g1541 (n1579, n1370, n1357, n1254, n1308);
or   g1542 (n1568, n1277, n1347, n1380, n1189);
xnor g1543 (n1424, n1377, n1314, n1280, n1271);
xnor g1544 (n1408, n1206, n1147, n1335, n1384);
xnor g1545 (n1561, n1316, n1359, n1404, n1331);
nand g1546 (n1512, n1322, n1263, n1265, n1355);
xnor g1547 (n1590, n1205, n1350, n1356, n1388);
nor  g1548 (n1586, n1320, n1304, n1256, n1176);
xnor g1549 (n1538, n1381, n1154, n1228, n1398);
and  g1550 (n1442, n1153, n1404, n1321, n1343);
nand g1551 (n1425, n1361, n1292, n1305, n1298);
or   g1552 (n1567, n1280, n1148, n1390, n1296);
nor  g1553 (n1548, n1360, n1341, n1300, n1284);
xnor g1554 (n1569, n1401, n1288, n1349, n1295);
nor  g1555 (n1482, n1284, n1255, n1288, n1375);
nor  g1556 (n1574, n1194, n1307, n1310, n1224);
nand g1557 (n1566, n125, n1326, n1274, n1384);
and  g1558 (n1452, n1375, n1278, n1274, n1347);
xnor g1559 (n1469, n1293, n1325, n1162, n1309);
xnor g1560 (n1588, n1163, n1326, n1338, n1328);
nor  g1561 (n1449, n1326, n1308, n1400, n1258);
xnor g1562 (n1519, n1317, n1356, n1285, n1342);
or   g1563 (n1527, n1273, n1294, n1391, n1283);
or   g1564 (n1542, n1264, n1344, n1177, n1358);
or   g1565 (n1483, n1334, n1300, n1166, n125);
xnor g1566 (n1506, n1338, n1393, n1328, n1261);
nand g1567 (n1464, n1297, n1368, n1283, n1174);
xor  g1568 (n1490, n1173, n1378, n1388, n1270);
or   g1569 (n1428, n1275, n1274, n1402, n1285);
xnor g1570 (n1564, n1401, n1321, n1284, n1268);
nand g1571 (n1504, n1279, n1303, n1386, n1317);
nor  g1572 (n1747, n1580, n1049, n1064, n1460);
and  g1573 (n1888, n1130, n1534, n1474, n1447);
xor  g1574 (n1669, n1071, n1476, n1117, n1459);
or   g1575 (n1644, n1418, n1477, n1505, n1475);
or   g1576 (n1831, n1545, n1118, n1100, n1133);
nand g1577 (n1723, n1109, n1460, n1115, n1598);
xor  g1578 (n1809, n1083, n1484, n1140, n1064);
xor  g1579 (n1879, n1592, n1125, n1117, n1575);
xnor g1580 (n1765, n1115, n1496, n1146, n1133);
and  g1581 (n1890, n1064, n1107, n1577, n1530);
and  g1582 (n1778, n1411, n1579, n1546, n1501);
nand g1583 (n1627, n1499, n1065, n1446, n1464);
or   g1584 (n1608, n1581, n1106, n1527, n1104);
nor  g1585 (n1647, n1559, n1084, n1457, n1075);
xnor g1586 (n1667, n1497, n1142, n1555, n1509);
xnor g1587 (n1850, n1408, n1464, n1056, n1117);
nand g1588 (n1740, n1513, n1044, n1135, n1497);
and  g1589 (n1726, n1489, n1573, n1110, n1514);
nor  g1590 (n1804, n1492, n1519, n1106, n1433);
nand g1591 (n1771, n1486, n1057, n1562, n1415);
and  g1592 (n1691, n1541, n1504, n1078, n1587);
xnor g1593 (n1611, n1116, n1493, n1521, n1057);
or   g1594 (n1792, n1422, n1491, n1468, n1547);
or   g1595 (n1736, n1550, n1597, n1127, n1123);
nand g1596 (n1696, n1588, n1481, n1083, n1047);
or   g1597 (n1683, n1411, n1044, n1577);
xnor g1598 (n1774, n1503, n1094, n1072, n1139);
nor  g1599 (n1613, n1058, n1599, n1511, n1053);
or   g1600 (n1815, n1078, n1104, n1073, n1111);
or   g1601 (n1766, n1419, n1146, n1055, n1494);
xor  g1602 (n1654, n1067, n1506, n1047, n1138);
or   g1603 (n1655, n1561, n1083, n1086, n1545);
xor  g1604 (n1833, n1059, n1444, n1466, n1533);
nand g1605 (n1794, n1481, n1584, n1088, n1107);
nor  g1606 (n1900, n1125, n1486, n1410, n1471);
nand g1607 (n1820, n1432, n1554, n1098, n1598);
and  g1608 (n1628, n1080, n1536, n1081, n1587);
and  g1609 (n1897, n1511, n1438, n1057, n1106);
nand g1610 (n1877, n1603, n1056, n1514, n1441);
and  g1611 (n1796, n1437, n1113, n1431, n1558);
xnor g1612 (n1818, n1490, n1484, n1591, n1588);
or   g1613 (n1769, n1585, n1493, n1114, n1482);
xor  g1614 (n1868, n1119, n1579, n1054, n1503);
nand g1615 (n1618, n1101, n1426, n1467, n1412);
xnor g1616 (n1832, n1568, n1443, n1487, n1052);
nand g1617 (n1713, n1551, n1474, n1480, n1544);
or   g1618 (n1684, n1539, n1496, n1121, n1535);
or   g1619 (n1821, n1503, n1060, n1130, n1134);
xor  g1620 (n1750, n1043, n1525, n1478, n1570);
nor  g1621 (n1673, n1508, n1500, n1589, n1529);
nand g1622 (n1870, n1556, n1413, n1075, n1597);
and  g1623 (n1836, n1131, n1452, n1434, n1101);
xor  g1624 (n1869, n1524, n1061, n1431, n1108);
nor  g1625 (n1715, n1142, n1093, n1085, n1453);
xor  g1626 (n1758, n1495, n1048, n1573, n1060);
nand g1627 (n1858, n1524, n1139, n1121, n1432);
xor  g1628 (n1635, n1542, n1506, n1124, n1534);
xor  g1629 (n1805, n1466, n1460, n1141, n1454);
or   g1630 (n1704, n1574, n1597, n1097, n1441);
nand g1631 (n1826, n1063, n1114, n1045, n1437);
nand g1632 (n1674, n1419, n1459, n1087, n1045);
and  g1633 (n1636, n1140, n1479, n1532, n1546);
nand g1634 (n1883, n1121, n1567, n1070, n1145);
xnor g1635 (n1884, n1505, n1512, n1116, n1530);
nand g1636 (n1873, n1552, n1063, n1553, n1067);
nor  g1637 (n1645, n1078, n1058, n1423, n1046);
nor  g1638 (n1642, n1446, n1092, n1484, n1491);
nor  g1639 (n1903, n1570, n1073, n1459, n1072);
nor  g1640 (n1775, n1427, n1065, n1098, n1455);
and  g1641 (n1767, n1451, n1453, n1146, n1493);
xnor g1642 (n1755, n1472, n1461, n1507, n1565);
xor  g1643 (n1901, n1595, n1089, n1117, n1502);
nand g1644 (n1632, n1479, n1561, n1527, n1430);
and  g1645 (n1716, n1048, n1072, n1067, n1085);
nor  g1646 (n1898, n1602, n1574, n1426, n1095);
xnor g1647 (n1663, n1563, n1061, n1458, n1126);
and  g1648 (n1799, n1116, n1532, n1572, n1482);
nor  g1649 (n1714, n1100, n1464, n1091, n1442);
xor  g1650 (n1902, n1092, n1466, n1128, n1453);
and  g1651 (n1670, n1138, n1123, n1596, n1044);
nand g1652 (n1759, n1535, n1143, n1046, n1090);
and  g1653 (n1822, n1542, n1565, n1097, n1074);
and  g1654 (n1641, n1548, n1518, n1603, n1496);
xor  g1655 (n1841, n1416, n1579, n1050, n1548);
or   g1656 (n1834, n1079, n1474, n1602, n1488);
xnor g1657 (n1709, n1422, n1412, n1568, n1068);
or   g1658 (n1702, n1575, n1448, n1492, n1510);
or   g1659 (n1745, n1595, n1526, n1518, n1449);
nand g1660 (n1904, n1052, n1518, n1504, n1120);
nor  g1661 (n1609, n1578, n1045, n1546, n1139);
xor  g1662 (n1708, n1051, n1058, n1563, n1517);
xor  g1663 (n1886, n1068, n1069, n1473, n1483);
xor  g1664 (n1606, n1080, n1469, n1425, n1087);
and  g1665 (n1612, n1542, n1537, n1525, n1430);
xnor g1666 (n1875, n1485, n1430, n1082, n1474);
or   g1667 (n1707, n1128, n1110, n1099, n1063);
or   g1668 (n1893, n1484, n1126, n1598, n1143);
nor  g1669 (n1827, n1584, n1508, n1415, n1554);
and  g1670 (n1777, n1422, n1598, n1463, n1424);
and  g1671 (n1692, n1447, n1590, n1540, n1134);
or   g1672 (n1867, n1429, n1409, n1445, n1071);
nor  g1673 (n1681, n1565, n1567, n1113, n1475);
xor  g1674 (n1800, n1597, n1458, n1094, n1539);
nor  g1675 (n1881, n1594, n1548, n1557, n1497);
xnor g1676 (n1737, n1550, n1549, n1070, n1063);
and  g1677 (n1677, n1580, n1521, n1103, n1444);
xnor g1678 (n1637, n1532, n1421, n1139, n1497);
and  g1679 (n1811, n1577, n1573, n1583, n1439);
nor  g1680 (n1729, n1544, n1434, n1593, n1425);
nor  g1681 (n1835, n1414, n1545, n1556, n1074);
or   g1682 (n1712, n1076, n1558, n1131, n1498);
nand g1683 (n1720, n1098, n1055, n1062, n1604);
nor  g1684 (n1754, n1115, n1076, n1425, n1415);
nand g1685 (n1852, n1549, n1437, n1519, n1052);
nand g1686 (n1807, n1567, n1512, n1436, n1600);
xnor g1687 (n1722, n1448, n1430, n1128, n1575);
xnor g1688 (n1651, n1480, n1090, n1112, n1512);
and  g1689 (n1843, n1508, n1455, n1119, n1538);
nand g1690 (n1741, n1458, n1568, n1470, n1560);
nand g1691 (n1752, n1429, n1059, n1127, n1091);
nand g1692 (n1662, n1472, n1581, n1531, n1127);
or   g1693 (n1810, n1141, n1457, n1575, n1520);
xnor g1694 (n1738, n1109, n1595, n1136);
xnor g1695 (n1860, n1554, n1550, n1130, n1109);
and  g1696 (n1838, n1588, n1543, n1553, n1526);
and  g1697 (n1788, n1126, n1448, n1527, n1461);
or   g1698 (n1676, n1135, n1488, n1433, n1594);
and  g1699 (n1744, n1080, n1435, n1581, n1538);
xnor g1700 (n1871, n1428, n1438, n1113, n1498);
xnor g1701 (n1790, n1523, n1513, n1518, n1463);
nor  g1702 (n1685, n1433, n1140, n1102, n1077);
xnor g1703 (n1607, n1089, n1492, n1467, n1599);
and  g1704 (n1625, n1554, n1112, n1471, n1133);
xor  g1705 (n1679, n1081, n1465, n1118, n1576);
xnor g1706 (n1630, n1409, n1134, n1539, n1090);
nand g1707 (n1801, n1476, n1138, n1523, n1502);
and  g1708 (n1862, n1461, n1489, n1129);
nand g1709 (n1751, n1419, n1053, n1132, n1075);
nor  g1710 (n1814, n1557, n1418, n1102, n1071);
and  g1711 (n1703, n1444, n1463, n1555, n1526);
xor  g1712 (n1837, n1466, n1070, n1410, n1132);
and  g1713 (n1847, n1424, n1467, n1091, n1076);
xnor g1714 (n1816, n1569, n1534, n1048, n1124);
xor  g1715 (n1733, n1540, n1100, n1462, n1110);
xnor g1716 (n1665, n1439, n1462, n1599, n1074);
or   g1717 (n1885, n1496, n1418, n1085, n1062);
and  g1718 (n1895, n1120, n1535, n1106, n1483);
or   g1719 (n1797, n1584, n1414, n1469, n1595);
nand g1720 (n1761, n1099, n1488, n1069, n1543);
and  g1721 (n1840, n1427, n1088, n1594, n1093);
and  g1722 (n1659, n1439, n1578, n1478, n1592);
and  g1723 (n1773, n1438, n1452, n1506, n1462);
xor  g1724 (n1633, n1513, n1053, n1082, n1583);
and  g1725 (n1671, n1585, n1048, n1137, n1094);
nor  g1726 (n1846, n1068, n1141, n1101, n1600);
nand g1727 (n1661, n1451, n1480, n1129, n1504);
xnor g1728 (n1764, n1082, n1440, n1428, n1105);
or   g1729 (n1664, n1449, n1445, n1077, n1521);
and  g1730 (n1855, n1470, n1446, n1487, n1435);
nor  g1731 (n1798, n1093, n1529, n1560, n1095);
nand g1732 (n1782, n1092, n1508, n1543, n1080);
and  g1733 (n1763, n1543, n1145, n1436, n1105);
nor  g1734 (n1734, n1525, n1050, n1566, n1533);
nand g1735 (n1678, n1423, n1481, n1498, n1046);
nor  g1736 (n1813, n1552, n1490, n1507, n1563);
nand g1737 (n1779, n1412, n1552, n1528);
nor  g1738 (n1682, n1585, n1524, n1483, n1600);
nand g1739 (n1689, n1105, n1571, n1565, n1564);
and  g1740 (n1694, n1084, n1136, n1437, n1600);
or   g1741 (n1863, n1506, n1601, n1564, n1066);
nand g1742 (n1719, n1544, n1515, n1146, n1440);
xnor g1743 (n1762, n1432, n1576, n1079, n1448);
nand g1744 (n1894, n1529, n1569, n1509, n1469);
or   g1745 (n1851, n1411, n1586, n1502, n1559);
or   g1746 (n1780, n1441, n1572, n1468, n1585);
nor  g1747 (n1878, n1135, n1072, n1604, n1418);
or   g1748 (n1739, n1593, n1586, n1594, n1051);
xor  g1749 (n1768, n1482, n1477, n1529, n1571);
or   g1750 (n1786, n1109, n1140, n1059, n1097);
or   g1751 (n1639, n1551, n1047, n1096, n1534);
xnor g1752 (n1817, n1530, n1054, n1059, n1451);
xnor g1753 (n1638, n1570, n1443, n1054, n1586);
xor  g1754 (n1849, n1549, n1564, n1125, n1416);
xor  g1755 (n1823, n1046, n1571, n1431, n1490);
nor  g1756 (n1892, n1111, n1131, n1522, n1473);
nor  g1757 (n1785, n1458, n1533, n1103, n1453);
xor  g1758 (n1643, n1083, n1411, n1503, n1089);
and  g1759 (n1666, n1467, n1105, n1100, n1442);
nand g1760 (n1728, n1409, n1516, n1462, n1572);
or   g1761 (n1622, n1494, n1425, n1132, n1584);
xnor g1762 (n1705, n1052, n1491, n1509, n1515);
nor  g1763 (n1760, n1452, n1429, n1082, n1541);
nand g1764 (n1830, n1535, n1439, n1112, n1424);
or   g1765 (n1657, n1464, n1519, n1553, n1094);
xor  g1766 (n1887, n1516, n1580, n1120, n1138);
and  g1767 (n1857, n1049, n1461, n1412, n1095);
or   g1768 (n1889, n1102, n1525, n1050, n1476);
nor  g1769 (n1652, n1524, n1469, n1051, n1447);
nand g1770 (n1808, n1522, n1500, n1056, n1108);
or   g1771 (n1710, n1520, n1433, n1478, n1429);
xor  g1772 (n1649, n1583, n1564, n1573, n1099);
or   g1773 (n1748, n1454, n1570, n1088, n1044);
or   g1774 (n1853, n1522, n1528, n1426, n1108);
xor  g1775 (n1789, n1487, n1485, n1576, n1549);
xor  g1776 (n1776, n1125, n1420, n1428, n1590);
nor  g1777 (n1791, n1486, n1556, n1417, n1582);
or   g1778 (n1730, n1587, n1057, n1592, n1542);
nand g1779 (n1653, n1546, n1533, n1131, n1091);
nand g1780 (n1687, n1592, n1421, n1110, n1416);
nor  g1781 (n1718, n1431, n1101, n1589, n1055);
and  g1782 (n1802, n1054, n1551, n1471, n1489);
nand g1783 (n1859, n1456, n1126, n1133, n1134);
xnor g1784 (n1819, n1114, n1122, n1561, n1479);
and  g1785 (n1880, n1591, n1143, n1574, n1435);
nand g1786 (n1727, n1050, n1531, n1555, n1485);
nand g1787 (n1700, n1413, n1562, n1589, n1127);
nand g1788 (n1806, n1540, n1571, n1096, n1113);
nor  g1789 (n1680, n1144, n1123, n1507, n1536);
nor  g1790 (n1848, n1123, n1058, n1450, n1587);
nor  g1791 (n1787, n1142, n1493, n1443, n1531);
or   g1792 (n1619, n1065, n1049, n1520, n1547);
or   g1793 (n1839, n1450, n1445, n1410, n1588);
nor  g1794 (n1614, n1098, n1604, n1075, n1500);
nand g1795 (n1845, n1558, n1129, n1513, n1413);
xor  g1796 (n1675, n1119, n1460, n1510, n1122);
xnor g1797 (n1784, n1465, n1053, n1515, n1562);
nand g1798 (n1724, n1536, n1144, n1066, n1578);
and  g1799 (n1783, n1599, n1559, n1563, n1096);
nand g1800 (n1620, n1591, n1145, n1555, n1086);
and  g1801 (n1795, n1071, n1086, n1528, n1423);
nand g1802 (n1781, n1512, n1499, n1043, n1445);
xor  g1803 (n1640, n1089, n1509, n1558, n1122);
xnor g1804 (n1693, n1079, n1556, n1421, n1077);
or   g1805 (n1731, n1586, n1130, n1062, n1591);
or   g1806 (n1742, n1472, n1104, n1471, n1135);
xor  g1807 (n1856, n1602, n1081, n1114, n1073);
nor  g1808 (n1757, n1442, n1103, n1455, n1498);
xnor g1809 (n1646, n1421, n1517, n1087, n1520);
and  g1810 (n1725, n1120, n1523, n1420, n1501);
nand g1811 (n1634, n1473, n1087, n1490, n1593);
or   g1812 (n1899, n1511, n1414, n1456, n1424);
xor  g1813 (n1803, n1590, n1468, n1581, n1507);
or   g1814 (n1866, n1081, n1436, n1116, n1486);
nand g1815 (n1624, n1073, n1444, n1567, n1510);
or   g1816 (n1864, n1435, n1530, n1061, n1449);
xnor g1817 (n1743, n1066, n1574, n1085, n1428);
xnor g1818 (n1610, n1060, n1092, n1069, n1077);
nor  g1819 (n1882, n1128, n1045, n1548, n1078);
and  g1820 (n1824, n1532, n1560, n1065, n1468);
and  g1821 (n1844, n1526, n1068, n1076, n1562);
nor  g1822 (n1829, n1521, n1099, n1601, n1423);
and  g1823 (n1825, n1495, n1118, n1516, n1455);
or   g1824 (n1842, n1505, n1410, n1463, n1136);
and  g1825 (n1699, n1132, n1141, n1569, n1137);
and  g1826 (n1717, n1434, n1145, n1580, n1523);
xnor g1827 (n1701, n1446, n1115, n1495, n1043);
xor  g1828 (n1672, n1495, n1596, n1578, n1511);
xor  g1829 (n1656, n1475, n1451, n1589, n1566);
or   g1830 (n1812, n1539, n1596, n1502, n1527);
xnor g1831 (n1648, n1544, n1420, n1480, n1545);
xnor g1832 (n1621, n1124, n1477, n1067, n1522);
and  g1833 (n1706, n1441, n1501, n1470, n1541);
nor  g1834 (n1650, n1449, n1436, n1062, n1144);
xor  g1835 (n1735, n1440, n1472, n1432, n1079);
xnor g1836 (n1861, n1553, n1447, n1066, n1557);
nand g1837 (n1854, n1452, n1500, n1454, n1601);
nand g1838 (n1658, n1124, n1074, n1568, n1514);
nor  g1839 (n1690, n1505, n1603, n1583, n1536);
or   g1840 (n1631, n1541, n1415, n1602, n1061);
or   g1841 (n1711, n1137, n1119, n1102, n1604);
nor  g1842 (n1746, n1475, n1488, n1442, n1047);
or   g1843 (n1626, n1084, n1064, n1104, n1510);
or   g1844 (n1891, n1481, n1538, n1528, n1470);
xnor g1845 (n1697, n1582, n1056, n1491, n1579);
or   g1846 (n1695, n1576, n1515, n1551, n1434);
nand g1847 (n1896, n1070, n1582, n1483, n1409);
xor  g1848 (n1660, n1427, n1118, n1450, n1414);
xor  g1849 (n1872, n1069, n1122, n1097, n1422);
nand g1850 (n1698, n1454, n1137, n1465, n1538);
and  g1851 (n1688, n1093, n1473, n1111, n1489);
nand g1852 (n1770, n1440, n1499, n1417, n1593);
nor  g1853 (n1721, n1557, n1547, n1112, n1090);
and  g1854 (n1865, n1456, n1590, n1107, n1413);
and  g1855 (n1732, n1596, n1049, n1479, n1142);
or   g1856 (n1615, n1121, n1560, n1540, n1517);
or   g1857 (n1686, n1566, n1514, n1516, n1519);
xnor g1858 (n1629, n1499, n1456, n1485, n1419);
xnor g1859 (n1753, n1550, n1443, n1084, n1477);
nor  g1860 (n1756, n1095, n1111, n1603, n1572);
xnor g1861 (n1617, n1547, n1478, n1537);
nor  g1862 (n1793, n1427, n1144, n1457, n1417);
nand g1863 (n1668, n1060, n1501, n1108, n1107);
or   g1864 (n1772, n1096, n1494, n1531, n1420);
xnor g1865 (n1874, n1569, n1582, n1465, n1055);
and  g1866 (n1828, n1459, n1426, n1601, n1517);
xnor g1867 (n1623, n1103, n1487, n1051, n1416);
xnor g1868 (n1616, n1504, n1494, n1417, n1086);
or   g1869 (n1749, n1559, n1566, n1457, n1537);
xnor g1870 (n1876, n1492, n1476, n1450, n1438);
nand g1871 (n1605, n1482, n1143, n1088, n1561);
xnor g1872 (n1985, n1757, n93, n1846, n159);
xor  g1873 (n1955, n1725, n1608, n1652, n1623);
nor  g1874 (n1987, n1830, n1792, n1716, n1682);
nand g1875 (n1984, n1699, n89, n93, n1849);
and  g1876 (n1960, n1615, n89, n1895, n1782);
xor  g1877 (n1905, n1727, n86, n1728, n1872);
nor  g1878 (n1916, n1638, n1804, n1651, n1660);
or   g1879 (n1953, n1676, n1761, n1625, n1663);
xnor g1880 (n1991, n1859, n1862, n92, n85);
nor  g1881 (n1946, n1719, n1882, n1669, n1711);
nand g1882 (n1911, n1824, n158, n86, n1702);
nand g1883 (n1925, n1794, n1730, n1735, n1693);
nor  g1884 (n1920, n1802, n1861, n1871, n1640);
nand g1885 (n1976, n1636, n1818, n157, n1783);
xor  g1886 (n1928, n1705, n93, n1808, n1677);
nor  g1887 (n1922, n1626, n88, n1826, n1856);
or   g1888 (n1977, n1724, n1875, n1646, n158);
or   g1889 (n1941, n1722, n1629, n1686, n1888);
xnor g1890 (n1993, n1854, n90, n1762, n1864);
and  g1891 (n1927, n1723, n1837, n1746, n1763);
and  g1892 (n1921, n1805, n1812, n91, n1834);
or   g1893 (n1950, n1685, n1879, n1795, n1852);
nand g1894 (n1972, n95, n1815, n1821, n1656);
xor  g1895 (n1978, n1809, n1659, n92, n1827);
or   g1896 (n1945, n1680, n1825, n1667, n1700);
xor  g1897 (n1923, n1624, n1733, n92, n1901);
xor  g1898 (n1961, n91, n1840, n1870, n1644);
nand g1899 (n1967, n1744, n1793, n1609, n1787);
and  g1900 (n1981, n89, n1694, n1807, n1833);
or   g1901 (n1964, n1838, n1679, n1769, n1813);
and  g1902 (n1936, n1823, n1828, n1880, n87);
nand g1903 (n1932, n90, n1731, n1616, n1892);
and  g1904 (n1958, n1732, n1890, n1622, n89);
nor  g1905 (n1908, n1832, n1621, n156, n1780);
xor  g1906 (n1929, n1695, n1884, n87, n1745);
nand g1907 (n1940, n1642, n1766, n95, n94);
or   g1908 (n1919, n1771, n1803, n1647, n1635);
or   g1909 (n1975, n1627, n1868, n92, n1831);
nand g1910 (n1980, n1631, n1639, n1721, n158);
and  g1911 (n1912, n1684, n1697, n1689, n1633);
xor  g1912 (n1944, n1810, n1877, n1666, n1873);
and  g1913 (n1971, n1798, n1632, n1747, n157);
xor  g1914 (n1966, n1754, n1740, n1714, n91);
and  g1915 (n1938, n1738, n1777, n1878, n1898);
nor  g1916 (n1963, n1710, n1696, n88, n1836);
or   g1917 (n1933, n1775, n1881, n1752, n1726);
or   g1918 (n1906, n1790, n1772, n1641, n228);
xor  g1919 (n1942, n91, n1749, n95, n1767);
xor  g1920 (n1917, n1897, n1683, n1791, n1800);
xor  g1921 (n1943, n88, n1774, n1876, n1743);
nor  g1922 (n1986, n1789, n1606, n1896, n1703);
nor  g1923 (n1915, n1670, n1649, n1902, n1886);
or   g1924 (n1935, n1799, n1891, n1894, n1681);
nor  g1925 (n1930, n1753, n1887, n1712, n1779);
or   g1926 (n1952, n1674, n86, n1758, n1842);
xnor g1927 (n1918, n90, n1869, n1867, n158);
xnor g1928 (n1934, n1701, n1778, n1657, n1729);
nand g1929 (n1947, n1816, n1691, n1841, n1707);
and  g1930 (n1957, n156, n159, n1687, n94);
and  g1931 (n1956, n93, n1607, n1610, n1672);
xor  g1932 (n1965, n1675, n1819, n1844, n1634);
nand g1933 (n1924, n1850, n157, n1643, n1858);
xor  g1934 (n1982, n1756, n1661, n94, n1688);
and  g1935 (n1968, n1889, n1765, n1734, n1899);
xor  g1936 (n1970, n1664, n1611, n88, n1900);
xor  g1937 (n1937, n1855, n1776, n1773, n1717);
xnor g1938 (n1926, n1742, n1648, n1863, n87);
and  g1939 (n1959, n1617, n1806, n1755, n1851);
nor  g1940 (n1992, n1883, n1709, n1650, n1704);
or   g1941 (n1909, n1768, n1665, n1801, n1796);
xnor g1942 (n1983, n1885, n1866, n1718, n1839);
or   g1943 (n1969, n1865, n1853, n1829, n1655);
or   g1944 (n1939, n1630, n1658, n1620, n1857);
xor  g1945 (n1910, n1822, n1760, n1784, n1848);
nand g1946 (n1914, n1788, n1811, n159, n1720);
or   g1947 (n1974, n95, n1706, n1673, n1637);
nand g1948 (n1949, n1713, n1843, n1698, n1736);
nand g1949 (n1913, n1662, n1860, n94, n1619);
nor  g1950 (n1962, n1613, n1814, n1618, n1605);
nor  g1951 (n1989, n1671, n1692, n1750, n1786);
nor  g1952 (n1931, n1614, n1653, n228, n1785);
nand g1953 (n1954, n1668, n1764, n1845, n1741);
or   g1954 (n1973, n159, n1739, n1612, n1654);
nor  g1955 (n1951, n1748, n1715, n1628, n1645);
or   g1956 (n1979, n86, n1835, n1759, n90);
or   g1957 (n1988, n1781, n1817, n157, n87);
nand g1958 (n1948, n1737, n156, n1874, n1797);
or   g1959 (n1990, n1893, n1678, n1708, n1847);
nand g1960 (n1907, n1751, n1690, n1820, n1770);
nor  g1961 (n2007, n1914, n1925, n1973, n1934);
xnor g1962 (n1994, n1956, n1905, n1970, n1982);
nor  g1963 (n2002, n1975, n1968, n1992, n1918);
and  g1964 (n2015, n1957, n1923, n1985, n1976);
nor  g1965 (n2006, n1962, n1915, n1912, n1966);
nor  g1966 (n2013, n1961, n1958, n1941, n1944);
xnor g1967 (n1995, n1949, n1964, n1929, n1917);
or   g1968 (n1998, n1971, n1955, n1935, n1928);
xnor g1969 (n2005, n1940, n1927, n1959, n1951);
xnor g1970 (n1997, n1978, n1943, n1986, n1952);
xnor g1971 (n2008, n1933, n1919, n1990, n1922);
nand g1972 (n2012, n1920, n1967, n1983, n1981);
or   g1973 (n2001, n1907, n1991, n1926, n1924);
nor  g1974 (n1999, n1987, n1909, n1977, n1947);
nor  g1975 (n2000, n1936, n1979, n1938, n1974);
or   g1976 (n2010, n1916, n1969, n1930, n1931);
nor  g1977 (n1996, n1913, n1953, n1932, n1946);
or   g1978 (n2004, n1980, n1988, n1910, n1942);
or   g1979 (n2011, n1963, n1950, n1954, n1908);
xor  g1980 (n2014, n1960, n1989, n1972, n1911);
and  g1981 (n2009, n1945, n1984, n1965, n1939);
and  g1982 (n2003, n1921, n1937, n1948, n1906);
not  g1983 (n2029, n2007);
not  g1984 (n2017, n2005);
buf  g1985 (n2025, n1998);
buf  g1986 (n2030, n1904);
not  g1987 (n2022, n1993);
buf  g1988 (n2027, n2003);
buf  g1989 (n2021, n2014);
not  g1990 (n2024, n2012);
not  g1991 (n2026, n2009);
buf  g1992 (n2020, n2006);
buf  g1993 (n2018, n2010);
not  g1994 (n2031, n1903);
not  g1995 (n2019, n2001);
not  g1996 (n2016, n2000);
buf  g1997 (n2028, n2013);
or   g1998 (n2032, n2011, n2015, n2004);
xor  g1999 (n2023, n2002, n2008, n1999, n1997);
endmodule
