

module Stat_2000_221
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1108,
  n1157,
  n1049,
  n1098,
  n1061,
  n1134,
  n1128,
  n1082,
  n1147,
  n1051,
  n1107,
  n1060,
  n1144,
  n1085,
  n1057,
  n1130,
  n1897,
  n1900,
  n2029,
  n2023,
  n2022,
  n2027,
  n2024,
  n2020,
  n2032,
  n2026,
  n2030,
  n2021,
  n2025,
  n2028,
  n2019,
  n2031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1108;output n1157;output n1049;output n1098;output n1061;output n1134;output n1128;output n1082;output n1147;output n1051;output n1107;output n1060;output n1144;output n1085;output n1057;output n1130;output n1897;output n1900;output n2029;output n2023;output n2022;output n2027;output n2024;output n2020;output n2032;output n2026;output n2030;output n2021;output n2025;output n2028;output n2019;output n2031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1050;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1058;wire n1059;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1083;wire n1084;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1129;wire n1131;wire n1132;wire n1133;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1145;wire n1146;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1898;wire n1899;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n70,
    n1
  );


  not
  g1
  (
    n46,
    n2
  );


  buf
  g2
  (
    n36,
    n26
  );


  buf
  g3
  (
    n154,
    n8
  );


  buf
  g4
  (
    n71,
    n28
  );


  buf
  g5
  (
    n34,
    n6
  );


  buf
  g6
  (
    n79,
    n8
  );


  not
  g7
  (
    n73,
    n29
  );


  not
  g8
  (
    n148,
    n23
  );


  buf
  g9
  (
    n142,
    n2
  );


  not
  g10
  (
    n44,
    n18
  );


  not
  g11
  (
    n85,
    n30
  );


  not
  g12
  (
    n65,
    n10
  );


  buf
  g13
  (
    n54,
    n22
  );


  buf
  g14
  (
    n156,
    n3
  );


  buf
  g15
  (
    n120,
    n19
  );


  buf
  g16
  (
    n151,
    n28
  );


  buf
  g17
  (
    n136,
    n5
  );


  not
  g18
  (
    n72,
    n26
  );


  not
  g19
  (
    n134,
    n29
  );


  not
  g20
  (
    n75,
    n28
  );


  not
  g21
  (
    n60,
    n1
  );


  not
  g22
  (
    n96,
    n2
  );


  buf
  g23
  (
    n121,
    n20
  );


  not
  g24
  (
    n41,
    n23
  );


  buf
  g25
  (
    n39,
    n11
  );


  buf
  g26
  (
    n78,
    n15
  );


  buf
  g27
  (
    n145,
    n30
  );


  not
  g28
  (
    n100,
    n11
  );


  buf
  g29
  (
    n115,
    n5
  );


  buf
  g30
  (
    n95,
    n7
  );


  buf
  g31
  (
    n66,
    n22
  );


  buf
  g32
  (
    n111,
    n5
  );


  buf
  g33
  (
    n118,
    n30
  );


  not
  g34
  (
    n74,
    n6
  );


  not
  g35
  (
    n90,
    n10
  );


  not
  g36
  (
    n119,
    n23
  );


  not
  g37
  (
    n124,
    n18
  );


  buf
  g38
  (
    n102,
    n19
  );


  not
  g39
  (
    n52,
    n13
  );


  not
  g40
  (
    n155,
    n10
  );


  not
  g41
  (
    n82,
    n27
  );


  buf
  g42
  (
    n101,
    n27
  );


  not
  g43
  (
    n125,
    n29
  );


  buf
  g44
  (
    n35,
    n17
  );


  not
  g45
  (
    n67,
    n9
  );


  not
  g46
  (
    n103,
    n4
  );


  not
  g47
  (
    n81,
    n5
  );


  buf
  g48
  (
    n114,
    n26
  );


  buf
  g49
  (
    n135,
    n9
  );


  not
  g50
  (
    n117,
    n4
  );


  not
  g51
  (
    n131,
    n29
  );


  not
  g52
  (
    n69,
    n26
  );


  not
  g53
  (
    n51,
    n24
  );


  buf
  g54
  (
    n86,
    n21
  );


  not
  g55
  (
    n133,
    n9
  );


  not
  g56
  (
    n53,
    n30
  );


  buf
  g57
  (
    n129,
    n12
  );


  buf
  g58
  (
    n62,
    n27
  );


  buf
  g59
  (
    n139,
    n1
  );


  not
  g60
  (
    n76,
    n16
  );


  buf
  g61
  (
    n150,
    n22
  );


  not
  g62
  (
    n61,
    n19
  );


  buf
  g63
  (
    n109,
    n12
  );


  not
  g64
  (
    n108,
    n14
  );


  not
  g65
  (
    n38,
    n6
  );


  not
  g66
  (
    n126,
    n3
  );


  not
  g67
  (
    n116,
    n22
  );


  not
  g68
  (
    n57,
    n27
  );


  buf
  g69
  (
    n50,
    n31
  );


  buf
  g70
  (
    n144,
    n20
  );


  buf
  g71
  (
    n37,
    n4
  );


  not
  g72
  (
    n48,
    n15
  );


  buf
  g73
  (
    n138,
    n16
  );


  not
  g74
  (
    n104,
    n13
  );


  not
  g75
  (
    n113,
    n25
  );


  not
  g76
  (
    n137,
    n25
  );


  buf
  g77
  (
    n128,
    n28
  );


  not
  g78
  (
    n105,
    n21
  );


  not
  g79
  (
    n80,
    n11
  );


  not
  g80
  (
    n123,
    n21
  );


  buf
  g81
  (
    n149,
    n31
  );


  not
  g82
  (
    n141,
    n31
  );


  not
  g83
  (
    n40,
    n10
  );


  buf
  g84
  (
    n63,
    n7
  );


  buf
  g85
  (
    n146,
    n18
  );


  buf
  g86
  (
    n127,
    n24
  );


  buf
  g87
  (
    n58,
    n19
  );


  not
  g88
  (
    n92,
    n6
  );


  buf
  g89
  (
    n45,
    n8
  );


  not
  g90
  (
    n107,
    n4
  );


  not
  g91
  (
    n49,
    n7
  );


  not
  g92
  (
    n106,
    n14
  );


  not
  g93
  (
    n153,
    n14
  );


  buf
  g94
  (
    n42,
    n25
  );


  buf
  g95
  (
    n43,
    n15
  );


  not
  g96
  (
    n77,
    n16
  );


  buf
  g97
  (
    n152,
    n2
  );


  not
  g98
  (
    n68,
    n18
  );


  not
  g99
  (
    n55,
    n17
  );


  not
  g100
  (
    n98,
    n20
  );


  buf
  g101
  (
    n83,
    n3
  );


  not
  g102
  (
    n94,
    n24
  );


  not
  g103
  (
    n110,
    n25
  );


  not
  g104
  (
    n99,
    n15
  );


  not
  g105
  (
    n130,
    n24
  );


  buf
  g106
  (
    n97,
    n12
  );


  buf
  g107
  (
    n122,
    n17
  );


  not
  g108
  (
    n132,
    n7
  );


  not
  g109
  (
    n91,
    n20
  );


  not
  g110
  (
    n47,
    n17
  );


  buf
  g111
  (
    n87,
    n21
  );


  not
  g112
  (
    n59,
    n8
  );


  buf
  g113
  (
    n93,
    n11
  );


  not
  g114
  (
    n56,
    n1
  );


  not
  g115
  (
    n88,
    n9
  );


  buf
  g116
  (
    n33,
    n12
  );


  buf
  g117
  (
    n64,
    n14
  );


  not
  g118
  (
    n147,
    n13
  );


  buf
  g119
  (
    n143,
    n23
  );


  not
  g120
  (
    n84,
    n31
  );


  not
  g121
  (
    n89,
    n16
  );


  buf
  g122
  (
    n140,
    n3
  );


  buf
  g123
  (
    n112,
    n13
  );


  buf
  g124
  (
    n181,
    n55
  );


  buf
  g125
  (
    n244,
    n59
  );


  buf
  g126
  (
    n161,
    n55
  );


  not
  g127
  (
    n388,
    n48
  );


  not
  g128
  (
    n280,
    n96
  );


  not
  g129
  (
    n376,
    n120
  );


  not
  g130
  (
    n507,
    n91
  );


  not
  g131
  (
    n534,
    n138
  );


  not
  g132
  (
    n583,
    n89
  );


  buf
  g133
  (
    n229,
    n107
  );


  not
  g134
  (
    n333,
    n51
  );


  not
  g135
  (
    n396,
    n130
  );


  not
  g136
  (
    n238,
    n60
  );


  not
  g137
  (
    n362,
    n72
  );


  not
  g138
  (
    n423,
    n140
  );


  not
  g139
  (
    n286,
    n100
  );


  not
  g140
  (
    n432,
    n37
  );


  buf
  g141
  (
    n468,
    n119
  );


  not
  g142
  (
    n446,
    n120
  );


  buf
  g143
  (
    n518,
    n78
  );


  not
  g144
  (
    n546,
    n46
  );


  buf
  g145
  (
    n278,
    n117
  );


  not
  g146
  (
    n565,
    n82
  );


  not
  g147
  (
    n542,
    n58
  );


  buf
  g148
  (
    n259,
    n99
  );


  buf
  g149
  (
    n459,
    n81
  );


  not
  g150
  (
    n581,
    n41
  );


  not
  g151
  (
    n342,
    n143
  );


  buf
  g152
  (
    n308,
    n133
  );


  not
  g153
  (
    n266,
    n147
  );


  buf
  g154
  (
    n326,
    n126
  );


  not
  g155
  (
    n558,
    n123
  );


  buf
  g156
  (
    n486,
    n102
  );


  buf
  g157
  (
    n568,
    n46
  );


  not
  g158
  (
    n281,
    n39
  );


  not
  g159
  (
    n576,
    n73
  );


  buf
  g160
  (
    n292,
    n77
  );


  not
  g161
  (
    n344,
    n150
  );


  not
  g162
  (
    n582,
    n71
  );


  not
  g163
  (
    n587,
    n140
  );


  buf
  g164
  (
    n254,
    n154
  );


  not
  g165
  (
    n214,
    n85
  );


  not
  g166
  (
    n276,
    n87
  );


  buf
  g167
  (
    n537,
    n95
  );


  buf
  g168
  (
    n305,
    n113
  );


  buf
  g169
  (
    n195,
    n152
  );


  not
  g170
  (
    n465,
    n42
  );


  buf
  g171
  (
    n427,
    n98
  );


  buf
  g172
  (
    n221,
    n102
  );


  buf
  g173
  (
    n398,
    n95
  );


  not
  g174
  (
    n393,
    n98
  );


  not
  g175
  (
    n458,
    n138
  );


  not
  g176
  (
    n517,
    n133
  );


  not
  g177
  (
    n401,
    n69
  );


  buf
  g178
  (
    n457,
    n62
  );


  buf
  g179
  (
    n339,
    n127
  );


  buf
  g180
  (
    n334,
    n66
  );


  not
  g181
  (
    n520,
    n149
  );


  not
  g182
  (
    n416,
    n141
  );


  buf
  g183
  (
    n338,
    n108
  );


  not
  g184
  (
    n544,
    n149
  );


  not
  g185
  (
    n588,
    n65
  );


  buf
  g186
  (
    n570,
    n62
  );


  not
  g187
  (
    n476,
    n114
  );


  buf
  g188
  (
    n370,
    n126
  );


  buf
  g189
  (
    n538,
    n131
  );


  buf
  g190
  (
    n553,
    n119
  );


  not
  g191
  (
    n348,
    n120
  );


  not
  g192
  (
    n400,
    n89
  );


  not
  g193
  (
    n352,
    n64
  );


  not
  g194
  (
    n212,
    n128
  );


  buf
  g195
  (
    n464,
    n34
  );


  buf
  g196
  (
    n523,
    n148
  );


  not
  g197
  (
    n360,
    n123
  );


  buf
  g198
  (
    n371,
    n112
  );


  not
  g199
  (
    n477,
    n105
  );


  not
  g200
  (
    n321,
    n137
  );


  not
  g201
  (
    n443,
    n121
  );


  not
  g202
  (
    n269,
    n139
  );


  not
  g203
  (
    n482,
    n109
  );


  not
  g204
  (
    n366,
    n92
  );


  not
  g205
  (
    n384,
    n72
  );


  not
  g206
  (
    n220,
    n56
  );


  buf
  g207
  (
    n255,
    n54
  );


  buf
  g208
  (
    n365,
    n33
  );


  not
  g209
  (
    n447,
    n127
  );


  buf
  g210
  (
    n347,
    n110
  );


  buf
  g211
  (
    n375,
    n88
  );


  not
  g212
  (
    n425,
    n101
  );


  buf
  g213
  (
    n324,
    n101
  );


  buf
  g214
  (
    n232,
    n49
  );


  buf
  g215
  (
    n336,
    n128
  );


  buf
  g216
  (
    n179,
    n154
  );


  not
  g217
  (
    n218,
    n64
  );


  not
  g218
  (
    n580,
    n37
  );


  buf
  g219
  (
    n584,
    n98
  );


  not
  g220
  (
    n204,
    n36
  );


  buf
  g221
  (
    n411,
    n125
  );


  not
  g222
  (
    n472,
    n134
  );


  not
  g223
  (
    n250,
    n43
  );


  buf
  g224
  (
    n562,
    n144
  );


  not
  g225
  (
    n183,
    n40
  );


  buf
  g226
  (
    n288,
    n136
  );


  buf
  g227
  (
    n402,
    n145
  );


  not
  g228
  (
    n252,
    n109
  );


  not
  g229
  (
    n448,
    n142
  );


  not
  g230
  (
    n378,
    n89
  );


  not
  g231
  (
    n258,
    n65
  );


  buf
  g232
  (
    n315,
    n100
  );


  buf
  g233
  (
    n386,
    n84
  );


  not
  g234
  (
    n412,
    n103
  );


  not
  g235
  (
    n199,
    n131
  );


  not
  g236
  (
    n555,
    n72
  );


  not
  g237
  (
    n474,
    n37
  );


  not
  g238
  (
    n529,
    n116
  );


  not
  g239
  (
    n391,
    n75
  );


  not
  g240
  (
    n484,
    n148
  );


  buf
  g241
  (
    n527,
    n109
  );


  buf
  g242
  (
    n551,
    n90
  );


  buf
  g243
  (
    n230,
    n42
  );


  not
  g244
  (
    n557,
    n58
  );


  not
  g245
  (
    n549,
    n68
  );


  not
  g246
  (
    n206,
    n53
  );


  buf
  g247
  (
    n403,
    n137
  );


  buf
  g248
  (
    n180,
    n127
  );


  buf
  g249
  (
    n475,
    n129
  );


  not
  g250
  (
    n247,
    n44
  );


  not
  g251
  (
    n417,
    n87
  );


  not
  g252
  (
    n579,
    n39
  );


  buf
  g253
  (
    n367,
    n132
  );


  buf
  g254
  (
    n535,
    n110
  );


  buf
  g255
  (
    n239,
    n53
  );


  buf
  g256
  (
    n256,
    n35
  );


  buf
  g257
  (
    n525,
    n104
  );


  buf
  g258
  (
    n577,
    n56
  );


  not
  g259
  (
    n355,
    n91
  );


  not
  g260
  (
    n424,
    n74
  );


  buf
  g261
  (
    n316,
    n128
  );


  not
  g262
  (
    n241,
    n95
  );


  not
  g263
  (
    n536,
    n96
  );


  not
  g264
  (
    n216,
    n122
  );


  not
  g265
  (
    n275,
    n73
  );


  not
  g266
  (
    n253,
    n108
  );


  buf
  g267
  (
    n585,
    n104
  );


  buf
  g268
  (
    n406,
    n59
  );


  buf
  g269
  (
    n550,
    n80
  );


  buf
  g270
  (
    n318,
    n137
  );


  not
  g271
  (
    n192,
    n74
  );


  not
  g272
  (
    n189,
    n154
  );


  buf
  g273
  (
    n298,
    n57
  );


  not
  g274
  (
    n506,
    n110
  );


  buf
  g275
  (
    n299,
    n63
  );


  buf
  g276
  (
    n283,
    n146
  );


  buf
  g277
  (
    n184,
    n83
  );


  not
  g278
  (
    n586,
    n155
  );


  not
  g279
  (
    n162,
    n135
  );


  buf
  g280
  (
    n510,
    n136
  );


  not
  g281
  (
    n373,
    n73
  );


  buf
  g282
  (
    n483,
    n146
  );


  not
  g283
  (
    n561,
    n113
  );


  buf
  g284
  (
    n478,
    n56
  );


  not
  g285
  (
    n235,
    n66
  );


  buf
  g286
  (
    n530,
    n140
  );


  not
  g287
  (
    n201,
    n154
  );


  buf
  g288
  (
    n480,
    n92
  );


  buf
  g289
  (
    n531,
    n96
  );


  not
  g290
  (
    n194,
    n63
  );


  buf
  g291
  (
    n290,
    n136
  );


  not
  g292
  (
    n395,
    n139
  );


  buf
  g293
  (
    n351,
    n84
  );


  buf
  g294
  (
    n320,
    n102
  );


  buf
  g295
  (
    n485,
    n67
  );


  not
  g296
  (
    n327,
    n50
  );


  buf
  g297
  (
    n173,
    n131
  );


  not
  g298
  (
    n452,
    n36
  );


  buf
  g299
  (
    n528,
    n54
  );


  buf
  g300
  (
    n503,
    n51
  );


  not
  g301
  (
    n307,
    n33
  );


  buf
  g302
  (
    n233,
    n123
  );


  buf
  g303
  (
    n501,
    n142
  );


  buf
  g304
  (
    n499,
    n48
  );


  not
  g305
  (
    n203,
    n79
  );


  not
  g306
  (
    n231,
    n148
  );


  buf
  g307
  (
    n571,
    n103
  );


  not
  g308
  (
    n418,
    n70
  );


  buf
  g309
  (
    n306,
    n101
  );


  buf
  g310
  (
    n431,
    n137
  );


  not
  g311
  (
    n569,
    n130
  );


  buf
  g312
  (
    n168,
    n85
  );


  buf
  g313
  (
    n169,
    n71
  );


  buf
  g314
  (
    n166,
    n49
  );


  buf
  g315
  (
    n493,
    n97
  );


  buf
  g316
  (
    n350,
    n130
  );


  buf
  g317
  (
    n157,
    n144
  );


  not
  g318
  (
    n332,
    n152
  );


  buf
  g319
  (
    n313,
    n121
  );


  buf
  g320
  (
    n242,
    n66
  );


  buf
  g321
  (
    n444,
    n84
  );


  buf
  g322
  (
    n441,
    n82
  );


  not
  g323
  (
    n190,
    n119
  );


  buf
  g324
  (
    n213,
    n46
  );


  buf
  g325
  (
    n383,
    n69
  );


  buf
  g326
  (
    n160,
    n90
  );


  not
  g327
  (
    n454,
    n52
  );


  not
  g328
  (
    n346,
    n63
  );


  not
  g329
  (
    n323,
    n105
  );


  buf
  g330
  (
    n548,
    n52
  );


  not
  g331
  (
    n374,
    n45
  );


  not
  g332
  (
    n267,
    n70
  );


  buf
  g333
  (
    n377,
    n143
  );


  buf
  g334
  (
    n337,
    n51
  );


  not
  g335
  (
    n270,
    n82
  );


  buf
  g336
  (
    n277,
    n115
  );


  not
  g337
  (
    n196,
    n91
  );


  buf
  g338
  (
    n422,
    n90
  );


  buf
  g339
  (
    n541,
    n106
  );


  buf
  g340
  (
    n361,
    n36
  );


  not
  g341
  (
    n291,
    n118
  );


  not
  g342
  (
    n567,
    n77
  );


  not
  g343
  (
    n165,
    n152
  );


  not
  g344
  (
    n543,
    n147
  );


  buf
  g345
  (
    n331,
    n92
  );


  not
  g346
  (
    n294,
    n144
  );


  buf
  g347
  (
    n413,
    n126
  );


  buf
  g348
  (
    n504,
    n67
  );


  not
  g349
  (
    n496,
    n57
  );


  buf
  g350
  (
    n574,
    n48
  );


  buf
  g351
  (
    n302,
    n76
  );


  not
  g352
  (
    n304,
    n77
  );


  buf
  g353
  (
    n442,
    n146
  );


  buf
  g354
  (
    n426,
    n34
  );


  buf
  g355
  (
    n394,
    n145
  );


  buf
  g356
  (
    n547,
    n134
  );


  not
  g357
  (
    n439,
    n43
  );


  not
  g358
  (
    n554,
    n38
  );


  not
  g359
  (
    n363,
    n78
  );


  buf
  g360
  (
    n261,
    n76
  );


  buf
  g361
  (
    n471,
    n149
  );


  buf
  g362
  (
    n430,
    n141
  );


  not
  g363
  (
    n158,
    n76
  );


  not
  g364
  (
    n462,
    n124
  );


  not
  g365
  (
    n193,
    n90
  );


  buf
  g366
  (
    n455,
    n140
  );


  not
  g367
  (
    n434,
    n78
  );


  buf
  g368
  (
    n564,
    n134
  );


  not
  g369
  (
    n237,
    n120
  );


  buf
  g370
  (
    n211,
    n134
  );


  buf
  g371
  (
    n264,
    n93
  );


  buf
  g372
  (
    n178,
    n91
  );


  not
  g373
  (
    n505,
    n82
  );


  not
  g374
  (
    n526,
    n60
  );


  not
  g375
  (
    n498,
    n71
  );


  not
  g376
  (
    n364,
    n36
  );


  buf
  g377
  (
    n479,
    n47
  );


  not
  g378
  (
    n245,
    n67
  );


  not
  g379
  (
    n589,
    n54
  );


  buf
  g380
  (
    n297,
    n43
  );


  buf
  g381
  (
    n248,
    n44
  );


  not
  g382
  (
    n488,
    n112
  );


  not
  g383
  (
    n215,
    n87
  );


  not
  g384
  (
    n197,
    n71
  );


  buf
  g385
  (
    n265,
    n33
  );


  buf
  g386
  (
    n481,
    n45
  );


  buf
  g387
  (
    n490,
    n58
  );


  not
  g388
  (
    n243,
    n147
  );


  not
  g389
  (
    n387,
    n93
  );


  not
  g390
  (
    n282,
    n153
  );


  buf
  g391
  (
    n210,
    n77
  );


  buf
  g392
  (
    n522,
    n69
  );


  buf
  g393
  (
    n575,
    n130
  );


  buf
  g394
  (
    n500,
    n127
  );


  not
  g395
  (
    n556,
    n115
  );


  buf
  g396
  (
    n227,
    n64
  );


  not
  g397
  (
    n524,
    n40
  );


  not
  g398
  (
    n407,
    n47
  );


  not
  g399
  (
    n198,
    n86
  );


  not
  g400
  (
    n389,
    n50
  );


  not
  g401
  (
    n311,
    n41
  );


  buf
  g402
  (
    n260,
    n92
  );


  buf
  g403
  (
    n219,
    n61
  );


  buf
  g404
  (
    n438,
    n56
  );


  not
  g405
  (
    n515,
    n150
  );


  buf
  g406
  (
    n272,
    n50
  );


  buf
  g407
  (
    n494,
    n93
  );


  not
  g408
  (
    n300,
    n101
  );


  buf
  g409
  (
    n236,
    n139
  );


  buf
  g410
  (
    n295,
    n118
  );


  buf
  g411
  (
    n353,
    n44
  );


  not
  g412
  (
    n289,
    n88
  );


  buf
  g413
  (
    n415,
    n125
  );


  not
  g414
  (
    n240,
    n114
  );


  buf
  g415
  (
    n519,
    n94
  );


  buf
  g416
  (
    n509,
    n48
  );


  not
  g417
  (
    n185,
    n39
  );


  buf
  g418
  (
    n382,
    n75
  );


  not
  g419
  (
    n172,
    n128
  );


  not
  g420
  (
    n285,
    n142
  );


  not
  g421
  (
    n263,
    n117
  );


  not
  g422
  (
    n343,
    n114
  );


  buf
  g423
  (
    n188,
    n145
  );


  buf
  g424
  (
    n390,
    n87
  );


  buf
  g425
  (
    n445,
    n64
  );


  not
  g426
  (
    n330,
    n143
  );


  buf
  g427
  (
    n419,
    n43
  );


  not
  g428
  (
    n284,
    n44
  );


  not
  g429
  (
    n303,
    n118
  );


  not
  g430
  (
    n222,
    n74
  );


  not
  g431
  (
    n202,
    n106
  );


  buf
  g432
  (
    n470,
    n86
  );


  buf
  g433
  (
    n514,
    n35
  );


  buf
  g434
  (
    n461,
    n60
  );


  buf
  g435
  (
    n246,
    n103
  );


  buf
  g436
  (
    n512,
    n53
  );


  not
  g437
  (
    n317,
    n141
  );


  not
  g438
  (
    n497,
    n141
  );


  not
  g439
  (
    n420,
    n51
  );


  buf
  g440
  (
    n249,
    n45
  );


  not
  g441
  (
    n453,
    n94
  );


  not
  g442
  (
    n492,
    n126
  );


  not
  g443
  (
    n175,
    n99
  );


  buf
  g444
  (
    n456,
    n146
  );


  buf
  g445
  (
    n223,
    n62
  );


  buf
  g446
  (
    n473,
    n132
  );


  buf
  g447
  (
    n354,
    n107
  );


  buf
  g448
  (
    n312,
    n144
  );


  not
  g449
  (
    n358,
    n74
  );


  buf
  g450
  (
    n207,
    n122
  );


  buf
  g451
  (
    n451,
    n151
  );


  not
  g452
  (
    n257,
    n83
  );


  not
  g453
  (
    n559,
    n111
  );


  buf
  g454
  (
    n186,
    n151
  );


  buf
  g455
  (
    n437,
    n55
  );


  not
  g456
  (
    n491,
    n63
  );


  not
  g457
  (
    n301,
    n80
  );


  not
  g458
  (
    n404,
    n50
  );


  buf
  g459
  (
    n385,
    n41
  );


  buf
  g460
  (
    n532,
    n49
  );


  buf
  g461
  (
    n159,
    n57
  );


  buf
  g462
  (
    n381,
    n73
  );


  buf
  g463
  (
    n440,
    n153
  );


  buf
  g464
  (
    n511,
    n129
  );


  buf
  g465
  (
    n224,
    n75
  );


  buf
  g466
  (
    n421,
    n37
  );


  buf
  g467
  (
    n209,
    n38
  );


  buf
  g468
  (
    n310,
    n95
  );


  not
  g469
  (
    n187,
    n133
  );


  not
  g470
  (
    n191,
    n68
  );


  buf
  g471
  (
    n380,
    n52
  );


  buf
  g472
  (
    n540,
    n97
  );


  not
  g473
  (
    n356,
    n138
  );


  not
  g474
  (
    n533,
    n35
  );


  buf
  g475
  (
    n309,
    n125
  );


  buf
  g476
  (
    n329,
    n81
  );


  buf
  g477
  (
    n345,
    n58
  );


  not
  g478
  (
    n408,
    n55
  );


  not
  g479
  (
    n487,
    n116
  );


  buf
  g480
  (
    n513,
    n122
  );


  not
  g481
  (
    n414,
    n70
  );


  not
  g482
  (
    n296,
    n117
  );


  buf
  g483
  (
    n262,
    n75
  );


  buf
  g484
  (
    n273,
    n96
  );


  not
  g485
  (
    n325,
    n45
  );


  buf
  g486
  (
    n409,
    n86
  );


  not
  g487
  (
    n552,
    n103
  );


  buf
  g488
  (
    n369,
    n98
  );


  not
  g489
  (
    n463,
    n65
  );


  buf
  g490
  (
    n578,
    n153
  );


  buf
  g491
  (
    n450,
    n111
  );


  buf
  g492
  (
    n379,
    n133
  );


  not
  g493
  (
    n274,
    n150
  );


  buf
  g494
  (
    n502,
    n142
  );


  not
  g495
  (
    n566,
    n105
  );


  buf
  g496
  (
    n521,
    n114
  );


  buf
  g497
  (
    n467,
    n72
  );


  buf
  g498
  (
    n174,
    n40
  );


  not
  g499
  (
    n163,
    n116
  );


  not
  g500
  (
    n489,
    n138
  );


  buf
  g501
  (
    n251,
    n145
  );


  buf
  g502
  (
    n590,
    n60
  );


  buf
  g503
  (
    n410,
    n83
  );


  buf
  g504
  (
    n335,
    n150
  );


  not
  g505
  (
    n271,
    n135
  );


  not
  g506
  (
    n372,
    n88
  );


  buf
  g507
  (
    n495,
    n61
  );


  not
  g508
  (
    n287,
    n131
  );


  buf
  g509
  (
    n539,
    n67
  );


  buf
  g510
  (
    n428,
    n35
  );


  not
  g511
  (
    n225,
    n129
  );


  buf
  g512
  (
    n545,
    n76
  );


  buf
  g513
  (
    n357,
    n132
  );


  buf
  g514
  (
    n563,
    n113
  );


  buf
  g515
  (
    n314,
    n151
  );


  buf
  g516
  (
    n170,
    n62
  );


  not
  g517
  (
    n516,
    n47
  );


  buf
  g518
  (
    n208,
    n97
  );


  buf
  g519
  (
    n279,
    n117
  );


  buf
  g520
  (
    n176,
    n151
  );


  buf
  g521
  (
    n433,
    n106
  );


  buf
  g522
  (
    n572,
    n68
  );


  buf
  g523
  (
    n293,
    n94
  );


  not
  g524
  (
    n573,
    n66
  );


  not
  g525
  (
    n466,
    n149
  );


  buf
  g526
  (
    n319,
    n79
  );


  not
  g527
  (
    n182,
    n34
  );


  buf
  g528
  (
    n340,
    n88
  );


  not
  g529
  (
    n328,
    n79
  );


  not
  g530
  (
    n429,
    n79
  );


  buf
  g531
  (
    n560,
    n81
  );


  not
  g532
  (
    n226,
    n85
  );


  not
  g533
  (
    n167,
    n34
  );


  buf
  g534
  (
    n268,
    n107
  );


  buf
  g535
  (
    n228,
    n108
  );


  buf
  g536
  (
    n368,
    n119
  );


  buf
  g537
  (
    n469,
    n84
  );


  not
  g538
  (
    n177,
    n121
  );


  and
  g539
  (
    n164,
    n104,
    n136
  );


  xor
  g540
  (
    n359,
    n110,
    n33,
    n107,
    n135
  );


  nand
  g541
  (
    n397,
    n116,
    n105,
    n86,
    n70
  );


  nor
  g542
  (
    n200,
    n112,
    n65,
    n124,
    n113
  );


  xor
  g543
  (
    n449,
    n83,
    n94,
    n42,
    n54
  );


  xor
  g544
  (
    n508,
    n118,
    n53,
    n99,
    n143
  );


  nor
  g545
  (
    n341,
    n129,
    n115,
    n42,
    n78
  );


  and
  g546
  (
    n205,
    n47,
    n152,
    n81,
    n125
  );


  nor
  g547
  (
    n171,
    n41,
    n115,
    n104,
    n85
  );


  or
  g548
  (
    n217,
    n46,
    n93,
    n97,
    n99
  );


  xor
  g549
  (
    n460,
    n111,
    n123,
    n132,
    n49
  );


  nor
  g550
  (
    n405,
    n57,
    n122,
    n124,
    n61
  );


  or
  g551
  (
    n392,
    n109,
    n69,
    n124,
    n68
  );


  and
  g552
  (
    n322,
    n59,
    n111,
    n61,
    n38
  );


  and
  g553
  (
    n399,
    n40,
    n38,
    n80,
    n106
  );


  xnor
  g554
  (
    n234,
    n59,
    n147,
    n102,
    n148
  );


  xnor
  g555
  (
    n435,
    n39,
    n139,
    n121,
    n135
  );


  nor
  g556
  (
    n436,
    n108,
    n52,
    n153,
    n80
  );


  or
  g557
  (
    n349,
    n100,
    n100,
    n112,
    n89
  );


  not
  g558
  (
    n715,
    n381
  );


  buf
  g559
  (
    n855,
    n238
  );


  buf
  g560
  (
    n748,
    n469
  );


  buf
  g561
  (
    n733,
    n390
  );


  buf
  g562
  (
    n685,
    n405
  );


  buf
  g563
  (
    n762,
    n32
  );


  buf
  g564
  (
    n606,
    n282
  );


  not
  g565
  (
    n757,
    n346
  );


  buf
  g566
  (
    n792,
    n323
  );


  not
  g567
  (
    n712,
    n362
  );


  not
  g568
  (
    n800,
    n217
  );


  buf
  g569
  (
    n775,
    n451
  );


  buf
  g570
  (
    n817,
    n459
  );


  not
  g571
  (
    n666,
    n441
  );


  buf
  g572
  (
    n761,
    n336
  );


  not
  g573
  (
    n839,
    n493
  );


  buf
  g574
  (
    n706,
    n364
  );


  not
  g575
  (
    n831,
    n375
  );


  not
  g576
  (
    n840,
    n383
  );


  buf
  g577
  (
    n773,
    n386
  );


  not
  g578
  (
    n822,
    n479
  );


  buf
  g579
  (
    n835,
    n406
  );


  not
  g580
  (
    n638,
    n264
  );


  not
  g581
  (
    n668,
    n203
  );


  buf
  g582
  (
    n816,
    n280
  );


  buf
  g583
  (
    n842,
    n190
  );


  not
  g584
  (
    n728,
    n420
  );


  not
  g585
  (
    n681,
    n418
  );


  buf
  g586
  (
    n841,
    n423
  );


  buf
  g587
  (
    n665,
    n455
  );


  buf
  g588
  (
    n592,
    n498
  );


  buf
  g589
  (
    n652,
    n517
  );


  buf
  g590
  (
    n722,
    n449
  );


  not
  g591
  (
    n672,
    n438
  );


  not
  g592
  (
    n673,
    n202
  );


  buf
  g593
  (
    n694,
    n456
  );


  buf
  g594
  (
    n716,
    n286
  );


  buf
  g595
  (
    n714,
    n510
  );


  not
  g596
  (
    n649,
    n427
  );


  buf
  g597
  (
    n600,
    n349
  );


  not
  g598
  (
    n812,
    n170
  );


  not
  g599
  (
    n594,
    n201
  );


  buf
  g600
  (
    n727,
    n341
  );


  buf
  g601
  (
    n660,
    n489
  );


  not
  g602
  (
    n732,
    n454
  );


  buf
  g603
  (
    n861,
    n178
  );


  not
  g604
  (
    n791,
    n539
  );


  buf
  g605
  (
    n749,
    n310
  );


  not
  g606
  (
    n785,
    n157
  );


  not
  g607
  (
    n752,
    n397
  );


  not
  g608
  (
    n726,
    n325
  );


  buf
  g609
  (
    n631,
    n446
  );


  buf
  g610
  (
    n782,
    n313
  );


  not
  g611
  (
    n744,
    n301
  );


  not
  g612
  (
    n736,
    n215
  );


  buf
  g613
  (
    n711,
    n251
  );


  not
  g614
  (
    n787,
    n347
  );


  buf
  g615
  (
    n696,
    n166
  );


  buf
  g616
  (
    n620,
    n532
  );


  buf
  g617
  (
    n635,
    n320
  );


  buf
  g618
  (
    n833,
    n32
  );


  buf
  g619
  (
    n760,
    n173
  );


  not
  g620
  (
    n676,
    n443
  );


  buf
  g621
  (
    n795,
    n165
  );


  not
  g622
  (
    n725,
    n351
  );


  buf
  g623
  (
    n717,
    n433
  );


  not
  g624
  (
    n664,
    n237
  );


  not
  g625
  (
    n648,
    n334
  );


  buf
  g626
  (
    n623,
    n542
  );


  buf
  g627
  (
    n700,
    n319
  );


  buf
  g628
  (
    n843,
    n512
  );


  not
  g629
  (
    n789,
    n276
  );


  not
  g630
  (
    n814,
    n186
  );


  not
  g631
  (
    n597,
    n533
  );


  buf
  g632
  (
    n758,
    n552
  );


  buf
  g633
  (
    n671,
    n354
  );


  not
  g634
  (
    n836,
    n348
  );


  buf
  g635
  (
    n679,
    n359
  );


  buf
  g636
  (
    n598,
    n249
  );


  not
  g637
  (
    n713,
    n486
  );


  buf
  g638
  (
    n615,
    n429
  );


  not
  g639
  (
    n846,
    n252
  );


  not
  g640
  (
    n820,
    n399
  );


  not
  g641
  (
    n810,
    n507
  );


  not
  g642
  (
    n844,
    n260
  );


  buf
  g643
  (
    n860,
    n345
  );


  not
  g644
  (
    n729,
    n470
  );


  buf
  g645
  (
    n610,
    n232
  );


  not
  g646
  (
    n826,
    n541
  );


  not
  g647
  (
    n639,
    n184
  );


  buf
  g648
  (
    n621,
    n234
  );


  buf
  g649
  (
    n680,
    n377
  );


  buf
  g650
  (
    n675,
    n544
  );


  not
  g651
  (
    n739,
    n283
  );


  not
  g652
  (
    n740,
    n548
  );


  not
  g653
  (
    n720,
    n374
  );


  not
  g654
  (
    n763,
    n285
  );


  not
  g655
  (
    n609,
    n478
  );


  not
  g656
  (
    n601,
    n227
  );


  buf
  g657
  (
    n663,
    n309
  );


  not
  g658
  (
    n695,
    n273
  );


  buf
  g659
  (
    n693,
    n226
  );


  buf
  g660
  (
    n779,
    n487
  );


  not
  g661
  (
    n599,
    n463
  );


  not
  g662
  (
    n625,
    n287
  );


  not
  g663
  (
    n818,
    n32
  );


  buf
  g664
  (
    n703,
    n550
  );


  not
  g665
  (
    n838,
    n216
  );


  not
  g666
  (
    n622,
    n236
  );


  not
  g667
  (
    n815,
    n317
  );


  not
  g668
  (
    n604,
    n316
  );


  not
  g669
  (
    n830,
    n272
  );


  not
  g670
  (
    n858,
    n247
  );


  not
  g671
  (
    n737,
    n530
  );


  buf
  g672
  (
    n677,
    n255
  );


  buf
  g673
  (
    n783,
    n222
  );


  buf
  g674
  (
    n661,
    n277
  );


  buf
  g675
  (
    n662,
    n240
  );


  not
  g676
  (
    n853,
    n307
  );


  not
  g677
  (
    n742,
    n332
  );


  not
  g678
  (
    n697,
    n492
  );


  buf
  g679
  (
    n778,
    n302
  );


  not
  g680
  (
    n845,
    n183
  );


  not
  g681
  (
    n643,
    n426
  );


  buf
  g682
  (
    n731,
    n461
  );


  not
  g683
  (
    n854,
    n466
  );


  not
  g684
  (
    n644,
    n164
  );


  buf
  g685
  (
    n756,
    n417
  );


  not
  g686
  (
    n786,
    n239
  );


  not
  g687
  (
    n650,
    n546
  );


  not
  g688
  (
    n658,
    n372
  );


  not
  g689
  (
    n847,
    n484
  );


  buf
  g690
  (
    n832,
    n180
  );


  buf
  g691
  (
    n751,
    n407
  );


  buf
  g692
  (
    n718,
    n502
  );


  buf
  g693
  (
    n755,
    n520
  );


  not
  g694
  (
    n708,
    n514
  );


  not
  g695
  (
    n851,
    n472
  );


  buf
  g696
  (
    n811,
    n174
  );


  buf
  g697
  (
    n595,
    n194
  );


  not
  g698
  (
    n852,
    n297
  );


  buf
  g699
  (
    n684,
    n160
  );


  not
  g700
  (
    n616,
    n181
  );


  buf
  g701
  (
    n784,
    n430
  );


  buf
  g702
  (
    n730,
    n248
  );


  buf
  g703
  (
    n655,
    n223
  );


  not
  g704
  (
    n827,
    n439
  );


  not
  g705
  (
    n799,
    n494
  );


  buf
  g706
  (
    n614,
    n196
  );


  not
  g707
  (
    n813,
    n501
  );


  not
  g708
  (
    n741,
    n523
  );


  not
  g709
  (
    n687,
    n367
  );


  buf
  g710
  (
    n634,
    n213
  );


  not
  g711
  (
    n856,
    n350
  );


  buf
  g712
  (
    n721,
    n321
  );


  buf
  g713
  (
    n669,
    n370
  );


  buf
  g714
  (
    n806,
    n527
  );


  not
  g715
  (
    n809,
    n534
  );


  buf
  g716
  (
    n774,
    n491
  );


  buf
  g717
  (
    n659,
    n169
  );


  not
  g718
  (
    n777,
    n495
  );


  not
  g719
  (
    n629,
    n480
  );


  buf
  g720
  (
    n608,
    n329
  );


  not
  g721
  (
    n704,
    n434
  );


  not
  g722
  (
    n764,
    n391
  );


  buf
  g723
  (
    n642,
    n192
  );


  buf
  g724
  (
    n654,
    n177
  );


  not
  g725
  (
    n735,
    n250
  );


  buf
  g726
  (
    n651,
    n214
  );


  buf
  g727
  (
    n793,
    n210
  );


  buf
  g728
  (
    n647,
    n398
  );


  buf
  g729
  (
    n724,
    n337
  );


  not
  g730
  (
    n596,
    n274
  );


  not
  g731
  (
    n801,
    n444
  );


  buf
  g732
  (
    n632,
    n328
  );


  not
  g733
  (
    n745,
    n483
  );


  not
  g734
  (
    n803,
    n355
  );


  not
  g735
  (
    n709,
    n296
  );


  not
  g736
  (
    n828,
    n424
  );


  not
  g737
  (
    n591,
    n208
  );


  not
  g738
  (
    n759,
    n342
  );


  not
  g739
  (
    n857,
    n545
  );


  buf
  g740
  (
    n674,
    n551
  );


  buf
  g741
  (
    n611,
    n508
  );


  not
  g742
  (
    n776,
    n188
  );


  not
  g743
  (
    n808,
    n299
  );


  buf
  g744
  (
    n807,
    n211
  );


  not
  g745
  (
    n699,
    n340
  );


  not
  g746
  (
    n626,
    n267
  );


  buf
  g747
  (
    n682,
    n318
  );


  buf
  g748
  (
    n689,
    n293
  );


  not
  g749
  (
    n657,
    n525
  );


  not
  g750
  (
    n710,
    n476
  );


  not
  g751
  (
    n825,
    n327
  );


  buf
  g752
  (
    n691,
    n360
  );


  buf
  g753
  (
    n678,
    n477
  );


  buf
  g754
  (
    n633,
    n504
  );


  buf
  g755
  (
    n805,
    n314
  );


  buf
  g756
  (
    n788,
    n195
  );


  buf
  g757
  (
    n824,
    n535
  );


  buf
  g758
  (
    n617,
    n246
  );


  not
  g759
  (
    n796,
    n197
  );


  not
  g760
  (
    n690,
    n528
  );


  not
  g761
  (
    n653,
    n531
  );


  not
  g762
  (
    n667,
    n338
  );


  not
  g763
  (
    n849,
    n256
  );


  not
  g764
  (
    n821,
    n220
  );


  not
  g765
  (
    n698,
    n228
  );


  not
  g766
  (
    n743,
    n428
  );


  buf
  g767
  (
    n771,
    n488
  );


  buf
  g768
  (
    n646,
    n305
  );


  buf
  g769
  (
    n640,
    n290
  );


  buf
  g770
  (
    n738,
    n524
  );


  buf
  g771
  (
    n754,
    n462
  );


  not
  g772
  (
    n819,
    n221
  );


  buf
  g773
  (
    n850,
    n505
  );


  not
  g774
  (
    n612,
    n416
  );


  buf
  g775
  (
    n848,
    n413
  );


  buf
  g776
  (
    n765,
    n294
  );


  not
  g777
  (
    n670,
    n475
  );


  not
  g778
  (
    n802,
    n450
  );


  buf
  g779
  (
    n734,
    n193
  );


  not
  g780
  (
    n781,
    n388
  );


  buf
  g781
  (
    n770,
    n402
  );


  not
  g782
  (
    n707,
    n233
  );


  not
  g783
  (
    n750,
    n243
  );


  not
  g784
  (
    n829,
    n404
  );


  not
  g785
  (
    n628,
    n179
  );


  not
  g786
  (
    n705,
    n437
  );


  buf
  g787
  (
    n766,
    n275
  );


  and
  g788
  (
    n768,
    n263,
    n261
  );


  or
  g789
  (
    n797,
    n254,
    n468,
    n421,
    n171
  );


  and
  g790
  (
    n603,
    n509,
    n209,
    n311,
    n266
  );


  xor
  g791
  (
    n862,
    n205,
    n547,
    n518,
    n284
  );


  xnor
  g792
  (
    n627,
    n380,
    n403,
    n212,
    n511
  );


  or
  g793
  (
    n686,
    n207,
    n185,
    n503,
    n32
  );


  nor
  g794
  (
    n746,
    n442,
    n315,
    n167,
    n522
  );


  nand
  g795
  (
    n637,
    n303,
    n432,
    n187,
    n312
  );


  xor
  g796
  (
    n859,
    n387,
    n271,
    n335,
    n435
  );


  nor
  g797
  (
    n798,
    n245,
    n447,
    n229,
    n369
  );


  xor
  g798
  (
    n863,
    n536,
    n224,
    n235,
    n457
  );


  nor
  g799
  (
    n804,
    n497,
    n445,
    n361,
    n358
  );


  nand
  g800
  (
    n656,
    n401,
    n230,
    n163,
    n425
  );


  xor
  g801
  (
    n767,
    n485,
    n490,
    n204,
    n253
  );


  nand
  g802
  (
    n624,
    n521,
    n191,
    n175,
    n265
  );


  and
  g803
  (
    n747,
    n343,
    n159,
    n396,
    n182
  );


  or
  g804
  (
    n723,
    n382,
    n161,
    n519,
    n356
  );


  and
  g805
  (
    n701,
    n409,
    n298,
    n378,
    n458
  );


  and
  g806
  (
    n772,
    n422,
    n330,
    n344,
    n288
  );


  xnor
  g807
  (
    n790,
    n411,
    n415,
    n482,
    n300
  );


  nand
  g808
  (
    n719,
    n291,
    n259,
    n331,
    n500
  );


  nand
  g809
  (
    n692,
    n242,
    n176,
    n389,
    n322
  );


  xor
  g810
  (
    n593,
    n464,
    n393,
    n394,
    n244
  );


  nor
  g811
  (
    n794,
    n219,
    n268,
    n326,
    n410
  );


  xnor
  g812
  (
    n702,
    n465,
    n308,
    n241,
    n189
  );


  and
  g813
  (
    n607,
    n385,
    n306,
    n278,
    n481
  );


  nor
  g814
  (
    n834,
    n162,
    n412,
    n440,
    n270
  );


  nand
  g815
  (
    n602,
    n198,
    n158,
    n540,
    n473
  );


  nand
  g816
  (
    n618,
    n371,
    n395,
    n172,
    n467
  );


  nand
  g817
  (
    n641,
    n352,
    n168,
    n526,
    n199
  );


  xor
  g818
  (
    n636,
    n353,
    n515,
    n258,
    n474
  );


  nand
  g819
  (
    n823,
    n448,
    n373,
    n513,
    n452
  );


  and
  g820
  (
    n837,
    n431,
    n376,
    n460,
    n262
  );


  nor
  g821
  (
    n769,
    n295,
    n419,
    n496,
    n218
  );


  xnor
  g822
  (
    n630,
    n436,
    n499,
    n231,
    n357
  );


  nor
  g823
  (
    n605,
    n453,
    n400,
    n366,
    n279
  );


  and
  g824
  (
    n683,
    n529,
    n365,
    n363,
    n506
  );


  xnor
  g825
  (
    n619,
    n339,
    n304,
    n549,
    n392
  );


  xnor
  g826
  (
    n753,
    n537,
    n333,
    n368,
    n292
  );


  or
  g827
  (
    n780,
    n206,
    n379,
    n516,
    n281
  );


  or
  g828
  (
    n688,
    n384,
    n324,
    n257,
    n289
  );


  xnor
  g829
  (
    n645,
    n225,
    n200,
    n538,
    n414
  );


  and
  g830
  (
    n613,
    n269,
    n471,
    n408,
    n543
  );


  buf
  g831
  (
    n865,
    n592
  );


  buf
  g832
  (
    n864,
    n591
  );


  and
  g833
  (
    n873,
    n563,
    n570,
    n571,
    n574
  );


  nor
  g834
  (
    n868,
    n575,
    n865,
    n566
  );


  xnor
  g835
  (
    n872,
    n864,
    n567,
    n560,
    n572
  );


  nand
  g836
  (
    n869,
    n568,
    n864,
    n562,
    n865
  );


  nor
  g837
  (
    n871,
    n573,
    n864,
    n565,
    n554
  );


  nor
  g838
  (
    n866,
    n576,
    n864,
    n558,
    n559
  );


  nor
  g839
  (
    n870,
    n555,
    n561,
    n569,
    n564
  );


  or
  g840
  (
    n867,
    n865,
    n556,
    n557,
    n553
  );


  buf
  g841
  (
    n880,
    n869
  );


  buf
  g842
  (
    n882,
    n866
  );


  not
  g843
  (
    n884,
    n867
  );


  buf
  g844
  (
    n889,
    n869
  );


  not
  g845
  (
    n876,
    n867
  );


  not
  g846
  (
    n887,
    n870
  );


  not
  g847
  (
    n888,
    n867
  );


  buf
  g848
  (
    n878,
    n866
  );


  not
  g849
  (
    n879,
    n867
  );


  not
  g850
  (
    n885,
    n868
  );


  not
  g851
  (
    n877,
    n868
  );


  not
  g852
  (
    n883,
    n869
  );


  not
  g853
  (
    n886,
    n869
  );


  buf
  g854
  (
    n875,
    n868
  );


  buf
  g855
  (
    n874,
    n868
  );


  not
  g856
  (
    n881,
    n870
  );


  xor
  g857
  (
    n929,
    n606,
    n688,
    n704,
    n878
  );


  nand
  g858
  (
    n920,
    n628,
    n629,
    n881,
    n880
  );


  nor
  g859
  (
    n923,
    n714,
    n709,
    n600,
    n877
  );


  or
  g860
  (
    n919,
    n676,
    n702,
    n715,
    n875
  );


  xor
  g861
  (
    n892,
    n875,
    n601,
    n708,
    n664
  );


  nand
  g862
  (
    n895,
    n882,
    n696,
    n712,
    n876
  );


  nand
  g863
  (
    n924,
    n630,
    n683,
    n717,
    n670
  );


  nand
  g864
  (
    n897,
    n597,
    n710,
    n678,
    n614
  );


  or
  g865
  (
    n917,
    n697,
    n632,
    n695,
    n875
  );


  xnor
  g866
  (
    n906,
    n653,
    n669,
    n883,
    n874
  );


  xnor
  g867
  (
    n930,
    n634,
    n883,
    n640,
    n713
  );


  or
  g868
  (
    n927,
    n593,
    n694,
    n685,
    n642
  );


  nor
  g869
  (
    n891,
    n668,
    n661,
    n880,
    n656
  );


  and
  g870
  (
    n899,
    n618,
    n626,
    n620,
    n663
  );


  and
  g871
  (
    n898,
    n648,
    n609,
    n631,
    n674
  );


  nand
  g872
  (
    n925,
    n619,
    n613,
    n881,
    n636
  );


  xor
  g873
  (
    n922,
    n875,
    n605,
    n687,
    n623
  );


  xnor
  g874
  (
    n903,
    n654,
    n877,
    n652,
    n878
  );


  xor
  g875
  (
    n913,
    n877,
    n686,
    n639,
    n658
  );


  nor
  g876
  (
    n918,
    n666,
    n647,
    n706,
    n655
  );


  nand
  g877
  (
    n894,
    n650,
    n879,
    n876,
    n667
  );


  xnor
  g878
  (
    n910,
    n874,
    n681,
    n701,
    n883
  );


  or
  g879
  (
    n915,
    n671,
    n603,
    n660,
    n675
  );


  xor
  g880
  (
    n916,
    n612,
    n662,
    n684,
    n635
  );


  xnor
  g881
  (
    n931,
    n596,
    n633,
    n637,
    n621
  );


  or
  g882
  (
    n928,
    n881,
    n698,
    n699,
    n716
  );


  and
  g883
  (
    n904,
    n884,
    n672,
    n881,
    n877
  );


  nor
  g884
  (
    n893,
    n665,
    n595,
    n682,
    n679
  );


  xnor
  g885
  (
    n912,
    n673,
    n625,
    n690,
    n645
  );


  nor
  g886
  (
    n911,
    n876,
    n649,
    n878,
    n705
  );


  nand
  g887
  (
    n921,
    n707,
    n882,
    n615,
    n622
  );


  nor
  g888
  (
    n896,
    n879,
    n599,
    n874,
    n624
  );


  xor
  g889
  (
    n909,
    n651,
    n608,
    n617,
    n644
  );


  xor
  g890
  (
    n926,
    n643,
    n882,
    n689,
    n703
  );


  nand
  g891
  (
    n901,
    n680,
    n638,
    n607,
    n594
  );


  or
  g892
  (
    n907,
    n700,
    n610,
    n693,
    n646
  );


  xor
  g893
  (
    n908,
    n883,
    n876,
    n878,
    n880
  );


  xor
  g894
  (
    n902,
    n677,
    n616,
    n641,
    n880
  );


  xnor
  g895
  (
    n900,
    n711,
    n611,
    n692,
    n657
  );


  or
  g896
  (
    n905,
    n598,
    n718,
    n627,
    n602
  );


  or
  g897
  (
    n890,
    n604,
    n884,
    n882,
    n659
  );


  nor
  g898
  (
    n914,
    n874,
    n879,
    n691
  );


  buf
  g899
  (
    n940,
    n896
  );


  buf
  g900
  (
    n937,
    n894
  );


  buf
  g901
  (
    n938,
    n897
  );


  not
  g902
  (
    n941,
    n898
  );


  not
  g903
  (
    n934,
    n892
  );


  not
  g904
  (
    n936,
    n899
  );


  not
  g905
  (
    n933,
    n890
  );


  buf
  g906
  (
    n939,
    n893
  );


  buf
  g907
  (
    n935,
    n895
  );


  not
  g908
  (
    n932,
    n891
  );


  or
  g909
  (
    n966,
    n939,
    n584
  );


  or
  g910
  (
    n967,
    n936,
    n730,
    n578,
    n724
  );


  nor
  g911
  (
    n958,
    n581,
    n935,
    n585,
    n909
  );


  and
  g912
  (
    n946,
    n885,
    n934,
    n156,
    n582
  );


  or
  g913
  (
    n964,
    n901,
    n889,
    n886,
    n937
  );


  xnor
  g914
  (
    n968,
    n940,
    n940,
    n885,
    n933
  );


  nand
  g915
  (
    n961,
    n579,
    n935,
    n886,
    n583
  );


  nand
  g916
  (
    n944,
    n934,
    n871,
    n728,
    n938
  );


  or
  g917
  (
    n952,
    n936,
    n902,
    n584,
    n720
  );


  nand
  g918
  (
    n956,
    n578,
    n578,
    n870,
    n903
  );


  nor
  g919
  (
    n943,
    n941,
    n887,
    n933,
    n938
  );


  xnor
  g920
  (
    n957,
    n585,
    n873,
    n722,
    n937
  );


  xnor
  g921
  (
    n953,
    n582,
    n577,
    n579,
    n155
  );


  nand
  g922
  (
    n960,
    n940,
    n937,
    n907,
    n908
  );


  xor
  g923
  (
    n963,
    n871,
    n887,
    n577,
    n884
  );


  or
  g924
  (
    n977,
    n932,
    n940,
    n581,
    n933
  );


  xor
  g925
  (
    n948,
    n585,
    n155,
    n900,
    n936
  );


  and
  g926
  (
    n954,
    n583,
    n873,
    n578,
    n581
  );


  or
  g927
  (
    n971,
    n580,
    n580,
    n939,
    n729
  );


  and
  g928
  (
    n950,
    n937,
    n932,
    n939,
    n871
  );


  xor
  g929
  (
    n978,
    n887,
    n577,
    n726,
    n582
  );


  xor
  g930
  (
    n949,
    n932,
    n584,
    n934,
    n586
  );


  and
  g931
  (
    n972,
    n905,
    n941,
    n873,
    n579
  );


  nand
  g932
  (
    n962,
    n889,
    n719,
    n583,
    n580
  );


  xnor
  g933
  (
    n955,
    n732,
    n886,
    n725,
    n936
  );


  nand
  g934
  (
    n959,
    n941,
    n932,
    n934,
    n939
  );


  nand
  g935
  (
    n969,
    n583,
    n585,
    n872,
    n871
  );


  xnor
  g936
  (
    n951,
    n586,
    n885,
    n872
  );


  or
  g937
  (
    n965,
    n579,
    n580,
    n872,
    n933
  );


  xnor
  g938
  (
    n975,
    n884,
    n584,
    n731,
    n938
  );


  xor
  g939
  (
    n947,
    n870,
    n889,
    n872,
    n577
  );


  nor
  g940
  (
    n970,
    n734,
    n888,
    n938,
    n911
  );


  or
  g941
  (
    n976,
    n889,
    n727,
    n888,
    n886
  );


  xor
  g942
  (
    n942,
    n935,
    n935,
    n910,
    n888
  );


  nand
  g943
  (
    n945,
    n904,
    n733,
    n723,
    n582
  );


  xnor
  g944
  (
    n973,
    n887,
    n941,
    n873,
    n906
  );


  nand
  g945
  (
    n974,
    n581,
    n155,
    n888,
    n721
  );


  not
  g946
  (
    n986,
    n912
  );


  buf
  g947
  (
    n979,
    n914
  );


  not
  g948
  (
    n983,
    n952
  );


  buf
  g949
  (
    n982,
    n917
  );


  not
  g950
  (
    n989,
    n951
  );


  not
  g951
  (
    n988,
    n917
  );


  buf
  g952
  (
    n984,
    n917
  );


  buf
  g953
  (
    n994,
    n954
  );


  buf
  g954
  (
    n990,
    n950
  );


  xnor
  g955
  (
    n992,
    n956,
    n915,
    n947
  );


  xor
  g956
  (
    n980,
    n955,
    n946,
    n949,
    n916
  );


  nor
  g957
  (
    n981,
    n916,
    n943,
    n913
  );


  xnor
  g958
  (
    n991,
    n944,
    n957,
    n915,
    n942
  );


  or
  g959
  (
    n993,
    n914,
    n953,
    n916,
    n917
  );


  or
  g960
  (
    n985,
    n914,
    n916,
    n913,
    n948
  );


  nor
  g961
  (
    n987,
    n945,
    n914,
    n915
  );


  not
  g962
  (
    n998,
    n918
  );


  buf
  g963
  (
    n1000,
    n979
  );


  buf
  g964
  (
    n996,
    n981
  );


  not
  g965
  (
    n997,
    n919
  );


  buf
  g966
  (
    n999,
    n979
  );


  or
  g967
  (
    n1003,
    n918,
    n979
  );


  xor
  g968
  (
    n995,
    n918,
    n980,
    n919
  );


  xor
  g969
  (
    n1001,
    n918,
    n980
  );


  xor
  g970
  (
    n1002,
    n979,
    n919,
    n980
  );


  not
  g971
  (
    n1036,
    n920
  );


  not
  g972
  (
    n1035,
    n922
  );


  buf
  g973
  (
    n1016,
    n1003
  );


  buf
  g974
  (
    n1015,
    n968
  );


  buf
  g975
  (
    n1022,
    n968
  );


  not
  g976
  (
    n1014,
    n921
  );


  not
  g977
  (
    n1021,
    n969
  );


  not
  g978
  (
    n1023,
    n1002
  );


  not
  g979
  (
    n1017,
    n1003
  );


  not
  g980
  (
    n1030,
    n997
  );


  buf
  g981
  (
    n1025,
    n922
  );


  not
  g982
  (
    n1009,
    n967
  );


  not
  g983
  (
    n1011,
    n998
  );


  buf
  g984
  (
    n1007,
    n961
  );


  buf
  g985
  (
    n1020,
    n1003
  );


  buf
  g986
  (
    n1005,
    n995
  );


  not
  g987
  (
    n1008,
    n964
  );


  not
  g988
  (
    n1038,
    n958
  );


  not
  g989
  (
    n1004,
    n969
  );


  buf
  g990
  (
    n1018,
    n921
  );


  not
  g991
  (
    n1031,
    n1002
  );


  not
  g992
  (
    n1019,
    n1001
  );


  and
  g993
  (
    n1026,
    n920,
    n1002
  );


  nor
  g994
  (
    n1032,
    n1001,
    n962,
    n997,
    n967
  );


  nor
  g995
  (
    n1033,
    n1003,
    n968,
    n960
  );


  xor
  g996
  (
    n1013,
    n920,
    n969,
    n1000,
    n996
  );


  or
  g997
  (
    n1027,
    n995,
    n963,
    n999,
    n996
  );


  nor
  g998
  (
    n1006,
    n998,
    n1000,
    n920,
    n997
  );


  and
  g999
  (
    n1010,
    n998,
    n967,
    n1001,
    n997
  );


  nor
  g1000
  (
    n1029,
    n995,
    n1002,
    n966,
    n970
  );


  xnor
  g1001
  (
    n1012,
    n969,
    n959,
    n998,
    n996
  );


  xor
  g1002
  (
    n1037,
    n922,
    n999,
    n1001
  );


  or
  g1003
  (
    n1028,
    n922,
    n970,
    n999,
    n1000
  );


  xor
  g1004
  (
    n1024,
    n996,
    n921,
    n1000,
    n919
  );


  and
  g1005
  (
    n1034,
    n970,
    n965,
    n967,
    n921
  );


  not
  g1006
  (
    n1110,
    n1025
  );


  not
  g1007
  (
    n1153,
    n1024
  );


  buf
  g1008
  (
    n1168,
    n1025
  );


  not
  g1009
  (
    n1117,
    n1033
  );


  not
  g1010
  (
    n1164,
    n974
  );


  not
  g1011
  (
    n1102,
    n1018
  );


  buf
  g1012
  (
    n1053,
    n1013
  );


  buf
  g1013
  (
    n1063,
    n1021
  );


  buf
  g1014
  (
    n1125,
    n984
  );


  not
  g1015
  (
    n1064,
    n981
  );


  buf
  g1016
  (
    n1104,
    n985
  );


  not
  g1017
  (
    n1041,
    n992
  );


  buf
  g1018
  (
    n1067,
    n1016
  );


  not
  g1019
  (
    n1145,
    n1034
  );


  not
  g1020
  (
    n1121,
    n1005
  );


  buf
  g1021
  (
    n1098,
    n1005
  );


  not
  g1022
  (
    n1144,
    n1014
  );


  buf
  g1023
  (
    n1149,
    n972
  );


  buf
  g1024
  (
    n1105,
    n1014
  );


  buf
  g1025
  (
    n1130,
    n1008
  );


  buf
  g1026
  (
    n1103,
    n1005
  );


  buf
  g1027
  (
    n1097,
    n982
  );


  not
  g1028
  (
    n1055,
    n1011
  );


  not
  g1029
  (
    n1079,
    n1012
  );


  not
  g1030
  (
    n1096,
    n1019
  );


  not
  g1031
  (
    n1113,
    n1015
  );


  not
  g1032
  (
    n1136,
    n1017
  );


  buf
  g1033
  (
    n1106,
    n988
  );


  not
  g1034
  (
    n1140,
    n1029
  );


  buf
  g1035
  (
    n1163,
    n1026
  );


  not
  g1036
  (
    n1135,
    n1008
  );


  not
  g1037
  (
    n1151,
    n991
  );


  not
  g1038
  (
    n1081,
    n976
  );


  buf
  g1039
  (
    n1085,
    n1017
  );


  not
  g1040
  (
    n1131,
    n1011
  );


  buf
  g1041
  (
    n1165,
    n976
  );


  buf
  g1042
  (
    n1040,
    n1020
  );


  buf
  g1043
  (
    n1083,
    n1032
  );


  buf
  g1044
  (
    n1047,
    n992
  );


  buf
  g1045
  (
    n1120,
    n1008
  );


  not
  g1046
  (
    n1076,
    n1024
  );


  buf
  g1047
  (
    n1075,
    n1007
  );


  not
  g1048
  (
    n1128,
    n990
  );


  not
  g1049
  (
    n1112,
    n987
  );


  not
  g1050
  (
    n1090,
    n1028
  );


  not
  g1051
  (
    n1074,
    n1027
  );


  not
  g1052
  (
    n1147,
    n1012
  );


  buf
  g1053
  (
    n1095,
    n1021
  );


  buf
  g1054
  (
    n1160,
    n1033
  );


  not
  g1055
  (
    n1062,
    n990
  );


  buf
  g1056
  (
    n1157,
    n989
  );


  not
  g1057
  (
    n1082,
    n985
  );


  not
  g1058
  (
    n1124,
    n1018
  );


  not
  g1059
  (
    n1167,
    n1031
  );


  not
  g1060
  (
    n1065,
    n1036
  );


  buf
  g1061
  (
    n1060,
    n735
  );


  not
  g1062
  (
    n1162,
    n1011
  );


  not
  g1063
  (
    n1143,
    n986
  );


  buf
  g1064
  (
    n1133,
    n1020
  );


  buf
  g1065
  (
    n1101,
    n974
  );


  not
  g1066
  (
    n1127,
    n990
  );


  buf
  g1067
  (
    n1089,
    n1018
  );


  not
  g1068
  (
    n1166,
    n1029
  );


  buf
  g1069
  (
    n1092,
    n982
  );


  buf
  g1070
  (
    n1066,
    n742
  );


  buf
  g1071
  (
    n1108,
    n971
  );


  not
  g1072
  (
    n1044,
    n988
  );


  buf
  g1073
  (
    n1078,
    n975
  );


  not
  g1074
  (
    n1156,
    n985
  );


  not
  g1075
  (
    n1154,
    n1004
  );


  not
  g1076
  (
    n1086,
    n972
  );


  not
  g1077
  (
    n1080,
    n987
  );


  buf
  g1078
  (
    n1132,
    n974
  );


  not
  g1079
  (
    n1057,
    n983
  );


  buf
  g1080
  (
    n1161,
    n1015
  );


  not
  g1081
  (
    n1094,
    n987
  );


  buf
  g1082
  (
    n1158,
    n1006
  );


  not
  g1083
  (
    n1146,
    n978
  );


  not
  g1084
  (
    n1087,
    n971
  );


  buf
  g1085
  (
    n1138,
    n1008
  );


  not
  g1086
  (
    n1126,
    n1007
  );


  not
  g1087
  (
    n1045,
    n989
  );


  buf
  g1088
  (
    n1139,
    n1019
  );


  buf
  g1089
  (
    n1071,
    n1035
  );


  buf
  g1090
  (
    n1039,
    n972
  );


  buf
  g1091
  (
    n1059,
    n984
  );


  buf
  g1092
  (
    n1046,
    n1033
  );


  buf
  g1093
  (
    n1114,
    n971
  );


  not
  g1094
  (
    n1116,
    n1026
  );


  buf
  g1095
  (
    n1155,
    n1035
  );


  not
  g1096
  (
    n1054,
    n740
  );


  not
  g1097
  (
    n1148,
    n984
  );


  not
  g1098
  (
    n1042,
    n983
  );


  buf
  g1099
  (
    n1122,
    n988
  );


  not
  g1100
  (
    n1118,
    n1032
  );


  not
  g1101
  (
    n1137,
    n974
  );


  buf
  g1102
  (
    n1119,
    n981
  );


  buf
  g1103
  (
    n1100,
    n741
  );


  nand
  g1104
  (
    n1123,
    n1028,
    n1022,
    n1031,
    n985
  );


  xnor
  g1105
  (
    n1043,
    n1023,
    n1014,
    n1013
  );


  or
  g1106
  (
    n1152,
    n1010,
    n1005,
    n1034,
    n738
  );


  or
  g1107
  (
    n1109,
    n1028,
    n992,
    n1012,
    n989
  );


  or
  g1108
  (
    n1058,
    n1036,
    n1030,
    n993,
    n1025
  );


  and
  g1109
  (
    n1134,
    n1030,
    n1023,
    n1010,
    n736
  );


  xor
  g1110
  (
    n1048,
    n983,
    n1028,
    n975,
    n1027
  );


  xnor
  g1111
  (
    n1141,
    n971,
    n1015,
    n977,
    n1023
  );


  xnor
  g1112
  (
    n1056,
    n986,
    n991,
    n973,
    n1007
  );


  and
  g1113
  (
    n1099,
    n1009,
    n1032,
    n981,
    n1016
  );


  nor
  g1114
  (
    n1115,
    n975,
    n1030,
    n1022,
    n982
  );


  nor
  g1115
  (
    n1111,
    n1034,
    n1016,
    n1006,
    n1007
  );


  nand
  g1116
  (
    n1072,
    n975,
    n994,
    n1009,
    n977
  );


  xnor
  g1117
  (
    n1061,
    n1021,
    n970,
    n1027,
    n1015
  );


  or
  g1118
  (
    n1150,
    n978,
    n1035,
    n983,
    n994
  );


  or
  g1119
  (
    n1049,
    n994,
    n993,
    n1021,
    n988
  );


  or
  g1120
  (
    n1084,
    n973,
    n1009,
    n1025,
    n1030
  );


  nand
  g1121
  (
    n1051,
    n984,
    n739,
    n1026,
    n990
  );


  xnor
  g1122
  (
    n1088,
    n1029,
    n1034,
    n1024
  );


  or
  g1123
  (
    n1107,
    n973,
    n993,
    n1010,
    n994
  );


  xor
  g1124
  (
    n1070,
    n976,
    n1019,
    n1012,
    n986
  );


  or
  g1125
  (
    n1077,
    n1004,
    n978,
    n1009,
    n1011
  );


  or
  g1126
  (
    n1068,
    n1017,
    n1022,
    n992,
    n1026
  );


  nand
  g1127
  (
    n1073,
    n1017,
    n1022,
    n1006,
    n986
  );


  xor
  g1128
  (
    n1159,
    n1013,
    n976,
    n737,
    n1006
  );


  nand
  g1129
  (
    n1129,
    n1035,
    n987,
    n972,
    n977
  );


  nand
  g1130
  (
    n1093,
    n978,
    n1032,
    n1027,
    n977
  );


  nor
  g1131
  (
    n1142,
    n989,
    n1029,
    n1031,
    n991
  );


  xnor
  g1132
  (
    n1091,
    n993,
    n1004,
    n1013
  );


  nand
  g1133
  (
    n1050,
    n1031,
    n982,
    n1020,
    n1019
  );


  or
  g1134
  (
    n1052,
    n1033,
    n1016,
    n991,
    n973
  );


  xor
  g1135
  (
    n1069,
    n1023,
    n1018,
    n1020,
    n1010
  );


  buf
  g1136
  (
    n1375,
    n1080
  );


  buf
  g1137
  (
    n1604,
    n1084
  );


  buf
  g1138
  (
    n1228,
    n1058
  );


  buf
  g1139
  (
    n1210,
    n1098
  );


  buf
  g1140
  (
    n1374,
    n1073
  );


  buf
  g1141
  (
    n1288,
    n1072
  );


  not
  g1142
  (
    n1420,
    n1110
  );


  buf
  g1143
  (
    n1551,
    n1155
  );


  not
  g1144
  (
    n1337,
    n1154
  );


  not
  g1145
  (
    n1538,
    n1133
  );


  buf
  g1146
  (
    n1359,
    n1052
  );


  buf
  g1147
  (
    n1186,
    n1166
  );


  not
  g1148
  (
    n1506,
    n1129
  );


  not
  g1149
  (
    n1434,
    n1079
  );


  not
  g1150
  (
    n1302,
    n1144
  );


  not
  g1151
  (
    n1250,
    n1120
  );


  buf
  g1152
  (
    n1325,
    n1095
  );


  buf
  g1153
  (
    n1297,
    n1130
  );


  not
  g1154
  (
    n1172,
    n1064
  );


  buf
  g1155
  (
    n1642,
    n1084
  );


  buf
  g1156
  (
    n1358,
    n1097
  );


  buf
  g1157
  (
    n1317,
    n1111
  );


  not
  g1158
  (
    n1328,
    n1052
  );


  buf
  g1159
  (
    n1666,
    n1085
  );


  not
  g1160
  (
    n1266,
    n1086
  );


  buf
  g1161
  (
    n1242,
    n1056
  );


  not
  g1162
  (
    n1380,
    n1120
  );


  buf
  g1163
  (
    n1277,
    n1076
  );


  not
  g1164
  (
    n1182,
    n1101
  );


  buf
  g1165
  (
    n1430,
    n1078
  );


  buf
  g1166
  (
    n1361,
    n1102
  );


  buf
  g1167
  (
    n1458,
    n1156
  );


  not
  g1168
  (
    n1413,
    n1128
  );


  buf
  g1169
  (
    n1638,
    n1094
  );


  buf
  g1170
  (
    n1577,
    n1137
  );


  buf
  g1171
  (
    n1282,
    n1090
  );


  buf
  g1172
  (
    n1540,
    n1061
  );


  buf
  g1173
  (
    n1402,
    n1057
  );


  buf
  g1174
  (
    n1294,
    n1127
  );


  buf
  g1175
  (
    n1527,
    n1082
  );


  not
  g1176
  (
    n1450,
    n1090
  );


  not
  g1177
  (
    n1425,
    n1087
  );


  buf
  g1178
  (
    n1409,
    n1094
  );


  buf
  g1179
  (
    n1646,
    n1117
  );


  buf
  g1180
  (
    n1481,
    n1142
  );


  buf
  g1181
  (
    n1447,
    n1105
  );


  not
  g1182
  (
    n1292,
    n1105
  );


  buf
  g1183
  (
    n1227,
    n1088
  );


  buf
  g1184
  (
    n1314,
    n1068
  );


  not
  g1185
  (
    n1239,
    n1099
  );


  not
  g1186
  (
    n1568,
    n1107
  );


  not
  g1187
  (
    n1443,
    n1104
  );


  not
  g1188
  (
    n1201,
    n1159
  );


  not
  g1189
  (
    n1609,
    n1089
  );


  not
  g1190
  (
    n1483,
    n1041
  );


  buf
  g1191
  (
    n1246,
    n1093
  );


  buf
  g1192
  (
    n1468,
    n1109
  );


  buf
  g1193
  (
    n1644,
    n1153
  );


  buf
  g1194
  (
    n1581,
    n1077
  );


  buf
  g1195
  (
    n1170,
    n1060
  );


  not
  g1196
  (
    n1514,
    n1138
  );


  buf
  g1197
  (
    n1377,
    n1073
  );


  buf
  g1198
  (
    n1441,
    n1049
  );


  not
  g1199
  (
    n1368,
    n1167
  );


  buf
  g1200
  (
    n1179,
    n1059
  );


  not
  g1201
  (
    n1629,
    n1149
  );


  not
  g1202
  (
    n1332,
    n1061
  );


  not
  g1203
  (
    n1516,
    n1075
  );


  not
  g1204
  (
    n1575,
    n1048
  );


  buf
  g1205
  (
    n1321,
    n1121
  );


  buf
  g1206
  (
    n1622,
    n1115
  );


  buf
  g1207
  (
    n1196,
    n1137
  );


  buf
  g1208
  (
    n1519,
    n1045
  );


  not
  g1209
  (
    n1549,
    n1054
  );


  buf
  g1210
  (
    n1611,
    n1111
  );


  not
  g1211
  (
    n1659,
    n1071
  );


  not
  g1212
  (
    n1370,
    n1066
  );


  not
  g1213
  (
    n1534,
    n1162
  );


  buf
  g1214
  (
    n1176,
    n1132
  );


  buf
  g1215
  (
    n1449,
    n1063
  );


  not
  g1216
  (
    n1346,
    n1065
  );


  buf
  g1217
  (
    n1316,
    n1163
  );


  not
  g1218
  (
    n1469,
    n1095
  );


  buf
  g1219
  (
    n1618,
    n1135
  );


  buf
  g1220
  (
    n1555,
    n1078
  );


  buf
  g1221
  (
    n1379,
    n1142
  );


  buf
  g1222
  (
    n1561,
    n1109
  );


  not
  g1223
  (
    n1268,
    n1148
  );


  not
  g1224
  (
    n1645,
    n1105
  );


  buf
  g1225
  (
    n1407,
    n1138
  );


  buf
  g1226
  (
    n1560,
    n1137
  );


  buf
  g1227
  (
    n1471,
    n1118
  );


  buf
  g1228
  (
    n1207,
    n1072
  );


  buf
  g1229
  (
    n1499,
    n1069
  );


  not
  g1230
  (
    n1366,
    n1124
  );


  buf
  g1231
  (
    n1605,
    n1139
  );


  buf
  g1232
  (
    n1442,
    n1099
  );


  not
  g1233
  (
    n1329,
    n1064
  );


  buf
  g1234
  (
    n1405,
    n1101
  );


  buf
  g1235
  (
    n1218,
    n1157
  );


  not
  g1236
  (
    n1465,
    n1141
  );


  not
  g1237
  (
    n1486,
    n1052
  );


  not
  g1238
  (
    n1427,
    n1116
  );


  buf
  g1239
  (
    n1665,
    n1114
  );


  buf
  g1240
  (
    n1459,
    n1167
  );


  buf
  g1241
  (
    n1464,
    n1097
  );


  not
  g1242
  (
    n1304,
    n1167
  );


  buf
  g1243
  (
    n1237,
    n1155
  );


  not
  g1244
  (
    n1640,
    n1073
  );


  buf
  g1245
  (
    n1617,
    n1138
  );


  buf
  g1246
  (
    n1383,
    n1082
  );


  not
  g1247
  (
    n1270,
    n1067
  );


  buf
  g1248
  (
    n1215,
    n1098
  );


  buf
  g1249
  (
    n1670,
    n1059
  );


  not
  g1250
  (
    n1570,
    n1049
  );


  not
  g1251
  (
    n1523,
    n1141
  );


  not
  g1252
  (
    n1320,
    n1163
  );


  not
  g1253
  (
    n1515,
    n1054
  );


  buf
  g1254
  (
    n1342,
    n1159
  );


  buf
  g1255
  (
    n1290,
    n1076
  );


  buf
  g1256
  (
    n1654,
    n1050
  );


  buf
  g1257
  (
    n1580,
    n1108
  );


  not
  g1258
  (
    n1457,
    n1118
  );


  not
  g1259
  (
    n1336,
    n1166
  );


  buf
  g1260
  (
    n1276,
    n1065
  );


  buf
  g1261
  (
    n1511,
    n1057
  );


  not
  g1262
  (
    n1259,
    n1162
  );


  buf
  g1263
  (
    n1590,
    n1054
  );


  not
  g1264
  (
    n1295,
    n1146
  );


  buf
  g1265
  (
    n1508,
    n1075
  );


  not
  g1266
  (
    n1626,
    n1116
  );


  not
  g1267
  (
    n1663,
    n1165
  );


  buf
  g1268
  (
    n1510,
    n1147
  );


  not
  g1269
  (
    n1403,
    n1062
  );


  buf
  g1270
  (
    n1344,
    n1050
  );


  not
  g1271
  (
    n1574,
    n1146
  );


  not
  g1272
  (
    n1619,
    n1061
  );


  buf
  g1273
  (
    n1197,
    n1103
  );


  not
  g1274
  (
    n1429,
    n1112
  );


  buf
  g1275
  (
    n1394,
    n1100
  );


  not
  g1276
  (
    n1621,
    n1154
  );


  buf
  g1277
  (
    n1661,
    n1119
  );


  buf
  g1278
  (
    n1173,
    n1141
  );


  not
  g1279
  (
    n1236,
    n1163
  );


  not
  g1280
  (
    n1298,
    n1087
  );


  buf
  g1281
  (
    n1253,
    n1048
  );


  not
  g1282
  (
    n1355,
    n1103
  );


  not
  g1283
  (
    n1426,
    n1067
  );


  not
  g1284
  (
    n1365,
    n1127
  );


  buf
  g1285
  (
    n1264,
    n1132
  );


  not
  g1286
  (
    n1198,
    n1145
  );


  not
  g1287
  (
    n1222,
    n1088
  );


  not
  g1288
  (
    n1423,
    n1163
  );


  buf
  g1289
  (
    n1669,
    n1101
  );


  buf
  g1290
  (
    n1520,
    n1131
  );


  not
  g1291
  (
    n1556,
    n1168
  );


  buf
  g1292
  (
    n1299,
    n1051
  );


  buf
  g1293
  (
    n1616,
    n1158
  );


  buf
  g1294
  (
    n1194,
    n1156
  );


  not
  g1295
  (
    n1440,
    n1110
  );


  not
  g1296
  (
    n1362,
    n1115
  );


  buf
  g1297
  (
    n1428,
    n1056
  );


  not
  g1298
  (
    n1562,
    n1159
  );


  not
  g1299
  (
    n1334,
    n1144
  );


  not
  g1300
  (
    n1489,
    n1100
  );


  not
  g1301
  (
    n1477,
    n1060
  );


  not
  g1302
  (
    n1241,
    n1166
  );


  buf
  g1303
  (
    n1456,
    n1070
  );


  not
  g1304
  (
    n1591,
    n1143
  );


  not
  g1305
  (
    n1279,
    n1086
  );


  buf
  g1306
  (
    n1630,
    n1132
  );


  not
  g1307
  (
    n1492,
    n1070
  );


  buf
  g1308
  (
    n1573,
    n1076
  );


  buf
  g1309
  (
    n1401,
    n1153
  );


  not
  g1310
  (
    n1658,
    n1117
  );


  buf
  g1311
  (
    n1649,
    n1069
  );


  buf
  g1312
  (
    n1522,
    n1058
  );


  buf
  g1313
  (
    n1204,
    n1096
  );


  not
  g1314
  (
    n1262,
    n1053
  );


  buf
  g1315
  (
    n1598,
    n1061
  );


  buf
  g1316
  (
    n1478,
    n1125
  );


  not
  g1317
  (
    n1498,
    n1059
  );


  buf
  g1318
  (
    n1437,
    n1158
  );


  not
  g1319
  (
    n1559,
    n1139
  );


  buf
  g1320
  (
    n1352,
    n1083
  );


  not
  g1321
  (
    n1491,
    n1064
  );


  buf
  g1322
  (
    n1582,
    n1057
  );


  not
  g1323
  (
    n1391,
    n1100
  );


  not
  g1324
  (
    n1267,
    n1055
  );


  not
  g1325
  (
    n1613,
    n1091
  );


  not
  g1326
  (
    n1461,
    n1164
  );


  buf
  g1327
  (
    n1417,
    n1126
  );


  buf
  g1328
  (
    n1623,
    n1151
  );


  buf
  g1329
  (
    n1552,
    n1068
  );


  buf
  g1330
  (
    n1341,
    n1131
  );


  not
  g1331
  (
    n1526,
    n1046
  );


  buf
  g1332
  (
    n1312,
    n1094
  );


  buf
  g1333
  (
    n1300,
    n1140
  );


  buf
  g1334
  (
    n1550,
    n1160
  );


  not
  g1335
  (
    n1376,
    n1050
  );


  not
  g1336
  (
    n1482,
    n1047
  );


  not
  g1337
  (
    n1301,
    n1072
  );


  not
  g1338
  (
    n1502,
    n1155
  );


  not
  g1339
  (
    n1184,
    n1066
  );


  buf
  g1340
  (
    n1202,
    n1149
  );


  buf
  g1341
  (
    n1180,
    n1099
  );


  buf
  g1342
  (
    n1495,
    n1143
  );


  buf
  g1343
  (
    n1205,
    n1122
  );


  buf
  g1344
  (
    n1479,
    n1106
  );


  buf
  g1345
  (
    n1517,
    n1096
  );


  buf
  g1346
  (
    n1233,
    n1149
  );


  buf
  g1347
  (
    n1177,
    n1142
  );


  not
  g1348
  (
    n1372,
    n1164
  );


  buf
  g1349
  (
    n1356,
    n1103
  );


  buf
  g1350
  (
    n1291,
    n1112
  );


  not
  g1351
  (
    n1397,
    n1085
  );


  not
  g1352
  (
    n1521,
    n1079
  );


  not
  g1353
  (
    n1615,
    n1113
  );


  buf
  g1354
  (
    n1608,
    n1081
  );


  buf
  g1355
  (
    n1306,
    n1125
  );


  not
  g1356
  (
    n1569,
    n1040
  );


  not
  g1357
  (
    n1271,
    n1057
  );


  buf
  g1358
  (
    n1548,
    n1168
  );


  buf
  g1359
  (
    n1281,
    n1078
  );


  buf
  g1360
  (
    n1283,
    n1138
  );


  not
  g1361
  (
    n1333,
    n1047
  );


  buf
  g1362
  (
    n1251,
    n1081
  );


  not
  g1363
  (
    n1178,
    n1109
  );


  not
  g1364
  (
    n1221,
    n1134
  );


  buf
  g1365
  (
    n1488,
    n1052
  );


  buf
  g1366
  (
    n1566,
    n1102
  );


  not
  g1367
  (
    n1331,
    n1166
  );


  buf
  g1368
  (
    n1354,
    n1147
  );


  not
  g1369
  (
    n1505,
    n1069
  );


  not
  g1370
  (
    n1214,
    n1131
  );


  not
  g1371
  (
    n1234,
    n1081
  );


  buf
  g1372
  (
    n1466,
    n1108
  );


  buf
  g1373
  (
    n1351,
    n1105
  );


  buf
  g1374
  (
    n1200,
    n1140
  );


  not
  g1375
  (
    n1545,
    n1079
  );


  not
  g1376
  (
    n1399,
    n1125
  );


  not
  g1377
  (
    n1596,
    n1098
  );


  not
  g1378
  (
    n1470,
    n1076
  );


  not
  g1379
  (
    n1480,
    n1134
  );


  buf
  g1380
  (
    n1289,
    n1104
  );


  buf
  g1381
  (
    n1188,
    n1160
  );


  buf
  g1382
  (
    n1187,
    n1077
  );


  not
  g1383
  (
    n1432,
    n1120
  );


  buf
  g1384
  (
    n1597,
    n1093
  );


  not
  g1385
  (
    n1650,
    n1069
  );


  buf
  g1386
  (
    n1530,
    n1070
  );


  buf
  g1387
  (
    n1175,
    n1162
  );


  buf
  g1388
  (
    n1503,
    n1088
  );


  not
  g1389
  (
    n1436,
    n1123
  );


  buf
  g1390
  (
    n1185,
    n1113
  );


  not
  g1391
  (
    n1633,
    n1092
  );


  buf
  g1392
  (
    n1199,
    n1114
  );


  not
  g1393
  (
    n1627,
    n1045
  );


  buf
  g1394
  (
    n1261,
    n1059
  );


  not
  g1395
  (
    n1607,
    n1111
  );


  buf
  g1396
  (
    n1558,
    n1091
  );


  buf
  g1397
  (
    n1586,
    n1127
  );


  not
  g1398
  (
    n1238,
    n1153
  );


  buf
  g1399
  (
    n1330,
    n1046
  );


  not
  g1400
  (
    n1315,
    n1127
  );


  not
  g1401
  (
    n1347,
    n1168
  );


  not
  g1402
  (
    n1260,
    n1082
  );


  buf
  g1403
  (
    n1369,
    n1055
  );


  buf
  g1404
  (
    n1232,
    n1074
  );


  not
  g1405
  (
    n1224,
    n1060
  );


  not
  g1406
  (
    n1311,
    n1111
  );


  buf
  g1407
  (
    n1191,
    n1062
  );


  buf
  g1408
  (
    n1373,
    n1092
  );


  not
  g1409
  (
    n1579,
    n1150
  );


  not
  g1410
  (
    n1664,
    n1165
  );


  not
  g1411
  (
    n1263,
    n1084
  );


  buf
  g1412
  (
    n1509,
    n1154
  );


  buf
  g1413
  (
    n1169,
    n1113
  );


  not
  g1414
  (
    n1257,
    n1143
  );


  not
  g1415
  (
    n1529,
    n1146
  );


  not
  g1416
  (
    n1512,
    n1151
  );


  buf
  g1417
  (
    n1418,
    n1165
  );


  buf
  g1418
  (
    n1648,
    n1128
  );


  buf
  g1419
  (
    n1431,
    n1091
  );


  buf
  g1420
  (
    n1193,
    n1106
  );


  not
  g1421
  (
    n1606,
    n1121
  );


  not
  g1422
  (
    n1252,
    n1097
  );


  not
  g1423
  (
    n1229,
    n1083
  );


  not
  g1424
  (
    n1406,
    n1046
  );


  not
  g1425
  (
    n1213,
    n1102
  );


  not
  g1426
  (
    n1274,
    n1095
  );


  not
  g1427
  (
    n1319,
    n1140
  );


  not
  g1428
  (
    n1285,
    n1106
  );


  not
  g1429
  (
    n1657,
    n1046
  );


  buf
  g1430
  (
    n1455,
    n1054
  );


  not
  g1431
  (
    n1392,
    n1051
  );


  not
  g1432
  (
    n1497,
    n1160
  );


  buf
  g1433
  (
    n1243,
    n1152
  );


  not
  g1434
  (
    n1303,
    n1123
  );


  buf
  g1435
  (
    n1594,
    n1067
  );


  buf
  g1436
  (
    n1553,
    n1102
  );


  not
  g1437
  (
    n1585,
    n1047
  );


  not
  g1438
  (
    n1554,
    n1161
  );


  not
  g1439
  (
    n1371,
    n1086
  );


  buf
  g1440
  (
    n1453,
    n1120
  );


  not
  g1441
  (
    n1208,
    n1128
  );


  not
  g1442
  (
    n1542,
    n1139
  );


  not
  g1443
  (
    n1181,
    n1072
  );


  not
  g1444
  (
    n1338,
    n1129
  );


  not
  g1445
  (
    n1536,
    n1075
  );


  not
  g1446
  (
    n1416,
    n1077
  );


  buf
  g1447
  (
    n1357,
    n1071
  );


  buf
  g1448
  (
    n1335,
    n1049
  );


  buf
  g1449
  (
    n1564,
    n1136
  );


  not
  g1450
  (
    n1452,
    n1142
  );


  not
  g1451
  (
    n1254,
    n1130
  );


  buf
  g1452
  (
    n1614,
    n1151
  );


  buf
  g1453
  (
    n1513,
    n1093
  );


  not
  g1454
  (
    n1326,
    n1129
  );


  buf
  g1455
  (
    n1602,
    n1074
  );


  not
  g1456
  (
    n1367,
    n1143
  );


  buf
  g1457
  (
    n1415,
    n1089
  );


  not
  g1458
  (
    n1635,
    n1080
  );


  not
  g1459
  (
    n1398,
    n1087
  );


  buf
  g1460
  (
    n1547,
    n1118
  );


  not
  g1461
  (
    n1286,
    n1150
  );


  not
  g1462
  (
    n1410,
    n1145
  );


  buf
  g1463
  (
    n1313,
    n1051
  );


  buf
  g1464
  (
    n1668,
    n1083
  );


  not
  g1465
  (
    n1433,
    n1161
  );


  not
  g1466
  (
    n1472,
    n1108
  );


  not
  g1467
  (
    n1445,
    n1161
  );


  buf
  g1468
  (
    n1340,
    n1107
  );


  buf
  g1469
  (
    n1305,
    n1093
  );


  not
  g1470
  (
    n1390,
    n1146
  );


  not
  g1471
  (
    n1240,
    n1104
  );


  buf
  g1472
  (
    n1275,
    n1051
  );


  not
  g1473
  (
    n1601,
    n1097
  );


  buf
  g1474
  (
    n1610,
    n1055
  );


  buf
  g1475
  (
    n1572,
    n1065
  );


  not
  g1476
  (
    n1475,
    n1136
  );


  buf
  g1477
  (
    n1400,
    n1085
  );


  not
  g1478
  (
    n1595,
    n1122
  );


  not
  g1479
  (
    n1223,
    n1063
  );


  not
  g1480
  (
    n1424,
    n1152
  );


  buf
  g1481
  (
    n1652,
    n1117
  );


  buf
  g1482
  (
    n1183,
    n1048
  );


  not
  g1483
  (
    n1421,
    n1100
  );


  not
  g1484
  (
    n1600,
    n1152
  );


  not
  g1485
  (
    n1226,
    n1066
  );


  not
  g1486
  (
    n1386,
    n1117
  );


  not
  g1487
  (
    n1565,
    n1092
  );


  not
  g1488
  (
    n1284,
    n1068
  );


  not
  g1489
  (
    n1280,
    n1083
  );


  not
  g1490
  (
    n1339,
    n1085
  );


  buf
  g1491
  (
    n1235,
    n1140
  );


  not
  g1492
  (
    n1592,
    n1119
  );


  not
  g1493
  (
    n1322,
    n1106
  );


  not
  g1494
  (
    n1360,
    n1058
  );


  buf
  g1495
  (
    n1576,
    n1091
  );


  not
  g1496
  (
    n1190,
    n1132
  );


  buf
  g1497
  (
    n1220,
    n1078
  );


  buf
  g1498
  (
    n1324,
    n1109
  );


  buf
  g1499
  (
    n1209,
    n1079
  );


  buf
  g1500
  (
    n1255,
    n1095
  );


  buf
  g1501
  (
    n1533,
    n1157
  );


  buf
  g1502
  (
    n1454,
    n1152
  );


  not
  g1503
  (
    n1381,
    n1101
  );


  not
  g1504
  (
    n1544,
    n1144
  );


  not
  g1505
  (
    n1460,
    n1047
  );


  not
  g1506
  (
    n1206,
    n1062
  );


  buf
  g1507
  (
    n1620,
    n1112
  );


  not
  g1508
  (
    n1578,
    n1116
  );


  buf
  g1509
  (
    n1171,
    n1124
  );


  not
  g1510
  (
    n1230,
    n1044
  );


  not
  g1511
  (
    n1448,
    n1141
  );


  buf
  g1512
  (
    n1451,
    n1135
  );


  not
  g1513
  (
    n1612,
    n1129
  );


  not
  g1514
  (
    n1189,
    n1133
  );


  not
  g1515
  (
    n1435,
    n1049
  );


  not
  g1516
  (
    n1219,
    n1065
  );


  not
  g1517
  (
    n1484,
    n1045
  );


  not
  g1518
  (
    n1388,
    n1053
  );


  buf
  g1519
  (
    n1414,
    n1124
  );


  not
  g1520
  (
    n1563,
    n1154
  );


  buf
  g1521
  (
    n1310,
    n1124
  );


  not
  g1522
  (
    n1588,
    n1089
  );


  not
  g1523
  (
    n1396,
    n1089
  );


  not
  g1524
  (
    n1382,
    n1165
  );


  buf
  g1525
  (
    n1203,
    n1133
  );


  not
  g1526
  (
    n1628,
    n1071
  );


  not
  g1527
  (
    n1496,
    n1103
  );


  not
  g1528
  (
    n1216,
    n1148
  );


  buf
  g1529
  (
    n1217,
    n1162
  );


  buf
  g1530
  (
    n1174,
    n1126
  );


  not
  g1531
  (
    n1593,
    n1096
  );


  not
  g1532
  (
    n1363,
    n1121
  );


  not
  g1533
  (
    n1287,
    n1118
  );


  buf
  g1534
  (
    n1389,
    n1159
  );


  buf
  g1535
  (
    n1422,
    n1060
  );


  not
  g1536
  (
    n1660,
    n1039
  );


  buf
  g1537
  (
    n1395,
    n1156
  );


  not
  g1538
  (
    n1273,
    n1148
  );


  not
  g1539
  (
    n1364,
    n1050
  );


  not
  g1540
  (
    n1528,
    n1115
  );


  buf
  g1541
  (
    n1476,
    n1096
  );


  not
  g1542
  (
    n1444,
    n1055
  );


  not
  g1543
  (
    n1518,
    n1080
  );


  not
  g1544
  (
    n1539,
    n1080
  );


  not
  g1545
  (
    n1408,
    n1107
  );


  not
  g1546
  (
    n1631,
    n1075
  );


  not
  g1547
  (
    n1535,
    n1168
  );


  buf
  g1548
  (
    n1247,
    n1149
  );


  buf
  g1549
  (
    n1632,
    n1164
  );


  not
  g1550
  (
    n1393,
    n1160
  );


  buf
  g1551
  (
    n1353,
    n1133
  );


  buf
  g1552
  (
    n1571,
    n1123
  );


  buf
  g1553
  (
    n1531,
    n1156
  );


  buf
  g1554
  (
    n1599,
    n1158
  );


  not
  g1555
  (
    n1462,
    n1150
  );


  buf
  g1556
  (
    n1524,
    n1094
  );


  not
  g1557
  (
    n1308,
    n1112
  );


  not
  g1558
  (
    n1473,
    n1064
  );


  buf
  g1559
  (
    n1525,
    n1070
  );


  buf
  g1560
  (
    n1537,
    n1110
  );


  not
  g1561
  (
    n1584,
    n1045
  );


  buf
  g1562
  (
    n1411,
    n1136
  );


  not
  g1563
  (
    n1504,
    n1135
  );


  not
  g1564
  (
    n1557,
    n1048
  );


  buf
  g1565
  (
    n1463,
    n1161
  );


  buf
  g1566
  (
    n1662,
    n1121
  );


  not
  g1567
  (
    n1378,
    n1114
  );


  buf
  g1568
  (
    n1494,
    n1153
  );


  buf
  g1569
  (
    n1643,
    n1150
  );


  buf
  g1570
  (
    n1412,
    n1056
  );


  not
  g1571
  (
    n1192,
    n1092
  );


  buf
  g1572
  (
    n1636,
    n1116
  );


  not
  g1573
  (
    n1485,
    n1088
  );


  buf
  g1574
  (
    n1248,
    n1148
  );


  buf
  g1575
  (
    n1384,
    n1073
  );


  buf
  g1576
  (
    n1487,
    n1134
  );


  not
  g1577
  (
    n1634,
    n1151
  );


  not
  g1578
  (
    n1500,
    n1126
  );


  buf
  g1579
  (
    n1256,
    n1115
  );


  buf
  g1580
  (
    n1493,
    n1067
  );


  buf
  g1581
  (
    n1350,
    n1119
  );


  not
  g1582
  (
    n1467,
    n1066
  );


  not
  g1583
  (
    n1318,
    n1134
  );


  not
  g1584
  (
    n1307,
    n1098
  );


  not
  g1585
  (
    n1269,
    n1086
  );


  not
  g1586
  (
    n1439,
    n1107
  );


  not
  g1587
  (
    n1507,
    n1058
  );


  buf
  g1588
  (
    n1474,
    n1145
  );


  buf
  g1589
  (
    n1587,
    n1157
  );


  buf
  g1590
  (
    n1446,
    n1082
  );


  not
  g1591
  (
    n1589,
    n1126
  );


  buf
  g1592
  (
    n1349,
    n1144
  );


  buf
  g1593
  (
    n1385,
    n1130
  );


  not
  g1594
  (
    n1501,
    n1164
  );


  buf
  g1595
  (
    n1387,
    n1063
  );


  buf
  g1596
  (
    n1323,
    n1167
  );


  not
  g1597
  (
    n1272,
    n1128
  );


  not
  g1598
  (
    n1245,
    n1063
  );


  not
  g1599
  (
    n1231,
    n1155
  );


  buf
  g1600
  (
    n1212,
    n1053
  );


  not
  g1601
  (
    n1309,
    n1056
  );


  buf
  g1602
  (
    n1655,
    n1136
  );


  buf
  g1603
  (
    n1348,
    n1099
  );


  not
  g1604
  (
    n1603,
    n1071
  );


  not
  g1605
  (
    n1296,
    n1147
  );


  not
  g1606
  (
    n1546,
    n1122
  );


  not
  g1607
  (
    n1583,
    n1147
  );


  buf
  g1608
  (
    n1667,
    n1131
  );


  not
  g1609
  (
    n1653,
    n1077
  );


  buf
  g1610
  (
    n1244,
    n1125
  );


  buf
  g1611
  (
    n1211,
    n1119
  );


  buf
  g1612
  (
    n1624,
    n1114
  );


  not
  g1613
  (
    n1345,
    n1043
  );


  not
  g1614
  (
    n1543,
    n1074
  );


  not
  g1615
  (
    n1343,
    n1145
  );


  buf
  g1616
  (
    n1639,
    n1139
  );


  not
  g1617
  (
    n1225,
    n1123
  );


  buf
  g1618
  (
    n1249,
    n1108
  );


  buf
  g1619
  (
    n1532,
    n1081
  );


  not
  g1620
  (
    n1419,
    n1090
  );


  not
  g1621
  (
    n1651,
    n1130
  );


  not
  g1622
  (
    n1293,
    n1158
  );


  buf
  g1623
  (
    n1647,
    n1090
  );


  not
  g1624
  (
    n1490,
    n1122
  );


  buf
  g1625
  (
    n1567,
    n1084
  );


  buf
  g1626
  (
    n1656,
    n1087
  );


  buf
  g1627
  (
    n1541,
    n1137
  );


  not
  g1628
  (
    n1641,
    n1110
  );


  buf
  g1629
  (
    n1625,
    n1062
  );


  not
  g1630
  (
    n1278,
    n1135
  );


  not
  g1631
  (
    n1258,
    n1074
  );


  not
  g1632
  (
    n1404,
    n1104
  );


  buf
  g1633
  (
    n1637,
    n1068
  );


  not
  g1634
  (
    n1438,
    n1042
  );


  not
  g1635
  (
    n1265,
    n1053
  );


  buf
  g1636
  (
    n1195,
    n1157
  );


  not
  g1637
  (
    n1327,
    n1113
  );


  xnor
  g1638
  (
    n1812,
    n1321,
    n1625,
    n1338,
    n1605
  );


  or
  g1639
  (
    n1793,
    n1187,
    n1419,
    n1560,
    n1444
  );


  and
  g1640
  (
    n1843,
    n1519,
    n1214,
    n1638,
    n1185
  );


  nand
  g1641
  (
    n1695,
    n1282,
    n1357,
    n1193,
    n1489
  );


  xnor
  g1642
  (
    n1813,
    n1615,
    n1645,
    n1595,
    n1184
  );


  nor
  g1643
  (
    n1830,
    n1382,
    n1619,
    n1652,
    n744
  );


  nor
  g1644
  (
    n1679,
    n1619,
    n1322,
    n1281,
    n1336
  );


  nand
  g1645
  (
    n1691,
    n1618,
    n1649,
    n1591,
    n1653
  );


  nand
  g1646
  (
    n1766,
    n1548,
    n1614,
    n1388,
    n1300
  );


  xnor
  g1647
  (
    n1709,
    n1189,
    n1638,
    n1566,
    n1642
  );


  xor
  g1648
  (
    n1693,
    n1596,
    n1475,
    n1374,
    n1654
  );


  xor
  g1649
  (
    n1850,
    n1250,
    n1288,
    n1548,
    n1635
  );


  xnor
  g1650
  (
    n1784,
    n1223,
    n746,
    n1633,
    n1169
  );


  nand
  g1651
  (
    n1862,
    n1530,
    n1646,
    n1639,
    n1343
  );


  nand
  g1652
  (
    n1833,
    n1658,
    n1550,
    n1628,
    n1533
  );


  nand
  g1653
  (
    n1689,
    n1037,
    n1607,
    n1311,
    n1557
  );


  nand
  g1654
  (
    n1686,
    n1038,
    n1307,
    n1426,
    n1387
  );


  xnor
  g1655
  (
    n1780,
    n1594,
    n1624,
    n1317,
    n1205
  );


  nor
  g1656
  (
    n1682,
    n1629,
    n1588,
    n1461,
    n1263
  );


  nand
  g1657
  (
    n1826,
    n1592,
    n1456,
    n1261,
    n1637
  );


  nand
  g1658
  (
    n1825,
    n1645,
    n1518,
    n1637,
    n1333
  );


  xnor
  g1659
  (
    n1782,
    n1608,
    n1278,
    n1490,
    n1552
  );


  nand
  g1660
  (
    n1749,
    n1173,
    n1298,
    n1538,
    n1431
  );


  or
  g1661
  (
    n1823,
    n1597,
    n1593,
    n1460,
    n1621
  );


  or
  g1662
  (
    n1772,
    n1527,
    n1291,
    n1436,
    n1526
  );


  xor
  g1663
  (
    n1714,
    n1640,
    n1468,
    n745,
    n1651
  );


  or
  g1664
  (
    n1753,
    n1340,
    n1285,
    n1478,
    n1409
  );


  nand
  g1665
  (
    n1719,
    n1454,
    n1549,
    n1645,
    n1545
  );


  nor
  g1666
  (
    n1799,
    n1326,
    n1641,
    n1512,
    n1463
  );


  nand
  g1667
  (
    n1864,
    n1659,
    n1540,
    n1628,
    n1416
  );


  nor
  g1668
  (
    n1715,
    n1654,
    n1439,
    n1247,
    n1582
  );


  xnor
  g1669
  (
    n1839,
    n1498,
    n1610,
    n1412,
    n1628
  );


  nor
  g1670
  (
    n1809,
    n1599,
    n1547,
    n1462,
    n1414
  );


  or
  g1671
  (
    n1814,
    n1289,
    n1334,
    n1579,
    n1458
  );


  nand
  g1672
  (
    n1855,
    n1348,
    n1440,
    n1546,
    n1598
  );


  and
  g1673
  (
    n1685,
    n1481,
    n1443,
    n1590,
    n1551
  );


  xor
  g1674
  (
    n1761,
    n1541,
    n1350,
    n1636,
    n1232
  );


  nor
  g1675
  (
    n1744,
    n743,
    n1178,
    n1556,
    n1611
  );


  nand
  g1676
  (
    n1854,
    n1643,
    n1647,
    n1639,
    n1400
  );


  nor
  g1677
  (
    n1676,
    n1655,
    n1544,
    n1601,
    n1612
  );


  nand
  g1678
  (
    n1722,
    n1379,
    n1598,
    n1323,
    n1487
  );


  nand
  g1679
  (
    n1771,
    n1260,
    n1599,
    n1591,
    n1623
  );


  or
  g1680
  (
    n1853,
    n1432,
    n1547,
    n1203,
    n1249
  );


  xnor
  g1681
  (
    n1846,
    n1628,
    n1658,
    n1647,
    n1631
  );


  and
  g1682
  (
    n1705,
    n1597,
    n1198,
    n1643,
    n1639
  );


  nand
  g1683
  (
    n1795,
    n1530,
    n1656,
    n1483,
    n1546
  );


  or
  g1684
  (
    n1802,
    n1634,
    n1356,
    n1616,
    n1425
  );


  xnor
  g1685
  (
    n1747,
    n1467,
    n1308,
    n1351,
    n1315
  );


  and
  g1686
  (
    n1828,
    n1614,
    n923,
    n1435,
    n1283
  );


  and
  g1687
  (
    n1687,
    n1459,
    n1620,
    n1637,
    n1252
  );


  nor
  g1688
  (
    n1713,
    n1320,
    n1617,
    n1452,
    n1623
  );


  xor
  g1689
  (
    n1848,
    n1625,
    n1306,
    n1601,
    n1624
  );


  and
  g1690
  (
    n1821,
    n1274,
    n1597,
    n1502,
    n1313
  );


  nor
  g1691
  (
    n1698,
    n1208,
    n1640,
    n1473,
    n1592
  );


  nor
  g1692
  (
    n1765,
    n1469,
    n1255,
    n1500,
    n1622
  );


  and
  g1693
  (
    n1789,
    n1610,
    n1623,
    n1375,
    n1328
  );


  nand
  g1694
  (
    n1824,
    n1537,
    n1588,
    n1606,
    n1579
  );


  nand
  g1695
  (
    n1851,
    n1591,
    n1305,
    n1606,
    n1428
  );


  xnor
  g1696
  (
    n1840,
    n1272,
    n1531,
    n1618,
    n1399
  );


  nor
  g1697
  (
    n1841,
    n1441,
    n1449,
    n1557,
    n1275
  );


  xnor
  g1698
  (
    n1684,
    n1174,
    n1396,
    n1190,
    n1341
  );


  xnor
  g1699
  (
    n1739,
    n1609,
    n1606,
    n1420,
    n1230
  );


  nand
  g1700
  (
    n1738,
    n1559,
    n1429,
    n1638,
    n1488
  );


  and
  g1701
  (
    n1680,
    n1615,
    n1571,
    n1542,
    n1629
  );


  nand
  g1702
  (
    n1822,
    n1268,
    n1371,
    n1572,
    n1355
  );


  nand
  g1703
  (
    n1733,
    n1632,
    n1604,
    n1642,
    n1365
  );


  xor
  g1704
  (
    n1806,
    n1257,
    n1633,
    n1612,
    n1603
  );


  xor
  g1705
  (
    n1712,
    n1404,
    n1614,
    n1657,
    n1626
  );


  xnor
  g1706
  (
    n1807,
    n1267,
    n1202,
    n1614,
    n1625
  );


  xor
  g1707
  (
    n1838,
    n1318,
    n1514,
    n1329,
    n1634
  );


  xnor
  g1708
  (
    n1792,
    n1352,
    n1276,
    n1453,
    n1418
  );


  and
  g1709
  (
    n1718,
    n1319,
    n1037,
    n1309,
    n1197
  );


  nor
  g1710
  (
    n1819,
    n1624,
    n1604,
    n1601,
    n1620
  );


  xor
  g1711
  (
    n1723,
    n1622,
    n1474,
    n1568,
    n1476
  );


  xor
  g1712
  (
    n1767,
    n1517,
    n1516,
    n1242,
    n1535
  );


  xor
  g1713
  (
    n1844,
    n1389,
    n1573,
    n1180,
    n1537
  );


  xor
  g1714
  (
    n1865,
    n1240,
    n1633,
    n1605,
    n1589
  );


  nor
  g1715
  (
    n1743,
    n1601,
    n1542,
    n1645,
    n1195
  );


  and
  g1716
  (
    n1675,
    n1221,
    n1640,
    n1621,
    n1646
  );


  xnor
  g1717
  (
    n1758,
    n1484,
    n1538,
    n1556,
    n1592
  );


  xor
  g1718
  (
    n1731,
    n1301,
    n1575,
    n1646,
    n1337
  );


  xnor
  g1719
  (
    n1820,
    n1204,
    n1580,
    n1658,
    n1655
  );


  xnor
  g1720
  (
    n1694,
    n1385,
    n1638,
    n1277,
    n1570
  );


  nand
  g1721
  (
    n1811,
    n1657,
    n1621,
    n1558,
    n1644
  );


  and
  g1722
  (
    n1717,
    n1363,
    n1482,
    n1619,
    n1493
  );


  and
  g1723
  (
    n1788,
    n1568,
    n1631,
    n1181,
    n1632
  );


  xor
  g1724
  (
    n1835,
    n1550,
    n1621,
    n1238,
    n1211
  );


  and
  g1725
  (
    n1781,
    n1312,
    n1581,
    n1324,
    n1327
  );


  xor
  g1726
  (
    n1681,
    n1345,
    n1590,
    n1598,
    n1224
  );


  nor
  g1727
  (
    n1775,
    n1629,
    n1265,
    n1529,
    n1603
  );


  nand
  g1728
  (
    n1740,
    n1273,
    n1491,
    n1391,
    n1591
  );


  xnor
  g1729
  (
    n1783,
    n1616,
    n1610,
    n1602,
    n1434
  );


  xor
  g1730
  (
    n1674,
    n1347,
    n1567,
    n1640,
    n1605
  );


  nor
  g1731
  (
    n1827,
    n1386,
    n1636,
    n1609,
    n1495
  );


  nor
  g1732
  (
    n1863,
    n1201,
    n1511,
    n1534,
    n1647
  );


  or
  g1733
  (
    n1829,
    n1362,
    n1617,
    n1569,
    n1616
  );


  or
  g1734
  (
    n1735,
    n1219,
    n1569,
    n1594,
    n1633
  );


  xor
  g1735
  (
    n1764,
    n1403,
    n1616,
    n1421,
    n1587
  );


  and
  g1736
  (
    n1690,
    n1531,
    n1286,
    n1532,
    n1631
  );


  xnor
  g1737
  (
    n1673,
    n1643,
    n1523,
    n1600,
    n1394
  );


  xor
  g1738
  (
    n1734,
    n1652,
    n1369,
    n1636,
    n1611
  );


  and
  g1739
  (
    n1688,
    n1186,
    n1566,
    n1656,
    n1422
  );


  nand
  g1740
  (
    n1845,
    n1641,
    n1544,
    n1606,
    n1608
  );


  or
  g1741
  (
    n1831,
    n1634,
    n1217,
    n1188,
    n1038
  );


  or
  g1742
  (
    n1710,
    n1503,
    n1210,
    n1564,
    n1036
  );


  and
  g1743
  (
    n1836,
    n1373,
    n1648,
    n1536,
    n1587
  );


  or
  g1744
  (
    n1796,
    n1358,
    n1553,
    n1225,
    n1641
  );


  xnor
  g1745
  (
    n1726,
    n1236,
    n1402,
    n1280,
    n1528
  );


  xnor
  g1746
  (
    n1790,
    n1574,
    n1597,
    n1643,
    n1406
  );


  xor
  g1747
  (
    n1737,
    n1573,
    n1237,
    n1522,
    n1368
  );


  nor
  g1748
  (
    n1859,
    n1526,
    n1520,
    n1622,
    n1554
  );


  nand
  g1749
  (
    n1741,
    n1182,
    n1611,
    n1423,
    n1209
  );


  xor
  g1750
  (
    n1776,
    n1651,
    n1653,
    n1626,
    n1585
  );


  nand
  g1751
  (
    n1757,
    n1593,
    n1631,
    n1603,
    n1600
  );


  or
  g1752
  (
    n1701,
    n1200,
    n1648
  );


  and
  g1753
  (
    n1778,
    n1172,
    n1630,
    n1485,
    n1038
  );


  xor
  g1754
  (
    n1837,
    n1586,
    n1630,
    n1656,
    n1554
  );


  or
  g1755
  (
    n1770,
    n1576,
    n1589,
    n1433,
    n1408
  );


  or
  g1756
  (
    n1774,
    n1594,
    n1175,
    n1206,
    n1398
  );


  nor
  g1757
  (
    n1702,
    n749,
    n1215,
    n1596,
    n1342
  );


  or
  g1758
  (
    n1816,
    n1413,
    n1596,
    n1644,
    n1248
  );


  nor
  g1759
  (
    n1817,
    n1619,
    n1578,
    n1234,
    n1479
  );


  xnor
  g1760
  (
    n1834,
    n1494,
    n1228,
    n1625,
    n1360
  );


  or
  g1761
  (
    n1746,
    n1471,
    n1294,
    n1377,
    n1525
  );


  xor
  g1762
  (
    n1805,
    n1509,
    n1270,
    n1299,
    n1578
  );


  nand
  g1763
  (
    n1791,
    n1584,
    n1302,
    n1577,
    n1316
  );


  and
  g1764
  (
    n1756,
    n1038,
    n1602,
    n1346,
    n1604
  );


  xor
  g1765
  (
    n1703,
    n1410,
    n1451,
    n1652,
    n1510
  );


  and
  g1766
  (
    n1728,
    n1220,
    n1627,
    n1615
  );


  and
  g1767
  (
    n1700,
    n923,
    n1613,
    n1605,
    n1588
  );


  or
  g1768
  (
    n1810,
    n1472,
    n1612,
    n1253,
    n1593
  );


  nor
  g1769
  (
    n1777,
    n1297,
    n1241,
    n1254,
    n1513
  );


  nor
  g1770
  (
    n1736,
    n1636,
    n1407,
    n1634,
    n1576
  );


  xnor
  g1771
  (
    n1760,
    n1555,
    n1657,
    n1653,
    n1650
  );


  nor
  g1772
  (
    n1720,
    n1521,
    n1611,
    n1364,
    n1246
  );


  and
  g1773
  (
    n1759,
    n1613,
    n1477,
    n1657,
    n1595
  );


  xor
  g1774
  (
    n1677,
    n1649,
    n1424,
    n1589,
    n1626
  );


  xor
  g1775
  (
    n1707,
    n1654,
    n1543,
    n1607,
    n1586
  );


  or
  g1776
  (
    n1762,
    n1384,
    n1447,
    n1590,
    n748
  );


  and
  g1777
  (
    n1867,
    n1641,
    n1620,
    n1411,
    n1266
  );


  nor
  g1778
  (
    n1815,
    n1380,
    n1466,
    n1612,
    n1244
  );


  or
  g1779
  (
    n1801,
    n1577,
    n1486,
    n1446,
    n1582
  );


  xor
  g1780
  (
    n1697,
    n1290,
    n1335,
    n1571,
    n1649
  );


  or
  g1781
  (
    n1727,
    n1437,
    n1383,
    n1499,
    n1635
  );


  nand
  g1782
  (
    n1725,
    n1595,
    n1196,
    n1563,
    n1194
  );


  and
  g1783
  (
    n1818,
    n1559,
    n1496,
    n1226,
    n1243
  );


  nand
  g1784
  (
    n1842,
    n1541,
    n1567,
    n1561,
    n1646
  );


  nand
  g1785
  (
    n1773,
    n1572,
    n1378,
    n1581,
    n1370
  );


  xor
  g1786
  (
    n1706,
    n1372,
    n1590,
    n1239,
    n1610
  );


  xnor
  g1787
  (
    n1857,
    n1652,
    n1271,
    n1199,
    n1251
  );


  and
  g1788
  (
    n1755,
    n1354,
    n1650,
    n1504,
    n1191
  );


  or
  g1789
  (
    n1716,
    n1213,
    n1608,
    n1262,
    n1264
  );


  nor
  g1790
  (
    n1748,
    n1415,
    n1367,
    n1617,
    n923
  );


  and
  g1791
  (
    n1763,
    n1231,
    n1654,
    n1555,
    n1624
  );


  nor
  g1792
  (
    n1721,
    n1216,
    n1269,
    n1332,
    n1553
  );


  or
  g1793
  (
    n1769,
    n1593,
    n1507,
    n1218,
    n1445
  );


  nor
  g1794
  (
    n1832,
    n1626,
    n1651,
    n1207,
    n1497
  );


  and
  g1795
  (
    n1711,
    n1533,
    n1325,
    n1349,
    n1212
  );


  nor
  g1796
  (
    n1742,
    n1607,
    n1630,
    n1233,
    n1583
  );


  xor
  g1797
  (
    n1860,
    n1599,
    n1658,
    n1303,
    n1630
  );


  xor
  g1798
  (
    n1678,
    n1256,
    n1596,
    n1245,
    n1529
  );


  nand
  g1799
  (
    n1849,
    n1465,
    n1618,
    n1417,
    n1575
  );


  nor
  g1800
  (
    n1866,
    n1304,
    n1642,
    n1361,
    n1310
  );


  nand
  g1801
  (
    n1808,
    n1644,
    n1508,
    n1604,
    n1563
  );


  and
  g1802
  (
    n1708,
    n1455,
    n1227,
    n1599,
    n1587
  );


  xnor
  g1803
  (
    n1797,
    n1565,
    n1279,
    n1480,
    n1545
  );


  nor
  g1804
  (
    n1672,
    n1635,
    n1258,
    n1589,
    n1492
  );


  or
  g1805
  (
    n1699,
    n1635,
    n1622,
    n1618,
    n1390
  );


  nor
  g1806
  (
    n1794,
    n1613,
    n1292,
    n1653,
    n1287
  );


  nand
  g1807
  (
    n1750,
    n1330,
    n1585,
    n1600,
    n1293
  );


  xnor
  g1808
  (
    n1861,
    n1649,
    n1427,
    n1620,
    n1442
  );


  nand
  g1809
  (
    n1732,
    n1650,
    n1229,
    n1515,
    n1551
  );


  nor
  g1810
  (
    n1800,
    n1592,
    n1570,
    n1651,
    n1170
  );


  xnor
  g1811
  (
    n1730,
    n1284,
    n1401,
    n1629,
    n1623
  );


  nand
  g1812
  (
    n1847,
    n1655,
    n1549,
    n1607,
    n1448
  );


  nand
  g1813
  (
    n1724,
    n1539,
    n1594,
    n1331,
    n1532
  );


  xor
  g1814
  (
    n1745,
    n1613,
    n1574,
    n1584,
    n1376
  );


  xnor
  g1815
  (
    n1683,
    n1171,
    n1430,
    n1650,
    n1192
  );


  xor
  g1816
  (
    n1704,
    n1339,
    n1438,
    n1235,
    n1036
  );


  and
  g1817
  (
    n1858,
    n1564,
    n1561,
    n1540,
    n1609
  );


  xor
  g1818
  (
    n1856,
    n1558,
    n1617,
    n1562,
    n1501
  );


  nor
  g1819
  (
    n1798,
    n1552,
    n1464,
    n1539,
    n1644
  );


  and
  g1820
  (
    n1671,
    n1598,
    n1627,
    n1588,
    n1222
  );


  and
  g1821
  (
    n1803,
    n1534,
    n1359,
    n1637,
    n1344
  );


  or
  g1822
  (
    n1852,
    n1183,
    n1647,
    n1450,
    n1037
  );


  nand
  g1823
  (
    n1754,
    n1353,
    n1176,
    n1656,
    n1524
  );


  xor
  g1824
  (
    n1787,
    n1528,
    n1602,
    n1627,
    n1295
  );


  and
  g1825
  (
    n1752,
    n1366,
    n1560,
    n1393,
    n1395
  );


  xor
  g1826
  (
    n1729,
    n1392,
    n1179,
    n1536,
    n1583
  );


  xnor
  g1827
  (
    n1779,
    n1642,
    n1595,
    n1639,
    n1506
  );


  xnor
  g1828
  (
    n1692,
    n1580,
    n1543,
    n1600,
    n1381
  );


  xnor
  g1829
  (
    n1786,
    n1405,
    n1608,
    n1615,
    n1587
  );


  xnor
  g1830
  (
    n1804,
    n747,
    n1037,
    n1603,
    n1314
  );


  or
  g1831
  (
    n1751,
    n1535,
    n1602,
    n1609,
    n1655
  );


  nand
  g1832
  (
    n1768,
    n1457,
    n1527,
    n1505,
    n1177
  );


  xor
  g1833
  (
    n1696,
    n1632,
    n1397,
    n1259,
    n1470
  );


  nand
  g1834
  (
    n1785,
    n1565,
    n1632,
    n1296,
    n1562
  );


  buf
  g1835
  (
    n1870,
    n1676
  );


  not
  g1836
  (
    n1872,
    n1672
  );


  buf
  g1837
  (
    n1868,
    n1675
  );


  nand
  g1838
  (
    n1871,
    n1678,
    n1680,
    n1671
  );


  nor
  g1839
  (
    n1869,
    n1673,
    n1679,
    n1677,
    n1674
  );


  nor
  g1840
  (
    n1876,
    n1869,
    n1662,
    n1669,
    n1663
  );


  or
  g1841
  (
    n1886,
    n1663,
    n1669,
    n1664,
    n1870
  );


  xor
  g1842
  (
    n1874,
    n1665,
    n1871,
    n587
  );


  nand
  g1843
  (
    n1879,
    n1662,
    n1666,
    n1872
  );


  xnor
  g1844
  (
    n1884,
    n1660,
    n586,
    n1870,
    n1868
  );


  nand
  g1845
  (
    n1873,
    n1669,
    n1668,
    n1871
  );


  and
  g1846
  (
    n1877,
    n1667,
    n1665,
    n1872,
    n1669
  );


  xor
  g1847
  (
    n1881,
    n586,
    n1668,
    n1661,
    n1667
  );


  nor
  g1848
  (
    n1890,
    n1871,
    n1663,
    n1664
  );


  nand
  g1849
  (
    n1885,
    n1668,
    n1661,
    n1659,
    n1868
  );


  xnor
  g1850
  (
    n1887,
    n1666,
    n1660,
    n1667
  );


  nand
  g1851
  (
    n1882,
    n1664,
    n1869,
    n1665,
    n588
  );


  xnor
  g1852
  (
    n1888,
    n1869,
    n1670,
    n1667,
    n1668
  );


  xor
  g1853
  (
    n1883,
    n587,
    n1872,
    n1670,
    n1659
  );


  xor
  g1854
  (
    n1875,
    n1664,
    n1869,
    n1659,
    n1870
  );


  nand
  g1855
  (
    n1880,
    n1661,
    n1670,
    n1870,
    n1666
  );


  nand
  g1856
  (
    n1878,
    n1670,
    n1666,
    n1660,
    n1662
  );


  nand
  g1857
  (
    n1889,
    n1662,
    n1661,
    n587,
    n1665
  );


  xor
  g1858
  (
    n1891,
    n1681,
    n1716,
    n1695,
    n1690
  );


  nand
  g1859
  (
    n1900,
    n1697,
    n1696,
    n1683,
    n1687
  );


  or
  g1860
  (
    n1897,
    n1880,
    n1708,
    n1704,
    n1699
  );


  and
  g1861
  (
    n1898,
    n1881,
    n1878,
    n1702,
    n1720
  );


  or
  g1862
  (
    n1904,
    n1711,
    n1694,
    n1714,
    n1684
  );


  or
  g1863
  (
    n1903,
    n1700,
    n1882,
    n1703,
    n1724
  );


  or
  g1864
  (
    n1893,
    n1713,
    n1721,
    n1874,
    n1688
  );


  xor
  g1865
  (
    n1901,
    n1698,
    n1877,
    n1879,
    n1717
  );


  xor
  g1866
  (
    n1902,
    n1701,
    n1883,
    n1882,
    n1725
  );


  xor
  g1867
  (
    n1899,
    n1881,
    n1883,
    n1705,
    n1685
  );


  or
  g1868
  (
    n1895,
    n1691,
    n1707,
    n1712,
    n1875
  );


  and
  g1869
  (
    n1905,
    n1706,
    n1709,
    n1873,
    n1718
  );


  nor
  g1870
  (
    n1892,
    n1723,
    n1715,
    n1693,
    n1719
  );


  or
  g1871
  (
    n1894,
    n1722,
    n1686,
    n1692,
    n1682
  );


  nand
  g1872
  (
    n1896,
    n1876,
    n1689,
    n1710,
    n1880
  );


  not
  g1873
  (
    n1912,
    n750
  );


  not
  g1874
  (
    n1915,
    n1896
  );


  not
  g1875
  (
    n1910,
    n1904
  );


  not
  g1876
  (
    n1906,
    n1902
  );


  buf
  g1877
  (
    n1914,
    n1905
  );


  buf
  g1878
  (
    n1908,
    n925
  );


  not
  g1879
  (
    n1913,
    n924
  );


  not
  g1880
  (
    n1918,
    n1729
  );


  nand
  g1881
  (
    n1907,
    n1899,
    n1894,
    n1727
  );


  xnor
  g1882
  (
    n1911,
    n923,
    n1893,
    n1903
  );


  nor
  g1883
  (
    n1917,
    n925,
    n1726,
    n1728,
    n924
  );


  xnor
  g1884
  (
    n1909,
    n925,
    n924,
    n1901,
    n1897
  );


  xor
  g1885
  (
    n1916,
    n1895,
    n1898,
    n1900,
    n924
  );


  xor
  g1886
  (
    n1931,
    n1768,
    n1846,
    n1888,
    n1912
  );


  or
  g1887
  (
    n1924,
    n1909,
    n1758,
    n1741,
    n1866
  );


  or
  g1888
  (
    n1928,
    n1742,
    n1914,
    n1908,
    n1917
  );


  nand
  g1889
  (
    n1943,
    n1856,
    n1749,
    n1744,
    n1909
  );


  xnor
  g1890
  (
    n1954,
    n1776,
    n1807,
    n1843,
    n1826
  );


  and
  g1891
  (
    n1944,
    n925,
    n1833,
    n1918,
    n1913
  );


  nor
  g1892
  (
    n1964,
    n1909,
    n1755,
    n1760,
    n1834
  );


  xor
  g1893
  (
    n1929,
    n1838,
    n1912,
    n1803,
    n1828
  );


  nand
  g1894
  (
    n1968,
    n1827,
    n1916,
    n1738,
    n1890
  );


  nor
  g1895
  (
    n1935,
    n1750,
    n1910,
    n1784,
    n1773
  );


  xor
  g1896
  (
    n1939,
    n1748,
    n1885,
    n1778,
    n1918
  );


  xor
  g1897
  (
    n1941,
    n1814,
    n1809,
    n1886,
    n1852
  );


  nand
  g1898
  (
    n1942,
    n1915,
    n1907,
    n1914,
    n1835
  );


  nor
  g1899
  (
    n1947,
    n1886,
    n1918,
    n1864,
    n1822
  );


  and
  g1900
  (
    n1936,
    n1820,
    n1796,
    n1788,
    n1860
  );


  nand
  g1901
  (
    n1920,
    n1819,
    n1910,
    n1837,
    n1911
  );


  xor
  g1902
  (
    n1966,
    n1915,
    n1823,
    n1766,
    n1888
  );


  nand
  g1903
  (
    n1967,
    n1732,
    n1801,
    n1906,
    n1911
  );


  xnor
  g1904
  (
    n1951,
    n1914,
    n926,
    n1763,
    n1917
  );


  xnor
  g1905
  (
    n1956,
    n1884,
    n1854,
    n1794,
    n1797
  );


  nor
  g1906
  (
    n1969,
    n1786,
    n1806,
    n1800,
    n1781
  );


  xnor
  g1907
  (
    n1934,
    n1858,
    n1885,
    n1911,
    n1845
  );


  nand
  g1908
  (
    n1945,
    n1769,
    n1916,
    n1913,
    n1802
  );


  xnor
  g1909
  (
    n1938,
    n1839,
    n1855,
    n1908,
    n1739
  );


  xor
  g1910
  (
    n1926,
    n1734,
    n1813,
    n1830,
    n1867
  );


  and
  g1911
  (
    n1963,
    n1765,
    n1916,
    n1842,
    n1829
  );


  xnor
  g1912
  (
    n1932,
    n1756,
    n1844,
    n1791,
    n1824
  );


  xor
  g1913
  (
    n1950,
    n1832,
    n1798,
    n1762,
    n1745
  );


  xor
  g1914
  (
    n1933,
    n1840,
    n1793,
    n1889,
    n1770
  );


  xor
  g1915
  (
    n1960,
    n1752,
    n1862,
    n1908,
    n1859
  );


  and
  g1916
  (
    n1919,
    n1916,
    n1863,
    n1907,
    n1757
  );


  xor
  g1917
  (
    n1961,
    n1861,
    n1747,
    n1774,
    n1799
  );


  or
  g1918
  (
    n1965,
    n1759,
    n1787,
    n1907,
    n1789
  );


  xnor
  g1919
  (
    n1970,
    n1736,
    n1910,
    n1913,
    n1847
  );


  xor
  g1920
  (
    n1948,
    n1906,
    n1853,
    n1767,
    n1825
  );


  xnor
  g1921
  (
    n1959,
    n1850,
    n1775,
    n1887,
    n1754
  );


  nor
  g1922
  (
    n1957,
    n1733,
    n1764,
    n1792,
    n1795
  );


  nor
  g1923
  (
    n1953,
    n751,
    n1782,
    n1810,
    n1771
  );


  or
  g1924
  (
    n1946,
    n1889,
    n1779,
    n1785,
    n1848
  );


  xnor
  g1925
  (
    n1940,
    n1836,
    n1817,
    n1818,
    n1913
  );


  nand
  g1926
  (
    n1925,
    n1917,
    n1884,
    n1841,
    n926
  );


  and
  g1927
  (
    n1923,
    n1865,
    n1912,
    n1746,
    n1731
  );


  xnor
  g1928
  (
    n1955,
    n1735,
    n1857,
    n1751,
    n1740
  );


  xnor
  g1929
  (
    n1958,
    n1907,
    n1831,
    n1780,
    n1849
  );


  xor
  g1930
  (
    n1949,
    n1918,
    n1811,
    n1917,
    n1914
  );


  xnor
  g1931
  (
    n1922,
    n1777,
    n1912,
    n1815,
    n1821
  );


  and
  g1932
  (
    n1927,
    n1772,
    n1910,
    n1911,
    n1783
  );


  xnor
  g1933
  (
    n1962,
    n1890,
    n1851,
    n1816,
    n1906
  );


  xnor
  g1934
  (
    n1921,
    n1915,
    n1743,
    n1808,
    n1887
  );


  and
  g1935
  (
    n1930,
    n1812,
    n1804,
    n1761,
    n1753
  );


  or
  g1936
  (
    n1952,
    n1730,
    n1906,
    n1908,
    n1805
  );


  xor
  g1937
  (
    n1937,
    n1790,
    n1909,
    n1737,
    n1915
  );


  nor
  g1938
  (
    n1984,
    n1924,
    n791,
    n1946,
    n156
  );


  xor
  g1939
  (
    n2010,
    n929,
    n1921,
    n1953,
    n840
  );


  nor
  g1940
  (
    n2013,
    n790,
    n1959,
    n1947,
    n855
  );


  xor
  g1941
  (
    n1996,
    n775,
    n1958,
    n765,
    n767
  );


  and
  g1942
  (
    n2018,
    n795,
    n841,
    n774,
    n837
  );


  or
  g1943
  (
    n2015,
    n839,
    n590,
    n833,
    n1954
  );


  nor
  g1944
  (
    n1987,
    n1948,
    n811,
    n926,
    n809
  );


  or
  g1945
  (
    n2017,
    n754,
    n1934,
    n768,
    n829
  );


  xor
  g1946
  (
    n1997,
    n929,
    n590,
    n849
  );


  nand
  g1947
  (
    n1976,
    n826,
    n1925,
    n928,
    n803
  );


  nand
  g1948
  (
    n1973,
    n777,
    n588,
    n815,
    n818
  );


  or
  g1949
  (
    n2012,
    n793,
    n1927,
    n1931,
    n1944
  );


  xor
  g1950
  (
    n1974,
    n1942,
    n821,
    n798,
    n823
  );


  xor
  g1951
  (
    n1971,
    n787,
    n847,
    n1940,
    n845
  );


  xnor
  g1952
  (
    n1989,
    n812,
    n1955,
    n1919,
    n804
  );


  nand
  g1953
  (
    n1986,
    n794,
    n792,
    n927,
    n824
  );


  xnor
  g1954
  (
    n2006,
    n832,
    n820,
    n1970,
    n788
  );


  nor
  g1955
  (
    n2014,
    n771,
    n1965,
    n806,
    n1961
  );


  and
  g1956
  (
    n1992,
    n856,
    n1943,
    n926,
    n1928
  );


  and
  g1957
  (
    n2009,
    n860,
    n755,
    n1920,
    n759
  );


  and
  g1958
  (
    n2011,
    n589,
    n828,
    n1962,
    n852
  );


  and
  g1959
  (
    n1988,
    n772,
    n1964,
    n834,
    n850
  );


  xnor
  g1960
  (
    n1990,
    n757,
    n782,
    n797,
    n1945
  );


  nand
  g1961
  (
    n1983,
    n1922,
    n783,
    n761,
    n1951
  );


  and
  g1962
  (
    n2000,
    n760,
    n1935,
    n827,
    n1950
  );


  nor
  g1963
  (
    n1982,
    n844,
    n588,
    n1968,
    n810
  );


  xor
  g1964
  (
    n1993,
    n1923,
    n589,
    n863,
    n928
  );


  nor
  g1965
  (
    n2002,
    n1929,
    n764,
    n1966,
    n780
  );


  nand
  g1966
  (
    n1980,
    n781,
    n752,
    n800,
    n763
  );


  and
  g1967
  (
    n1979,
    n156,
    n854,
    n842,
    n779
  );


  xor
  g1968
  (
    n2016,
    n1932,
    n928,
    n1960,
    n784
  );


  xnor
  g1969
  (
    n1999,
    n758,
    n853,
    n819,
    n1941
  );


  xnor
  g1970
  (
    n2001,
    n1956,
    n846,
    n1926,
    n590
  );


  or
  g1971
  (
    n2005,
    n776,
    n927,
    n766,
    n778
  );


  nand
  g1972
  (
    n1995,
    n1937,
    n858,
    n1969,
    n1930
  );


  xnor
  g1973
  (
    n2004,
    n799,
    n1952,
    n770,
    n762
  );


  nand
  g1974
  (
    n1998,
    n862,
    n851,
    n927,
    n805
  );


  nand
  g1975
  (
    n1991,
    n843,
    n929,
    n835,
    n836
  );


  xor
  g1976
  (
    n1994,
    n807,
    n813,
    n1963,
    n838
  );


  or
  g1977
  (
    n2003,
    n816,
    n1949,
    n861,
    n1939
  );


  xor
  g1978
  (
    n1972,
    n589,
    n1933,
    n927,
    n831
  );


  nor
  g1979
  (
    n2008,
    n756,
    n928,
    n1967,
    n789
  );


  or
  g1980
  (
    n1985,
    n589,
    n830,
    n929,
    n588
  );


  xor
  g1981
  (
    n1975,
    n802,
    n825,
    n822,
    n753
  );


  nor
  g1982
  (
    n2007,
    n769,
    n817,
    n857,
    n1957
  );


  nand
  g1983
  (
    n1978,
    n814,
    n156,
    n1938,
    n848
  );


  nand
  g1984
  (
    n1981,
    n1936,
    n796,
    n859,
    n808
  );


  nand
  g1985
  (
    n1977,
    n786,
    n801,
    n785,
    n773
  );


  or
  g1986
  (
    AntiSAT_key_wire,
    n2014,
    n1995,
    n1974,
    n1986
  );


  nand
  g1987
  (
    n2025,
    n2015,
    n931,
    n2004,
    n1989
  );


  and
  g1988
  (
    n2030,
    n1997,
    n1990,
    n1992,
    n1976
  );


  nand
  g1989
  (
    n2027,
    n1979,
    n1999,
    n930,
    n2001
  );


  nand
  g1990
  (
    n2028,
    n1987,
    n931,
    n1981
  );


  or
  g1991
  (
    n2019,
    n1984,
    n2016,
    n2012,
    n2006
  );


  nand
  g1992
  (
    n2026,
    n2008,
    n930,
    n2005,
    n1983
  );


  xnor
  g1993
  (
    n2022,
    n2017,
    n930,
    n1991
  );


  and
  g1994
  (
    n2029,
    n1975,
    n1977,
    n2011,
    n1988
  );


  xor
  g1995
  (
    n2021,
    n2000,
    n2013,
    n931,
    n2003
  );


  and
  g1996
  (
    n2023,
    n1994,
    n1982,
    n2018,
    n1971
  );


  xor
  g1997
  (
    n2020,
    n1985,
    n2010,
    n1993,
    n2002
  );


  xnor
  g1998
  (
    n2032,
    n2009,
    n1980,
    n1998,
    n1996
  );


  and
  g1999
  (
    n2024,
    n2007,
    n1973,
    n1972,
    n1978
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n2031,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

