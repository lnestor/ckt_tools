

module Stat_100_69
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n123,
  n117,
  n103,
  n109,
  n115,
  n116,
  n118,
  n98,
  n104,
  n108,
  n106,
  n120,
  n107,
  n101,
  n102,
  n97,
  n122,
  n119,
  n100,
  n110,
  n111,
  n99,
  n114,
  n121,
  n129,
  n128,
  n126,
  n131,
  n130,
  n125,
  n127,
  n132
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n123;output n117;output n103;output n109;output n115;output n116;output n118;output n98;output n104;output n108;output n106;output n120;output n107;output n101;output n102;output n97;output n122;output n119;output n100;output n110;output n111;output n99;output n114;output n121;output n129;output n128;output n126;output n131;output n130;output n125;output n127;output n132;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n105;wire n112;wire n113;wire n124;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;

  buf
  g0
  (
    KeyWire_0_15,
    n22
  );


  buf
  g1
  (
    KeyWire_0_3,
    n3
  );


  buf
  g2
  (
    KeyWire_0_61,
    n17
  );


  buf
  g3
  (
    n34,
    n20
  );


  nor
  g4
  (
    n38,
    n11,
    n15,
    n16
  );


  nand
  g5
  (
    n40,
    n8,
    n1,
    n19,
    n18
  );


  or
  g6
  (
    KeyWire_0_52,
    n9,
    n5,
    n10,
    n2
  );


  nor
  g7
  (
    n33,
    n4,
    n21,
    n23,
    n6
  );


  xor
  g8
  (
    KeyWire_0_20,
    n7,
    n12,
    n13,
    n14
  );


  buf
  g9
  (
    n47,
    n40
  );


  not
  g10
  (
    KeyWire_0_63,
    n37
  );


  buf
  g11
  (
    KeyWire_0_59,
    n36
  );


  not
  g12
  (
    n42,
    n34
  );


  not
  g13
  (
    KeyWire_0_60,
    n33
  );


  buf
  g14
  (
    KeyWire_0_32,
    n39
  );


  not
  g15
  (
    n43,
    n38
  );


  buf
  g16
  (
    KeyWire_0_51,
    n35
  );


  not
  g17
  (
    KeyWire_0_23,
    n46
  );


  buf
  g18
  (
    KeyWire_0_22,
    n44
  );


  buf
  g19
  (
    n61,
    n43
  );


  not
  g20
  (
    KeyWire_0_38,
    n48
  );


  not
  g21
  (
    KeyWire_0_48,
    n49
  );


  not
  g22
  (
    KeyWire_0_36,
    n42
  );


  buf
  g23
  (
    KeyWire_0_42,
    n46
  );


  buf
  g24
  (
    KeyWire_0_8,
    n44
  );


  not
  g25
  (
    n69,
    n45
  );


  not
  g26
  (
    KeyWire_0_46,
    n45
  );


  not
  g27
  (
    KeyWire_0_18,
    n47
  );


  not
  g28
  (
    n66,
    n43
  );


  not
  g29
  (
    n76,
    n43
  );


  not
  g30
  (
    KeyWire_0_26,
    n46
  );


  not
  g31
  (
    KeyWire_0_44,
    n43
  );


  buf
  g32
  (
    KeyWire_0_0,
    n48
  );


  buf
  g33
  (
    KeyWire_0_47,
    n48
  );


  not
  g34
  (
    KeyWire_0_34,
    n47
  );


  buf
  g35
  (
    KeyWire_0_7,
    n48
  );


  not
  g36
  (
    n74,
    n45
  );


  not
  g37
  (
    KeyWire_0_21,
    n46
  );


  buf
  g38
  (
    KeyWire_0_40,
    n42
  );


  not
  g39
  (
    KeyWire_0_17,
    n47
  );


  not
  g40
  (
    KeyWire_0_53,
    n47
  );


  not
  g41
  (
    KeyWire_0_12,
    n49
  );


  buf
  g42
  (
    KeyWire_0_54,
    n44
  );


  buf
  g43
  (
    n67,
    n44
  );


  nor
  g44
  (
    n65,
    n49,
    n45,
    n41
  );


  not
  g45
  (
    KeyWire_0_11,
    n50
  );


  buf
  g46
  (
    KeyWire_0_6,
    n54
  );


  not
  g47
  (
    n93,
    n29
  );


  not
  g48
  (
    KeyWire_0_28,
    n55
  );


  not
  g49
  (
    KeyWire_0_16,
    n53
  );


  buf
  g50
  (
    n83,
    n55
  );


  not
  g51
  (
    KeyWire_0_4,
    n53
  );


  buf
  g52
  (
    KeyWire_0_50,
    n32
  );


  not
  g53
  (
    KeyWire_0_14,
    n26
  );


  buf
  g54
  (
    n89,
    n25
  );


  buf
  g55
  (
    n95,
    n31
  );


  buf
  g56
  (
    n92,
    n53
  );


  not
  g57
  (
    KeyWire_0_33,
    n28
  );


  nor
  g58
  (
    KeyWire_0_58,
    n55,
    n24,
    n49
  );


  xor
  g59
  (
    KeyWire_0_49,
    n27,
    n54,
    n55
  );


  xor
  g60
  (
    KeyWire_0_62,
    n54,
    n56,
    n30
  );


  xnor
  g61
  (
    n84,
    n53,
    n51,
    n52
  );


  xnor
  g62
  (
    n94,
    n54,
    n52,
    n51
  );


  nand
  g63
  (
    KeyWire_0_41,
    n67,
    n68,
    n74,
    n84
  );


  xnor
  g64
  (
    n118,
    n70,
    n72,
    n93
  );


  or
  g65
  (
    n110,
    n70,
    n68,
    n69,
    n63
  );


  xor
  g66
  (
    KeyWire_0_25,
    n90,
    n76,
    n64,
    n80
  );


  and
  g67
  (
    n112,
    n56,
    n93,
    n74
  );


  nor
  g68
  (
    KeyWire_0_1,
    n77,
    n68,
    n61,
    n83
  );


  xor
  g69
  (
    n108,
    n65,
    n76,
    n57,
    n61
  );


  xor
  g70
  (
    n114,
    n60,
    n91,
    n70,
    n57
  );


  and
  g71
  (
    KeyWire_0_24,
    n61,
    n66,
    n75,
    n89
  );


  and
  g72
  (
    KeyWire_0_31,
    n90,
    n71,
    n67,
    n88
  );


  and
  g73
  (
    KeyWire_0_5,
    n77,
    n73,
    n89,
    n57
  );


  nand
  g74
  (
    KeyWire_0_43,
    n63,
    n73,
    n81
  );


  nand
  g75
  (
    KeyWire_0_57,
    n92,
    n69,
    n74,
    n91
  );


  nor
  g76
  (
    KeyWire_0_30,
    n63,
    n65,
    n72
  );


  nor
  g77
  (
    n111,
    n82,
    n58,
    n60
  );


  or
  g78
  (
    KeyWire_0_37,
    n58,
    n85,
    n61,
    n67
  );


  xnor
  g79
  (
    n124,
    n91,
    n72,
    n68,
    n78
  );


  nand
  g80
  (
    KeyWire_0_13,
    n62,
    n79,
    n73,
    n57
  );


  nand
  g81
  (
    KeyWire_0_56,
    n86,
    n59,
    n71
  );


  xnor
  g82
  (
    KeyWire_0_27,
    n91,
    n92,
    n66
  );


  xor
  g83
  (
    n100,
    n75,
    n62,
    n90,
    n77
  );


  or
  g84
  (
    KeyWire_0_2,
    n64,
    n71,
    n70,
    n65
  );


  xor
  g85
  (
    n119,
    n69,
    n64,
    n89,
    n60
  );


  nand
  g86
  (
    n113,
    n75,
    n62,
    n69,
    n87
  );


  or
  g87
  (
    KeyWire_0_39,
    n89,
    n56,
    n67,
    n66
  );


  nand
  g88
  (
    KeyWire_0_9,
    n76,
    n64,
    n60,
    n75
  );


  xnor
  g89
  (
    n121,
    n92,
    n62,
    n77,
    n59
  );


  nand
  g90
  (
    KeyWire_0_45,
    n59,
    n71,
    n63,
    n90
  );


  nor
  g91
  (
    n104,
    n58,
    n76,
    n56,
    n66
  );


  buf
  g92
  (
    KeyWire_0_19,
    n94
  );


  buf
  g93
  (
    KeyWire_0_10,
    n117
  );


  buf
  g94
  (
    KeyWire_0_35,
    n115
  );


  xnor
  g95
  (
    KeyWire_0_55,
    n118,
    n123,
    n94
  );


  nand
  g96
  (
    n129,
    n94,
    n95
  );


  xnor
  g97
  (
    KeyWire_0_29,
    n120,
    n114,
    n95,
    n93
  );


  nand
  g98
  (
    n131,
    n93,
    n122,
    n95,
    n124
  );


  xnor
  g99
  (
    n128,
    n119,
    n116,
    n113,
    n121
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n72,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n117,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n107,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n39,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n86,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n123,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n78,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n77,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n54,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n98,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n125,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n82,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n59,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n115,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n90,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n35,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n91,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n64,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n52,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n127,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n36,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n53,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n56,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n55,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n122,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n106,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n68,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n120,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n88,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n130,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n96,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n109,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n45,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n79,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n62,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n132,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n70,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n97,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n51,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n101,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n73,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n103,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n57,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n102,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n63,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n105,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n75,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n50,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n60,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n80,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n87,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n46,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n37,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n71,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n58,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n126,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n99,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n116,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n85,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n48,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n44,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n41,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n81,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n49,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


