

module Stat_114_49
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n130,
  n118,
  n131,
  n123,
  n115,
  n117,
  n114,
  n120,
  n128,
  n121,
  n119,
  n126,
  n129,
  n124,
  n116,
  n125,
  n127,
  n122,
  n113,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n130;
  output n118;
  output n131;
  output n123;
  output n115;
  output n117;
  output n114;
  output n120;
  output n128;
  output n121;
  output n119;
  output n126;
  output n129;
  output n124;
  output n116;
  output n125;
  output n127;
  output n122;
  output n113;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    KeyWire_0_50,
    n17
  );


  buf
  g1
  (
    n26,
    n7
  );


  buf
  g2
  (
    n20,
    n11
  );


  not
  g3
  (
    n24,
    n6
  );


  not
  g4
  (
    n18,
    n9
  );


  buf
  g5
  (
    n25,
    n17
  );


  buf
  g6
  (
    n23,
    n12
  );


  buf
  g7
  (
    n28,
    n15
  );


  buf
  g8
  (
    n30,
    n14
  );


  not
  g9
  (
    n35,
    n13
  );


  buf
  g10
  (
    n27,
    n10
  );


  not
  g11
  (
    KeyWire_0_58,
    n16
  );


  buf
  g12
  (
    KeyWire_0_45,
    n5
  );


  not
  g13
  (
    KeyWire_0_54,
    n3
  );


  buf
  g14
  (
    n21,
    n1
  );


  buf
  g15
  (
    KeyWire_0_37,
    n4
  );


  buf
  g16
  (
    KeyWire_0_6,
    n2
  );


  buf
  g17
  (
    KeyWire_0_11,
    n8
  );


  not
  g18
  (
    KeyWire_0_53,
    n31
  );


  buf
  g19
  (
    KeyWire_0_63,
    n34
  );


  not
  g20
  (
    KeyWire_0_24,
    n24
  );


  not
  g21
  (
    n65,
    n20
  );


  buf
  g22
  (
    KeyWire_0_31,
    n27
  );


  not
  g23
  (
    KeyWire_0_48,
    n35
  );


  not
  g24
  (
    n64,
    n19
  );


  buf
  g25
  (
    KeyWire_0_18,
    n26
  );


  not
  g26
  (
    n42,
    n24
  );


  buf
  g27
  (
    KeyWire_0_0,
    n35
  );


  not
  g28
  (
    KeyWire_0_39,
    n27
  );


  not
  g29
  (
    KeyWire_0_47,
    n29
  );


  not
  g30
  (
    n72,
    n30
  );


  buf
  g31
  (
    KeyWire_0_8,
    n35
  );


  not
  g32
  (
    KeyWire_0_60,
    n31
  );


  not
  g33
  (
    n70,
    n33
  );


  buf
  g34
  (
    KeyWire_0_27,
    n22
  );


  not
  g35
  (
    n44,
    n18
  );


  not
  g36
  (
    n66,
    n29
  );


  not
  g37
  (
    n61,
    n23
  );


  not
  g38
  (
    n37,
    n22
  );


  buf
  g39
  (
    KeyWire_0_5,
    n18
  );


  not
  g40
  (
    n40,
    n34
  );


  not
  g41
  (
    n47,
    n28
  );


  not
  g42
  (
    KeyWire_0_57,
    n34
  );


  buf
  g43
  (
    KeyWire_0_46,
    n25
  );


  not
  g44
  (
    n38,
    n30
  );


  buf
  g45
  (
    n58,
    n20
  );


  buf
  g46
  (
    KeyWire_0_3,
    n19
  );


  buf
  g47
  (
    KeyWire_0_33,
    n33
  );


  buf
  g48
  (
    KeyWire_0_51,
    n28
  );


  buf
  g49
  (
    KeyWire_0_22,
    n23
  );


  buf
  g50
  (
    KeyWire_0_30,
    n32
  );


  not
  g51
  (
    n46,
    n21
  );


  not
  g52
  (
    KeyWire_0_4,
    n26
  );


  not
  g53
  (
    KeyWire_0_1,
    n21
  );


  buf
  g54
  (
    KeyWire_0_40,
    n32
  );


  not
  g55
  (
    KeyWire_0_32,
    n25
  );


  not
  g56
  (
    KeyWire_0_55,
    n49
  );


  not
  g57
  (
    KeyWire_0_42,
    n68
  );


  buf
  g58
  (
    n100,
    n39
  );


  buf
  g59
  (
    KeyWire_0_38,
    n38
  );


  buf
  g60
  (
    n74,
    n55
  );


  buf
  g61
  (
    KeyWire_0_17,
    n43
  );


  not
  g62
  (
    KeyWire_0_21,
    n37
  );


  buf
  g63
  (
    KeyWire_0_49,
    n42
  );


  buf
  g64
  (
    KeyWire_0_7,
    n51
  );


  not
  g65
  (
    n75,
    n65
  );


  buf
  g66
  (
    KeyWire_0_16,
    n66
  );


  not
  g67
  (
    KeyWire_0_41,
    n60
  );


  not
  g68
  (
    n103,
    n64
  );


  buf
  g69
  (
    KeyWire_0_52,
    n53
  );


  buf
  g70
  (
    KeyWire_0_56,
    n69
  );


  not
  g71
  (
    KeyWire_0_2,
    n40
  );


  buf
  g72
  (
    n97,
    n72
  );


  not
  g73
  (
    KeyWire_0_34,
    n36
  );


  buf
  g74
  (
    n85,
    n46
  );


  buf
  g75
  (
    KeyWire_0_20,
    n48
  );


  not
  g76
  (
    n79,
    n71
  );


  buf
  g77
  (
    KeyWire_0_15,
    n57
  );


  buf
  g78
  (
    KeyWire_0_10,
    n73
  );


  buf
  g79
  (
    KeyWire_0_44,
    n58
  );


  not
  g80
  (
    n99,
    n61
  );


  buf
  g81
  (
    n101,
    n41
  );


  buf
  g82
  (
    n102,
    n54
  );


  not
  g83
  (
    KeyWire_0_29,
    n59
  );


  not
  g84
  (
    KeyWire_0_25,
    n52
  );


  not
  g85
  (
    KeyWire_0_28,
    n67
  );


  not
  g86
  (
    n110,
    n73
  );


  not
  g87
  (
    KeyWire_0_36,
    n63
  );


  buf
  g88
  (
    n87,
    n62
  );


  buf
  g89
  (
    KeyWire_0_61,
    n56
  );


  buf
  g90
  (
    KeyWire_0_35,
    n50
  );


  not
  g91
  (
    n111,
    n70
  );


  not
  g92
  (
    n108,
    n44
  );


  buf
  g93
  (
    n81,
    n45
  );


  not
  g94
  (
    KeyWire_0_9,
    n47
  );


  not
  g95
  (
    KeyWire_0_62,
    n88
  );


  buf
  g96
  (
    KeyWire_0_59,
    n108
  );


  not
  g97
  (
    n129,
    n107
  );


  buf
  g98
  (
    KeyWire_0_14,
    n106
  );


  buf
  g99
  (
    n119,
    n75
  );


  buf
  g100
  (
    KeyWire_0_13,
    n100
  );


  buf
  g101
  (
    n126,
    n98
  );


  buf
  g102
  (
    n131,
    n78
  );


  not
  g103
  (
    KeyWire_0_12,
    n82
  );


  not
  g104
  (
    KeyWire_0_19,
    n93
  );


  not
  g105
  (
    n127,
    n110
  );


  not
  g106
  (
    KeyWire_0_23,
    n94
  );


  xnor
  g107
  (
    n116,
    n105,
    n101,
    n92
  );


  xor
  g108
  (
    n130,
    n102,
    n109,
    n87,
    n96
  );


  and
  g109
  (
    n118,
    n91,
    n97,
    n77,
    n99
  );


  xor
  g110
  (
    n114,
    n80,
    n90,
    n76,
    n79
  );


  nor
  g111
  (
    n117,
    n74,
    n111,
    n95,
    n83
  );


  nand
  g112
  (
    KeyWire_0_26,
    n81,
    n104,
    n112,
    n86
  );


  or
  g113
  (
    KeyWire_0_43,
    n84,
    n103,
    n89,
    n85
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n45,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n71,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n93,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n51,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n67,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n68,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n31,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n90,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n50,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n95,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n105,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n29,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n125,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n128,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n124,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n88,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n83,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n106,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n49,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n120,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n98,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n94,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n62,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n121,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n43,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n77,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n113,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n55,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n84,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n86,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n54,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n52,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n59,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n57,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n96,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n82,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n80,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n19,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n107,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n36,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n53,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n112,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n104,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n122,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n89,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n34,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n69,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n48,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n39,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n92,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n32,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n73,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n91,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n41,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n33,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n76,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n78,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n56,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n22,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n123,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n60,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n109,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n115,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n63,
    KeyNOTWire_0_63
  );


endmodule

