

module Stat_100_49
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n96,
  n107,
  n118,
  n110,
  n98,
  n106,
  n113,
  n121,
  n99,
  n111,
  n109,
  n97,
  n114,
  n93,
  n88,
  n119,
  n116,
  n101,
  n120,
  n103,
  n87,
  n108,
  n104,
  n115,
  n123,
  n128,
  n127,
  n129,
  n126,
  n124,
  n132,
  n131
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n96;output n107;output n118;output n110;output n98;output n106;output n113;output n121;output n99;output n111;output n109;output n97;output n114;output n93;output n88;output n119;output n116;output n101;output n120;output n103;output n87;output n108;output n104;output n115;output n123;output n128;output n127;output n129;output n126;output n124;output n132;output n131;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n89;wire n90;wire n91;wire n92;wire n94;wire n95;wire n100;wire n102;wire n105;wire n112;wire n117;wire n122;wire n125;wire n130;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;

  buf
  g0
  (
    KeyWire_0_8,
    n19
  );


  not
  g1
  (
    n49,
    n27
  );


  buf
  g2
  (
    n59,
    n5
  );


  buf
  g3
  (
    KeyWire_0_3,
    n32
  );


  buf
  g4
  (
    n42,
    n28
  );


  buf
  g5
  (
    KeyWire_0_5,
    n31
  );


  not
  g6
  (
    KeyWire_0_6,
    n21
  );


  not
  g7
  (
    n33,
    n10
  );


  not
  g8
  (
    n46,
    n15
  );


  buf
  g9
  (
    n76,
    n2
  );


  buf
  g10
  (
    n53,
    n3
  );


  buf
  g11
  (
    KeyWire_0_0,
    n26
  );


  buf
  g12
  (
    n69,
    n29
  );


  buf
  g13
  (
    n35,
    n20
  );


  not
  g14
  (
    n36,
    n26
  );


  buf
  g15
  (
    n45,
    n16
  );


  buf
  g16
  (
    KeyWire_0_15,
    n26
  );


  buf
  g17
  (
    n61,
    n24
  );


  not
  g18
  (
    n70,
    n13
  );


  buf
  g19
  (
    n78,
    n8
  );


  not
  g20
  (
    n52,
    n25
  );


  buf
  g21
  (
    n73,
    n17
  );


  not
  g22
  (
    n58,
    n24
  );


  buf
  g23
  (
    n72,
    n18
  );


  not
  g24
  (
    n68,
    n28
  );


  not
  g25
  (
    n43,
    n29
  );


  buf
  g26
  (
    n66,
    n27
  );


  not
  g27
  (
    n60,
    n11
  );


  buf
  g28
  (
    n67,
    n14
  );


  not
  g29
  (
    n62,
    n12
  );


  buf
  g30
  (
    n54,
    n25
  );


  buf
  g31
  (
    KeyWire_0_13,
    n4
  );


  buf
  g32
  (
    KeyWire_0_2,
    n31
  );


  not
  g33
  (
    n80,
    n23
  );


  buf
  g34
  (
    n64,
    n30
  );


  buf
  g35
  (
    n56,
    n27
  );


  buf
  g36
  (
    n82,
    n30
  );


  not
  g37
  (
    n79,
    n25
  );


  not
  g38
  (
    n77,
    n22
  );


  not
  g39
  (
    n41,
    n32
  );


  buf
  g40
  (
    n48,
    n29
  );


  buf
  g41
  (
    n71,
    n32
  );


  not
  g42
  (
    n57,
    n28
  );


  buf
  g43
  (
    n74,
    n1
  );


  buf
  g44
  (
    n44,
    n6
  );


  not
  g45
  (
    n40,
    n7
  );


  buf
  g46
  (
    KeyWire_0_14,
    n31
  );


  not
  g47
  (
    KeyWire_0_9,
    n24
  );


  not
  g48
  (
    n37,
    n9
  );


  not
  g49
  (
    n38,
    n30
  );


  or
  g50
  (
    n100,
    n61,
    n47,
    n36,
    n37
  );


  nand
  g51
  (
    n114,
    n53,
    n55,
    n78,
    n75
  );


  or
  g52
  (
    n86,
    n73,
    n50,
    n65,
    n51
  );


  nand
  g53
  (
    n93,
    n39,
    n56,
    n51,
    n37
  );


  xnor
  g54
  (
    n84,
    n79,
    n50,
    n70,
    n39
  );


  nand
  g55
  (
    n104,
    n35,
    n63,
    n33,
    n68
  );


  or
  g56
  (
    KeyWire_0_4,
    n40,
    n80,
    n72,
    n39
  );


  nor
  g57
  (
    n106,
    n73,
    n74,
    n77,
    n38
  );


  nand
  g58
  (
    n116,
    n44,
    n67,
    n66
  );


  nor
  g59
  (
    KeyWire_0_10,
    n65,
    n45,
    n79,
    n35
  );


  xnor
  g60
  (
    n121,
    n42,
    n59,
    n60,
    n77
  );


  and
  g61
  (
    n117,
    n55,
    n33,
    n67,
    n58
  );


  or
  g62
  (
    n120,
    n72,
    n58,
    n56,
    n79
  );


  or
  g63
  (
    n91,
    n75,
    n66,
    n37,
    n47
  );


  or
  g64
  (
    n97,
    n62,
    n78,
    n48,
    n41
  );


  nor
  g65
  (
    n119,
    n67,
    n52,
    n78
  );


  nand
  g66
  (
    n94,
    n65,
    n70,
    n71
  );


  xor
  g67
  (
    n105,
    n57,
    n59,
    n68,
    n62
  );


  xnor
  g68
  (
    n113,
    n53,
    n74,
    n63,
    n35
  );


  and
  g69
  (
    n107,
    n61,
    n50,
    n75,
    n76
  );


  and
  g70
  (
    n89,
    n68,
    n44,
    n71,
    n69
  );


  or
  g71
  (
    n98,
    n46,
    n68,
    n67,
    n36
  );


  nand
  g72
  (
    n109,
    n64,
    n76,
    n34
  );


  nor
  g73
  (
    n95,
    n57,
    n44,
    n46,
    n41
  );


  or
  g74
  (
    n118,
    n54,
    n45,
    n41,
    n74
  );


  xor
  g75
  (
    n85,
    n49,
    n71,
    n46,
    n43
  );


  nand
  g76
  (
    KeyWire_0_1,
    n78,
    n45,
    n40,
    n65
  );


  xnor
  g77
  (
    n90,
    n76,
    n42,
    n74
  );


  xor
  g78
  (
    KeyWire_0_12,
    n54,
    n49,
    n64,
    n53
  );


  nor
  g79
  (
    n122,
    n66,
    n48,
    n56,
    n70
  );


  nand
  g80
  (
    n96,
    n60,
    n69,
    n77,
    n52
  );


  or
  g81
  (
    n115,
    n73,
    n38,
    n75,
    n69
  );


  xnor
  g82
  (
    n87,
    n69,
    n71,
    n60,
    n64
  );


  xnor
  g83
  (
    n103,
    n72,
    n58,
    n64,
    n54
  );


  or
  g84
  (
    n83,
    n34,
    n36,
    n63,
    n55
  );


  nor
  g85
  (
    KeyWire_0_7,
    n61,
    n73,
    n51,
    n38
  );


  xnor
  g86
  (
    n112,
    n48,
    n72,
    n77,
    n43
  );


  xnor
  g87
  (
    n111,
    n63,
    n43,
    n79,
    n40
  );


  xor
  g88
  (
    KeyWire_0_11,
    n62,
    n57,
    n49,
    n47
  );


  xnor
  g89
  (
    n99,
    n59,
    n34,
    n80,
    n33
  );


  or
  g90
  (
    n125,
    n81,
    n115,
    n82
  );


  xnor
  g91
  (
    n127,
    n82,
    n110,
    n117
  );


  xor
  g92
  (
    n123,
    n120,
    n119,
    n121
  );


  nand
  g93
  (
    n126,
    n81,
    n122,
    n116
  );


  nor
  g94
  (
    n128,
    n113,
    n80,
    n82
  );


  xor
  g95
  (
    n124,
    n81,
    n114,
    n109
  );


  xor
  g96
  (
    n130,
    n81,
    n82,
    n80,
    n108
  );


  or
  g97
  (
    n129,
    n112,
    n118,
    n107,
    n111
  );


  buf
  g98
  (
    n132,
    n130
  );


  buf
  g99
  (
    n131,
    n129
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n81,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n88,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n65,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n55,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n101,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n34,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n51,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n108,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n39,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n50,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n102,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n92,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n110,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n47,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n63,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n75,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


