// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_186_441 written by SynthGen on 2021/05/24 19:47:14
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_186_441 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31,
 n210, n217, n212, n213, n215, n207, n208, n209,
 n211, n204, n203, n214, n206, n202, n216, n205,
 n201);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31;

output n210, n217, n212, n213, n215, n207, n208, n209,
 n211, n204, n203, n214, n206, n202, n216, n205,
 n201;

wire n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200;

not  g0 (n72, n15);
not  g1 (n54, n14);
not  g2 (n79, n13);
buf  g3 (n60, n14);
not  g4 (n68, n1);
not  g5 (n39, n7);
not  g6 (n69, n19);
buf  g7 (n52, n20);
not  g8 (n81, n6);
not  g9 (n64, n20);
not  g10 (n87, n13);
buf  g11 (n80, n10);
not  g12 (n63, n2);
buf  g13 (n62, n10);
not  g14 (n85, n3);
not  g15 (n33, n11);
buf  g16 (n67, n21);
not  g17 (n66, n6);
not  g18 (n83, n5);
buf  g19 (n53, n10);
buf  g20 (n82, n5);
buf  g21 (n55, n18);
not  g22 (n58, n3);
buf  g23 (n57, n8);
buf  g24 (n43, n14);
buf  g25 (n61, n20);
not  g26 (n35, n4);
not  g27 (n90, n9);
buf  g28 (n47, n11);
buf  g29 (n34, n19);
not  g30 (n59, n13);
buf  g31 (n42, n12);
not  g32 (n94, n17);
buf  g33 (n50, n8);
buf  g34 (n40, n4);
not  g35 (n92, n16);
not  g36 (n71, n7);
not  g37 (n91, n17);
buf  g38 (n56, n11);
buf  g39 (n32, n5);
not  g40 (n49, n2);
not  g41 (n44, n21);
not  g42 (n48, n6);
buf  g43 (n89, n7);
buf  g44 (n74, n16);
buf  g45 (n41, n4);
buf  g46 (n70, n8);
not  g47 (n51, n9);
not  g48 (n86, n12);
not  g49 (n36, n16);
buf  g50 (n73, n9);
buf  g51 (n38, n12);
buf  g52 (n88, n3);
buf  g53 (n78, n19);
not  g54 (n46, n1);
not  g55 (n65, n18);
not  g56 (n76, n15);
not  g57 (n75, n18);
not  g58 (n45, n1);
buf  g59 (n84, n21);
not  g60 (n77, n2);
buf  g61 (n93, n15);
not  g62 (n37, n17);
buf  g63 (n100, n43);
not  g64 (n115, n37);
not  g65 (n122, n36);
buf  g66 (n130, n39);
not  g67 (n116, n37);
buf  g68 (n127, n34);
buf  g69 (n97, n42);
buf  g70 (n105, n43);
buf  g71 (n107, n32);
not  g72 (n118, n32);
not  g73 (n106, n42);
not  g74 (n99, n36);
buf  g75 (n98, n37);
not  g76 (n117, n39);
not  g77 (n104, n38);
not  g78 (n96, n33);
not  g79 (n128, n40);
buf  g80 (n113, n33);
not  g81 (n129, n33);
buf  g82 (n103, n41);
not  g83 (n120, n44);
not  g84 (n126, n32);
not  g85 (n109, n41);
not  g86 (n132, n34);
not  g87 (n119, n36);
not  g88 (n101, n35);
not  g89 (n110, n40);
buf  g90 (n121, n41);
not  g91 (n95, n35);
not  g92 (n111, n39);
not  g93 (n131, n34);
buf  g94 (n102, n40);
not  g95 (n108, n42);
buf  g96 (n124, n44);
buf  g97 (n114, n35);
not  g98 (n123, n38);
not  g99 (n125, n43);
not  g100 (n112, n38);
and  g101 (n182, n125, n130, n106);
nor  g102 (n141, n64, n65, n113);
and  g103 (n144, n86, n124, n100);
xnor g104 (n147, n124, n92);
and  g105 (n167, n66, n84);
nand g106 (n187, n27, n51, n26);
nand g107 (n161, n57, n83, n72);
nand g108 (n159, n66, n82, n93);
or   g109 (n143, n28, n72, n69);
and  g110 (n150, n116, n121, n85);
xnor g111 (n195, n85, n91, n67);
xnor g112 (n190, n25, n30, n24);
nor  g113 (n181, n125, n31, n126);
xnor g114 (n135, n119, n50, n130);
or   g115 (n173, n45, n48, n61);
and  g116 (n200, n74, n47, n88);
nor  g117 (n151, n124, n79, n76);
nor  g118 (n192, n77, n125, n52);
nand g119 (n169, n128, n64, n89);
and  g120 (n189, n80, n29, n107);
nand g121 (n138, n62, n26, n86);
and  g122 (n148, n117, n55, n109);
xnor g123 (n186, n24, n131, n67);
or   g124 (n133, n54, n118, n93, n22);
or   g125 (n164, n59, n27, n91, n128);
nand g126 (n142, n79, n97, n61, n129);
or   g127 (n156, n71, n26, n57, n48);
and  g128 (n154, n47, n56, n126, n55);
nor  g129 (n179, n63, n89, n120, n45);
xnor g130 (n145, n25, n51, n73, n102);
and  g131 (n180, n132, n62, n50, n25);
nand g132 (n146, n55, n69, n128, n58);
xor  g133 (n155, n90, n58, n28);
and  g134 (n196, n110, n89, n94, n84);
nor  g135 (n166, n60, n81, n119, n27);
xor  g136 (n175, n105, n24, n29, n98);
or   g137 (n198, n52, n75, n118, n90);
nand g138 (n171, n72, n85, n94, n46);
xor  g139 (n165, n81, n53, n83, n63);
and  g140 (n157, n101, n87, n28, n70);
xor  g141 (n178, n87, n76, n78, n96);
xnor g142 (n152, n114, n60, n71, n126);
or   g143 (n188, n80, n76, n49, n62);
xnor g144 (n149, n92, n70, n22, n60);
nand g145 (n136, n99, n95, n91, n77);
or   g146 (n170, n83, n53, n49, n75);
xor  g147 (n191, n81, n69, n23, n82);
or   g148 (n177, n118, n31, n127, n54);
or   g149 (n163, n74, n68, n50, n61);
xor  g150 (n162, n121, n65, n123, n108);
xor  g151 (n139, n74, n79, n87, n64);
and  g152 (n172, n119, n123, n94, n77);
and  g153 (n184, n73, n112, n51, n131);
and  g154 (n193, n22, n127, n80, n88);
nand g155 (n197, n93, n129, n46, n66);
or   g156 (n137, n103, n75, n23, n120);
nand g157 (n153, n56, n122, n59, n53);
and  g158 (n134, n90, n78, n56, n132);
nor  g159 (n176, n122, n29, n57, n54);
nand g160 (n183, n121, n46, n65, n82);
xnor g161 (n194, n78, n63, n30, n123);
nor  g162 (n185, n68, n130, n122, n127);
xor  g163 (n174, n132, n111, n70, n131);
xnor g164 (n168, n88, n47, n45, n104);
nand g165 (n199, n49, n129, n68, n48);
nand g166 (n158, n31, n52, n67, n23);
nor  g167 (n140, n30, n44, n120, n73);
nand g168 (n160, n59, n86, n71, n115);
xor  g169 (n210, n156, n190, n165, n171);
or   g170 (n208, n177, n155, n135, n137);
and  g171 (n206, n144, n138, n186, n136);
or   g172 (n207, n147, n154, n134, n157);
and  g173 (n211, n163, n170, n182, n193);
nand g174 (n201, n168, n162, n183, n166);
nor  g175 (n209, n185, n188, n181, n194);
xor  g176 (n215, n172, n152, n191, n141);
xor  g177 (n213, n169, n184, n133, n200);
or   g178 (n214, n150, n195, n189, n196);
nor  g179 (n212, n198, n173, n151, n160);
and  g180 (n216, n179, n149, n153, n174);
or   g181 (n203, n192, n175, n139, n159);
or   g182 (n217, n164, n145, n161, n178);
nand g183 (n205, n143, n146, n167, n148);
xor  g184 (n202, n176, n187, n142, n180);
and  g185 (n204, n197, n199, n140, n158);
endmodule
