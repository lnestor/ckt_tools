

module Stat_1000_205
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n174,
  n148,
  n179,
  n165,
  n178,
  n151,
  n168,
  n139,
  n194,
  n150,
  n186,
  n124,
  n181,
  n147,
  n135,
  n182,
  n601,
  n613,
  n610,
  n611,
  n598,
  n608,
  n623,
  n605,
  n621,
  n602,
  n620,
  n606,
  n617,
  n622,
  n1031,
  n1032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n174;
  output n148;
  output n179;
  output n165;
  output n178;
  output n151;
  output n168;
  output n139;
  output n194;
  output n150;
  output n186;
  output n124;
  output n181;
  output n147;
  output n135;
  output n182;
  output n601;
  output n613;
  output n610;
  output n611;
  output n598;
  output n608;
  output n623;
  output n605;
  output n621;
  output n602;
  output n620;
  output n606;
  output n617;
  output n622;
  output n1031;
  output n1032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n136;
  wire n137;
  wire n138;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n149;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n166;
  wire n167;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n175;
  wire n176;
  wire n177;
  wire n180;
  wire n183;
  wire n184;
  wire n185;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n599;
  wire n600;
  wire n603;
  wire n604;
  wire n607;
  wire n609;
  wire n612;
  wire n614;
  wire n615;
  wire n616;
  wire n618;
  wire n619;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n87,
    n14
  );


  buf
  g1
  (
    n68,
    n17
  );


  not
  g2
  (
    n103,
    n14
  );


  not
  g3
  (
    n62,
    n2
  );


  not
  g4
  (
    n56,
    n21
  );


  not
  g5
  (
    n34,
    n20
  );


  buf
  g6
  (
    n49,
    n9
  );


  not
  g7
  (
    n53,
    n20
  );


  not
  g8
  (
    n72,
    n18
  );


  not
  g9
  (
    n117,
    n16
  );


  not
  g10
  (
    KeyWire_0_42,
    n6
  );


  buf
  g11
  (
    n79,
    n19
  );


  not
  g12
  (
    n71,
    n21
  );


  not
  g13
  (
    n108,
    n13
  );


  buf
  g14
  (
    n69,
    n9
  );


  buf
  g15
  (
    n102,
    n6
  );


  buf
  g16
  (
    n74,
    n5
  );


  buf
  g17
  (
    n38,
    n8
  );


  buf
  g18
  (
    n80,
    n10
  );


  buf
  g19
  (
    n43,
    n15
  );


  buf
  g20
  (
    n41,
    n13
  );


  buf
  g21
  (
    n110,
    n22
  );


  buf
  g22
  (
    n46,
    n23
  );


  buf
  g23
  (
    n115,
    n11
  );


  not
  g24
  (
    n113,
    n4
  );


  not
  g25
  (
    n70,
    n6
  );


  buf
  g26
  (
    n47,
    n3
  );


  buf
  g27
  (
    n109,
    n4
  );


  not
  g28
  (
    n54,
    n23
  );


  not
  g29
  (
    n86,
    n15
  );


  buf
  g30
  (
    n84,
    n23
  );


  not
  g31
  (
    n52,
    n6
  );


  not
  g32
  (
    n101,
    n7
  );


  not
  g33
  (
    n111,
    n7
  );


  buf
  g34
  (
    n104,
    n21
  );


  not
  g35
  (
    n78,
    n15
  );


  buf
  g36
  (
    n100,
    n17
  );


  not
  g37
  (
    n37,
    n11
  );


  buf
  g38
  (
    n67,
    n8
  );


  buf
  g39
  (
    n61,
    n15
  );


  not
  g40
  (
    n94,
    n17
  );


  not
  g41
  (
    n95,
    n9
  );


  not
  g42
  (
    n96,
    n5
  );


  not
  g43
  (
    n57,
    n12
  );


  not
  g44
  (
    n90,
    n24
  );


  not
  g45
  (
    n33,
    n9
  );


  not
  g46
  (
    n58,
    n13
  );


  buf
  g47
  (
    n98,
    n22
  );


  buf
  g48
  (
    n83,
    n19
  );


  not
  g49
  (
    n92,
    n20
  );


  buf
  g50
  (
    n105,
    n5
  );


  buf
  g51
  (
    n35,
    n10
  );


  not
  g52
  (
    n114,
    n16
  );


  not
  g53
  (
    n44,
    n10
  );


  buf
  g54
  (
    n75,
    n23
  );


  not
  g55
  (
    n89,
    n7
  );


  buf
  g56
  (
    n76,
    n17
  );


  buf
  g57
  (
    n106,
    n12
  );


  not
  g58
  (
    n59,
    n14
  );


  not
  g59
  (
    n107,
    n4
  );


  not
  g60
  (
    n55,
    n11
  );


  buf
  g61
  (
    n60,
    n18
  );


  buf
  g62
  (
    n42,
    n18
  );


  not
  g63
  (
    n77,
    n19
  );


  not
  g64
  (
    n88,
    n1
  );


  buf
  g65
  (
    n39,
    n21
  );


  not
  g66
  (
    n66,
    n12
  );


  not
  g67
  (
    n64,
    n14
  );


  not
  g68
  (
    n48,
    n22
  );


  not
  g69
  (
    KeyWire_0_30,
    n11
  );


  buf
  g70
  (
    n45,
    n4
  );


  buf
  g71
  (
    n51,
    n8
  );


  not
  g72
  (
    n85,
    n24
  );


  not
  g73
  (
    n93,
    n8
  );


  buf
  g74
  (
    n63,
    n13
  );


  not
  g75
  (
    n116,
    n10
  );


  not
  g76
  (
    n81,
    n16
  );


  not
  g77
  (
    n73,
    n19
  );


  not
  g78
  (
    n112,
    n20
  );


  not
  g79
  (
    n65,
    n22
  );


  buf
  g80
  (
    n36,
    n5
  );


  buf
  g81
  (
    n97,
    n7
  );


  buf
  g82
  (
    n82,
    n12
  );


  buf
  g83
  (
    n99,
    n16
  );


  not
  g84
  (
    n50,
    n18
  );


  not
  g85
  (
    n168,
    n63
  );


  not
  g86
  (
    n165,
    n75
  );


  buf
  g87
  (
    n150,
    n73
  );


  buf
  g88
  (
    n123,
    n72
  );


  not
  g89
  (
    n185,
    n56
  );


  buf
  g90
  (
    n162,
    n48
  );


  buf
  g91
  (
    n158,
    n56
  );


  buf
  g92
  (
    n147,
    n46
  );


  not
  g93
  (
    n166,
    n53
  );


  buf
  g94
  (
    n181,
    n56
  );


  not
  g95
  (
    n132,
    n65
  );


  not
  g96
  (
    n159,
    n68
  );


  buf
  g97
  (
    n167,
    n54
  );


  not
  g98
  (
    n155,
    n41
  );


  buf
  g99
  (
    n153,
    n59
  );


  not
  g100
  (
    n136,
    n75
  );


  not
  g101
  (
    n143,
    n52
  );


  not
  g102
  (
    n175,
    n63
  );


  not
  g103
  (
    n188,
    n53
  );


  buf
  g104
  (
    KeyWire_0_26,
    n63
  );


  not
  g105
  (
    n157,
    n74
  );


  buf
  g106
  (
    n196,
    n62
  );


  buf
  g107
  (
    n137,
    n53
  );


  buf
  g108
  (
    n124,
    n75
  );


  not
  g109
  (
    n141,
    n64
  );


  not
  g110
  (
    n135,
    n70
  );


  buf
  g111
  (
    n133,
    n61
  );


  not
  g112
  (
    n118,
    n55
  );


  not
  g113
  (
    n179,
    n67
  );


  buf
  g114
  (
    n160,
    n68
  );


  buf
  g115
  (
    KeyWire_0_33,
    n42
  );


  buf
  g116
  (
    n184,
    n50
  );


  buf
  g117
  (
    n134,
    n74
  );


  buf
  g118
  (
    n126,
    n35
  );


  buf
  g119
  (
    n120,
    n53
  );


  not
  g120
  (
    n163,
    n61
  );


  not
  g121
  (
    n170,
    n77
  );


  buf
  g122
  (
    n194,
    n67
  );


  not
  g123
  (
    n145,
    n70
  );


  not
  g124
  (
    n177,
    n45
  );


  not
  g125
  (
    n142,
    n46
  );


  buf
  g126
  (
    n169,
    n57
  );


  not
  g127
  (
    n139,
    n57
  );


  buf
  g128
  (
    n171,
    n50
  );


  buf
  g129
  (
    n195,
    n36
  );


  not
  g130
  (
    n154,
    n49
  );


  buf
  g131
  (
    n122,
    n50
  );


  buf
  g132
  (
    n149,
    n52
  );


  not
  g133
  (
    n173,
    n61
  );


  buf
  g134
  (
    n144,
    n76
  );


  not
  g135
  (
    n176,
    n64
  );


  buf
  g136
  (
    n183,
    n47
  );


  buf
  g137
  (
    n131,
    n59
  );


  buf
  g138
  (
    n191,
    n72
  );


  not
  g139
  (
    n182,
    n59
  );


  buf
  g140
  (
    n121,
    n60
  );


  buf
  g141
  (
    n125,
    n50
  );


  not
  g142
  (
    n129,
    n60
  );


  buf
  g143
  (
    n128,
    n58
  );


  nand
  g144
  (
    n192,
    n58,
    n55,
    n76,
    n74
  );


  nor
  g145
  (
    n146,
    n40,
    n62,
    n54,
    n77
  );


  or
  g146
  (
    n127,
    n73,
    n72,
    n51,
    n54
  );


  and
  g147
  (
    n172,
    n51,
    n65,
    n57,
    n70
  );


  nor
  g148
  (
    n164,
    n62,
    n66,
    n67,
    n46
  );


  or
  g149
  (
    n180,
    n65,
    n37,
    n69,
    n44
  );


  and
  g150
  (
    n174,
    n70,
    n51,
    n72,
    n65
  );


  nor
  g151
  (
    n189,
    n62,
    n49,
    n74,
    n46
  );


  or
  g152
  (
    KeyWire_0_48,
    n68,
    n68,
    n73,
    n33
  );


  or
  g153
  (
    KeyWire_0_49,
    n52,
    n55,
    n39,
    n48
  );


  nand
  g154
  (
    n151,
    n59,
    n71,
    n64,
    n38
  );


  nor
  g155
  (
    n152,
    n49,
    n47,
    n76,
    n58
  );


  xor
  g156
  (
    n161,
    n73,
    n71,
    n66,
    n43
  );


  xnor
  g157
  (
    n190,
    n48,
    n54,
    n60,
    n75
  );


  or
  g158
  (
    n178,
    n48,
    n66,
    n58,
    n47
  );


  nor
  g159
  (
    n187,
    n67,
    n76,
    n69,
    n60
  );


  xor
  g160
  (
    n130,
    n57,
    n71,
    n56,
    n63
  );


  or
  g161
  (
    n186,
    n49,
    n66,
    n69,
    n34
  );


  nor
  g162
  (
    n138,
    n52,
    n69,
    n47,
    n61
  );


  xor
  g163
  (
    KeyWire_0_23,
    n55,
    n71,
    n64,
    n51
  );


  not
  g164
  (
    n217,
    n162
  );


  buf
  g165
  (
    n212,
    n28
  );


  not
  g166
  (
    n221,
    n29
  );


  buf
  g167
  (
    n199,
    n79
  );


  not
  g168
  (
    n252,
    n158
  );


  buf
  g169
  (
    n232,
    n25
  );


  not
  g170
  (
    n234,
    n194
  );


  buf
  g171
  (
    KeyWire_0_12,
    n79
  );


  not
  g172
  (
    n250,
    n177
  );


  not
  g173
  (
    n254,
    n129
  );


  not
  g174
  (
    n211,
    n182
  );


  buf
  g175
  (
    n264,
    n178
  );


  not
  g176
  (
    n244,
    n146
  );


  buf
  g177
  (
    KeyWire_0_14,
    n30
  );


  buf
  g178
  (
    n262,
    n148
  );


  not
  g179
  (
    n245,
    n77
  );


  not
  g180
  (
    n243,
    n183
  );


  not
  g181
  (
    n201,
    n153
  );


  buf
  g182
  (
    KeyWire_0_24,
    n125
  );


  buf
  g183
  (
    n225,
    n144
  );


  not
  g184
  (
    n215,
    n124
  );


  not
  g185
  (
    n213,
    n136
  );


  buf
  g186
  (
    n220,
    n163
  );


  buf
  g187
  (
    n228,
    n152
  );


  not
  g188
  (
    n236,
    n128
  );


  not
  g189
  (
    n266,
    n195
  );


  buf
  g190
  (
    n202,
    n137
  );


  buf
  g191
  (
    n198,
    n150
  );


  not
  g192
  (
    n257,
    n26
  );


  buf
  g193
  (
    n261,
    n78
  );


  buf
  g194
  (
    n248,
    n196
  );


  not
  g195
  (
    n241,
    n142
  );


  buf
  g196
  (
    n223,
    n30
  );


  buf
  g197
  (
    n269,
    n191
  );


  not
  g198
  (
    n230,
    n31
  );


  not
  g199
  (
    n226,
    n186
  );


  buf
  g200
  (
    n246,
    n30
  );


  not
  g201
  (
    n216,
    n24
  );


  buf
  g202
  (
    n203,
    n161
  );


  buf
  g203
  (
    n222,
    n176
  );


  buf
  g204
  (
    n204,
    n138
  );


  buf
  g205
  (
    n206,
    n31
  );


  buf
  g206
  (
    n259,
    n25
  );


  buf
  g207
  (
    n210,
    n30
  );


  buf
  g208
  (
    n209,
    n78
  );


  not
  g209
  (
    n238,
    n193
  );


  buf
  g210
  (
    KeyWire_0_36,
    n132
  );


  not
  g211
  (
    n258,
    n80
  );


  not
  g212
  (
    n242,
    n31
  );


  buf
  g213
  (
    n205,
    n164
  );


  buf
  g214
  (
    n208,
    n160
  );


  not
  g215
  (
    n255,
    n156
  );


  or
  g216
  (
    KeyWire_0_28,
    n174,
    n135,
    n143
  );


  nor
  g217
  (
    n227,
    n26,
    n27,
    n79
  );


  nand
  g218
  (
    n197,
    n78,
    n175,
    n145
  );


  or
  g219
  (
    n267,
    n187,
    n184,
    n181
  );


  nor
  g220
  (
    n256,
    n170,
    n185,
    n31
  );


  xnor
  g221
  (
    n268,
    n192,
    n141,
    n28
  );


  and
  g222
  (
    n249,
    n189,
    n126,
    n32
  );


  nand
  g223
  (
    n200,
    n127,
    n78,
    n80
  );


  xor
  g224
  (
    n218,
    n26,
    n155,
    n168
  );


  and
  g225
  (
    n207,
    n171,
    n29
  );


  xnor
  g226
  (
    n237,
    n159,
    n180,
    n147
  );


  nor
  g227
  (
    n239,
    n134,
    n25,
    n139
  );


  or
  g228
  (
    n224,
    n133,
    n77,
    n190
  );


  xnor
  g229
  (
    n253,
    n29,
    n28,
    n79
  );


  xnor
  g230
  (
    n260,
    n27,
    n130,
    n165
  );


  nand
  g231
  (
    n219,
    n26,
    n140,
    n172
  );


  xnor
  g232
  (
    n233,
    n166,
    n167,
    n27
  );


  nor
  g233
  (
    n247,
    n157,
    n169,
    n173
  );


  nand
  g234
  (
    n235,
    n123,
    n28,
    n179
  );


  xor
  g235
  (
    n231,
    n32,
    n131,
    n154
  );


  nor
  g236
  (
    n265,
    n27,
    n149,
    n24
  );


  nor
  g237
  (
    n214,
    n188,
    n151,
    n25
  );


  not
  g238
  (
    n438,
    n99
  );


  buf
  g239
  (
    n393,
    n253
  );


  not
  g240
  (
    n428,
    n98
  );


  buf
  g241
  (
    n374,
    n242
  );


  not
  g242
  (
    KeyWire_0_25,
    n236
  );


  not
  g243
  (
    n354,
    n248
  );


  buf
  g244
  (
    n353,
    n229
  );


  not
  g245
  (
    n467,
    n84
  );


  buf
  g246
  (
    KeyWire_0_15,
    n90
  );


  buf
  g247
  (
    KeyWire_0_58,
    n234
  );


  buf
  g248
  (
    n494,
    n101
  );


  not
  g249
  (
    n462,
    n199
  );


  not
  g250
  (
    n471,
    n94
  );


  buf
  g251
  (
    n477,
    n222
  );


  not
  g252
  (
    n420,
    n208
  );


  buf
  g253
  (
    n454,
    n234
  );


  not
  g254
  (
    n280,
    n235
  );


  not
  g255
  (
    n401,
    n97
  );


  not
  g256
  (
    n434,
    n86
  );


  buf
  g257
  (
    n414,
    n109
  );


  not
  g258
  (
    n271,
    n227
  );


  buf
  g259
  (
    n491,
    n228
  );


  buf
  g260
  (
    n440,
    n264
  );


  buf
  g261
  (
    n368,
    n250
  );


  buf
  g262
  (
    n415,
    n200
  );


  not
  g263
  (
    KeyWire_0_41,
    n242
  );


  not
  g264
  (
    KeyWire_0_54,
    n84
  );


  not
  g265
  (
    n335,
    n253
  );


  buf
  g266
  (
    n442,
    n95
  );


  not
  g267
  (
    n389,
    n224
  );


  not
  g268
  (
    n383,
    n229
  );


  buf
  g269
  (
    n480,
    n102
  );


  not
  g270
  (
    n476,
    n233
  );


  buf
  g271
  (
    n326,
    n105
  );


  not
  g272
  (
    n288,
    n81
  );


  buf
  g273
  (
    n452,
    n198
  );


  buf
  g274
  (
    n427,
    n202
  );


  not
  g275
  (
    n329,
    n226
  );


  not
  g276
  (
    n364,
    n82
  );


  not
  g277
  (
    n313,
    n104
  );


  buf
  g278
  (
    KeyWire_0_19,
    n241
  );


  not
  g279
  (
    n449,
    n262
  );


  not
  g280
  (
    n277,
    n243
  );


  buf
  g281
  (
    n330,
    n209
  );


  not
  g282
  (
    n299,
    n242
  );


  buf
  g283
  (
    n404,
    n245
  );


  buf
  g284
  (
    KeyWire_0_6,
    n99
  );


  not
  g285
  (
    n387,
    n109
  );


  buf
  g286
  (
    n338,
    n213
  );


  not
  g287
  (
    n465,
    n262
  );


  buf
  g288
  (
    n334,
    n241
  );


  buf
  g289
  (
    n390,
    n99
  );


  not
  g290
  (
    n314,
    n251
  );


  not
  g291
  (
    n296,
    n239
  );


  buf
  g292
  (
    n429,
    n231
  );


  buf
  g293
  (
    n402,
    n259
  );


  not
  g294
  (
    n397,
    n248
  );


  not
  g295
  (
    n304,
    n207
  );


  not
  g296
  (
    n370,
    n270
  );


  not
  g297
  (
    n424,
    n106
  );


  buf
  g298
  (
    n305,
    n256
  );


  not
  g299
  (
    n486,
    n110
  );


  not
  g300
  (
    n351,
    n239
  );


  not
  g301
  (
    n275,
    n243
  );


  buf
  g302
  (
    n413,
    n266
  );


  buf
  g303
  (
    n483,
    n265
  );


  not
  g304
  (
    n484,
    n255
  );


  not
  g305
  (
    n380,
    n218
  );


  not
  g306
  (
    n410,
    n101
  );


  buf
  g307
  (
    KeyWire_0_8,
    n85
  );


  not
  g308
  (
    KeyWire_0_22,
    n232
  );


  not
  g309
  (
    n391,
    n211
  );


  buf
  g310
  (
    n367,
    n230
  );


  not
  g311
  (
    KeyWire_0_43,
    n254
  );


  not
  g312
  (
    n307,
    n265
  );


  buf
  g313
  (
    n319,
    n232
  );


  not
  g314
  (
    n336,
    n257
  );


  not
  g315
  (
    n388,
    n219
  );


  buf
  g316
  (
    n282,
    n103
  );


  not
  g317
  (
    n355,
    n263
  );


  not
  g318
  (
    n312,
    n233
  );


  buf
  g319
  (
    n430,
    n264
  );


  not
  g320
  (
    n488,
    n100
  );


  not
  g321
  (
    n362,
    n237
  );


  not
  g322
  (
    n448,
    n233
  );


  buf
  g323
  (
    n371,
    n214
  );


  buf
  g324
  (
    n341,
    n261
  );


  buf
  g325
  (
    n495,
    n90
  );


  buf
  g326
  (
    n392,
    n221
  );


  not
  g327
  (
    n381,
    n258
  );


  buf
  g328
  (
    n283,
    n93
  );


  buf
  g329
  (
    n363,
    n252
  );


  buf
  g330
  (
    n350,
    n241
  );


  not
  g331
  (
    n375,
    n87
  );


  not
  g332
  (
    n399,
    n208
  );


  not
  g333
  (
    n287,
    n206
  );


  buf
  g334
  (
    n366,
    n239
  );


  not
  g335
  (
    n333,
    n260
  );


  not
  g336
  (
    n411,
    n247
  );


  not
  g337
  (
    n400,
    n228
  );


  buf
  g338
  (
    n455,
    n110
  );


  buf
  g339
  (
    n479,
    n244
  );


  not
  g340
  (
    n281,
    n96
  );


  buf
  g341
  (
    n446,
    n94
  );


  not
  g342
  (
    n472,
    n265
  );


  not
  g343
  (
    n365,
    n213
  );


  buf
  g344
  (
    n290,
    n254
  );


  not
  g345
  (
    n273,
    n204
  );


  buf
  g346
  (
    n496,
    n224
  );


  buf
  g347
  (
    n426,
    n106
  );


  buf
  g348
  (
    n403,
    n204
  );


  buf
  g349
  (
    n385,
    n86
  );


  not
  g350
  (
    KeyWire_0_27,
    n229
  );


  buf
  g351
  (
    n318,
    n247
  );


  not
  g352
  (
    KeyWire_0_17,
    n249
  );


  not
  g353
  (
    n456,
    n230
  );


  buf
  g354
  (
    n379,
    n253
  );


  not
  g355
  (
    n396,
    n102
  );


  not
  g356
  (
    n492,
    n103
  );


  buf
  g357
  (
    n487,
    n109
  );


  buf
  g358
  (
    KeyWire_0_9,
    n106
  );


  not
  g359
  (
    n316,
    n205
  );


  not
  g360
  (
    n382,
    n108
  );


  not
  g361
  (
    n289,
    n92
  );


  buf
  g362
  (
    n322,
    n232
  );


  not
  g363
  (
    n278,
    n251
  );


  buf
  g364
  (
    n466,
    n212
  );


  buf
  g365
  (
    n356,
    n100
  );


  not
  g366
  (
    n418,
    n261
  );


  buf
  g367
  (
    n344,
    n97
  );


  not
  g368
  (
    n447,
    n84
  );


  buf
  g369
  (
    n272,
    n268
  );


  not
  g370
  (
    n464,
    n265
  );


  not
  g371
  (
    n274,
    n89
  );


  buf
  g372
  (
    n310,
    n108
  );


  buf
  g373
  (
    n470,
    n270
  );


  buf
  g374
  (
    n332,
    n105
  );


  not
  g375
  (
    n433,
    n223
  );


  buf
  g376
  (
    n352,
    n215
  );


  not
  g377
  (
    n419,
    n89
  );


  buf
  g378
  (
    n405,
    n106
  );


  not
  g379
  (
    n317,
    n227
  );


  buf
  g380
  (
    n417,
    n215
  );


  not
  g381
  (
    n302,
    n235
  );


  not
  g382
  (
    n489,
    n97
  );


  not
  g383
  (
    n345,
    n232
  );


  buf
  g384
  (
    n359,
    n110
  );


  buf
  g385
  (
    KeyWire_0_39,
    n259
  );


  buf
  g386
  (
    n327,
    n246
  );


  not
  g387
  (
    KeyWire_0_37,
    n95
  );


  buf
  g388
  (
    n349,
    n255
  );


  not
  g389
  (
    n279,
    n86
  );


  not
  g390
  (
    n340,
    n268
  );


  not
  g391
  (
    n298,
    n85
  );


  buf
  g392
  (
    KeyWire_0_62,
    n81
  );


  not
  g393
  (
    n445,
    n91
  );


  not
  g394
  (
    KeyWire_0_21,
    n217
  );


  not
  g395
  (
    n478,
    n248
  );


  buf
  g396
  (
    n421,
    n235
  );


  buf
  g397
  (
    n301,
    n107
  );


  not
  g398
  (
    n431,
    n230
  );


  not
  g399
  (
    n311,
    n269
  );


  not
  g400
  (
    n407,
    n205
  );


  buf
  g401
  (
    n451,
    n262
  );


  buf
  g402
  (
    n343,
    n105
  );


  buf
  g403
  (
    n463,
    n236
  );


  buf
  g404
  (
    n291,
    n210
  );


  buf
  g405
  (
    KeyWire_0_47,
    n231
  );


  not
  g406
  (
    n315,
    n266
  );


  not
  g407
  (
    n384,
    n97
  );


  not
  g408
  (
    n457,
    n212
  );


  buf
  g409
  (
    n303,
    n258
  );


  not
  g410
  (
    n460,
    n240
  );


  not
  g411
  (
    n328,
    n85
  );


  not
  g412
  (
    n453,
    n228
  );


  not
  g413
  (
    n450,
    n92
  );


  buf
  g414
  (
    n300,
    n95
  );


  not
  g415
  (
    n323,
    n94
  );


  buf
  g416
  (
    n295,
    n201
  );


  buf
  g417
  (
    n376,
    n259
  );


  not
  g418
  (
    n475,
    n237
  );


  buf
  g419
  (
    n294,
    n256
  );


  buf
  g420
  (
    n468,
    n216
  );


  buf
  g421
  (
    n412,
    n245
  );


  not
  g422
  (
    n276,
    n108
  );


  buf
  g423
  (
    n409,
    n90
  );


  and
  g424
  (
    n459,
    n84,
    n222
  );


  nor
  g425
  (
    n439,
    n82,
    n98,
    n250,
    n260
  );


  nand
  g426
  (
    n432,
    n268,
    n236,
    n251,
    n233
  );


  nand
  g427
  (
    n284,
    n107,
    n259,
    n231,
    n267
  );


  xor
  g428
  (
    n378,
    n255,
    n85,
    n80,
    n269
  );


  nor
  g429
  (
    n360,
    n226,
    n254,
    n266
  );


  and
  g430
  (
    n493,
    n100,
    n245,
    n257,
    n95
  );


  and
  g431
  (
    n297,
    n83,
    n82,
    n87,
    n91
  );


  and
  g432
  (
    n425,
    n255,
    n107,
    n240,
    n92
  );


  nand
  g433
  (
    n285,
    n98,
    n108,
    n238,
    n223
  );


  nor
  g434
  (
    n416,
    n234,
    n96,
    n237,
    n264
  );


  nor
  g435
  (
    n320,
    n104,
    n245,
    n218,
    n225
  );


  xnor
  g436
  (
    n481,
    n239,
    n241,
    n105,
    n92
  );


  xnor
  g437
  (
    n342,
    n96,
    n104,
    n263,
    n94
  );


  or
  g438
  (
    n293,
    n261,
    n250,
    n257,
    n91
  );


  or
  g439
  (
    n461,
    n98,
    n89,
    n263,
    n221
  );


  xor
  g440
  (
    n325,
    n249,
    n269,
    n246,
    n253
  );


  and
  g441
  (
    n485,
    n100,
    n83,
    n90,
    n88
  );


  or
  g442
  (
    n443,
    n209,
    n99,
    n249,
    n88
  );


  xor
  g443
  (
    n398,
    n268,
    n87,
    n235,
    n230
  );


  and
  g444
  (
    n358,
    n263,
    n270,
    n81,
    n210
  );


  or
  g445
  (
    n339,
    n219,
    n93,
    n91,
    n270
  );


  or
  g446
  (
    n394,
    n248,
    n261,
    n211,
    n249
  );


  nor
  g447
  (
    n406,
    n254,
    n238,
    n203,
    n243
  );


  or
  g448
  (
    n482,
    n267,
    n225,
    n238,
    n103
  );


  and
  g449
  (
    n458,
    n220,
    n247,
    n206,
    n229
  );


  xor
  g450
  (
    n331,
    n246,
    n217,
    n260,
    n236
  );


  or
  g451
  (
    n357,
    n247,
    n197,
    n82,
    n252
  );


  nand
  g452
  (
    n369,
    n101,
    n252,
    n244,
    n264
  );


  and
  g453
  (
    n337,
    n81,
    n207,
    n258,
    n256
  );


  and
  g454
  (
    n435,
    n267,
    n214,
    n252,
    n107
  );


  nor
  g455
  (
    n473,
    n267,
    n251,
    n87,
    n88
  );


  nor
  g456
  (
    n347,
    n240,
    n101,
    n244,
    n109
  );


  or
  g457
  (
    n437,
    n220,
    n244,
    n269,
    n93
  );


  nand
  g458
  (
    n292,
    n256,
    n83,
    n250,
    n231
  );


  or
  g459
  (
    n373,
    n243,
    n88,
    n102,
    n260
  );


  nor
  g460
  (
    n309,
    n103,
    n89,
    n83,
    n234
  );


  or
  g461
  (
    n474,
    n262,
    n104,
    n240,
    n228
  );


  nand
  g462
  (
    n469,
    n242,
    n216,
    n96,
    n257
  );


  xor
  g463
  (
    n348,
    n238,
    n93,
    n80,
    n237
  );


  and
  g464
  (
    n286,
    n246,
    n258,
    n86,
    n102
  );


  buf
  g465
  (
    n527,
    n275
  );


  not
  g466
  (
    n511,
    n291
  );


  buf
  g467
  (
    n528,
    n285
  );


  not
  g468
  (
    n522,
    n283
  );


  buf
  g469
  (
    n512,
    n300
  );


  not
  g470
  (
    n521,
    n279
  );


  buf
  g471
  (
    n506,
    n293
  );


  buf
  g472
  (
    n513,
    n276
  );


  buf
  g473
  (
    n504,
    n278
  );


  not
  g474
  (
    n499,
    n286
  );


  not
  g475
  (
    KeyWire_0_20,
    n296
  );


  buf
  g476
  (
    n503,
    n290
  );


  not
  g477
  (
    n523,
    n284
  );


  not
  g478
  (
    n520,
    n274
  );


  buf
  g479
  (
    n517,
    n271
  );


  not
  g480
  (
    n500,
    n280
  );


  not
  g481
  (
    n507,
    n287
  );


  not
  g482
  (
    n501,
    n298
  );


  buf
  g483
  (
    n519,
    n282
  );


  not
  g484
  (
    n518,
    n277
  );


  not
  g485
  (
    n505,
    n288
  );


  buf
  g486
  (
    n515,
    n289
  );


  buf
  g487
  (
    n526,
    n302
  );


  buf
  g488
  (
    n508,
    n297
  );


  not
  g489
  (
    n525,
    n281
  );


  not
  g490
  (
    n498,
    n292
  );


  buf
  g491
  (
    n509,
    n272
  );


  buf
  g492
  (
    n524,
    n294
  );


  buf
  g493
  (
    n502,
    n273
  );


  not
  g494
  (
    n514,
    n299
  );


  buf
  g495
  (
    n529,
    n301
  );


  buf
  g496
  (
    n510,
    n295
  );


  not
  g497
  (
    n566,
    n501
  );


  not
  g498
  (
    n558,
    n514
  );


  buf
  g499
  (
    KeyWire_0_35,
    n506
  );


  buf
  g500
  (
    n544,
    n505
  );


  not
  g501
  (
    n569,
    n499
  );


  buf
  g502
  (
    n568,
    n498
  );


  not
  g503
  (
    n563,
    n508
  );


  not
  g504
  (
    n545,
    n508
  );


  buf
  g505
  (
    n553,
    n511
  );


  not
  g506
  (
    n530,
    n498
  );


  not
  g507
  (
    n540,
    n512
  );


  not
  g508
  (
    n531,
    n506
  );


  not
  g509
  (
    n535,
    n502
  );


  not
  g510
  (
    n561,
    n506
  );


  buf
  g511
  (
    n549,
    n111
  );


  buf
  g512
  (
    n552,
    n499
  );


  buf
  g513
  (
    n536,
    n512
  );


  buf
  g514
  (
    KeyWire_0_2,
    n510
  );


  not
  g515
  (
    n548,
    n506
  );


  not
  g516
  (
    n550,
    n511
  );


  buf
  g517
  (
    n538,
    n505
  );


  buf
  g518
  (
    n537,
    n510
  );


  buf
  g519
  (
    n560,
    n503
  );


  not
  g520
  (
    n554,
    n498
  );


  buf
  g521
  (
    n567,
    n503
  );


  not
  g522
  (
    n562,
    n500
  );


  nand
  g523
  (
    n556,
    n513,
    n503
  );


  xor
  g524
  (
    n557,
    n515,
    n513
  );


  and
  g525
  (
    n555,
    n511,
    n514,
    n508,
    n515
  );


  or
  g526
  (
    n534,
    n515,
    n507,
    n511,
    n508
  );


  or
  g527
  (
    n547,
    n502,
    n507,
    n110,
    n505
  );


  nor
  g528
  (
    n533,
    n500,
    n509,
    n502,
    n501
  );


  nor
  g529
  (
    n564,
    n516,
    n498,
    n510,
    n505
  );


  or
  g530
  (
    n546,
    n507,
    n509,
    n514,
    n512
  );


  or
  g531
  (
    n565,
    n510,
    n507,
    n499,
    n512
  );


  or
  g532
  (
    n551,
    n509,
    n500,
    n504
  );


  nand
  g533
  (
    n539,
    n501,
    n502,
    n516,
    n513
  );


  nand
  g534
  (
    KeyWire_0_18,
    n509,
    n504,
    n499,
    n501
  );


  nand
  g535
  (
    n542,
    n513,
    n111,
    n516,
    n500
  );


  nand
  g536
  (
    n532,
    n514,
    n515,
    n503,
    n504
  );


  not
  g537
  (
    n570,
    n542
  );


  buf
  g538
  (
    n578,
    n532
  );


  buf
  g539
  (
    n583,
    n531
  );


  not
  g540
  (
    n575,
    n535
  );


  not
  g541
  (
    n572,
    n530
  );


  not
  g542
  (
    n584,
    n536
  );


  not
  g543
  (
    n574,
    n541
  );


  not
  g544
  (
    n571,
    n537
  );


  buf
  g545
  (
    n573,
    n543
  );


  not
  g546
  (
    n576,
    n533
  );


  not
  g547
  (
    n585,
    n534
  );


  buf
  g548
  (
    n579,
    n539
  );


  buf
  g549
  (
    n581,
    n545
  );


  buf
  g550
  (
    KeyWire_0_29,
    n544
  );


  not
  g551
  (
    n580,
    n540
  );


  not
  g552
  (
    KeyWire_0_16,
    n538
  );


  buf
  g553
  (
    n587,
    n304
  );


  buf
  g554
  (
    n594,
    n576
  );


  buf
  g555
  (
    n595,
    n305
  );


  not
  g556
  (
    n588,
    n578
  );


  nor
  g557
  (
    n591,
    n573,
    n303
  );


  xor
  g558
  (
    n589,
    n306,
    n570
  );


  and
  g559
  (
    n593,
    n571,
    n572
  );


  and
  g560
  (
    n586,
    n575,
    n579
  );


  xnor
  g561
  (
    n592,
    n577,
    n111
  );


  nor
  g562
  (
    n590,
    n574,
    n111
  );


  not
  g563
  (
    n608,
    n516
  );


  not
  g564
  (
    n599,
    n590
  );


  not
  g565
  (
    n613,
    n592
  );


  not
  g566
  (
    n612,
    n588
  );


  not
  g567
  (
    n601,
    n587
  );


  not
  g568
  (
    n606,
    n590
  );


  buf
  g569
  (
    n609,
    n587
  );


  not
  g570
  (
    n617,
    n590
  );


  buf
  g571
  (
    n623,
    n593
  );


  not
  g572
  (
    n596,
    n591
  );


  not
  g573
  (
    n610,
    n589
  );


  buf
  g574
  (
    n598,
    n588
  );


  buf
  g575
  (
    n614,
    n589
  );


  not
  g576
  (
    n615,
    n586
  );


  buf
  g577
  (
    n604,
    n586
  );


  not
  g578
  (
    n616,
    n591
  );


  not
  g579
  (
    n620,
    n592
  );


  buf
  g580
  (
    n619,
    n589
  );


  not
  g581
  (
    n602,
    n593
  );


  buf
  g582
  (
    n618,
    n587
  );


  buf
  g583
  (
    n605,
    n587
  );


  not
  g584
  (
    n622,
    n588
  );


  buf
  g585
  (
    n624,
    n517
  );


  buf
  g586
  (
    n625,
    n591
  );


  not
  g587
  (
    n597,
    n590
  );


  buf
  g588
  (
    n621,
    n588
  );


  buf
  g589
  (
    n603,
    n586
  );


  buf
  g590
  (
    n607,
    n586
  );


  buf
  g591
  (
    n600,
    n592
  );


  nor
  g592
  (
    n611,
    n591,
    n592,
    n589
  );


  buf
  g593
  (
    n631,
    n313
  );


  buf
  g594
  (
    n637,
    n551
  );


  buf
  g595
  (
    n629,
    n552
  );


  buf
  g596
  (
    n636,
    n563
  );


  or
  g597
  (
    n630,
    n564,
    n615,
    n549,
    n613
  );


  and
  g598
  (
    n627,
    n311,
    n557,
    n610,
    n618
  );


  or
  g599
  (
    n632,
    n619,
    n585,
    n622,
    n546
  );


  xor
  g600
  (
    n634,
    n556,
    n555,
    n580,
    n560
  );


  nand
  g601
  (
    n638,
    n620,
    n582,
    n307,
    n616
  );


  xor
  g602
  (
    n628,
    n553,
    n562,
    n315,
    n581
  );


  or
  g603
  (
    KeyWire_0_57,
    n617,
    n312,
    n316,
    n317
  );


  and
  g604
  (
    n633,
    n314,
    n561,
    n548,
    n624
  );


  nor
  g605
  (
    KeyWire_0_56,
    n583,
    n547,
    n612,
    n310
  );


  xnor
  g606
  (
    n640,
    n614,
    n584,
    n550,
    n621
  );


  nor
  g607
  (
    n639,
    n309,
    n559,
    n623,
    n554
  );


  nand
  g608
  (
    n641,
    n611,
    n308,
    n558,
    n625
  );


  not
  g609
  (
    n644,
    n631
  );


  buf
  g610
  (
    n647,
    n630
  );


  buf
  g611
  (
    n643,
    n629
  );


  buf
  g612
  (
    n650,
    n628
  );


  buf
  g613
  (
    n649,
    n323
  );


  buf
  g614
  (
    n646,
    n632
  );


  not
  g615
  (
    n651,
    n320
  );


  not
  g616
  (
    n642,
    n322
  );


  and
  g617
  (
    n645,
    n319,
    n626,
    n318,
    n629
  );


  or
  g618
  (
    n648,
    n630,
    n627,
    n631,
    n321
  );


  not
  g619
  (
    n661,
    n648
  );


  buf
  g620
  (
    n654,
    n646
  );


  nor
  g621
  (
    n653,
    n645,
    n326,
    n651,
    n334
  );


  xnor
  g622
  (
    n656,
    n333,
    n642,
    n644,
    n518
  );


  and
  g623
  (
    n657,
    n332,
    n325,
    n517
  );


  nor
  g624
  (
    n655,
    n335,
    n329,
    n520,
    n519
  );


  nand
  g625
  (
    n652,
    n328,
    n519,
    n518,
    n651
  );


  and
  g626
  (
    n658,
    n647,
    n643,
    n650,
    n519
  );


  or
  g627
  (
    n660,
    n518,
    n518,
    n331,
    n520
  );


  xor
  g628
  (
    n662,
    n520,
    n519,
    n324,
    n327
  );


  nand
  g629
  (
    n659,
    n517,
    n520,
    n330,
    n649
  );


  buf
  g630
  (
    n667,
    n638
  );


  buf
  g631
  (
    n673,
    n568
  );


  buf
  g632
  (
    KeyWire_0_40,
    n633
  );


  not
  g633
  (
    n697,
    n659
  );


  not
  g634
  (
    n703,
    n344
  );


  not
  g635
  (
    n688,
    n566
  );


  not
  g636
  (
    KeyWire_0_38,
    n639
  );


  buf
  g637
  (
    n666,
    n113
  );


  buf
  g638
  (
    n680,
    n657
  );


  buf
  g639
  (
    n699,
    n662
  );


  buf
  g640
  (
    n692,
    n656
  );


  buf
  g641
  (
    n690,
    n653
  );


  not
  g642
  (
    n681,
    n654
  );


  not
  g643
  (
    n685,
    n112
  );


  buf
  g644
  (
    n686,
    n112
  );


  buf
  g645
  (
    n678,
    n654
  );


  not
  g646
  (
    n689,
    n652
  );


  not
  g647
  (
    n705,
    n658
  );


  buf
  g648
  (
    n693,
    n660
  );


  buf
  g649
  (
    n683,
    n640
  );


  buf
  g650
  (
    n675,
    n113
  );


  not
  g651
  (
    n665,
    n637
  );


  buf
  g652
  (
    KeyWire_0_1,
    n660
  );


  buf
  g653
  (
    n701,
    n635
  );


  not
  g654
  (
    n679,
    n634
  );


  buf
  g655
  (
    n663,
    n636
  );


  and
  g656
  (
    n695,
    n658,
    n347,
    n661,
    n345
  );


  nand
  g657
  (
    n698,
    n338,
    n343,
    n662
  );


  nor
  g658
  (
    KeyWire_0_50,
    n112,
    n653,
    n641
  );


  xor
  g659
  (
    n669,
    n639,
    n661,
    n635,
    n640
  );


  or
  g660
  (
    n691,
    n636,
    n348,
    n653,
    n654
  );


  nand
  g661
  (
    n706,
    n652,
    n354,
    n353,
    n340
  );


  nand
  g662
  (
    n676,
    n656,
    n652,
    n339,
    n352
  );


  nor
  g663
  (
    n664,
    n641,
    n351,
    n652,
    n569
  );


  xnor
  g664
  (
    n671,
    n341,
    n659,
    n655,
    n657
  );


  and
  g665
  (
    n672,
    n656,
    n634,
    n655
  );


  and
  g666
  (
    KeyWire_0_55,
    n637,
    n114,
    n342,
    n349
  );


  nor
  g667
  (
    n696,
    n337,
    n657,
    n658
  );


  and
  g668
  (
    n670,
    n350,
    n654,
    n632,
    n656
  );


  or
  g669
  (
    n668,
    n638,
    n355,
    n659,
    n567
  );


  nor
  g670
  (
    n674,
    n346,
    n662,
    n565,
    n660
  );


  xor
  g671
  (
    n700,
    n336,
    n655,
    n661,
    n113
  );


  nor
  g672
  (
    n684,
    n113,
    n660,
    n114,
    n633
  );


  and
  g673
  (
    n687,
    n657,
    n661,
    n659,
    n112
  );


  nor
  g674
  (
    n747,
    n464,
    n436,
    n473,
    n684
  );


  and
  g675
  (
    n744,
    n474,
    n454,
    n448,
    n463
  );


  xnor
  g676
  (
    n746,
    n389,
    n481,
    n356,
    n415
  );


  and
  g677
  (
    n728,
    n467,
    n685,
    n452,
    n381
  );


  and
  g678
  (
    n709,
    n453,
    n481,
    n458,
    n444
  );


  and
  g679
  (
    n754,
    n479,
    n663,
    n373,
    n482
  );


  xor
  g680
  (
    n712,
    n486,
    n694,
    n469,
    n693
  );


  and
  g681
  (
    n742,
    n363,
    n691,
    n382,
    n686
  );


  xor
  g682
  (
    n768,
    n688,
    n455,
    n458,
    n478
  );


  nor
  g683
  (
    n745,
    n457,
    n476,
    n695,
    n452
  );


  nand
  g684
  (
    n753,
    n481,
    n685,
    n466,
    n693
  );


  and
  g685
  (
    KeyWire_0_44,
    n372,
    n683,
    n692,
    n481
  );


  nor
  g686
  (
    n785,
    n446,
    n687,
    n406,
    n423
  );


  or
  g687
  (
    n711,
    n429,
    n681,
    n689,
    n470
  );


  nor
  g688
  (
    n765,
    n485,
    n487,
    n455,
    n365
  );


  and
  g689
  (
    n735,
    n433,
    n469,
    n487,
    n402
  );


  xor
  g690
  (
    n770,
    n439,
    n370,
    n443,
    n690
  );


  xnor
  g691
  (
    n707,
    n412,
    n692,
    n394,
    n671
  );


  or
  g692
  (
    n763,
    n366,
    n479,
    n453,
    n386
  );


  xor
  g693
  (
    n760,
    n692,
    n420,
    n427,
    n694
  );


  nand
  g694
  (
    n714,
    n688,
    n404,
    n418,
    n486
  );


  and
  g695
  (
    KeyWire_0_59,
    n459,
    n688,
    n457,
    n484
  );


  and
  g696
  (
    n741,
    n424,
    n673,
    n685,
    n475
  );


  or
  g697
  (
    n776,
    n422,
    n395,
    n474,
    n469
  );


  or
  g698
  (
    n772,
    n466,
    n689,
    n442,
    n683
  );


  or
  g699
  (
    n736,
    n425,
    n387,
    n460,
    n691
  );


  xor
  g700
  (
    n748,
    n447,
    n693,
    n465,
    n455
  );


  xnor
  g701
  (
    n771,
    n397,
    n441,
    n377,
    n446
  );


  and
  g702
  (
    n758,
    n362,
    n456,
    n470,
    n467
  );


  nor
  g703
  (
    n780,
    n693,
    n694,
    n376,
    n477
  );


  or
  g704
  (
    n775,
    n449,
    n476,
    n459,
    n695
  );


  xnor
  g705
  (
    n731,
    n385,
    n676,
    n691,
    n480
  );


  xor
  g706
  (
    n730,
    n485,
    n692,
    n465,
    n411
  );


  or
  g707
  (
    n749,
    n465,
    n485,
    n471,
    n478
  );


  xor
  g708
  (
    n743,
    n468,
    n456,
    n681,
    n460
  );


  nand
  g709
  (
    n764,
    n407,
    n694,
    n487,
    n484
  );


  xor
  g710
  (
    n724,
    n431,
    n450,
    n674,
    n413
  );


  and
  g711
  (
    n729,
    n438,
    n446,
    n368,
    n448
  );


  xor
  g712
  (
    n738,
    n393,
    n419,
    n483,
    n461
  );


  xor
  g713
  (
    n786,
    n375,
    n447,
    n474,
    n484
  );


  xor
  g714
  (
    n727,
    n401,
    n690,
    n450,
    n379
  );


  nand
  g715
  (
    n719,
    n471,
    n687,
    n417,
    n400
  );


  or
  g716
  (
    n721,
    n440,
    n677,
    n408,
    n484
  );


  xnor
  g717
  (
    n722,
    n460,
    n468,
    n388,
    n467
  );


  nand
  g718
  (
    n732,
    n466,
    n472,
    n688
  );


  xnor
  g719
  (
    n781,
    n434,
    n696,
    n390,
    n462
  );


  nand
  g720
  (
    n774,
    n474,
    n432,
    n680,
    n687
  );


  xnor
  g721
  (
    n710,
    n462,
    n684,
    n454,
    n686
  );


  and
  g722
  (
    n769,
    n384,
    n480,
    n478,
    n471
  );


  nor
  g723
  (
    n756,
    n466,
    n683,
    n396,
    n691
  );


  or
  g724
  (
    n761,
    n416,
    n695,
    n479,
    n469
  );


  xnor
  g725
  (
    n708,
    n409,
    n430,
    n684,
    n453
  );


  xor
  g726
  (
    n767,
    n398,
    n482,
    n463,
    n451
  );


  xnor
  g727
  (
    n726,
    n454,
    n451,
    n445,
    n480
  );


  xnor
  g728
  (
    n750,
    n449,
    n479,
    n360,
    n472
  );


  nor
  g729
  (
    n762,
    n477,
    n374,
    n681,
    n403
  );


  or
  g730
  (
    n725,
    n696,
    n392,
    n668,
    n447
  );


  and
  g731
  (
    n733,
    n486,
    n686,
    n359,
    n480
  );


  xor
  g732
  (
    n766,
    n378,
    n468,
    n391,
    n690
  );


  xnor
  g733
  (
    n720,
    n421,
    n670,
    n483,
    n459
  );


  or
  g734
  (
    n734,
    n426,
    n364,
    n461,
    n678
  );


  nand
  g735
  (
    n784,
    n399,
    n369,
    n477,
    n682
  );


  xor
  g736
  (
    n715,
    n451,
    n471,
    n665,
    n683
  );


  xnor
  g737
  (
    n752,
    n465,
    n666,
    n357,
    n695
  );


  and
  g738
  (
    n723,
    n667,
    n468,
    n470,
    n696
  );


  nand
  g739
  (
    n779,
    n669,
    n358,
    n482,
    n684
  );


  nor
  g740
  (
    n759,
    n690,
    n682,
    n475
  );


  xnor
  g741
  (
    n777,
    n414,
    n467,
    n696,
    n470
  );


  xor
  g742
  (
    n782,
    n458,
    n380,
    n435,
    n685
  );


  or
  g743
  (
    n718,
    n371,
    n475,
    n473,
    n449
  );


  xor
  g744
  (
    KeyWire_0_0,
    n672,
    n452,
    n461,
    n457
  );


  xor
  g745
  (
    n713,
    n463,
    n464,
    n478,
    n361
  );


  and
  g746
  (
    n739,
    n448,
    n689,
    n383
  );


  and
  g747
  (
    n737,
    n456,
    n428,
    n487,
    n686
  );


  xnor
  g748
  (
    n716,
    n473,
    n477,
    n464,
    n367
  );


  or
  g749
  (
    n751,
    n405,
    n464,
    n664,
    n462
  );


  and
  g750
  (
    n783,
    n482,
    n483,
    n472,
    n675
  );


  xor
  g751
  (
    n717,
    n679,
    n476,
    n485,
    n450
  );


  and
  g752
  (
    n778,
    n437,
    n473,
    n483,
    n410
  );


  nand
  g753
  (
    n757,
    n486,
    n475,
    n687,
    n476
  );


  buf
  g754
  (
    n842,
    n758
  );


  not
  g755
  (
    KeyWire_0_61,
    n114
  );


  not
  g756
  (
    n797,
    n723
  );


  not
  g757
  (
    n942,
    n728
  );


  buf
  g758
  (
    n795,
    n747
  );


  buf
  g759
  (
    n863,
    n725
  );


  not
  g760
  (
    n798,
    n785
  );


  not
  g761
  (
    n843,
    n523
  );


  not
  g762
  (
    n883,
    n117
  );


  not
  g763
  (
    n933,
    n715
  );


  not
  g764
  (
    n849,
    n716
  );


  not
  g765
  (
    n817,
    n521
  );


  buf
  g766
  (
    n917,
    n527
  );


  buf
  g767
  (
    n877,
    n769
  );


  buf
  g768
  (
    n929,
    n741
  );


  not
  g769
  (
    n836,
    n731
  );


  not
  g770
  (
    n846,
    n784
  );


  not
  g771
  (
    n810,
    n732
  );


  not
  g772
  (
    n901,
    n720
  );


  not
  g773
  (
    n946,
    n528
  );


  not
  g774
  (
    n805,
    n762
  );


  not
  g775
  (
    n879,
    n521
  );


  not
  g776
  (
    n923,
    n773
  );


  not
  g777
  (
    n804,
    n710
  );


  not
  g778
  (
    n918,
    n595
  );


  not
  g779
  (
    n889,
    n528
  );


  buf
  g780
  (
    n848,
    n760
  );


  buf
  g781
  (
    KeyWire_0_45,
    n753
  );


  not
  g782
  (
    n893,
    n525
  );


  not
  g783
  (
    n847,
    n758
  );


  not
  g784
  (
    n818,
    n748
  );


  not
  g785
  (
    n807,
    n723
  );


  buf
  g786
  (
    n854,
    n785
  );


  not
  g787
  (
    n834,
    n756
  );


  buf
  g788
  (
    n788,
    n770
  );


  not
  g789
  (
    n868,
    n765
  );


  not
  g790
  (
    n808,
    n116
  );


  buf
  g791
  (
    n799,
    n761
  );


  not
  g792
  (
    n900,
    n734
  );


  buf
  g793
  (
    n855,
    n724
  );


  buf
  g794
  (
    n878,
    n709
  );


  buf
  g795
  (
    KeyWire_0_46,
    n718
  );


  not
  g796
  (
    n895,
    n780
  );


  not
  g797
  (
    n794,
    n751
  );


  buf
  g798
  (
    n914,
    n752
  );


  not
  g799
  (
    n845,
    n736
  );


  not
  g800
  (
    KeyWire_0_34,
    n742
  );


  buf
  g801
  (
    n857,
    n743
  );


  not
  g802
  (
    n821,
    n709
  );


  buf
  g803
  (
    n884,
    n755
  );


  buf
  g804
  (
    n861,
    n526
  );


  nor
  g805
  (
    n856,
    n766,
    n724,
    n593
  );


  nand
  g806
  (
    n882,
    n747,
    n730,
    n710
  );


  xnor
  g807
  (
    n787,
    n736,
    n525,
    n732
  );


  nor
  g808
  (
    n947,
    n766,
    n744,
    n738
  );


  nor
  g809
  (
    n791,
    n708,
    n722,
    n733
  );


  nor
  g810
  (
    n892,
    n748,
    n765,
    n784
  );


  xor
  g811
  (
    n824,
    n779,
    n755,
    n708
  );


  xnor
  g812
  (
    n871,
    n786,
    n526,
    n726
  );


  xor
  g813
  (
    n819,
    n786,
    n782,
    n719
  );


  xnor
  g814
  (
    n922,
    n716,
    n734,
    n743
  );


  nor
  g815
  (
    n872,
    n748,
    n529,
    n751
  );


  and
  g816
  (
    n812,
    n712,
    n771,
    n707
  );


  and
  g817
  (
    n909,
    n711,
    n783,
    n772
  );


  nand
  g818
  (
    n809,
    n774,
    n767,
    n735
  );


  nor
  g819
  (
    n875,
    n714,
    n716,
    n776
  );


  and
  g820
  (
    n865,
    n594,
    n726,
    n773
  );


  xnor
  g821
  (
    n858,
    n768,
    n780,
    n734
  );


  xnor
  g822
  (
    n935,
    n725,
    n764,
    n752
  );


  xor
  g823
  (
    n938,
    n715,
    n594,
    n523
  );


  nand
  g824
  (
    n862,
    n760,
    n719,
    n529
  );


  and
  g825
  (
    n851,
    n786,
    n779,
    n526
  );


  nand
  g826
  (
    KeyWire_0_3,
    n738,
    n737,
    n707
  );


  and
  g827
  (
    n860,
    n763,
    n757,
    n713
  );


  nor
  g828
  (
    KeyWire_0_51,
    n778,
    n116,
    n763
  );


  and
  g829
  (
    n925,
    n729,
    n524,
    n750
  );


  xor
  g830
  (
    n880,
    n780,
    n767,
    n521
  );


  xnor
  g831
  (
    n859,
    n739,
    n748,
    n728
  );


  xnor
  g832
  (
    n790,
    n718,
    n713,
    n759
  );


  or
  g833
  (
    n850,
    n766,
    n781,
    n711
  );


  xnor
  g834
  (
    n939,
    n735,
    n762,
    n754
  );


  or
  g835
  (
    n853,
    n744,
    n773,
    n761
  );


  or
  g836
  (
    n913,
    n711,
    n732,
    n766
  );


  xnor
  g837
  (
    n800,
    n115,
    n729,
    n720
  );


  nand
  g838
  (
    n873,
    n746,
    n744,
    n736
  );


  and
  g839
  (
    n911,
    n708,
    n733,
    n709
  );


  and
  g840
  (
    n813,
    n741,
    n528,
    n746
  );


  and
  g841
  (
    n910,
    n727,
    n742,
    n751
  );


  nor
  g842
  (
    n874,
    n750,
    n32,
    n761
  );


  or
  g843
  (
    n932,
    n760,
    n749,
    n719
  );


  xor
  g844
  (
    n915,
    n117,
    n728,
    n716
  );


  nor
  g845
  (
    n830,
    n764,
    n755
  );


  nand
  g846
  (
    n891,
    n771,
    n739,
    n707
  );


  or
  g847
  (
    KeyWire_0_52,
    n731,
    n753,
    n757
  );


  xnor
  g848
  (
    n890,
    n722,
    n115,
    n727
  );


  nor
  g849
  (
    n886,
    n115,
    n739,
    n754
  );


  and
  g850
  (
    n927,
    n594,
    n752,
    n730
  );


  xor
  g851
  (
    n803,
    n743,
    n774,
    n778
  );


  xor
  g852
  (
    n814,
    n785,
    n723,
    n777
  );


  and
  g853
  (
    n820,
    n721,
    n525,
    n723
  );


  or
  g854
  (
    n904,
    n775,
    n529,
    n759
  );


  xor
  g855
  (
    n796,
    n763,
    n773,
    n751
  );


  and
  g856
  (
    n816,
    n749,
    n772,
    n725
  );


  nand
  g857
  (
    KeyWire_0_11,
    n744,
    n522,
    n732
  );


  or
  g858
  (
    n907,
    n117,
    n762,
    n743
  );


  xor
  g859
  (
    n888,
    n730,
    n754,
    n722
  );


  xor
  g860
  (
    n827,
    n756,
    n772,
    n738
  );


  xor
  g861
  (
    n792,
    n786,
    n781,
    n718
  );


  xnor
  g862
  (
    n941,
    n726,
    n775,
    n720
  );


  nor
  g863
  (
    n898,
    n775,
    n729,
    n745
  );


  or
  g864
  (
    n839,
    n771,
    n774,
    n772
  );


  nand
  g865
  (
    n815,
    n720,
    n721,
    n768
  );


  xnor
  g866
  (
    n885,
    n767,
    n746,
    n770
  );


  and
  g867
  (
    n934,
    n595,
    n760,
    n741
  );


  nor
  g868
  (
    n829,
    n717,
    n759,
    n710
  );


  xor
  g869
  (
    n823,
    n768,
    n745,
    n737
  );


  nor
  g870
  (
    n926,
    n528,
    n724,
    n524
  );


  nand
  g871
  (
    n806,
    n781,
    n777,
    n769
  );


  nand
  g872
  (
    n930,
    n776,
    n737,
    n750
  );


  xor
  g873
  (
    n887,
    n758,
    n594,
    n721
  );


  or
  g874
  (
    n905,
    n764,
    n742,
    n747
  );


  nor
  g875
  (
    n825,
    n741,
    n115,
    n725
  );


  and
  g876
  (
    n896,
    n527,
    n783,
    n522
  );


  nor
  g877
  (
    n940,
    n708,
    n521,
    n117
  );


  and
  g878
  (
    n936,
    n722,
    n759,
    n526
  );


  and
  g879
  (
    n833,
    n761,
    n775,
    n770
  );


  nand
  g880
  (
    n919,
    n595,
    n739,
    n782
  );


  xnor
  g881
  (
    n944,
    n758,
    n713,
    n523
  );


  nand
  g882
  (
    n831,
    n740,
    n769,
    n733
  );


  and
  g883
  (
    n876,
    n745,
    n779,
    n774
  );


  nand
  g884
  (
    n864,
    n756,
    n529,
    n731
  );


  xnor
  g885
  (
    n943,
    n746,
    n740,
    n724
  );


  xor
  g886
  (
    n826,
    n707,
    n714,
    n522
  );


  and
  g887
  (
    n822,
    n765,
    n735,
    n727
  );


  or
  g888
  (
    n881,
    n777,
    n778,
    n769
  );


  and
  g889
  (
    n852,
    n733,
    n753,
    n757
  );


  xnor
  g890
  (
    n921,
    n771,
    n765,
    n747
  );


  xor
  g891
  (
    n899,
    n784,
    n735,
    n742
  );


  nor
  g892
  (
    n866,
    n523,
    n712
  );


  nand
  g893
  (
    n903,
    n736,
    n715,
    n721
  );


  and
  g894
  (
    n924,
    n776,
    n731,
    n734
  );


  xor
  g895
  (
    n916,
    n726,
    n527,
    n714
  );


  nand
  g896
  (
    n912,
    n525,
    n776,
    n768
  );


  and
  g897
  (
    n908,
    n709,
    n756,
    n752
  );


  xnor
  g898
  (
    n867,
    n737,
    n717,
    n783
  );


  xnor
  g899
  (
    n841,
    n712,
    n782,
    n717
  );


  xor
  g900
  (
    n837,
    n116,
    n715,
    n714
  );


  xnor
  g901
  (
    n838,
    n729,
    n749,
    n753
  );


  nor
  g902
  (
    n811,
    n719,
    n767,
    n717
  );


  and
  g903
  (
    n793,
    n738,
    n764,
    n749
  );


  xnor
  g904
  (
    n840,
    n711,
    n740,
    n763
  );


  xor
  g905
  (
    n802,
    n783,
    n730,
    n785
  );


  or
  g906
  (
    n844,
    n116,
    n778,
    n524
  );


  nand
  g907
  (
    n789,
    n114,
    n784,
    n728
  );


  nand
  g908
  (
    n828,
    n757,
    n740,
    n782
  );


  nor
  g909
  (
    n835,
    n595,
    n780,
    n754
  );


  nor
  g910
  (
    n937,
    n524,
    n777,
    n522
  );


  nand
  g911
  (
    KeyWire_0_31,
    n593,
    n781,
    n718
  );


  or
  g912
  (
    KeyWire_0_7,
    n762,
    n770,
    n779
  );


  and
  g913
  (
    n920,
    n727,
    n710,
    n750
  );


  xor
  g914
  (
    KeyWire_0_10,
    n527,
    n713,
    n745
  );


  xor
  g915
  (
    KeyWire_0_5,
    n808,
    n832,
    n793,
    n799
  );


  or
  g916
  (
    n950,
    n792,
    n787,
    n813,
    n836
  );


  xnor
  g917
  (
    n960,
    n830,
    n820,
    n842,
    n841
  );


  xor
  g918
  (
    n965,
    n816,
    n851,
    n814,
    n803
  );


  nor
  g919
  (
    n952,
    n806,
    n801,
    n800,
    n797
  );


  xnor
  g920
  (
    n956,
    n837,
    n789,
    n818,
    n809
  );


  or
  g921
  (
    n961,
    n810,
    n858,
    n833,
    n825
  );


  xor
  g922
  (
    n964,
    n850,
    n848,
    n802,
    n839
  );


  xnor
  g923
  (
    n963,
    n791,
    n828,
    n854,
    n855
  );


  xnor
  g924
  (
    n949,
    n852,
    n788,
    n821,
    n815
  );


  and
  g925
  (
    n957,
    n845,
    n838,
    n844,
    n847
  );


  xnor
  g926
  (
    n951,
    n846,
    n811,
    n795,
    n831
  );


  and
  g927
  (
    n959,
    n840,
    n857,
    n796,
    n849
  );


  and
  g928
  (
    n955,
    n819,
    n804,
    n817,
    n843
  );


  or
  g929
  (
    n958,
    n822,
    n790,
    n835,
    n827
  );


  xor
  g930
  (
    n962,
    n829,
    n826,
    n853,
    n834
  );


  and
  g931
  (
    n954,
    n824,
    n807,
    n805,
    n856
  );


  or
  g932
  (
    n948,
    n812,
    n798,
    n823,
    n794
  );


  nor
  g933
  (
    n979,
    n698,
    n965,
    n699,
    n701
  );


  or
  g934
  (
    n980,
    n948,
    n701,
    n495,
    n489
  );


  nor
  g935
  (
    n975,
    n497,
    n492,
    n704,
    n960
  );


  or
  g936
  (
    n976,
    n953,
    n488,
    n961,
    n702
  );


  or
  g937
  (
    n972,
    n699,
    n964,
    n493,
    n494
  );


  xnor
  g938
  (
    n984,
    n698,
    n496,
    n963,
    n700
  );


  xor
  g939
  (
    n966,
    n491,
    n495,
    n961,
    n706
  );


  and
  g940
  (
    n991,
    n697,
    n963,
    n706,
    n960
  );


  nand
  g941
  (
    n978,
    n706,
    n495,
    n700,
    n704
  );


  xor
  g942
  (
    n967,
    n698,
    n702,
    n959,
    n496
  );


  nor
  g943
  (
    KeyWire_0_4,
    n494,
    n703,
    n962,
    n497
  );


  nor
  g944
  (
    KeyWire_0_60,
    n699,
    n962,
    n955,
    n704
  );


  xnor
  g945
  (
    KeyWire_0_32,
    n700,
    n702,
    n494,
    n705
  );


  nand
  g946
  (
    n970,
    n957,
    n490,
    n962,
    n956
  );


  nor
  g947
  (
    n974,
    n490,
    n697,
    n965
  );


  nand
  g948
  (
    n983,
    n706,
    n491,
    n959,
    n497
  );


  xnor
  g949
  (
    n993,
    n494,
    n949,
    n488,
    n493
  );


  nor
  g950
  (
    n977,
    n951,
    n497,
    n963,
    n699
  );


  xnor
  g951
  (
    n985,
    n493,
    n952,
    n964,
    n488
  );


  nand
  g952
  (
    n986,
    n492,
    n496,
    n488,
    n701
  );


  xnor
  g953
  (
    n988,
    n950,
    n961,
    n489,
    n700
  );


  or
  g954
  (
    n982,
    n964,
    n965,
    n489,
    n490
  );


  xnor
  g955
  (
    n969,
    n492,
    n958,
    n705,
    n703
  );


  nand
  g956
  (
    n968,
    n960,
    n954,
    n701,
    n496
  );


  and
  g957
  (
    n973,
    n493,
    n703,
    n705,
    n698
  );


  or
  g958
  (
    n981,
    n704,
    n492,
    n702,
    n958
  );


  nand
  g959
  (
    n971,
    n697,
    n703,
    n490,
    n495
  );


  xor
  g960
  (
    n990,
    n489,
    n705,
    n491
  );


  nand
  g961
  (
    KeyWire_0_13,
    n922,
    n897,
    n918,
    n875
  );


  nand
  g962
  (
    n1010,
    n990,
    n879,
    n930,
    n914
  );


  nand
  g963
  (
    KeyWire_0_63,
    n873,
    n887,
    n920,
    n933
  );


  or
  g964
  (
    n999,
    n970,
    n945,
    n984,
    n971
  );


  nand
  g965
  (
    n1017,
    n862,
    n924,
    n928,
    n888
  );


  or
  g966
  (
    n996,
    n934,
    n940,
    n869,
    n890
  );


  or
  g967
  (
    n998,
    n884,
    n892,
    n880,
    n923
  );


  xnor
  g968
  (
    n1012,
    n909,
    n885,
    n966,
    n896
  );


  or
  g969
  (
    n1021,
    n878,
    n931,
    n944,
    n900
  );


  or
  g970
  (
    n1005,
    n993,
    n906,
    n988,
    n893
  );


  xnor
  g971
  (
    n1008,
    n883,
    n886,
    n937,
    n908
  );


  nand
  g972
  (
    n1016,
    n912,
    n904,
    n927,
    n972
  );


  or
  g973
  (
    n1014,
    n867,
    n877,
    n868,
    n973
  );


  and
  g974
  (
    n1022,
    n982,
    n943,
    n939,
    n986
  );


  nand
  g975
  (
    n1006,
    n874,
    n974,
    n917,
    n864
  );


  or
  g976
  (
    n1004,
    n872,
    n921,
    n975,
    n901
  );


  xnor
  g977
  (
    n1009,
    n915,
    n905,
    n898,
    n895
  );


  xor
  g978
  (
    n1001,
    n891,
    n882,
    n976,
    n938
  );


  xnor
  g979
  (
    KeyWire_0_53,
    n910,
    n981,
    n870,
    n942
  );


  nand
  g980
  (
    n1013,
    n993,
    n983,
    n935,
    n916
  );


  and
  g981
  (
    n997,
    n936,
    n866,
    n894,
    n978
  );


  or
  g982
  (
    n1007,
    n989,
    n863,
    n871,
    n926
  );


  and
  g983
  (
    n1002,
    n987,
    n903,
    n876,
    n977
  );


  xor
  g984
  (
    n1020,
    n985,
    n980,
    n865,
    n899
  );


  xnor
  g985
  (
    n995,
    n979,
    n889,
    n992,
    n907
  );


  nor
  g986
  (
    n1011,
    n991,
    n929,
    n859,
    n860
  );


  or
  g987
  (
    n1019,
    n881,
    n969,
    n941,
    n919
  );


  nor
  g988
  (
    n1018,
    n967,
    n913,
    n932,
    n968
  );


  nor
  g989
  (
    n994,
    n911,
    n902,
    n861,
    n925
  );


  nor
  g990
  (
    n1028,
    n1019,
    n1013,
    n1006,
    n1002
  );


  nor
  g991
  (
    n1026,
    n1001,
    n1014,
    n999,
    n1015
  );


  or
  g992
  (
    n1024,
    n998,
    n996,
    n1022,
    n1000
  );


  xnor
  g993
  (
    n1029,
    n1008,
    n1021,
    n995,
    n1017
  );


  nor
  g994
  (
    n1023,
    n1007,
    n1003,
    n1018,
    n997
  );


  or
  g995
  (
    n1027,
    n1005,
    n32,
    n994,
    n1010
  );


  and
  g996
  (
    n1030,
    n1016,
    n1012,
    n947,
    n1009
  );


  xor
  g997
  (
    n1025,
    n1020,
    n946,
    n1004,
    n1011
  );


  nor
  g998
  (
    n1032,
    n1030,
    n1027,
    n1028,
    n1024
  );


  xnor
  g999
  (
    n1031,
    n1029,
    n1025,
    n1026,
    n1023
  );


  xnor
  KeyGate_0_0
  (
    n755,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n677,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n541,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n801,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n987,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n953,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n490,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n897,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n306,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n441,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n870,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n869,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n229,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1000,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n240,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n497,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n577,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n422,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n543,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n423,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n516,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n308,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n436,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n140,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n270,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n408,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n193,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n372,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n263,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n582,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n91,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n928,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n989,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n119,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n894,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n559,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n251,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n321,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n704,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n386,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n702,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n444,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n40,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n324,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n740,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n945,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n902,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n346,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n156,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n148,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n694,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n832,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n931,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1015,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n395,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n682,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n626,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n635,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n361,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n773,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n992,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n906,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n377,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n1003,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

