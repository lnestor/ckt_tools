

module Stat_114_49
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n130,
  n118,
  n131,
  n123,
  n115,
  n117,
  n114,
  n120,
  n128,
  n121,
  n119,
  n126,
  n129,
  n124,
  n116,
  n125,
  n127,
  n122,
  n113,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;
  output n130;output n118;output n131;output n123;output n115;output n117;output n114;output n120;output n128;output n121;output n119;output n126;output n129;output n124;output n116;output n125;output n127;output n122;output n113;
  wire n18;wire n19;wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n32,
    n17
  );


  buf
  g1
  (
    n26,
    n7
  );


  buf
  g2
  (
    n20,
    n11
  );


  not
  g3
  (
    n24,
    n6
  );


  not
  g4
  (
    n18,
    n9
  );


  buf
  g5
  (
    n25,
    n17
  );


  buf
  g6
  (
    n23,
    n12
  );


  buf
  g7
  (
    n28,
    n15
  );


  buf
  g8
  (
    n30,
    n14
  );


  not
  g9
  (
    n35,
    n13
  );


  buf
  g10
  (
    n27,
    n10
  );


  not
  g11
  (
    n22,
    n16
  );


  buf
  g12
  (
    n34,
    n5
  );


  not
  g13
  (
    n33,
    n3
  );


  buf
  g14
  (
    n21,
    n1
  );


  buf
  g15
  (
    n19,
    n4
  );


  buf
  g16
  (
    n31,
    n2
  );


  buf
  g17
  (
    n29,
    n8
  );


  not
  g18
  (
    n41,
    n31
  );


  buf
  g19
  (
    n63,
    n34
  );


  not
  g20
  (
    n43,
    n24
  );


  not
  g21
  (
    n65,
    n20
  );


  buf
  g22
  (
    n52,
    n27
  );


  not
  g23
  (
    n39,
    n35
  );


  not
  g24
  (
    n64,
    n19
  );


  buf
  g25
  (
    n49,
    n26
  );


  not
  g26
  (
    n42,
    n24
  );


  buf
  g27
  (
    n45,
    n35
  );


  not
  g28
  (
    n36,
    n27
  );


  not
  g29
  (
    n48,
    n29
  );


  not
  g30
  (
    n72,
    n30
  );


  buf
  g31
  (
    n50,
    n35
  );


  not
  g32
  (
    n60,
    n31
  );


  not
  g33
  (
    n70,
    n33
  );


  buf
  g34
  (
    n55,
    n22
  );


  not
  g35
  (
    n44,
    n18
  );


  not
  g36
  (
    n66,
    n29
  );


  not
  g37
  (
    n61,
    n23
  );


  not
  g38
  (
    n37,
    n22
  );


  buf
  g39
  (
    n68,
    n18
  );


  not
  g40
  (
    n40,
    n34
  );


  not
  g41
  (
    n47,
    n28
  );


  not
  g42
  (
    n56,
    n34
  );


  buf
  g43
  (
    n69,
    n25
  );


  not
  g44
  (
    n38,
    n30
  );


  buf
  g45
  (
    n58,
    n20
  );


  buf
  g46
  (
    n51,
    n19
  );


  buf
  g47
  (
    n57,
    n33
  );


  buf
  g48
  (
    n73,
    n28
  );


  buf
  g49
  (
    n62,
    n23
  );


  buf
  g50
  (
    n54,
    n32
  );


  not
  g51
  (
    n46,
    n21
  );


  not
  g52
  (
    n67,
    n26
  );


  not
  g53
  (
    n71,
    n21
  );


  buf
  g54
  (
    n53,
    n32
  );


  not
  g55
  (
    n59,
    n25
  );


  not
  g56
  (
    n76,
    n49
  );


  not
  g57
  (
    n104,
    n68
  );


  buf
  g58
  (
    n100,
    n39
  );


  buf
  g59
  (
    n107,
    n38
  );


  buf
  g60
  (
    n74,
    n55
  );


  buf
  g61
  (
    n106,
    n43
  );


  not
  g62
  (
    n94,
    n37
  );


  buf
  g63
  (
    n92,
    n42
  );


  buf
  g64
  (
    n90,
    n51
  );


  not
  g65
  (
    n75,
    n65
  );


  buf
  g66
  (
    n83,
    n66
  );


  not
  g67
  (
    n112,
    n60
  );


  not
  g68
  (
    n103,
    n64
  );


  buf
  g69
  (
    n91,
    n53
  );


  buf
  g70
  (
    n78,
    n69
  );


  not
  g71
  (
    n93,
    n40
  );


  buf
  g72
  (
    n97,
    n72
  );


  not
  g73
  (
    n96,
    n36
  );


  buf
  g74
  (
    n85,
    n46
  );


  buf
  g75
  (
    n98,
    n48
  );


  not
  g76
  (
    n79,
    n71
  );


  buf
  g77
  (
    n88,
    n57
  );


  buf
  g78
  (
    n105,
    n73
  );


  buf
  g79
  (
    n89,
    n58
  );


  not
  g80
  (
    n99,
    n61
  );


  buf
  g81
  (
    n101,
    n41
  );


  buf
  g82
  (
    n102,
    n54
  );


  not
  g83
  (
    n86,
    n59
  );


  not
  g84
  (
    n77,
    n52
  );


  not
  g85
  (
    n84,
    n67
  );


  not
  g86
  (
    n110,
    n73
  );


  not
  g87
  (
    n80,
    n63
  );


  buf
  g88
  (
    n87,
    n62
  );


  buf
  g89
  (
    n109,
    n56
  );


  buf
  g90
  (
    n82,
    n50
  );


  not
  g91
  (
    n111,
    n70
  );


  not
  g92
  (
    n108,
    n44
  );


  buf
  g93
  (
    n81,
    n45
  );


  not
  g94
  (
    n95,
    n47
  );


  not
  g95
  (
    n115,
    n88
  );


  buf
  g96
  (
    n123,
    n108
  );


  not
  g97
  (
    n129,
    n107
  );


  buf
  g98
  (
    n124,
    n106
  );


  buf
  g99
  (
    n119,
    n75
  );


  buf
  g100
  (
    n128,
    n100
  );


  buf
  g101
  (
    n126,
    n98
  );


  buf
  g102
  (
    n131,
    n78
  );


  not
  g103
  (
    n125,
    n82
  );


  not
  g104
  (
    AntiSAT_key_wire,
    n93
  );


  not
  g105
  (
    n127,
    n110
  );


  not
  g106
  (
    n121,
    n94
  );


  xnor
  g107
  (
    n116,
    n105,
    n101,
    n92
  );


  xor
  g108
  (
    n130,
    n102,
    n109,
    n87,
    n96
  );


  and
  g109
  (
    n118,
    n91,
    n97,
    n77,
    n99
  );


  xor
  g110
  (
    n114,
    n80,
    n90,
    n76,
    n79
  );


  nor
  g111
  (
    n117,
    n74,
    n111,
    n95,
    n83
  );


  nand
  g112
  (
    n113,
    n81,
    n104,
    n112,
    n86
  );


  or
  g113
  (
    n122,
    n84,
    n103,
    n89,
    n85
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_17
  (
    gbar_input_0_0,
    keyIn_0_17,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_18
  (
    gbar_input_0_1,
    keyIn_0_18,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_19
  (
    gbar_input_0_2,
    keyIn_0_19,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_20
  (
    gbar_input_0_3,
    keyIn_0_20,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_21
  (
    gbar_input_0_4,
    keyIn_0_21,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_22
  (
    gbar_input_0_5,
    keyIn_0_22,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_23
  (
    gbar_input_0_6,
    keyIn_0_23,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_24
  (
    gbar_input_0_7,
    keyIn_0_24,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_25
  (
    gbar_input_0_8,
    keyIn_0_25,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_9,
    keyIn_0_26,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_10,
    keyIn_0_27,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_11,
    keyIn_0_28,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_12,
    keyIn_0_29,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_13,
    keyIn_0_30,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_14,
    keyIn_0_31,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_15,
    keyIn_0_32,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_16,
    keyIn_0_33,
    n17
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n120,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

