

module Stat_100_52
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n62,
  n48,
  n126,
  n122,
  n129,
  n104,
  n113,
  n117,
  n123,
  n115,
  n110,
  n111,
  n116,
  n105,
  n112,
  n132,
  n118,
  n120,
  n125,
  n103,
  n128,
  n109,
  n127,
  n121,
  n107,
  n130,
  n106,
  n124,
  n114,
  n119,
  n131,
  n108
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n62;output n48;output n126;output n122;output n129;output n104;output n113;output n117;output n123;output n115;output n110;output n111;output n116;output n105;output n112;output n132;output n118;output n120;output n125;output n103;output n128;output n109;output n127;output n121;output n107;output n130;output n106;output n124;output n114;output n119;output n131;output n108;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;

  buf
  g0
  (
    n41,
    n2
  );


  buf
  g1
  (
    KeyWire_0_56,
    n2
  );


  not
  g2
  (
    n38,
    n3
  );


  not
  g3
  (
    KeyWire_0_21,
    n1
  );


  buf
  g4
  (
    n39,
    n2
  );


  not
  g5
  (
    KeyWire_0_53,
    n1
  );


  not
  g6
  (
    KeyWire_0_55,
    n1
  );


  buf
  g7
  (
    KeyWire_0_3,
    n2
  );


  not
  g8
  (
    n42,
    n1
  );


  buf
  g9
  (
    n33,
    n3
  );


  xnor
  g10
  (
    KeyWire_0_36,
    n32,
    n10
  );


  and
  g11
  (
    KeyWire_0_28,
    n36,
    n39,
    n14,
    n25
  );


  and
  g12
  (
    KeyWire_0_11,
    n17,
    n7,
    n32,
    n28
  );


  xor
  g13
  (
    n62,
    n30,
    n14,
    n13,
    n4
  );


  xor
  g14
  (
    KeyWire_0_63,
    n18,
    n8,
    n31,
    n42
  );


  xnor
  g15
  (
    n66,
    n22,
    n26,
    n23,
    n20
  );


  nor
  g16
  (
    n73,
    n5,
    n33,
    n16,
    n22
  );


  xnor
  g17
  (
    KeyWire_0_48,
    n10,
    n31,
    n11,
    n12
  );


  xnor
  g18
  (
    KeyWire_0_54,
    n11,
    n25,
    n32,
    n35
  );


  or
  g19
  (
    n57,
    n6,
    n15,
    n29,
    n10
  );


  and
  g20
  (
    n52,
    n11,
    n28,
    n36,
    n15
  );


  nand
  g21
  (
    n61,
    n4,
    n19,
    n21
  );


  nor
  g22
  (
    KeyWire_0_26,
    n31,
    n11,
    n23,
    n42
  );


  or
  g23
  (
    n71,
    n38,
    n35,
    n3,
    n25
  );


  and
  g24
  (
    KeyWire_0_12,
    n23,
    n24,
    n15,
    n34
  );


  nand
  g25
  (
    n79,
    n30,
    n21,
    n28,
    n34
  );


  xor
  g26
  (
    KeyWire_0_44,
    n39,
    n6,
    n22,
    n14
  );


  and
  g27
  (
    KeyWire_0_39,
    n33,
    n26,
    n18,
    n6
  );


  or
  g28
  (
    KeyWire_0_35,
    n30,
    n20,
    n23,
    n26
  );


  or
  g29
  (
    n68,
    n42,
    n12,
    n9,
    n20
  );


  nor
  g30
  (
    n82,
    n19,
    n36,
    n18,
    n8
  );


  xnor
  g31
  (
    KeyWire_0_37,
    n17,
    n8,
    n18,
    n38
  );


  xnor
  g32
  (
    n74,
    n19,
    n13,
    n22,
    n5
  );


  nand
  g33
  (
    n45,
    n17,
    n40,
    n16
  );


  nand
  g34
  (
    n70,
    n28,
    n39,
    n13,
    n26
  );


  xor
  g35
  (
    KeyWire_0_17,
    n7,
    n31,
    n6,
    n24
  );


  nand
  g36
  (
    KeyWire_0_13,
    n20,
    n33,
    n3,
    n27
  );


  or
  g37
  (
    KeyWire_0_43,
    n19,
    n5,
    n41,
    n24
  );


  and
  g38
  (
    KeyWire_0_19,
    n37,
    n39,
    n4,
    n41
  );


  and
  g39
  (
    KeyWire_0_45,
    n16,
    n7,
    n42,
    n35
  );


  nor
  g40
  (
    KeyWire_0_20,
    n9,
    n37,
    n32,
    n34
  );


  or
  g41
  (
    n65,
    n37,
    n9,
    n29,
    n35
  );


  and
  g42
  (
    KeyWire_0_9,
    n24,
    n4,
    n17,
    n12
  );


  nand
  g43
  (
    KeyWire_0_34,
    n8,
    n33,
    n15,
    n16
  );


  xor
  g44
  (
    n50,
    n29,
    n27,
    n38
  );


  xnor
  g45
  (
    KeyWire_0_15,
    n36,
    n9,
    n5,
    n25
  );


  nand
  g46
  (
    KeyWire_0_30,
    n14,
    n37,
    n40,
    n10
  );


  xnor
  g47
  (
    KeyWire_0_29,
    n27,
    n40,
    n30,
    n34
  );


  nand
  g48
  (
    n59,
    n38,
    n29,
    n13,
    n21
  );


  xnor
  g49
  (
    KeyWire_0_32,
    n12,
    n7,
    n41
  );


  buf
  g50
  (
    KeyWire_0_33,
    n45
  );


  buf
  g51
  (
    KeyWire_0_1,
    n46
  );


  not
  g52
  (
    KeyWire_0_52,
    n47
  );


  buf
  g53
  (
    KeyWire_0_14,
    n48
  );


  nor
  g54
  (
    n92,
    n58,
    n56,
    n50,
    n53
  );


  and
  g55
  (
    KeyWire_0_59,
    n50,
    n60,
    n52
  );


  or
  g56
  (
    n90,
    n84,
    n58,
    n51,
    n83
  );


  and
  g57
  (
    KeyWire_0_51,
    n50,
    n53,
    n55,
    n52
  );


  or
  g58
  (
    KeyWire_0_16,
    n85,
    n59,
    n55
  );


  xor
  g59
  (
    KeyWire_0_31,
    n58,
    n86,
    n52,
    n56
  );


  xnor
  g60
  (
    KeyWire_0_41,
    n59,
    n51,
    n60,
    n54
  );


  xnor
  g61
  (
    KeyWire_0_61,
    n53,
    n54,
    n55,
    n57
  );


  and
  g62
  (
    n102,
    n86,
    n52,
    n83,
    n59
  );


  xnor
  g63
  (
    KeyWire_0_60,
    n84,
    n85,
    n56,
    n57
  );


  xor
  g64
  (
    n97,
    n54,
    n84,
    n51
  );


  xor
  g65
  (
    KeyWire_0_47,
    n83,
    n53,
    n58,
    n54
  );


  nand
  g66
  (
    n94,
    n86,
    n85,
    n49
  );


  xor
  g67
  (
    KeyWire_0_7,
    n59,
    n57,
    n49,
    n60
  );


  xor
  g68
  (
    KeyWire_0_46,
    n50,
    n51,
    n56,
    n49
  );


  and
  g69
  (
    n91,
    n86,
    n85,
    n57,
    n83
  );


  nand
  g70
  (
    KeyWire_0_2,
    n81,
    n63,
    n66,
    n96
  );


  nand
  g71
  (
    n115,
    n81,
    n101,
    n66,
    n69
  );


  nor
  g72
  (
    n110,
    n62,
    n100,
    n71,
    n69
  );


  xnor
  g73
  (
    KeyWire_0_42,
    n68,
    n100,
    n74,
    n99
  );


  nand
  g74
  (
    KeyWire_0_8,
    n98,
    n99,
    n82,
    n101
  );


  nand
  g75
  (
    KeyWire_0_58,
    n72,
    n61,
    n102,
    n78
  );


  and
  g76
  (
    KeyWire_0_5,
    n68,
    n100,
    n82,
    n64
  );


  nor
  g77
  (
    n107,
    n74,
    n67,
    n75,
    n98
  );


  or
  g78
  (
    n117,
    n71,
    n65,
    n99,
    n80
  );


  or
  g79
  (
    KeyWire_0_50,
    n74,
    n75,
    n91,
    n87
  );


  xor
  g80
  (
    KeyWire_0_0,
    n95,
    n68,
    n63,
    n73
  );


  nand
  g81
  (
    n109,
    n94,
    n77,
    n89,
    n102
  );


  xnor
  g82
  (
    KeyWire_0_27,
    n69,
    n71,
    n79,
    n65
  );


  xnor
  g83
  (
    KeyWire_0_24,
    n93,
    n100,
    n102,
    n61
  );


  nor
  g84
  (
    KeyWire_0_4,
    n80,
    n76,
    n98,
    n90
  );


  xnor
  g85
  (
    KeyWire_0_38,
    n68,
    n76,
    n65
  );


  xnor
  g86
  (
    n125,
    n72,
    n66,
    n98,
    n77
  );


  nand
  g87
  (
    KeyWire_0_22,
    n80,
    n82,
    n73,
    n71
  );


  xor
  g88
  (
    n128,
    n74,
    n79,
    n70,
    n88
  );


  xnor
  g89
  (
    KeyWire_0_40,
    n72,
    n73,
    n75,
    n76
  );


  xnor
  g90
  (
    n124,
    n78,
    n70,
    n101,
    n72
  );


  xnor
  g91
  (
    KeyWire_0_49,
    n92,
    n64,
    n67
  );


  xnor
  g92
  (
    KeyWire_0_23,
    n67,
    n63,
    n79,
    n65
  );


  xor
  g93
  (
    KeyWire_0_10,
    n62,
    n78,
    n99,
    n70
  );


  xnor
  g94
  (
    KeyWire_0_57,
    n82,
    n63,
    n62,
    n73
  );


  and
  g95
  (
    KeyWire_0_18,
    n97,
    n62,
    n77,
    n81
  );


  xnor
  g96
  (
    KeyWire_0_6,
    n79,
    n102,
    n66,
    n80
  );


  xnor
  g97
  (
    KeyWire_0_25,
    n101,
    n81,
    n97,
    n61
  );


  xor
  g98
  (
    n129,
    n70,
    n67,
    n64,
    n61
  );


  nand
  g99
  (
    KeyWire_0_62,
    n77,
    n78,
    n69,
    n75
  );


  xnor
  KeyGate_0_0
  (
    n123,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n86,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n126,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n40,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n113,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n118,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n127,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n87,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n119,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n47,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n114,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n46,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n43,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n69,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n84,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n54,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n99,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n58,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n121,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n60,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n51,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n35,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n111,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n105,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n104,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n116,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n67,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n112,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n63,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n77,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n49,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n88,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n64,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n85,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n80,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n48,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n56,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n78,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n131,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n72,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n106,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n95,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n103,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n75,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n55,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n53,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n101,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n89,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n76,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n130,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n120,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n100,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n83,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n34,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n81,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n36,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n37,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n122,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n132,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n96,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n98,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n93,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n108,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n44,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


