

module Stat_1000_206
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n415,
  n417,
  n1027,
  n1008,
  n1003,
  n1025,
  n1004,
  n1010,
  n1032,
  n1023,
  n1016,
  n1024,
  n1009,
  n1028,
  n1022,
  n1031,
  n1006,
  n1011,
  n1021,
  n1014,
  n1015,
  n1013,
  n1012,
  n1018,
  n1017,
  n1029,
  n1005,
  n1026,
  n1030,
  n1007,
  n1020,
  n1019,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n415;output n417;output n1027;output n1008;output n1003;output n1025;output n1004;output n1010;output n1032;output n1023;output n1016;output n1024;output n1009;output n1028;output n1022;output n1031;output n1006;output n1011;output n1021;output n1014;output n1015;output n1013;output n1012;output n1018;output n1017;output n1029;output n1005;output n1026;output n1030;output n1007;output n1020;output n1019;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n416;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n49,
    n17
  );


  buf
  g1
  (
    n134,
    n8
  );


  not
  g2
  (
    n85,
    n18
  );


  not
  g3
  (
    n145,
    n1
  );


  not
  g4
  (
    n153,
    n12
  );


  not
  g5
  (
    n143,
    n13
  );


  not
  g6
  (
    n34,
    n28
  );


  not
  g7
  (
    n140,
    n28
  );


  not
  g8
  (
    n142,
    n19
  );


  not
  g9
  (
    n36,
    n7
  );


  not
  g10
  (
    n107,
    n11
  );


  not
  g11
  (
    n117,
    n2
  );


  not
  g12
  (
    n38,
    n19
  );


  not
  g13
  (
    n52,
    n9
  );


  not
  g14
  (
    n148,
    n27
  );


  not
  g15
  (
    n64,
    n11
  );


  not
  g16
  (
    n46,
    n3
  );


  buf
  g17
  (
    n35,
    n24
  );


  not
  g18
  (
    n86,
    n1
  );


  buf
  g19
  (
    n56,
    n9
  );


  buf
  g20
  (
    n151,
    n6
  );


  buf
  g21
  (
    n100,
    n22
  );


  not
  g22
  (
    n108,
    n25
  );


  buf
  g23
  (
    n115,
    n16
  );


  not
  g24
  (
    n103,
    n3
  );


  buf
  g25
  (
    n91,
    n17
  );


  buf
  g26
  (
    n104,
    n4
  );


  not
  g27
  (
    n39,
    n22
  );


  buf
  g28
  (
    n126,
    n18
  );


  buf
  g29
  (
    n132,
    n25
  );


  not
  g30
  (
    n51,
    n29
  );


  not
  g31
  (
    n138,
    n29
  );


  not
  g32
  (
    n106,
    n30
  );


  buf
  g33
  (
    n99,
    n23
  );


  buf
  g34
  (
    n72,
    n31
  );


  buf
  g35
  (
    n123,
    n3
  );


  buf
  g36
  (
    n120,
    n26
  );


  buf
  g37
  (
    n124,
    n28
  );


  not
  g38
  (
    n77,
    n24
  );


  buf
  g39
  (
    n88,
    n20
  );


  not
  g40
  (
    n139,
    n17
  );


  not
  g41
  (
    n48,
    n16
  );


  buf
  g42
  (
    n121,
    n10
  );


  buf
  g43
  (
    n42,
    n18
  );


  not
  g44
  (
    n112,
    n13
  );


  not
  g45
  (
    n61,
    n16
  );


  not
  g46
  (
    n147,
    n24
  );


  buf
  g47
  (
    n69,
    n20
  );


  buf
  g48
  (
    n92,
    n23
  );


  not
  g49
  (
    n81,
    n14
  );


  buf
  g50
  (
    n131,
    n21
  );


  not
  g51
  (
    n89,
    n25
  );


  not
  g52
  (
    n156,
    n7
  );


  not
  g53
  (
    n129,
    n1
  );


  not
  g54
  (
    n111,
    n23
  );


  not
  g55
  (
    n109,
    n2
  );


  not
  g56
  (
    n90,
    n8
  );


  not
  g57
  (
    n67,
    n26
  );


  buf
  g58
  (
    n58,
    n22
  );


  not
  g59
  (
    n40,
    n6
  );


  not
  g60
  (
    n33,
    n26
  );


  not
  g61
  (
    n119,
    n2
  );


  buf
  g62
  (
    n66,
    n15
  );


  buf
  g63
  (
    n75,
    n13
  );


  not
  g64
  (
    n74,
    n28
  );


  not
  g65
  (
    n80,
    n15
  );


  not
  g66
  (
    n57,
    n14
  );


  not
  g67
  (
    n68,
    n4
  );


  buf
  g68
  (
    n135,
    n21
  );


  buf
  g69
  (
    n60,
    n26
  );


  buf
  g70
  (
    n84,
    n2
  );


  not
  g71
  (
    n47,
    n31
  );


  buf
  g72
  (
    n141,
    n19
  );


  not
  g73
  (
    n110,
    n4
  );


  not
  g74
  (
    n136,
    n5
  );


  buf
  g75
  (
    n95,
    n15
  );


  buf
  g76
  (
    n144,
    n24
  );


  buf
  g77
  (
    n118,
    n21
  );


  buf
  g78
  (
    n114,
    n6
  );


  not
  g79
  (
    n63,
    n31
  );


  not
  g80
  (
    n97,
    n29
  );


  buf
  g81
  (
    n127,
    n13
  );


  buf
  g82
  (
    n43,
    n30
  );


  not
  g83
  (
    n93,
    n3
  );


  not
  g84
  (
    n53,
    n11
  );


  not
  g85
  (
    n65,
    n9
  );


  not
  g86
  (
    n59,
    n10
  );


  buf
  g87
  (
    n44,
    n12
  );


  buf
  g88
  (
    n78,
    n1
  );


  not
  g89
  (
    n87,
    n14
  );


  buf
  g90
  (
    n45,
    n30
  );


  buf
  g91
  (
    n150,
    n27
  );


  not
  g92
  (
    n154,
    n6
  );


  buf
  g93
  (
    n102,
    n16
  );


  buf
  g94
  (
    n73,
    n9
  );


  buf
  g95
  (
    n41,
    n11
  );


  not
  g96
  (
    n155,
    n5
  );


  not
  g97
  (
    n137,
    n10
  );


  buf
  g98
  (
    n94,
    n25
  );


  buf
  g99
  (
    n70,
    n8
  );


  not
  g100
  (
    n125,
    n29
  );


  buf
  g101
  (
    n152,
    n5
  );


  buf
  g102
  (
    n101,
    n12
  );


  buf
  g103
  (
    n71,
    n20
  );


  buf
  g104
  (
    n76,
    n15
  );


  not
  g105
  (
    n54,
    n17
  );


  buf
  g106
  (
    n96,
    n31
  );


  buf
  g107
  (
    n146,
    n4
  );


  buf
  g108
  (
    n62,
    n18
  );


  not
  g109
  (
    n105,
    n5
  );


  buf
  g110
  (
    n149,
    n10
  );


  not
  g111
  (
    n130,
    n8
  );


  buf
  g112
  (
    n37,
    n21
  );


  not
  g113
  (
    n98,
    n27
  );


  buf
  g114
  (
    n128,
    n22
  );


  buf
  g115
  (
    n133,
    n14
  );


  not
  g116
  (
    n50,
    n30
  );


  buf
  g117
  (
    n55,
    n19
  );


  buf
  g118
  (
    n116,
    n20
  );


  not
  g119
  (
    n79,
    n23
  );


  buf
  g120
  (
    n82,
    n12
  );


  not
  g121
  (
    n83,
    n7
  );


  buf
  g122
  (
    n113,
    n7
  );


  not
  g123
  (
    n122,
    n27
  );


  not
  g124
  (
    n181,
    n91
  );


  and
  g125
  (
    n267,
    n136,
    n124,
    n133,
    n121
  );


  nor
  g126
  (
    n210,
    n94,
    n33,
    n77,
    n70
  );


  xor
  g127
  (
    n185,
    n147,
    n91,
    n82,
    n72
  );


  xnor
  g128
  (
    n162,
    n36,
    n98,
    n60,
    n105
  );


  and
  g129
  (
    n165,
    n103,
    n61,
    n44,
    n118
  );


  nor
  g130
  (
    n174,
    n85,
    n120,
    n118,
    n101
  );


  nor
  g131
  (
    n253,
    n39,
    n153,
    n130,
    n90
  );


  xor
  g132
  (
    n173,
    n150,
    n56,
    n70,
    n119
  );


  nand
  g133
  (
    n261,
    n78,
    n37,
    n64,
    n91
  );


  xnor
  g134
  (
    n214,
    n151,
    n123,
    n148,
    n65
  );


  nand
  g135
  (
    n260,
    n138,
    n112,
    n151,
    n82
  );


  or
  g136
  (
    n266,
    n70,
    n39,
    n129,
    n35
  );


  xor
  g137
  (
    n172,
    n81,
    n152,
    n87,
    n95
  );


  or
  g138
  (
    n243,
    n127,
    n134,
    n128,
    n150
  );


  xnor
  g139
  (
    n238,
    n151,
    n41,
    n94,
    n116
  );


  nand
  g140
  (
    n259,
    n149,
    n117,
    n56,
    n143
  );


  and
  g141
  (
    n203,
    n34,
    n75,
    n152,
    n61
  );


  nor
  g142
  (
    n250,
    n113,
    n146,
    n131,
    n132
  );


  nor
  g143
  (
    n202,
    n42,
    n102,
    n113,
    n116
  );


  nand
  g144
  (
    n158,
    n37,
    n149,
    n124,
    n58
  );


  xnor
  g145
  (
    n182,
    n60,
    n146,
    n95,
    n73
  );


  nand
  g146
  (
    n268,
    n133,
    n139,
    n119,
    n92
  );


  and
  g147
  (
    n236,
    n64,
    n106,
    n65,
    n111
  );


  xnor
  g148
  (
    n157,
    n95,
    n44,
    n81,
    n104
  );


  nor
  g149
  (
    n257,
    n58,
    n57,
    n123,
    n81
  );


  xnor
  g150
  (
    n263,
    n57,
    n146,
    n110,
    n46
  );


  xor
  g151
  (
    n277,
    n118,
    n57,
    n122,
    n80
  );


  nor
  g152
  (
    n239,
    n89,
    n46,
    n139,
    n79
  );


  and
  g153
  (
    n254,
    n93,
    n43,
    n100,
    n127
  );


  xnor
  g154
  (
    n228,
    n132,
    n117,
    n54,
    n70
  );


  and
  g155
  (
    n195,
    n42,
    n35,
    n57,
    n75
  );


  xor
  g156
  (
    n190,
    n114,
    n41,
    n55,
    n44
  );


  and
  g157
  (
    n159,
    n91,
    n53,
    n48,
    n141
  );


  nor
  g158
  (
    n184,
    n97,
    n138,
    n37,
    n77
  );


  nand
  g159
  (
    n186,
    n134,
    n137,
    n74
  );


  nand
  g160
  (
    n245,
    n133,
    n142,
    n117,
    n61
  );


  nand
  g161
  (
    n167,
    n143,
    n92,
    n77,
    n96
  );


  and
  g162
  (
    n265,
    n92,
    n125,
    n141,
    n153
  );


  and
  g163
  (
    n166,
    n47,
    n62,
    n52,
    n50
  );


  xor
  g164
  (
    n216,
    n108,
    n41,
    n144,
    n55
  );


  xor
  g165
  (
    n248,
    n74,
    n152,
    n80,
    n128
  );


  nor
  g166
  (
    n215,
    n69,
    n83,
    n49,
    n110
  );


  and
  g167
  (
    n237,
    n141,
    n64,
    n89,
    n67
  );


  nand
  g168
  (
    n196,
    n115,
    n135,
    n78,
    n139
  );


  nand
  g169
  (
    n234,
    n144,
    n121,
    n114,
    n108
  );


  xor
  g170
  (
    n218,
    n125,
    n122,
    n152,
    n102
  );


  nand
  g171
  (
    n249,
    n99,
    n135,
    n39,
    n38
  );


  or
  g172
  (
    n272,
    n93,
    n146,
    n104,
    n67
  );


  nand
  g173
  (
    n251,
    n34,
    n86,
    n58,
    n127
  );


  nand
  g174
  (
    n269,
    n140,
    n51,
    n80,
    n145
  );


  nand
  g175
  (
    n170,
    n145,
    n49,
    n102,
    n87
  );


  or
  g176
  (
    n232,
    n94,
    n78,
    n53,
    n114
  );


  xnor
  g177
  (
    n231,
    n76,
    n97,
    n90,
    n142
  );


  xor
  g178
  (
    n189,
    n145,
    n115,
    n63,
    n71
  );


  xnor
  g179
  (
    n255,
    n89,
    n108,
    n104,
    n116
  );


  xnor
  g180
  (
    n229,
    n90,
    n43,
    n82,
    n36
  );


  xnor
  g181
  (
    n178,
    n73,
    n89,
    n88
  );


  xnor
  g182
  (
    n168,
    n47,
    n85,
    n87,
    n48
  );


  and
  g183
  (
    n246,
    n150,
    n107,
    n113,
    n38
  );


  nor
  g184
  (
    n206,
    n100,
    n131,
    n59,
    n51
  );


  nor
  g185
  (
    n199,
    n96,
    n66,
    n61,
    n148
  );


  xnor
  g186
  (
    n188,
    n34,
    n85,
    n148,
    n45
  );


  or
  g187
  (
    n258,
    n52,
    n133,
    n127,
    n58
  );


  and
  g188
  (
    n183,
    n142,
    n84,
    n66,
    n33
  );


  nor
  g189
  (
    n274,
    n150,
    n62,
    n63,
    n53
  );


  nand
  g190
  (
    n200,
    n113,
    n52,
    n103,
    n130
  );


  xor
  g191
  (
    n193,
    n69,
    n129,
    n144,
    n122
  );


  and
  g192
  (
    n211,
    n132,
    n55,
    n66,
    n84
  );


  xor
  g193
  (
    n219,
    n106,
    n115,
    n149,
    n54
  );


  nor
  g194
  (
    n171,
    n110,
    n85,
    n121,
    n69
  );


  nand
  g195
  (
    n207,
    n99,
    n141,
    n66,
    n131
  );


  nand
  g196
  (
    n271,
    n111,
    n105,
    n114,
    n103
  );


  or
  g197
  (
    n220,
    n45,
    n102,
    n79,
    n56
  );


  xnor
  g198
  (
    n270,
    n67,
    n92,
    n97,
    n63
  );


  nor
  g199
  (
    n278,
    n81,
    n112,
    n72
  );


  nand
  g200
  (
    n227,
    n86,
    n116,
    n131,
    n111
  );


  nand
  g201
  (
    n160,
    n107,
    n132,
    n49,
    n51
  );


  or
  g202
  (
    n213,
    n104,
    n60,
    n112,
    n43
  );


  nand
  g203
  (
    n221,
    n50,
    n62,
    n51,
    n147
  );


  xor
  g204
  (
    n247,
    n68,
    n60,
    n44,
    n142
  );


  and
  g205
  (
    n273,
    n137,
    n98,
    n75
  );


  nand
  g206
  (
    n226,
    n45,
    n118,
    n154,
    n82
  );


  xor
  g207
  (
    n187,
    n48,
    n40,
    n137,
    n33
  );


  nor
  g208
  (
    n191,
    n48,
    n78,
    n55,
    n83
  );


  nor
  g209
  (
    n180,
    n46,
    n59,
    n97,
    n72
  );


  nor
  g210
  (
    n252,
    n76,
    n112,
    n107,
    n68
  );


  xor
  g211
  (
    n204,
    n148,
    n59,
    n136,
    n40
  );


  xnor
  g212
  (
    n161,
    n77,
    n86,
    n124,
    n111
  );


  and
  g213
  (
    n275,
    n45,
    n71,
    n125,
    n138
  );


  nand
  g214
  (
    n242,
    n143,
    n119,
    n39,
    n135
  );


  xnor
  g215
  (
    n194,
    n109,
    n93,
    n56,
    n43
  );


  or
  g216
  (
    n175,
    n120,
    n40,
    n125
  );


  xor
  g217
  (
    n177,
    n88,
    n47,
    n120,
    n99
  );


  xnor
  g218
  (
    n256,
    n41,
    n76,
    n100,
    n120
  );


  and
  g219
  (
    n217,
    n105,
    n107,
    n138,
    n71
  );


  and
  g220
  (
    n176,
    n126,
    n64,
    n147,
    n103
  );


  xnor
  g221
  (
    n240,
    n126,
    n115,
    n54,
    n117
  );


  xor
  g222
  (
    n197,
    n126,
    n47,
    n52,
    n119
  );


  nor
  g223
  (
    n223,
    n86,
    n101,
    n50
  );


  and
  g224
  (
    n212,
    n80,
    n84,
    n129,
    n42
  );


  nand
  g225
  (
    n222,
    n74,
    n134,
    n136,
    n59
  );


  xnor
  g226
  (
    n224,
    n149,
    n68,
    n65,
    n147
  );


  or
  g227
  (
    n264,
    n130,
    n35,
    n126,
    n37
  );


  xor
  g228
  (
    n164,
    n83,
    n71,
    n109,
    n65
  );


  nor
  g229
  (
    n235,
    n140,
    n79,
    n67,
    n36
  );


  or
  g230
  (
    n163,
    n38,
    n94,
    n54,
    n122
  );


  nand
  g231
  (
    n192,
    n130,
    n96,
    n128,
    n123
  );


  xor
  g232
  (
    n205,
    n53,
    n46,
    n90,
    n144
  );


  xnor
  g233
  (
    n233,
    n62,
    n83,
    n76,
    n108
  );


  nand
  g234
  (
    n276,
    n38,
    n128,
    n87,
    n36
  );


  xor
  g235
  (
    n179,
    n79,
    n34,
    n135,
    n42
  );


  xor
  g236
  (
    n169,
    n124,
    n110,
    n105,
    n136
  );


  or
  g237
  (
    n209,
    n95,
    n139,
    n101,
    n73
  );


  nor
  g238
  (
    n198,
    n109,
    n93,
    n35,
    n106
  );


  nor
  g239
  (
    n208,
    n68,
    n153,
    n99,
    n49
  );


  nand
  g240
  (
    n225,
    n100,
    n69,
    n88,
    n143
  );


  nand
  g241
  (
    n244,
    n98,
    n121,
    n109,
    n106
  );


  nand
  g242
  (
    n262,
    n50,
    n140,
    n134,
    n73
  );


  nand
  g243
  (
    n230,
    n75,
    n63,
    n151,
    n145
  );


  and
  g244
  (
    n241,
    n33,
    n153,
    n84,
    n74
  );


  xor
  g245
  (
    n201,
    n96,
    n123,
    n140,
    n129
  );


  or
  g246
  (
    n289,
    n179,
    n160,
    n181,
    n183
  );


  xor
  g247
  (
    n284,
    n173,
    n188,
    n184,
    n186
  );


  xnor
  g248
  (
    n281,
    n174,
    n176,
    n190,
    n185
  );


  xor
  g249
  (
    n292,
    n176,
    n169,
    n187,
    n168
  );


  xor
  g250
  (
    n282,
    n160,
    n158,
    n166
  );


  or
  g251
  (
    n294,
    n169,
    n164,
    n175,
    n183
  );


  xor
  g252
  (
    n287,
    n157,
    n159,
    n163,
    n179
  );


  xor
  g253
  (
    n279,
    n187,
    n178,
    n172,
    n165
  );


  xor
  g254
  (
    n285,
    n182,
    n180,
    n184,
    n186
  );


  xnor
  g255
  (
    n290,
    n173,
    n181,
    n162
  );


  nor
  g256
  (
    n288,
    n188,
    n182,
    n171,
    n167
  );


  nor
  g257
  (
    n280,
    n161,
    n161,
    n165,
    n171
  );


  and
  g258
  (
    n291,
    n177,
    n174,
    n170,
    n168
  );


  and
  g259
  (
    n293,
    n163,
    n175,
    n172,
    n164
  );


  xnor
  g260
  (
    n286,
    n180,
    n189,
    n185,
    n177
  );


  nor
  g261
  (
    n283,
    n189,
    n178,
    n170,
    n167
  );


  buf
  g262
  (
    n304,
    n280
  );


  buf
  g263
  (
    n296,
    n281
  );


  not
  g264
  (
    n299,
    n282
  );


  not
  g265
  (
    n295,
    n288
  );


  buf
  g266
  (
    n302,
    n284
  );


  buf
  g267
  (
    n297,
    n287
  );


  not
  g268
  (
    n301,
    n283
  );


  not
  g269
  (
    n300,
    n286
  );


  buf
  g270
  (
    n298,
    n279
  );


  not
  g271
  (
    n303,
    n285
  );


  nor
  g272
  (
    n335,
    n297,
    n301,
    n209,
    n193
  );


  and
  g273
  (
    n327,
    n302,
    n220,
    n234,
    n200
  );


  and
  g274
  (
    n307,
    n234,
    n228,
    n296,
    n302
  );


  nand
  g275
  (
    n325,
    n223,
    n206,
    n194,
    n302
  );


  xnor
  g276
  (
    n317,
    n205,
    n296,
    n228,
    n295
  );


  or
  g277
  (
    n316,
    n235,
    n231,
    n208,
    n219
  );


  or
  g278
  (
    n306,
    n298,
    n233,
    n207,
    n194
  );


  xor
  g279
  (
    n326,
    n298,
    n205,
    n216,
    n203
  );


  and
  g280
  (
    n315,
    n218,
    n230,
    n191,
    n301
  );


  xnor
  g281
  (
    n334,
    n222,
    n235,
    n199,
    n231
  );


  and
  g282
  (
    n323,
    n214,
    n218,
    n217,
    n224
  );


  or
  g283
  (
    n305,
    n224,
    n204,
    n214,
    n300
  );


  and
  g284
  (
    n329,
    n202,
    n302,
    n212,
    n217
  );


  nor
  g285
  (
    n312,
    n223,
    n232,
    n199,
    n215
  );


  xor
  g286
  (
    n324,
    n206,
    n301,
    n211,
    n296
  );


  nand
  g287
  (
    n318,
    n225,
    n236,
    n297,
    n219
  );


  nor
  g288
  (
    n311,
    n195,
    n299,
    n300,
    n297
  );


  nand
  g289
  (
    n331,
    n300,
    n299,
    n196,
    n204
  );


  nand
  g290
  (
    n319,
    n200,
    n220,
    n209,
    n230
  );


  and
  g291
  (
    n320,
    n232,
    n216,
    n196,
    n229
  );


  nor
  g292
  (
    n330,
    n210,
    n227,
    n299
  );


  and
  g293
  (
    n332,
    n190,
    n208,
    n201,
    n221
  );


  xor
  g294
  (
    n328,
    n295,
    n300,
    n221,
    n213
  );


  xnor
  g295
  (
    n310,
    n297,
    n299,
    n193,
    n212
  );


  nor
  g296
  (
    n313,
    n197,
    n295,
    n229,
    n215
  );


  or
  g297
  (
    n309,
    n211,
    n203,
    n301,
    n233
  );


  nand
  g298
  (
    n314,
    n226,
    n236,
    n201,
    n191
  );


  xnor
  g299
  (
    n333,
    n197,
    n198,
    n298
  );


  or
  g300
  (
    n322,
    n296,
    n225,
    n222,
    n298
  );


  or
  g301
  (
    n321,
    n213,
    n192,
    n210,
    n195
  );


  xnor
  g302
  (
    n308,
    n226,
    n202,
    n192,
    n207
  );


  buf
  g303
  (
    n343,
    n305
  );


  buf
  g304
  (
    n344,
    n306
  );


  buf
  g305
  (
    n338,
    n307
  );


  buf
  g306
  (
    n339,
    n307
  );


  not
  g307
  (
    n337,
    n306
  );


  buf
  g308
  (
    n340,
    n306
  );


  buf
  g309
  (
    n345,
    n307
  );


  buf
  g310
  (
    n336,
    n305
  );


  not
  g311
  (
    n342,
    n307
  );


  not
  g312
  (
    n341,
    n306
  );


  and
  g313
  (
    n351,
    n338,
    n248,
    n239,
    n242
  );


  or
  g314
  (
    n353,
    n341,
    n244,
    n245,
    n248
  );


  xor
  g315
  (
    n347,
    n245,
    n246,
    n237,
    n241
  );


  nor
  g316
  (
    n350,
    n247,
    n340,
    n243,
    n342
  );


  xnor
  g317
  (
    n348,
    n343,
    n241,
    n246,
    n247
  );


  or
  g318
  (
    n346,
    n337,
    n240,
    n244
  );


  xnor
  g319
  (
    n352,
    n336,
    n242,
    n243,
    n237
  );


  and
  g320
  (
    n349,
    n239,
    n238,
    n339
  );


  not
  g321
  (
    n363,
    n346
  );


  not
  g322
  (
    n362,
    n348
  );


  buf
  g323
  (
    n355,
    n349
  );


  buf
  g324
  (
    n356,
    n349
  );


  not
  g325
  (
    n357,
    n347
  );


  not
  g326
  (
    n359,
    n346
  );


  buf
  g327
  (
    n358,
    n347
  );


  buf
  g328
  (
    n360,
    n349
  );


  not
  g329
  (
    n354,
    n349
  );


  not
  g330
  (
    n361,
    n348
  );


  buf
  g331
  (
    n396,
    n356
  );


  not
  g332
  (
    n365,
    n352
  );


  buf
  g333
  (
    n379,
    n356
  );


  not
  g334
  (
    n369,
    n263
  );


  nand
  g335
  (
    n393,
    n314,
    n309
  );


  nor
  g336
  (
    n400,
    n263,
    n314,
    n361,
    n259
  );


  and
  g337
  (
    n375,
    n356,
    n249,
    n355,
    n308
  );


  xnor
  g338
  (
    n383,
    n251,
    n361,
    n350,
    n354
  );


  xor
  g339
  (
    n373,
    n312,
    n255,
    n303,
    n304
  );


  xnor
  g340
  (
    n370,
    n350,
    n360,
    n361,
    n352
  );


  nor
  g341
  (
    n403,
    n357,
    n265,
    n355,
    n317
  );


  nor
  g342
  (
    n386,
    n356,
    n358,
    n254,
    n362
  );


  nor
  g343
  (
    n401,
    n363,
    n264,
    n358,
    n357
  );


  xnor
  g344
  (
    n377,
    n359,
    n309,
    n350,
    n303
  );


  and
  g345
  (
    n392,
    n257,
    n363,
    n252,
    n315
  );


  nor
  g346
  (
    n399,
    n154,
    n308,
    n262,
    n257
  );


  or
  g347
  (
    n387,
    n250,
    n351,
    n357,
    n254
  );


  xnor
  g348
  (
    n374,
    n358,
    n311,
    n355,
    n359
  );


  and
  g349
  (
    n380,
    n260,
    n313,
    n312,
    n310
  );


  xnor
  g350
  (
    n385,
    n304,
    n309,
    n312,
    n310
  );


  xnor
  g351
  (
    n364,
    n251,
    n363,
    n318,
    n265
  );


  or
  g352
  (
    n371,
    n267,
    n319,
    n314,
    n313
  );


  or
  g353
  (
    n395,
    n304,
    n267,
    n354,
    n310
  );


  nand
  g354
  (
    n389,
    n316,
    n253,
    n303,
    n317
  );


  xnor
  g355
  (
    n367,
    n313,
    n351,
    n310,
    n319
  );


  xnor
  g356
  (
    n390,
    n256,
    n266,
    n357,
    n311
  );


  or
  g357
  (
    n384,
    n350,
    n352,
    n354,
    n316
  );


  nor
  g358
  (
    n378,
    n359,
    n309,
    n351,
    n360
  );


  and
  g359
  (
    n382,
    n311,
    n313,
    n253,
    n351
  );


  nand
  g360
  (
    n391,
    n304,
    n266,
    n316,
    n264
  );


  or
  g361
  (
    n402,
    n354,
    n311,
    n261,
    n249
  );


  nor
  g362
  (
    n381,
    n255,
    n250,
    n308,
    n362
  );


  xor
  g363
  (
    n366,
    n315,
    n315,
    n256,
    n363
  );


  xor
  g364
  (
    n376,
    n318,
    n362,
    n314,
    n358
  );


  and
  g365
  (
    n368,
    n362,
    n318,
    n359,
    n308
  );


  or
  g366
  (
    n388,
    n252,
    n260,
    n312,
    n258
  );


  nor
  g367
  (
    n394,
    n360,
    n303,
    n318,
    n262
  );


  xnor
  g368
  (
    n398,
    n259,
    n315,
    n258,
    n361
  );


  xor
  g369
  (
    n397,
    n154,
    n360,
    n261,
    n316
  );


  nor
  g370
  (
    n372,
    n355,
    n317,
    n352
  );


  not
  g371
  (
    n419,
    n364
  );


  not
  g372
  (
    n404,
    n322
  );


  buf
  g373
  (
    n416,
    n323
  );


  buf
  g374
  (
    n411,
    n320
  );


  buf
  g375
  (
    n409,
    n370
  );


  buf
  g376
  (
    n413,
    n367
  );


  buf
  g377
  (
    n408,
    n320
  );


  not
  g378
  (
    n420,
    n370
  );


  or
  g379
  (
    n407,
    n368,
    n365,
    n322,
    n321
  );


  xor
  g380
  (
    n405,
    n319,
    n366,
    n365
  );


  and
  g381
  (
    n406,
    n367,
    n368,
    n372,
    n320
  );


  nand
  g382
  (
    n415,
    n370,
    n369,
    n367,
    n322
  );


  nor
  g383
  (
    n410,
    n365,
    n371,
    n369,
    n364
  );


  nor
  g384
  (
    n412,
    n319,
    n366,
    n321
  );


  and
  g385
  (
    n422,
    n367,
    n321,
    n369
  );


  xnor
  g386
  (
    n421,
    n371,
    n371,
    n323,
    n372
  );


  or
  g387
  (
    n417,
    n322,
    n368,
    n364,
    n320
  );


  xnor
  g388
  (
    n414,
    n372,
    n369,
    n370,
    n368
  );


  nor
  g389
  (
    n418,
    n364,
    n371,
    n365,
    n372
  );


  and
  g390
  (
    n437,
    n154,
    n345,
    n293
  );


  nand
  g391
  (
    n439,
    n415,
    n324,
    n323
  );


  nor
  g392
  (
    n438,
    n155,
    n417,
    n325
  );


  xnor
  g393
  (
    n427,
    n414,
    n292,
    n324
  );


  or
  g394
  (
    n434,
    n271,
    n155,
    n32
  );


  xor
  g395
  (
    n433,
    n406,
    n420,
    n270
  );


  nand
  g396
  (
    n436,
    n409,
    n268,
    n32
  );


  or
  g397
  (
    n425,
    n419,
    n325
  );


  and
  g398
  (
    n429,
    n294,
    n293,
    n324,
    n411
  );


  and
  g399
  (
    n432,
    n323,
    n155,
    n421,
    n413
  );


  xnor
  g400
  (
    n423,
    n292,
    n408,
    n156,
    n416
  );


  or
  g401
  (
    n424,
    n344,
    n156,
    n155,
    n326
  );


  xor
  g402
  (
    n431,
    n294,
    n422,
    n407,
    n418
  );


  and
  g403
  (
    n435,
    n289,
    n268,
    n156,
    n269
  );


  xnor
  g404
  (
    n426,
    n269,
    n324,
    n32,
    n290
  );


  and
  g405
  (
    n428,
    n270,
    n412,
    n291
  );


  nand
  g406
  (
    n430,
    n325,
    n410,
    n271,
    n32
  );


  not
  g407
  (
    n460,
    n391
  );


  not
  g408
  (
    n452,
    n373
  );


  buf
  g409
  (
    n457,
    n428
  );


  not
  g410
  (
    n474,
    n402
  );


  and
  g411
  (
    n473,
    n439,
    n434,
    n403
  );


  nor
  g412
  (
    n443,
    n391,
    n353,
    n379
  );


  nor
  g413
  (
    n446,
    n399,
    n375,
    n429
  );


  or
  g414
  (
    n502,
    n392,
    n376,
    n381
  );


  and
  g415
  (
    n506,
    n398,
    n438,
    n402
  );


  nor
  g416
  (
    n495,
    n374,
    n394,
    n380
  );


  or
  g417
  (
    n476,
    n403,
    n377,
    n386
  );


  nor
  g418
  (
    n479,
    n395,
    n386,
    n431
  );


  xnor
  g419
  (
    n455,
    n432,
    n385,
    n376
  );


  or
  g420
  (
    n441,
    n401,
    n377,
    n400
  );


  and
  g421
  (
    n498,
    n384,
    n438,
    n398
  );


  or
  g422
  (
    n464,
    n374,
    n396,
    n395
  );


  xor
  g423
  (
    n470,
    n394,
    n397,
    n401
  );


  or
  g424
  (
    n492,
    n382,
    n383,
    n432
  );


  nor
  g425
  (
    n445,
    n433,
    n400,
    n429
  );


  xnor
  g426
  (
    n496,
    n374,
    n403,
    n425
  );


  xnor
  g427
  (
    n480,
    n382,
    n439,
    n383
  );


  nand
  g428
  (
    n450,
    n384,
    n438,
    n381
  );


  xnor
  g429
  (
    n504,
    n430,
    n426,
    n434
  );


  and
  g430
  (
    n493,
    n377,
    n436,
    n427
  );


  nand
  g431
  (
    n490,
    n427,
    n435,
    n385
  );


  xor
  g432
  (
    n468,
    n399,
    n429,
    n403
  );


  xor
  g433
  (
    n488,
    n433,
    n390
  );


  nand
  g434
  (
    n459,
    n426,
    n439,
    n393
  );


  nand
  g435
  (
    n442,
    n424,
    n433,
    n437
  );


  nor
  g436
  (
    n481,
    n393,
    n397,
    n437
  );


  and
  g437
  (
    n478,
    n398,
    n378,
    n431
  );


  or
  g438
  (
    n500,
    n398,
    n401,
    n382
  );


  nand
  g439
  (
    n453,
    n423,
    n388,
    n379
  );


  and
  g440
  (
    n491,
    n382,
    n374,
    n437
  );


  or
  g441
  (
    n507,
    n389,
    n400,
    n378
  );


  xnor
  g442
  (
    n449,
    n387,
    n380,
    n428
  );


  xnor
  g443
  (
    n467,
    n396,
    n373,
    n426
  );


  nand
  g444
  (
    n466,
    n397,
    n428,
    n378
  );


  nor
  g445
  (
    n503,
    n385,
    n425,
    n432
  );


  xor
  g446
  (
    n469,
    n426,
    n392,
    n402
  );


  nor
  g447
  (
    n461,
    n381,
    n389,
    n388
  );


  nor
  g448
  (
    n440,
    n439,
    n423,
    n385
  );


  nand
  g449
  (
    n489,
    n395,
    n384,
    n427
  );


  xnor
  g450
  (
    n485,
    n400,
    n387
  );


  xor
  g451
  (
    n487,
    n376,
    n393,
    n391
  );


  nand
  g452
  (
    n475,
    n353,
    n424,
    n388
  );


  and
  g453
  (
    n444,
    n389,
    n392,
    n434
  );


  and
  g454
  (
    n486,
    n392,
    n431,
    n399
  );


  nand
  g455
  (
    n477,
    n375,
    n424,
    n380
  );


  nand
  g456
  (
    n482,
    n425,
    n427,
    n402
  );


  or
  g457
  (
    n465,
    n436,
    n353,
    n394
  );


  xor
  g458
  (
    n447,
    n425,
    n436,
    n431
  );


  xor
  g459
  (
    n451,
    n401,
    n428,
    n399
  );


  nor
  g460
  (
    n483,
    n389,
    n353,
    n379
  );


  and
  g461
  (
    n494,
    n433,
    n397,
    n390
  );


  nor
  g462
  (
    n501,
    n381,
    n430,
    n396
  );


  nand
  g463
  (
    n497,
    n388,
    n378,
    n437
  );


  nand
  g464
  (
    n472,
    n423,
    n429,
    n436
  );


  xor
  g465
  (
    n462,
    n435,
    n423,
    n432
  );


  nand
  g466
  (
    n456,
    n373,
    n424,
    n383
  );


  nor
  g467
  (
    n454,
    n396,
    n395,
    n375
  );


  xor
  g468
  (
    n463,
    n380,
    n383,
    n390
  );


  nand
  g469
  (
    n484,
    n435,
    n377,
    n384
  );


  xnor
  g470
  (
    n505,
    n379,
    n375,
    n434
  );


  or
  g471
  (
    n458,
    n394,
    n430,
    n393
  );


  xor
  g472
  (
    n499,
    n386,
    n430,
    n435
  );


  nand
  g473
  (
    n448,
    n438,
    n373,
    n376
  );


  or
  g474
  (
    n471,
    n387,
    n391,
    n386
  );


  buf
  g475
  (
    n667,
    n276
  );


  not
  g476
  (
    n537,
    n478
  );


  buf
  g477
  (
    n629,
    n481
  );


  buf
  g478
  (
    n527,
    n484
  );


  not
  g479
  (
    n626,
    n272
  );


  buf
  g480
  (
    n540,
    n486
  );


  buf
  g481
  (
    n614,
    n453
  );


  not
  g482
  (
    n607,
    n503
  );


  buf
  g483
  (
    n528,
    n503
  );


  not
  g484
  (
    n551,
    n489
  );


  buf
  g485
  (
    n612,
    n497
  );


  buf
  g486
  (
    n587,
    n480
  );


  buf
  g487
  (
    n678,
    n472
  );


  not
  g488
  (
    n682,
    n477
  );


  not
  g489
  (
    n617,
    n487
  );


  not
  g490
  (
    n592,
    n440
  );


  not
  g491
  (
    n636,
    n447
  );


  not
  g492
  (
    n568,
    n481
  );


  buf
  g493
  (
    n590,
    n471
  );


  buf
  g494
  (
    n611,
    n471
  );


  buf
  g495
  (
    n526,
    n489
  );


  not
  g496
  (
    n642,
    n479
  );


  buf
  g497
  (
    n685,
    n479
  );


  not
  g498
  (
    n579,
    n473
  );


  not
  g499
  (
    n634,
    n476
  );


  buf
  g500
  (
    n599,
    n466
  );


  not
  g501
  (
    n597,
    n460
  );


  not
  g502
  (
    n673,
    n456
  );


  buf
  g503
  (
    n512,
    n474
  );


  not
  g504
  (
    n660,
    n483
  );


  not
  g505
  (
    n534,
    n475
  );


  buf
  g506
  (
    n606,
    n493
  );


  buf
  g507
  (
    n652,
    n453
  );


  buf
  g508
  (
    n675,
    n458
  );


  buf
  g509
  (
    n595,
    n479
  );


  not
  g510
  (
    n603,
    n450
  );


  not
  g511
  (
    n516,
    n465
  );


  not
  g512
  (
    n571,
    n440
  );


  not
  g513
  (
    n596,
    n442
  );


  buf
  g514
  (
    n657,
    n444
  );


  buf
  g515
  (
    n572,
    n506
  );


  not
  g516
  (
    n600,
    n469
  );


  not
  g517
  (
    n649,
    n488
  );


  buf
  g518
  (
    n525,
    n483
  );


  not
  g519
  (
    n594,
    n481
  );


  not
  g520
  (
    n570,
    n457
  );


  not
  g521
  (
    n542,
    n457
  );


  buf
  g522
  (
    n591,
    n450
  );


  not
  g523
  (
    n664,
    n504
  );


  buf
  g524
  (
    n661,
    n475
  );


  buf
  g525
  (
    n680,
    n507
  );


  buf
  g526
  (
    n647,
    n455
  );


  not
  g527
  (
    n628,
    n442
  );


  not
  g528
  (
    n582,
    n485
  );


  buf
  g529
  (
    n622,
    n460
  );


  not
  g530
  (
    n604,
    n276
  );


  buf
  g531
  (
    n651,
    n498
  );


  not
  g532
  (
    n548,
    n497
  );


  buf
  g533
  (
    n535,
    n273
  );


  buf
  g534
  (
    n643,
    n443
  );


  not
  g535
  (
    n566,
    n494
  );


  not
  g536
  (
    n635,
    n483
  );


  buf
  g537
  (
    n674,
    n441
  );


  buf
  g538
  (
    n646,
    n503
  );


  not
  g539
  (
    n586,
    n464
  );


  not
  g540
  (
    n532,
    n490
  );


  buf
  g541
  (
    n556,
    n447
  );


  not
  g542
  (
    n513,
    n461
  );


  buf
  g543
  (
    n521,
    n461
  );


  not
  g544
  (
    n509,
    n504
  );


  not
  g545
  (
    n633,
    n440
  );


  not
  g546
  (
    n624,
    n481
  );


  buf
  g547
  (
    n580,
    n471
  );


  not
  g548
  (
    n631,
    n272
  );


  buf
  g549
  (
    n519,
    n493
  );


  buf
  g550
  (
    n658,
    n462
  );


  not
  g551
  (
    n613,
    n445
  );


  not
  g552
  (
    n524,
    n498
  );


  not
  g553
  (
    n511,
    n507
  );


  not
  g554
  (
    n621,
    n500
  );


  not
  g555
  (
    n533,
    n451
  );


  buf
  g556
  (
    n619,
    n480
  );


  buf
  g557
  (
    n560,
    n495
  );


  buf
  g558
  (
    n554,
    n494
  );


  buf
  g559
  (
    n546,
    n443
  );


  not
  g560
  (
    n605,
    n448
  );


  buf
  g561
  (
    n565,
    n444
  );


  buf
  g562
  (
    n645,
    n490
  );


  buf
  g563
  (
    n615,
    n278
  );


  buf
  g564
  (
    n508,
    n460
  );


  not
  g565
  (
    n545,
    n473
  );


  not
  g566
  (
    n574,
    n454
  );


  buf
  g567
  (
    n549,
    n274
  );


  not
  g568
  (
    n536,
    n466
  );


  not
  g569
  (
    n514,
    n504
  );


  not
  g570
  (
    n541,
    n451
  );


  not
  g571
  (
    n539,
    n502
  );


  buf
  g572
  (
    n558,
    n469
  );


  not
  g573
  (
    n547,
    n275
  );


  not
  g574
  (
    n553,
    n484
  );


  buf
  g575
  (
    n585,
    n456
  );


  not
  g576
  (
    n679,
    n467
  );


  not
  g577
  (
    n569,
    n462
  );


  buf
  g578
  (
    n602,
    n475
  );


  buf
  g579
  (
    n518,
    n496
  );


  buf
  g580
  (
    n627,
    n465
  );


  not
  g581
  (
    n561,
    n505
  );


  not
  g582
  (
    n623,
    n501
  );


  not
  g583
  (
    n567,
    n457
  );


  not
  g584
  (
    n632,
    n469
  );


  not
  g585
  (
    n659,
    n463
  );


  buf
  g586
  (
    n637,
    n494
  );


  buf
  g587
  (
    n529,
    n464
  );


  buf
  g588
  (
    n559,
    n447
  );


  not
  g589
  (
    n653,
    n449
  );


  not
  g590
  (
    n543,
    n451
  );


  buf
  g591
  (
    n638,
    n482
  );


  not
  g592
  (
    n644,
    n487
  );


  buf
  g593
  (
    n650,
    n493
  );


  not
  g594
  (
    n550,
    n462
  );


  buf
  g595
  (
    n557,
    n501
  );


  not
  g596
  (
    n578,
    n492
  );


  not
  g597
  (
    n630,
    n480
  );


  buf
  g598
  (
    n583,
    n274
  );


  buf
  g599
  (
    n608,
    n494
  );


  buf
  g600
  (
    n655,
    n476
  );


  buf
  g601
  (
    n610,
    n442
  );


  buf
  g602
  (
    n620,
    n456
  );


  buf
  g603
  (
    n640,
    n486
  );


  buf
  g604
  (
    n588,
    n493
  );


  buf
  g605
  (
    n593,
    n465
  );


  buf
  g606
  (
    n517,
    n463
  );


  not
  g607
  (
    n601,
    n456
  );


  buf
  g608
  (
    n510,
    n454
  );


  buf
  g609
  (
    n677,
    n485
  );


  buf
  g610
  (
    n625,
    n497
  );


  not
  g611
  (
    n564,
    n440
  );


  buf
  g612
  (
    n589,
    n487
  );


  buf
  g613
  (
    n573,
    n505
  );


  buf
  g614
  (
    n648,
    n455
  );


  buf
  g615
  (
    n666,
    n273
  );


  not
  g616
  (
    n654,
    n504
  );


  and
  g617
  (
    n552,
    n278,
    n484,
    n458,
    n445
  );


  or
  g618
  (
    n662,
    n446,
    n463,
    n501,
    n459
  );


  xnor
  g619
  (
    n616,
    n506,
    n495,
    n480,
    n499
  );


  or
  g620
  (
    n522,
    n503,
    n486,
    n495,
    n489
  );


  xnor
  g621
  (
    n555,
    n501,
    n506,
    n499,
    n453
  );


  or
  g622
  (
    n669,
    n498,
    n452,
    n491,
    n275
  );


  xor
  g623
  (
    n515,
    n444,
    n442,
    n277,
    n450
  );


  xor
  g624
  (
    n663,
    n491,
    n495,
    n277,
    n454
  );


  xnor
  g625
  (
    n656,
    n476,
    n453,
    n465,
    n464
  );


  xnor
  g626
  (
    n538,
    n476,
    n472,
    n497,
    n496
  );


  nor
  g627
  (
    n670,
    n459,
    n463,
    n449,
    n468
  );


  or
  g628
  (
    n641,
    n483,
    n482,
    n500,
    n478
  );


  nand
  g629
  (
    n672,
    n492,
    n470,
    n477,
    n496
  );


  nand
  g630
  (
    n520,
    n488,
    n470,
    n474,
    n461
  );


  nand
  g631
  (
    n665,
    n490,
    n446,
    n445,
    n485
  );


  and
  g632
  (
    n575,
    n474,
    n507,
    n454,
    n485
  );


  nand
  g633
  (
    n683,
    n443,
    n490,
    n479,
    n492
  );


  xor
  g634
  (
    n584,
    n455,
    n468,
    n478,
    n488
  );


  xor
  g635
  (
    n563,
    n467,
    n446,
    n482,
    n469
  );


  xnor
  g636
  (
    n681,
    n473,
    n448,
    n468,
    n462
  );


  xnor
  g637
  (
    n671,
    n472,
    n449,
    n447,
    n441
  );


  xnor
  g638
  (
    n523,
    n461,
    n484,
    n472,
    n451
  );


  and
  g639
  (
    n576,
    n455,
    n502,
    n500,
    n446
  );


  nand
  g640
  (
    n531,
    n482,
    n468,
    n499,
    n459
  );


  nor
  g641
  (
    n562,
    n478,
    n470,
    n452
  );


  nor
  g642
  (
    n530,
    n505,
    n460,
    n477,
    n498
  );


  nand
  g643
  (
    n544,
    n458,
    n448,
    n488,
    n491
  );


  or
  g644
  (
    n609,
    n470,
    n452,
    n499,
    n500
  );


  and
  g645
  (
    n668,
    n443,
    n458,
    n445,
    n477
  );


  or
  g646
  (
    n581,
    n475,
    n505,
    n448,
    n449
  );


  xor
  g647
  (
    n618,
    n491,
    n496,
    n441,
    n502
  );


  or
  g648
  (
    n676,
    n502,
    n471,
    n467,
    n441
  );


  xnor
  g649
  (
    n684,
    n444,
    n466,
    n450,
    n489
  );


  xnor
  g650
  (
    n598,
    n457,
    n507,
    n473,
    n506
  );


  xnor
  g651
  (
    n577,
    n464,
    n466,
    n492,
    n487
  );


  or
  g652
  (
    n639,
    n467,
    n474,
    n459,
    n486
  );


  not
  g653
  (
    n692,
    n526
  );


  not
  g654
  (
    n697,
    n573
  );


  not
  g655
  (
    n740,
    n543
  );


  not
  g656
  (
    n762,
    n549
  );


  buf
  g657
  (
    n789,
    n658
  );


  buf
  g658
  (
    n787,
    n572
  );


  buf
  g659
  (
    n793,
    n567
  );


  buf
  g660
  (
    n706,
    n624
  );


  not
  g661
  (
    n713,
    n647
  );


  not
  g662
  (
    n721,
    n601
  );


  not
  g663
  (
    n730,
    n614
  );


  not
  g664
  (
    n743,
    n530
  );


  buf
  g665
  (
    n695,
    n563
  );


  not
  g666
  (
    n699,
    n519
  );


  buf
  g667
  (
    n711,
    n667
  );


  buf
  g668
  (
    n788,
    n615
  );


  not
  g669
  (
    n712,
    n646
  );


  buf
  g670
  (
    n716,
    n629
  );


  buf
  g671
  (
    n754,
    n599
  );


  buf
  g672
  (
    n742,
    n634
  );


  not
  g673
  (
    n705,
    n589
  );


  not
  g674
  (
    n767,
    n566
  );


  buf
  g675
  (
    n792,
    n625
  );


  buf
  g676
  (
    n720,
    n616
  );


  buf
  g677
  (
    n778,
    n568
  );


  not
  g678
  (
    n717,
    n626
  );


  not
  g679
  (
    n756,
    n565
  );


  not
  g680
  (
    n783,
    n553
  );


  not
  g681
  (
    n727,
    n657
  );


  not
  g682
  (
    n689,
    n636
  );


  buf
  g683
  (
    n770,
    n575
  );


  buf
  g684
  (
    n696,
    n580
  );


  buf
  g685
  (
    n748,
    n564
  );


  not
  g686
  (
    n761,
    n534
  );


  buf
  g687
  (
    n715,
    n555
  );


  buf
  g688
  (
    n759,
    n529
  );


  buf
  g689
  (
    n734,
    n535
  );


  not
  g690
  (
    n776,
    n641
  );


  or
  g691
  (
    n726,
    n645,
    n548
  );


  xor
  g692
  (
    n702,
    n657,
    n604,
    n627,
    n584
  );


  nand
  g693
  (
    n786,
    n522,
    n641,
    n574,
    n520
  );


  xnor
  g694
  (
    n703,
    n606,
    n551,
    n573,
    n652
  );


  nor
  g695
  (
    n686,
    n612,
    n562,
    n664,
    n632
  );


  nand
  g696
  (
    n714,
    n618,
    n637,
    n629,
    n600
  );


  nor
  g697
  (
    n766,
    n660,
    n517,
    n638,
    n539
  );


  nand
  g698
  (
    n731,
    n530,
    n571,
    n592,
    n585
  );


  and
  g699
  (
    n691,
    n560,
    n642,
    n654,
    n603
  );


  nand
  g700
  (
    n760,
    n633,
    n602,
    n580,
    n556
  );


  and
  g701
  (
    n701,
    n528,
    n547,
    n524,
    n577
  );


  or
  g702
  (
    n750,
    n563,
    n610,
    n606,
    n626
  );


  xnor
  g703
  (
    n777,
    n533,
    n514,
    n590,
    n509
  );


  xor
  g704
  (
    n718,
    n605,
    n659,
    n612,
    n599
  );


  and
  g705
  (
    n790,
    n564,
    n637,
    n551,
    n545
  );


  or
  g706
  (
    n764,
    n644,
    n555,
    n639,
    n533
  );


  nand
  g707
  (
    n735,
    n582,
    n666,
    n662,
    n515
  );


  nor
  g708
  (
    n769,
    n609,
    n588,
    n647,
    n600
  );


  nor
  g709
  (
    n707,
    n589,
    n579,
    n594,
    n591
  );


  xor
  g710
  (
    n773,
    n552,
    n649,
    n651,
    n594
  );


  xor
  g711
  (
    n708,
    n661,
    n616,
    n518,
    n613
  );


  nor
  g712
  (
    n694,
    n618,
    n545,
    n602,
    n652
  );


  nor
  g713
  (
    n771,
    n575,
    n546,
    n550,
    n646
  );


  nand
  g714
  (
    n739,
    n508,
    n597,
    n542,
    n515
  );


  xnor
  g715
  (
    n736,
    n620,
    n559,
    n649,
    n548
  );


  or
  g716
  (
    n749,
    n571,
    n664,
    n579,
    n523
  );


  xor
  g717
  (
    n700,
    n632,
    n525,
    n565,
    n584
  );


  and
  g718
  (
    n690,
    n511,
    n621,
    n623,
    n550
  );


  nor
  g719
  (
    n782,
    n537,
    n538,
    n510,
    n514
  );


  xnor
  g720
  (
    n772,
    n521,
    n607,
    n622,
    n537
  );


  nor
  g721
  (
    n688,
    n661,
    n510,
    n509,
    n631
  );


  nor
  g722
  (
    n775,
    n558,
    n627,
    n523,
    n593
  );


  nor
  g723
  (
    n693,
    n663,
    n539,
    n528,
    n665
  );


  or
  g724
  (
    n774,
    n663,
    n557,
    n651,
    n608
  );


  nand
  g725
  (
    n791,
    n547,
    n520,
    n560,
    n569
  );


  and
  g726
  (
    n794,
    n645,
    n581,
    n643,
    n586
  );


  xor
  g727
  (
    n755,
    n662,
    n656,
    n595,
    n519
  );


  xnor
  g728
  (
    n728,
    n570,
    n540,
    n513,
    n525
  );


  or
  g729
  (
    n710,
    n609,
    n513,
    n534,
    n544
  );


  and
  g730
  (
    n704,
    n532,
    n622,
    n656,
    n531
  );


  nor
  g731
  (
    n709,
    n516,
    n596,
    n634,
    n592
  );


  and
  g732
  (
    n719,
    n572,
    n586,
    n608,
    n558
  );


  nand
  g733
  (
    n753,
    n593,
    n587,
    n659,
    n535
  );


  and
  g734
  (
    n781,
    n557,
    n620,
    n648,
    n568
  );


  or
  g735
  (
    n725,
    n531,
    n625,
    n522,
    n655
  );


  xor
  g736
  (
    n729,
    n615,
    n576,
    n587,
    n598
  );


  xnor
  g737
  (
    n687,
    n597,
    n590,
    n605,
    n544
  );


  nor
  g738
  (
    n744,
    n508,
    n577,
    n624,
    n607
  );


  xor
  g739
  (
    n763,
    n532,
    n552,
    n553,
    n617
  );


  nand
  g740
  (
    n751,
    n650,
    n526,
    n619,
    n585
  );


  nor
  g741
  (
    n757,
    n517,
    n578,
    n566,
    n518
  );


  and
  g742
  (
    n758,
    n581,
    n559,
    n540,
    n527
  );


  xnor
  g743
  (
    n768,
    n583,
    n512,
    n621,
    n561
  );


  nand
  g744
  (
    n722,
    n598,
    n643,
    n542,
    n603
  );


  xnor
  g745
  (
    n765,
    n613,
    n546,
    n611,
    n536
  );


  or
  g746
  (
    n723,
    n619,
    n583,
    n614,
    n569
  );


  nand
  g747
  (
    n745,
    n640,
    n529,
    n554,
    n631
  );


  xnor
  g748
  (
    n733,
    n556,
    n640,
    n667,
    n601
  );


  xnor
  g749
  (
    n752,
    n511,
    n567,
    n596,
    n512
  );


  xor
  g750
  (
    n746,
    n541,
    n604,
    n660,
    n549
  );


  nand
  g751
  (
    n784,
    n623,
    n638,
    n630,
    n666
  );


  or
  g752
  (
    n785,
    n648,
    n536,
    n595,
    n653
  );


  nor
  g753
  (
    n779,
    n582,
    n636,
    n570,
    n665
  );


  xor
  g754
  (
    n738,
    n578,
    n562,
    n576,
    n653
  );


  xnor
  g755
  (
    n698,
    n588,
    n538,
    n639,
    n561
  );


  nand
  g756
  (
    n724,
    n521,
    n650,
    n574,
    n628
  );


  and
  g757
  (
    n780,
    n527,
    n611,
    n541,
    n633
  );


  xnor
  g758
  (
    n732,
    n554,
    n635,
    n655,
    n543
  );


  or
  g759
  (
    n741,
    n628,
    n658,
    n642,
    n610
  );


  and
  g760
  (
    n747,
    n617,
    n516,
    n591,
    n654
  );


  xnor
  g761
  (
    n737,
    n524,
    n630,
    n644,
    n635
  );


  not
  g762
  (
    n796,
    n687
  );


  buf
  g763
  (
    n797,
    n687
  );


  not
  g764
  (
    n795,
    n686
  );


  buf
  g765
  (
    n798,
    n686
  );


  xor
  g766
  (
    n805,
    n798,
    n326,
    n674
  );


  xnor
  g767
  (
    n806,
    n672,
    n327,
    n796,
    n677
  );


  nor
  g768
  (
    n802,
    n796,
    n675,
    n671,
    n795
  );


  xor
  g769
  (
    n800,
    n668,
    n673,
    n798,
    n669
  );


  or
  g770
  (
    n804,
    n797,
    n670,
    n669,
    n795
  );


  or
  g771
  (
    n801,
    n675,
    n668,
    n671,
    n798
  );


  nor
  g772
  (
    n799,
    n327,
    n673,
    n672,
    n676
  );


  xnor
  g773
  (
    n803,
    n326,
    n677,
    n797,
    n674
  );


  nand
  g774
  (
    n807,
    n678,
    n678,
    n670,
    n676
  );


  buf
  g775
  (
    n808,
    n804
  );


  buf
  g776
  (
    n809,
    n802
  );


  buf
  g777
  (
    n810,
    n689
  );


  buf
  g778
  (
    n817,
    n799
  );


  buf
  g779
  (
    n821,
    n802
  );


  not
  g780
  (
    n816,
    n804
  );


  buf
  g781
  (
    n815,
    n807
  );


  not
  g782
  (
    n820,
    n688
  );


  buf
  g783
  (
    n812,
    n807
  );


  buf
  g784
  (
    n819,
    n805
  );


  buf
  g785
  (
    n822,
    n801
  );


  not
  g786
  (
    n818,
    n805
  );


  nand
  g787
  (
    n811,
    n806,
    n688
  );


  and
  g788
  (
    n813,
    n800,
    n803
  );


  or
  g789
  (
    n814,
    n803,
    n806
  );


  buf
  g790
  (
    n825,
    n820
  );


  not
  g791
  (
    n867,
    n333
  );


  not
  g792
  (
    n870,
    n817
  );


  buf
  g793
  (
    n841,
    n821
  );


  buf
  g794
  (
    n826,
    n817
  );


  buf
  g795
  (
    n868,
    n811
  );


  buf
  g796
  (
    n834,
    n683
  );


  buf
  g797
  (
    n830,
    n817
  );


  not
  g798
  (
    n882,
    n334
  );


  buf
  g799
  (
    n860,
    n815
  );


  buf
  g800
  (
    n849,
    n814
  );


  not
  g801
  (
    n837,
    n818
  );


  buf
  g802
  (
    n835,
    n683
  );


  buf
  g803
  (
    n842,
    n335
  );


  not
  g804
  (
    n824,
    n814
  );


  buf
  g805
  (
    n833,
    n683
  );


  buf
  g806
  (
    n854,
    n819
  );


  not
  g807
  (
    n845,
    n822
  );


  buf
  g808
  (
    n827,
    n819
  );


  buf
  g809
  (
    n855,
    n329
  );


  not
  g810
  (
    n877,
    n821
  );


  not
  g811
  (
    n843,
    n819
  );


  not
  g812
  (
    n852,
    n820
  );


  buf
  g813
  (
    n865,
    n808
  );


  not
  g814
  (
    n881,
    n815
  );


  buf
  g815
  (
    n828,
    n822
  );


  not
  g816
  (
    n832,
    n812
  );


  not
  g817
  (
    n863,
    n818
  );


  buf
  g818
  (
    n873,
    n816
  );


  buf
  g819
  (
    n840,
    n684
  );


  not
  g820
  (
    n836,
    n331
  );


  buf
  g821
  (
    n861,
    n333
  );


  not
  g822
  (
    n879,
    n810
  );


  buf
  g823
  (
    n858,
    n811
  );


  buf
  g824
  (
    n878,
    n335
  );


  not
  g825
  (
    n831,
    n334
  );


  buf
  g826
  (
    n839,
    n329
  );


  buf
  g827
  (
    n838,
    n816
  );


  buf
  g828
  (
    n866,
    n812
  );


  buf
  g829
  (
    n874,
    n679
  );


  buf
  g830
  (
    n872,
    n328
  );


  xnor
  g831
  (
    n875,
    n327,
    n822,
    n810
  );


  nand
  g832
  (
    n850,
    n685,
    n333,
    n813,
    n821
  );


  nor
  g833
  (
    n851,
    n335,
    n809,
    n685,
    n681
  );


  nand
  g834
  (
    n846,
    n332,
    n821,
    n681,
    n811
  );


  or
  g835
  (
    n829,
    n328,
    n819,
    n334,
    n808
  );


  nor
  g836
  (
    n844,
    n684,
    n814,
    n813,
    n822
  );


  xor
  g837
  (
    n869,
    n335,
    n808,
    n809,
    n810
  );


  or
  g838
  (
    n853,
    n680,
    n329,
    n331,
    n815
  );


  or
  g839
  (
    n876,
    n328,
    n684,
    n330,
    n682
  );


  xor
  g840
  (
    n856,
    n816,
    n683,
    n815,
    n331
  );


  nor
  g841
  (
    n857,
    n328,
    n330,
    n816,
    n818
  );


  nand
  g842
  (
    n880,
    n327,
    n680,
    n809,
    n330
  );


  nor
  g843
  (
    n859,
    n685,
    n817,
    n333,
    n811
  );


  and
  g844
  (
    n864,
    n809,
    n820,
    n332,
    n334
  );


  xnor
  g845
  (
    n848,
    n685,
    n813,
    n812
  );


  nor
  g846
  (
    n871,
    n818,
    n679,
    n682,
    n814
  );


  and
  g847
  (
    n862,
    n810,
    n820,
    n331,
    n684
  );


  nand
  g848
  (
    n847,
    n808,
    n329,
    n682,
    n332
  );


  or
  g849
  (
    n823,
    n813,
    n330,
    n682,
    n332
  );


  xor
  g850
  (
    n973,
    n771,
    n836,
    n751,
    n835
  );


  and
  g851
  (
    n959,
    n827,
    n856,
    n872,
    n841
  );


  or
  g852
  (
    n979,
    n849,
    n834,
    n836,
    n865
  );


  or
  g853
  (
    n963,
    n788,
    n850,
    n782,
    n731
  );


  or
  g854
  (
    n978,
    n739,
    n772,
    n740,
    n784
  );


  xnor
  g855
  (
    n1000,
    n876,
    n705,
    n699,
    n843
  );


  xor
  g856
  (
    n972,
    n738,
    n794,
    n778,
    n786
  );


  nand
  g857
  (
    n934,
    n690,
    n777,
    n827,
    n711
  );


  nand
  g858
  (
    n908,
    n833,
    n850,
    n788,
    n853
  );


  or
  g859
  (
    n945,
    n878,
    n851,
    n874,
    n862
  );


  xnor
  g860
  (
    n933,
    n703,
    n877,
    n782,
    n759
  );


  nor
  g861
  (
    n922,
    n867,
    n842,
    n741
  );


  nor
  g862
  (
    n988,
    n767,
    n752,
    n730,
    n877
  );


  and
  g863
  (
    n957,
    n729,
    n876,
    n834,
    n857
  );


  xor
  g864
  (
    n937,
    n771,
    n773,
    n848,
    n850
  );


  nand
  g865
  (
    n955,
    n878,
    n766,
    n842,
    n692
  );


  xor
  g866
  (
    n903,
    n730,
    n747,
    n768,
    n828
  );


  nand
  g867
  (
    n991,
    n843,
    n879,
    n824,
    n856
  );


  or
  g868
  (
    n917,
    n848,
    n752,
    n861,
    n864
  );


  xnor
  g869
  (
    n929,
    n725,
    n776,
    n865,
    n879
  );


  xor
  g870
  (
    n896,
    n831,
    n707,
    n701,
    n791
  );


  nor
  g871
  (
    n986,
    n773,
    n793,
    n858,
    n786
  );


  xor
  g872
  (
    n952,
    n777,
    n744,
    n852,
    n749
  );


  xor
  g873
  (
    n975,
    n781,
    n718,
    n872,
    n836
  );


  nor
  g874
  (
    n916,
    n720,
    n784,
    n745,
    n716
  );


  xnor
  g875
  (
    n906,
    n848,
    n783,
    n719,
    n876
  );


  nand
  g876
  (
    n890,
    n882,
    n877,
    n792,
    n857
  );


  nand
  g877
  (
    n976,
    n760,
    n695,
    n829,
    n869
  );


  nor
  g878
  (
    n927,
    n840,
    n873,
    n765,
    n878
  );


  nor
  g879
  (
    n981,
    n863,
    n702,
    n697,
    n826
  );


  xnor
  g880
  (
    n983,
    n775,
    n726,
    n856,
    n860
  );


  or
  g881
  (
    n898,
    n831,
    n834,
    n850,
    n848
  );


  and
  g882
  (
    n967,
    n703,
    n826,
    n877,
    n880
  );


  and
  g883
  (
    n962,
    n881,
    n766,
    n764,
    n691
  );


  nand
  g884
  (
    n935,
    n868,
    n872,
    n851,
    n831
  );


  xor
  g885
  (
    n899,
    n865,
    n832,
    n753,
    n723
  );


  xor
  g886
  (
    n909,
    n841,
    n854,
    n852
  );


  or
  g887
  (
    n900,
    n774,
    n767,
    n718,
    n843
  );


  or
  g888
  (
    n966,
    n762,
    n725,
    n869,
    n710
  );


  and
  g889
  (
    n965,
    n742,
    n835,
    n861,
    n862
  );


  nor
  g890
  (
    n987,
    n828,
    n852,
    n861,
    n849
  );


  nor
  g891
  (
    n907,
    n844,
    n706,
    n776,
    n754
  );


  or
  g892
  (
    n939,
    n756,
    n701,
    n825,
    n759
  );


  nor
  g893
  (
    n914,
    n840,
    n715,
    n860,
    n830
  );


  nand
  g894
  (
    n994,
    n881,
    n853,
    n710,
    n788
  );


  nor
  g895
  (
    n883,
    n845,
    n769,
    n700,
    n859
  );


  nor
  g896
  (
    n947,
    n858,
    n772,
    n774,
    n770
  );


  nor
  g897
  (
    n940,
    n707,
    n858,
    n722,
    n753
  );


  and
  g898
  (
    n923,
    n766,
    n837,
    n831,
    n712
  );


  and
  g899
  (
    n995,
    n740,
    n794,
    n840,
    n781
  );


  nor
  g900
  (
    n912,
    n790,
    n862,
    n700,
    n879
  );


  or
  g901
  (
    n989,
    n694,
    n870,
    n783,
    n830
  );


  nor
  g902
  (
    n911,
    n825,
    n747,
    n867,
    n774
  );


  nor
  g903
  (
    n924,
    n838,
    n846,
    n863,
    n763
  );


  or
  g904
  (
    n928,
    n750,
    n874,
    n824,
    n868
  );


  nand
  g905
  (
    n897,
    n734,
    n704,
    n857,
    n879
  );


  nand
  g906
  (
    n938,
    n741,
    n709,
    n833,
    n875
  );


  nand
  g907
  (
    n889,
    n875,
    n882,
    n743,
    n871
  );


  nor
  g908
  (
    n932,
    n841,
    n874,
    n829,
    n830
  );


  xnor
  g909
  (
    n931,
    n882,
    n758,
    n794,
    n789
  );


  xor
  g910
  (
    n887,
    n780,
    n760,
    n737,
    n842
  );


  or
  g911
  (
    n998,
    n769,
    n875,
    n869,
    n733
  );


  nand
  g912
  (
    n895,
    n726,
    n768,
    n764,
    n855
  );


  xor
  g913
  (
    n936,
    n696,
    n853,
    n785,
    n832
  );


  nand
  g914
  (
    n905,
    n704,
    n868,
    n876,
    n835
  );


  or
  g915
  (
    n950,
    n845,
    n698,
    n863,
    n713
  );


  nand
  g916
  (
    n920,
    n787,
    n853,
    n864,
    n836
  );


  xor
  g917
  (
    n971,
    n837,
    n882,
    n693,
    n780
  );


  nor
  g918
  (
    n913,
    n847,
    n698,
    n715,
    n690
  );


  and
  g919
  (
    n892,
    n783,
    n708,
    n695,
    n880
  );


  or
  g920
  (
    n958,
    n692,
    n792,
    n872,
    n845
  );


  nor
  g921
  (
    n970,
    n755,
    n778,
    n733,
    n874
  );


  xor
  g922
  (
    n953,
    n728,
    n855,
    n787,
    n840
  );


  nand
  g923
  (
    n1001,
    n712,
    n750,
    n827,
    n771
  );


  nor
  g924
  (
    n993,
    n855,
    n770,
    n763
  );


  xnor
  g925
  (
    n951,
    n866,
    n793,
    n779,
    n846
  );


  and
  g926
  (
    n974,
    n765,
    n773,
    n878,
    n706
  );


  xnor
  g927
  (
    n964,
    n720,
    n735,
    n843,
    n786
  );


  xnor
  g928
  (
    n992,
    n727,
    n722,
    n828,
    n867
  );


  or
  g929
  (
    n901,
    n825,
    n847,
    n832,
    n790
  );


  xnor
  g930
  (
    n960,
    n769,
    n835,
    n734,
    n778
  );


  xor
  g931
  (
    n926,
    n761,
    n855,
    n851,
    n871
  );


  and
  g932
  (
    n969,
    n827,
    n772,
    n860,
    n708
  );


  xor
  g933
  (
    n949,
    n870,
    n844,
    n866,
    n781
  );


  and
  g934
  (
    n999,
    n696,
    n789,
    n854,
    n791
  );


  xor
  g935
  (
    n919,
    n723,
    n844,
    n732,
    n777
  );


  xor
  g936
  (
    n943,
    n880,
    n867,
    n775,
    n849
  );


  xnor
  g937
  (
    n1002,
    n864,
    n869,
    n851,
    n724
  );


  nand
  g938
  (
    n980,
    n824,
    n852,
    n745,
    n866
  );


  xnor
  g939
  (
    n885,
    n834,
    n826,
    n757,
    n779
  );


  xnor
  g940
  (
    n921,
    n724,
    n699,
    n791,
    n714
  );


  or
  g941
  (
    n918,
    n838,
    n748,
    n839,
    n784
  );


  and
  g942
  (
    n904,
    n780,
    n846,
    n775,
    n839
  );


  xnor
  g943
  (
    n944,
    n871,
    n756,
    n873,
    n838
  );


  or
  g944
  (
    n956,
    n776,
    n751,
    n782,
    n758
  );


  nand
  g945
  (
    n946,
    n728,
    n709,
    n863,
    n719
  );


  xnor
  g946
  (
    n984,
    n854,
    n787,
    n736,
    n880
  );


  nor
  g947
  (
    n982,
    n702,
    n711,
    n761,
    n742
  );


  nand
  g948
  (
    n990,
    n737,
    n792,
    n779,
    n825
  );


  xor
  g949
  (
    n942,
    n714,
    n721,
    n694,
    n738
  );


  or
  g950
  (
    n886,
    n824,
    n859,
    n767,
    n856
  );


  or
  g951
  (
    n915,
    n716,
    n849,
    n845,
    n757
  );


  xor
  g952
  (
    n891,
    n729,
    n864,
    n823,
    n881
  );


  nand
  g953
  (
    n985,
    n156,
    n833,
    n868,
    n846
  );


  nor
  g954
  (
    n930,
    n785,
    n705,
    n858,
    n789
  );


  and
  g955
  (
    n948,
    n857,
    n881,
    n859,
    n829
  );


  xor
  g956
  (
    n894,
    n689,
    n743,
    n754,
    n713
  );


  xor
  g957
  (
    n977,
    n837,
    n717,
    n859,
    n744
  );


  and
  g958
  (
    n925,
    n861,
    n832,
    n717,
    n860
  );


  or
  g959
  (
    n888,
    n828,
    n833,
    n732,
    n871
  );


  nor
  g960
  (
    n893,
    n841,
    n866,
    n736,
    n838
  );


  nand
  g961
  (
    n902,
    n721,
    n762,
    n793,
    n748
  );


  nand
  g962
  (
    n968,
    n839,
    n765,
    n847,
    n862
  );


  xnor
  g963
  (
    n941,
    n844,
    n746,
    n865,
    n873
  );


  xor
  g964
  (
    n961,
    n873,
    n790,
    n785,
    n768
  );


  nand
  g965
  (
    n996,
    n727,
    n755,
    n829,
    n870
  );


  nor
  g966
  (
    n910,
    n830,
    n837,
    n826,
    n749
  );


  and
  g967
  (
    n884,
    n735,
    n847,
    n839,
    n746
  );


  nand
  g968
  (
    n954,
    n739,
    n697,
    n691,
    n731
  );


  or
  g969
  (
    n997,
    n823,
    n693,
    n870,
    n875
  );


  or
  g970
  (
    n1024,
    n944,
    n899,
    n886,
    n913
  );


  xnor
  g971
  (
    n1031,
    n965,
    n927,
    n948,
    n990
  );


  xnor
  g972
  (
    n1025,
    n932,
    n978,
    n986,
    n963
  );


  xnor
  g973
  (
    n1022,
    n928,
    n969,
    n961,
    n895
  );


  nor
  g974
  (
    n1016,
    n933,
    n979,
    n968,
    n959
  );


  xnor
  g975
  (
    n1013,
    n946,
    n929,
    n966,
    n994
  );


  nor
  g976
  (
    n1027,
    n983,
    n911,
    n991,
    n917
  );


  nor
  g977
  (
    n1005,
    n937,
    n988,
    n922,
    n952
  );


  nor
  g978
  (
    n1006,
    n920,
    n1000,
    n973,
    n992
  );


  xor
  g979
  (
    n1004,
    n935,
    n940,
    n941,
    n892
  );


  nor
  g980
  (
    n1008,
    n947,
    n890,
    n897,
    n993
  );


  nor
  g981
  (
    n1032,
    n997,
    n962,
    n902,
    n938
  );


  and
  g982
  (
    n1029,
    n955,
    n883,
    n985,
    n945
  );


  and
  g983
  (
    n1030,
    n915,
    n905,
    n910,
    n998
  );


  xnor
  g984
  (
    n1015,
    n943,
    n907,
    n896,
    n974
  );


  and
  g985
  (
    n1012,
    n1001,
    n916,
    n924,
    n887
  );


  and
  g986
  (
    n1019,
    n964,
    n989,
    n918,
    n906
  );


  xor
  g987
  (
    n1018,
    n987,
    n908,
    n967,
    n960
  );


  or
  g988
  (
    n1017,
    n923,
    n894,
    n936,
    n939
  );


  xnor
  g989
  (
    n1010,
    n996,
    n1002,
    n977,
    n984
  );


  nor
  g990
  (
    n1007,
    n900,
    n970,
    n953,
    n980
  );


  and
  g991
  (
    n1021,
    n950,
    n975,
    n972,
    n995
  );


  and
  g992
  (
    n1020,
    n885,
    n901,
    n971,
    n919
  );


  and
  g993
  (
    n1026,
    n981,
    n925,
    n921,
    n934
  );


  xor
  g994
  (
    n1023,
    n914,
    n957,
    n904,
    n893
  );


  nor
  g995
  (
    n1003,
    n884,
    n889,
    n976,
    n888
  );


  and
  g996
  (
    n1009,
    n930,
    n891,
    n931,
    n912
  );


  xnor
  g997
  (
    n1014,
    n951,
    n958,
    n954,
    n926
  );


  xor
  g998
  (
    n1011,
    n956,
    n903,
    n898,
    n909
  );


  or
  g999
  (
    AntiSAT_key_wire,
    n999,
    n982,
    n949,
    n942
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n1028,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

