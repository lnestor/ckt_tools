// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1619_32_1 written by SynthGen on 2021/06/15 15:04:53
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1619_32_1 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39,
 n1525, n1539, n1537, n1538, n1610, n1619, n1620, n1612,
 n1611, n1614, n1628, n1637, n1632, n1643, n1634, n1630,
 n1636, n1642, n1635, n1638, n1640, n1639, n1641, n1631,
 n1629, n1651, n1650, n1653, n1649, n1658, n1654, n1657,
 n1652, n1655, n1656);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39;

output n1525, n1539, n1537, n1538, n1610, n1619, n1620, n1612,
 n1611, n1614, n1628, n1637, n1632, n1643, n1634, n1630,
 n1636, n1642, n1635, n1638, n1640, n1639, n1641, n1631,
 n1629, n1651, n1650, n1653, n1649, n1658, n1654, n1657,
 n1652, n1655, n1656;

wire n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n402, n403, n404, n405, n406, n407,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n425, n426, n427, n428, n429, n430, n431,
 n432, n433, n434, n435, n436, n437, n438, n439,
 n440, n441, n442, n443, n444, n445, n446, n447,
 n448, n449, n450, n451, n452, n453, n454, n455,
 n456, n457, n458, n459, n460, n461, n462, n463,
 n464, n465, n466, n467, n468, n469, n470, n471,
 n472, n473, n474, n475, n476, n477, n478, n479,
 n480, n481, n482, n483, n484, n485, n486, n487,
 n488, n489, n490, n491, n492, n493, n494, n495,
 n496, n497, n498, n499, n500, n501, n502, n503,
 n504, n505, n506, n507, n508, n509, n510, n511,
 n512, n513, n514, n515, n516, n517, n518, n519,
 n520, n521, n522, n523, n524, n525, n526, n527,
 n528, n529, n530, n531, n532, n533, n534, n535,
 n536, n537, n538, n539, n540, n541, n542, n543,
 n544, n545, n546, n547, n548, n549, n550, n551,
 n552, n553, n554, n555, n556, n557, n558, n559,
 n560, n561, n562, n563, n564, n565, n566, n567,
 n568, n569, n570, n571, n572, n573, n574, n575,
 n576, n577, n578, n579, n580, n581, n582, n583,
 n584, n585, n586, n587, n588, n589, n590, n591,
 n592, n593, n594, n595, n596, n597, n598, n599,
 n600, n601, n602, n603, n604, n605, n606, n607,
 n608, n609, n610, n611, n612, n613, n614, n615,
 n616, n617, n618, n619, n620, n621, n622, n623,
 n624, n625, n626, n627, n628, n629, n630, n631,
 n632, n633, n634, n635, n636, n637, n638, n639,
 n640, n641, n642, n643, n644, n645, n646, n647,
 n648, n649, n650, n651, n652, n653, n654, n655,
 n656, n657, n658, n659, n660, n661, n662, n663,
 n664, n665, n666, n667, n668, n669, n670, n671,
 n672, n673, n674, n675, n676, n677, n678, n679,
 n680, n681, n682, n683, n684, n685, n686, n687,
 n688, n689, n690, n691, n692, n693, n694, n695,
 n696, n697, n698, n699, n700, n701, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735,
 n736, n737, n738, n739, n740, n741, n742, n743,
 n744, n745, n746, n747, n748, n749, n750, n751,
 n752, n753, n754, n755, n756, n757, n758, n759,
 n760, n761, n762, n763, n764, n765, n766, n767,
 n768, n769, n770, n771, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n794, n795, n796, n797, n798, n799,
 n800, n801, n802, n803, n804, n805, n806, n807,
 n808, n809, n810, n811, n812, n813, n814, n815,
 n816, n817, n818, n819, n820, n821, n822, n823,
 n824, n825, n826, n827, n828, n829, n830, n831,
 n832, n833, n834, n835, n836, n837, n838, n839,
 n840, n841, n842, n843, n844, n845, n846, n847,
 n848, n849, n850, n851, n852, n853, n854, n855,
 n856, n857, n858, n859, n860, n861, n862, n863,
 n864, n865, n866, n867, n868, n869, n870, n871,
 n872, n873, n874, n875, n876, n877, n878, n879,
 n880, n881, n882, n883, n884, n885, n886, n887,
 n888, n889, n890, n891, n892, n893, n894, n895,
 n896, n897, n898, n899, n900, n901, n902, n903,
 n904, n905, n906, n907, n908, n909, n910, n911,
 n912, n913, n914, n915, n916, n917, n918, n919,
 n920, n921, n922, n923, n924, n925, n926, n927,
 n928, n929, n930, n931, n932, n933, n934, n935,
 n936, n937, n938, n939, n940, n941, n942, n943,
 n944, n945, n946, n947, n948, n949, n950, n951,
 n952, n953, n954, n955, n956, n957, n958, n959,
 n960, n961, n962, n963, n964, n965, n966, n967,
 n968, n969, n970, n971, n972, n973, n974, n975,
 n976, n977, n978, n979, n980, n981, n982, n983,
 n984, n985, n986, n987, n988, n989, n990, n991,
 n992, n993, n994, n995, n996, n997, n998, n999,
 n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
 n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
 n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
 n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
 n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
 n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
 n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
 n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
 n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
 n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
 n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
 n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
 n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
 n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
 n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
 n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
 n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
 n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
 n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
 n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
 n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
 n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
 n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
 n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
 n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
 n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
 n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
 n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
 n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
 n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
 n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
 n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
 n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
 n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
 n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
 n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
 n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
 n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
 n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
 n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
 n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
 n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
 n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
 n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
 n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
 n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
 n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
 n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
 n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
 n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
 n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
 n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
 n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
 n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
 n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
 n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
 n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
 n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
 n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
 n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
 n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
 n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
 n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
 n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
 n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
 n1520, n1521, n1522, n1523, n1524, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
 n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
 n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
 n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
 n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
 n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
 n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
 n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
 n1604, n1605, n1606, n1607, n1608, n1609, n1613, n1615,
 n1616, n1617, n1618, n1621, n1622, n1623, n1624, n1625,
 n1626, n1627, n1633, n1644, n1645, n1646, n1647, n1648;

not  g0 (n47, n32);
not  g1 (n45, n16);
not  g2 (n168, n4);
buf  g3 (n143, n31);
not  g4 (n161, n31);
buf  g5 (n80, n31);
not  g6 (n84, n13);
buf  g7 (n60, n5);
buf  g8 (n171, n35);
buf  g9 (n91, n6);
buf  g10 (n89, n36);
not  g11 (n131, n2);
buf  g12 (n147, n12);
not  g13 (n132, n30);
not  g14 (n90, n22);
not  g15 (n102, n27);
not  g16 (n148, n13);
buf  g17 (n93, n18);
not  g18 (n74, n14);
not  g19 (n153, n10);
buf  g20 (n55, n12);
not  g21 (n160, n7);
not  g22 (n77, n37);
buf  g23 (n92, n29);
buf  g24 (n70, n8);
buf  g25 (n69, n21);
buf  g26 (n157, n5);
buf  g27 (n62, n15);
buf  g28 (n56, n28);
buf  g29 (n122, n27);
buf  g30 (n75, n14);
not  g31 (n96, n15);
not  g32 (n126, n20);
buf  g33 (n94, n24);
buf  g34 (n169, n27);
buf  g35 (n152, n25);
not  g36 (n53, n26);
not  g37 (n124, n29);
not  g38 (n127, n19);
buf  g39 (n177, n33);
not  g40 (n142, n20);
buf  g41 (n64, n8);
not  g42 (n82, n24);
buf  g43 (n117, n28);
buf  g44 (n111, n33);
not  g45 (n166, n31);
not  g46 (n167, n32);
buf  g47 (n46, n11);
not  g48 (n158, n13);
not  g49 (n65, n23);
not  g50 (n57, n17);
not  g51 (n43, n26);
buf  g52 (n134, n7);
not  g53 (n83, n30);
buf  g54 (n86, n4);
buf  g55 (n49, n36);
buf  g56 (n130, n16);
not  g57 (n100, n34);
not  g58 (n144, n23);
buf  g59 (n163, n35);
not  g60 (n165, n6);
not  g61 (n72, n19);
buf  g62 (n50, n18);
buf  g63 (n121, n10);
not  g64 (n112, n14);
buf  g65 (n155, n20);
not  g66 (n42, n25);
buf  g67 (n170, n33);
buf  g68 (n78, n7);
buf  g69 (n99, n23);
not  g70 (n120, n9);
buf  g71 (n145, n9);
not  g72 (n61, n22);
buf  g73 (n41, n10);
not  g74 (n175, n4);
not  g75 (n71, n37);
buf  g76 (n51, n8);
not  g77 (n151, n12);
not  g78 (n140, n15);
not  g79 (n159, n28);
not  g80 (n137, n19);
not  g81 (n114, n5);
not  g82 (n81, n28);
not  g83 (n44, n16);
buf  g84 (n150, n15);
buf  g85 (n59, n26);
buf  g86 (n164, n35);
buf  g87 (n101, n25);
buf  g88 (n156, n23);
not  g89 (n136, n17);
buf  g90 (n76, n21);
buf  g91 (n67, n14);
not  g92 (n129, n19);
buf  g93 (n107, n32);
not  g94 (n146, n8);
buf  g95 (n118, n36);
buf  g96 (n97, n5);
not  g97 (n104, n11);
buf  g98 (n48, n32);
buf  g99 (n162, n33);
not  g100 (n110, n3);
buf  g101 (n172, n17);
buf  g102 (n154, n27);
not  g103 (n68, n24);
not  g104 (n52, n13);
buf  g105 (n103, n34);
buf  g106 (n40, n34);
not  g107 (n58, n16);
buf  g108 (n79, n34);
buf  g109 (n125, n21);
buf  g110 (n135, n9);
buf  g111 (n173, n7);
not  g112 (n63, n22);
not  g113 (n133, n37);
not  g114 (n141, n20);
buf  g115 (n115, n21);
buf  g116 (n54, n18);
not  g117 (n106, n6);
buf  g118 (n119, n11);
not  g119 (n88, n29);
not  g120 (n128, n12);
not  g121 (n108, n30);
not  g122 (n149, n11);
not  g123 (n105, n4);
not  g124 (n116, n17);
buf  g125 (n123, n22);
buf  g126 (n139, n10);
buf  g127 (n174, n6);
buf  g128 (n138, n1);
not  g129 (n98, n24);
not  g130 (n73, n29);
not  g131 (n109, n25);
buf  g132 (n87, n26);
not  g133 (n66, n36);
not  g134 (n113, n35);
not  g135 (n95, n9);
not  g136 (n176, n30);
not  g137 (n85, n18);
buf  g138 (n396, n148);
buf  g139 (n392, n58);
buf  g140 (n362, n120);
not  g141 (n370, n135);
buf  g142 (n301, n92);
not  g143 (n277, n46);
buf  g144 (n343, n94);
buf  g145 (n389, n149);
not  g146 (n286, n49);
not  g147 (n347, n156);
buf  g148 (n247, n48);
buf  g149 (n278, n95);
buf  g150 (n195, n42);
buf  g151 (n365, n159);
buf  g152 (n284, n122);
not  g153 (n314, n164);
buf  g154 (n271, n74);
not  g155 (n291, n160);
not  g156 (n242, n91);
not  g157 (n225, n163);
buf  g158 (n191, n136);
buf  g159 (n305, n142);
buf  g160 (n182, n133);
not  g161 (n267, n169);
not  g162 (n212, n158);
not  g163 (n299, n172);
not  g164 (n334, n170);
not  g165 (n315, n153);
buf  g166 (n394, n128);
not  g167 (n214, n173);
not  g168 (n356, n96);
buf  g169 (n261, n146);
not  g170 (n378, n154);
not  g171 (n197, n61);
not  g172 (n223, n72);
not  g173 (n241, n68);
not  g174 (n181, n139);
not  g175 (n338, n93);
buf  g176 (n279, n137);
not  g177 (n254, n117);
not  g178 (n335, n100);
buf  g179 (n388, n162);
buf  g180 (n207, n173);
buf  g181 (n228, n81);
not  g182 (n302, n112);
buf  g183 (n262, n157);
not  g184 (n339, n102);
buf  g185 (n382, n90);
not  g186 (n189, n89);
buf  g187 (n219, n43);
buf  g188 (n344, n173);
buf  g189 (n321, n153);
not  g190 (n239, n111);
buf  g191 (n198, n131);
buf  g192 (n329, n40);
buf  g193 (n345, n163);
buf  g194 (n250, n41);
buf  g195 (n381, n126);
not  g196 (n213, n54);
buf  g197 (n310, n162);
not  g198 (n357, n156);
not  g199 (n243, n147);
buf  g200 (n322, n110);
buf  g201 (n319, n80);
not  g202 (n235, n51);
buf  g203 (n289, n108);
buf  g204 (n324, n151);
not  g205 (n386, n154);
not  g206 (n205, n158);
not  g207 (n202, n87);
not  g208 (n393, n167);
buf  g209 (n367, n151);
not  g210 (n185, n167);
not  g211 (n255, n168);
not  g212 (n265, n144);
buf  g213 (n385, n171);
not  g214 (n320, n162);
buf  g215 (n318, n116);
not  g216 (n337, n73);
not  g217 (n366, n157);
buf  g218 (n309, n164);
buf  g219 (n358, n147);
not  g220 (n364, n154);
not  g221 (n273, n159);
buf  g222 (n300, n129);
not  g223 (n375, n150);
buf  g224 (n374, n145);
not  g225 (n192, n99);
buf  g226 (n208, n146);
not  g227 (n257, n121);
buf  g228 (n281, n148);
buf  g229 (n333, n169);
not  g230 (n361, n155);
not  g231 (n326, n167);
not  g232 (n221, n84);
buf  g233 (n179, n155);
buf  g234 (n360, n70);
buf  g235 (n316, n134);
not  g236 (n246, n162);
not  g237 (n293, n165);
buf  g238 (n288, n153);
buf  g239 (n311, n124);
not  g240 (n351, n149);
buf  g241 (n236, n138);
buf  g242 (n353, n152);
buf  g243 (n234, n165);
not  g244 (n264, n161);
not  g245 (n204, n170);
buf  g246 (n184, n82);
not  g247 (n331, n119);
not  g248 (n325, n159);
not  g249 (n290, n168);
not  g250 (n248, n167);
buf  g251 (n283, n160);
buf  g252 (n256, n149);
buf  g253 (n298, n63);
not  g254 (n317, n169);
not  g255 (n187, n163);
buf  g256 (n194, n85);
buf  g257 (n216, n141);
not  g258 (n210, n64);
not  g259 (n354, n148);
buf  g260 (n297, n165);
buf  g261 (n183, n79);
buf  g262 (n359, n107);
not  g263 (n259, n168);
not  g264 (n231, n161);
buf  g265 (n227, n161);
not  g266 (n268, n114);
buf  g267 (n330, n171);
buf  g268 (n276, n154);
buf  g269 (n395, n166);
not  g270 (n270, n113);
buf  g271 (n296, n150);
buf  g272 (n178, n161);
buf  g273 (n391, n148);
buf  g274 (n253, n145);
not  g275 (n229, n171);
buf  g276 (n368, n140);
buf  g277 (n222, n147);
buf  g278 (n346, n150);
not  g279 (n280, n130);
buf  g280 (n232, n155);
not  g281 (n252, n76);
not  g282 (n312, n160);
not  g283 (n215, n147);
buf  g284 (n307, n101);
not  g285 (n237, n86);
not  g286 (n352, n103);
not  g287 (n275, n105);
not  g288 (n327, n127);
not  g289 (n211, n78);
buf  g290 (n199, n71);
not  g291 (n372, n67);
buf  g292 (n387, n160);
not  g293 (n295, n125);
buf  g294 (n383, n146);
buf  g295 (n218, n146);
buf  g296 (n379, n166);
not  g297 (n233, n97);
buf  g298 (n282, n171);
buf  g299 (n292, n173);
buf  g300 (n203, n45);
buf  g301 (n209, n83);
buf  g302 (n188, n59);
not  g303 (n244, n98);
buf  g304 (n220, n152);
not  g305 (n313, n55);
buf  g306 (n274, n169);
not  g307 (n303, n44);
not  g308 (n190, n164);
not  g309 (n251, n123);
not  g310 (n272, n168);
not  g311 (n349, n164);
not  g312 (n240, n56);
buf  g313 (n348, n66);
buf  g314 (n230, n143);
not  g315 (n224, n149);
buf  g316 (n308, n115);
buf  g317 (n371, n172);
not  g318 (n390, n104);
not  g319 (n269, n65);
buf  g320 (n200, n69);
not  g321 (n186, n62);
buf  g322 (n397, n109);
not  g323 (n376, n75);
buf  g324 (n332, n52);
not  g325 (n323, n155);
buf  g326 (n369, n174);
not  g327 (n355, n88);
buf  g328 (n380, n158);
buf  g329 (n263, n172);
not  g330 (n363, n170);
buf  g331 (n180, n158);
buf  g332 (n238, n163);
buf  g333 (n193, n157);
buf  g334 (n306, n153);
not  g335 (n350, n132);
not  g336 (n206, n166);
not  g337 (n266, n156);
not  g338 (n196, n166);
buf  g339 (n341, n165);
buf  g340 (n294, n150);
buf  g341 (n249, n57);
not  g342 (n342, n152);
not  g343 (n260, n118);
buf  g344 (n336, n152);
buf  g345 (n226, n172);
buf  g346 (n328, n159);
buf  g347 (n258, n47);
buf  g348 (n377, n106);
not  g349 (n245, n151);
buf  g350 (n287, n151);
buf  g351 (n304, n156);
buf  g352 (n384, n157);
not  g353 (n340, n50);
not  g354 (n217, n77);
buf  g355 (n201, n53);
buf  g356 (n373, n60);
not  g357 (n285, n170);
not  g358 (n715, n301);
buf  g359 (n779, n193);
not  g360 (n590, n263);
buf  g361 (n667, n292);
not  g362 (n569, n197);
not  g363 (n625, n349);
buf  g364 (n520, n350);
not  g365 (n553, n271);
buf  g366 (n435, n296);
not  g367 (n506, n192);
not  g368 (n444, n298);
not  g369 (n863, n265);
buf  g370 (n813, n386);
not  g371 (n727, n312);
buf  g372 (n1041, n315);
buf  g373 (n414, n192);
not  g374 (n424, n392);
buf  g375 (n833, n184);
not  g376 (n891, n259);
not  g377 (n769, n297);
not  g378 (n649, n364);
buf  g379 (n743, n367);
not  g380 (n449, n179);
not  g381 (n431, n211);
buf  g382 (n1042, n239);
buf  g383 (n636, n390);
buf  g384 (n1027, n260);
buf  g385 (n918, n183);
not  g386 (n934, n248);
buf  g387 (n1014, n178);
buf  g388 (n1015, n256);
not  g389 (n429, n202);
buf  g390 (n648, n302);
buf  g391 (n706, n352);
buf  g392 (n895, n367);
not  g393 (n1021, n257);
not  g394 (n577, n243);
not  g395 (n407, n306);
buf  g396 (n1005, n316);
buf  g397 (n929, n254);
not  g398 (n794, n277);
not  g399 (n678, n284);
buf  g400 (n995, n327);
buf  g401 (n511, n238);
not  g402 (n958, n335);
not  g403 (n997, n254);
not  g404 (n627, n391);
not  g405 (n544, n306);
not  g406 (n482, n243);
buf  g407 (n527, n207);
buf  g408 (n723, n197);
buf  g409 (n475, n264);
buf  g410 (n879, n389);
buf  g411 (n717, n206);
buf  g412 (n748, n246);
not  g413 (n543, n263);
not  g414 (n848, n217);
buf  g415 (n865, n396);
not  g416 (n498, n295);
not  g417 (n658, n231);
buf  g418 (n812, n212);
not  g419 (n936, n227);
not  g420 (n808, n305);
buf  g421 (n824, n252);
not  g422 (n840, n251);
buf  g423 (n857, n178);
buf  g424 (n476, n341);
buf  g425 (n460, n205);
buf  g426 (n613, n308);
not  g427 (n508, n279);
not  g428 (n841, n383);
not  g429 (n835, n319);
not  g430 (n777, n310);
buf  g431 (n898, n268);
not  g432 (n878, n397);
buf  g433 (n797, n383);
buf  g434 (n581, n283);
buf  g435 (n599, n229);
not  g436 (n602, n330);
buf  g437 (n849, n367);
not  g438 (n593, n267);
buf  g439 (n826, n228);
buf  g440 (n643, n240);
not  g441 (n908, n247);
not  g442 (n564, n256);
buf  g443 (n888, n250);
not  g444 (n696, n219);
buf  g445 (n802, n319);
not  g446 (n418, n393);
buf  g447 (n950, n353);
not  g448 (n796, n234);
not  g449 (n529, n315);
not  g450 (n585, n391);
not  g451 (n647, n392);
not  g452 (n746, n373);
not  g453 (n709, n237);
buf  g454 (n839, n273);
buf  g455 (n832, n378);
not  g456 (n959, n269);
not  g457 (n881, n238);
not  g458 (n909, n239);
not  g459 (n586, n321);
not  g460 (n1046, n356);
buf  g461 (n838, n282);
buf  g462 (n622, n275);
not  g463 (n971, n366);
not  g464 (n1010, n251);
not  g465 (n740, n240);
buf  g466 (n415, n185);
not  g467 (n861, n363);
buf  g468 (n720, n274);
buf  g469 (n912, n314);
buf  g470 (n547, n333);
buf  g471 (n651, n376);
buf  g472 (n836, n324);
not  g473 (n922, n301);
not  g474 (n781, n275);
buf  g475 (n852, n189);
not  g476 (n1056, n237);
buf  g477 (n565, n226);
not  g478 (n481, n386);
buf  g479 (n489, n181);
buf  g480 (n983, n320);
buf  g481 (n919, n397);
buf  g482 (n722, n199);
buf  g483 (n1020, n253);
not  g484 (n550, n379);
not  g485 (n731, n222);
not  g486 (n539, n199);
not  g487 (n528, n214);
not  g488 (n710, n388);
not  g489 (n906, n205);
buf  g490 (n662, n376);
not  g491 (n1007, n209);
not  g492 (n1053, n250);
not  g493 (n533, n323);
buf  g494 (n799, n325);
not  g495 (n583, n288);
buf  g496 (n432, n191);
not  g497 (n611, n393);
not  g498 (n792, n372);
buf  g499 (n608, n278);
buf  g500 (n981, n233);
not  g501 (n1019, n340);
buf  g502 (n409, n178);
not  g503 (n1052, n295);
buf  g504 (n855, n360);
buf  g505 (n1045, n286);
not  g506 (n567, n230);
buf  g507 (n926, n244);
buf  g508 (n921, n270);
buf  g509 (n478, n342);
not  g510 (n523, n283);
not  g511 (n494, n394);
not  g512 (n614, n188);
not  g513 (n411, n230);
not  g514 (n837, n219);
buf  g515 (n516, n259);
buf  g516 (n561, n369);
not  g517 (n576, n292);
buf  g518 (n862, n180);
buf  g519 (n421, n320);
buf  g520 (n700, n331);
not  g521 (n635, n322);
buf  g522 (n461, n372);
buf  g523 (n521, n224);
not  g524 (n964, n300);
buf  g525 (n470, n284);
not  g526 (n616, n395);
not  g527 (n745, n178);
buf  g528 (n509, n191);
not  g529 (n440, n357);
not  g530 (n446, n222);
not  g531 (n448, n275);
buf  g532 (n1044, n320);
not  g533 (n554, n217);
not  g534 (n619, n257);
buf  g535 (n659, n302);
buf  g536 (n398, n199);
buf  g537 (n988, n365);
buf  g538 (n970, n319);
not  g539 (n692, n321);
buf  g540 (n897, n341);
buf  g541 (n853, n208);
not  g542 (n755, n396);
not  g543 (n699, n337);
not  g544 (n677, n304);
buf  g545 (n1000, n285);
not  g546 (n454, n356);
buf  g547 (n707, n305);
not  g548 (n491, n289);
buf  g549 (n675, n355);
not  g550 (n977, n193);
not  g551 (n534, n243);
buf  g552 (n1058, n366);
not  g553 (n526, n186);
buf  g554 (n883, n395);
not  g555 (n472, n372);
buf  g556 (n473, n233);
not  g557 (n428, n241);
buf  g558 (n546, n384);
buf  g559 (n1036, n377);
buf  g560 (n538, n255);
buf  g561 (n1009, n265);
buf  g562 (n517, n311);
not  g563 (n789, n377);
not  g564 (n673, n223);
not  g565 (n525, n209);
buf  g566 (n617, n302);
not  g567 (n400, n358);
not  g568 (n633, n342);
not  g569 (n917, n246);
not  g570 (n939, n289);
not  g571 (n920, n347);
not  g572 (n656, n252);
buf  g573 (n911, n299);
buf  g574 (n626, n280);
buf  g575 (n930, n295);
not  g576 (n637, n260);
buf  g577 (n856, n194);
buf  g578 (n902, n332);
buf  g579 (n828, n282);
not  g580 (n843, n380);
not  g581 (n782, n389);
not  g582 (n1011, n212);
not  g583 (n725, n220);
not  g584 (n864, n338);
not  g585 (n992, n379);
buf  g586 (n890, n328);
not  g587 (n702, n228);
buf  g588 (n447, n286);
buf  g589 (n767, n179);
buf  g590 (n773, n339);
buf  g591 (n969, n219);
not  g592 (n598, n371);
not  g593 (n882, n273);
buf  g594 (n660, n340);
not  g595 (n935, n222);
not  g596 (n972, n314);
buf  g597 (n805, n312);
not  g598 (n504, n218);
not  g599 (n697, n240);
buf  g600 (n798, n349);
buf  g601 (n433, n285);
buf  g602 (n910, n378);
buf  g603 (n962, n307);
not  g604 (n500, n235);
buf  g605 (n928, n273);
not  g606 (n787, n204);
buf  g607 (n994, n221);
not  g608 (n750, n290);
buf  g609 (n519, n224);
not  g610 (n795, n182);
buf  g611 (n819, n352);
not  g612 (n445, n204);
buf  g613 (n587, n232);
buf  g614 (n807, n334);
not  g615 (n427, n393);
not  g616 (n634, n264);
not  g617 (n718, n267);
buf  g618 (n416, n388);
buf  g619 (n495, n311);
not  g620 (n987, n180);
buf  g621 (n595, n370);
not  g622 (n542, n245);
buf  g623 (n899, n213);
not  g624 (n548, n346);
not  g625 (n701, n336);
not  g626 (n758, n208);
not  g627 (n893, n332);
not  g628 (n744, n243);
buf  g629 (n557, n272);
not  g630 (n681, n270);
buf  g631 (n483, n303);
buf  g632 (n570, n211);
buf  g633 (n632, n228);
buf  g634 (n698, n203);
buf  g635 (n612, n246);
buf  g636 (n621, n354);
not  g637 (n628, n337);
not  g638 (n484, n252);
not  g639 (n674, n350);
buf  g640 (n721, n263);
buf  g641 (n426, n353);
not  g642 (n954, n264);
buf  g643 (n846, n303);
not  g644 (n873, n206);
not  g645 (n676, n215);
buf  g646 (n610, n278);
buf  g647 (n584, n242);
buf  g648 (n956, n310);
not  g649 (n1034, n223);
buf  g650 (n640, n287);
buf  g651 (n459, n273);
not  g652 (n502, n269);
buf  g653 (n563, n371);
buf  g654 (n984, n195);
not  g655 (n742, n220);
buf  g656 (n551, n357);
buf  g657 (n1012, n198);
not  g658 (n671, n323);
buf  g659 (n624, n258);
not  g660 (n940, n208);
buf  g661 (n747, n382);
buf  g662 (n901, n277);
buf  g663 (n993, n362);
not  g664 (n916, n278);
buf  g665 (n809, n231);
not  g666 (n961, n235);
buf  g667 (n947, n328);
not  g668 (n847, n271);
not  g669 (n804, n264);
buf  g670 (n915, n224);
not  g671 (n402, n193);
buf  g672 (n594, n358);
not  g673 (n1002, n335);
buf  g674 (n949, n358);
buf  g675 (n403, n186);
not  g676 (n946, n271);
not  g677 (n726, n368);
buf  g678 (n457, n306);
not  g679 (n914, n293);
not  g680 (n1028, n229);
buf  g681 (n800, n332);
not  g682 (n765, n306);
buf  g683 (n412, n307);
buf  g684 (n859, n342);
not  g685 (n965, n310);
buf  g686 (n844, n386);
not  g687 (n686, n221);
not  g688 (n401, n203);
not  g689 (n762, n336);
buf  g690 (n752, n348);
not  g691 (n514, n336);
not  g692 (n945, n345);
buf  g693 (n575, n388);
not  g694 (n1035, n262);
not  g695 (n596, n274);
not  g696 (n605, n233);
buf  g697 (n406, n359);
buf  g698 (n405, n378);
not  g699 (n708, n211);
not  g700 (n501, n326);
buf  g701 (n486, n385);
not  g702 (n803, n255);
not  g703 (n763, n298);
buf  g704 (n786, n195);
buf  g705 (n711, n234);
not  g706 (n927, n225);
buf  g707 (n887, n247);
buf  g708 (n513, n384);
not  g709 (n704, n314);
not  g710 (n810, n387);
not  g711 (n785, n232);
not  g712 (n738, n308);
buf  g713 (n858, n371);
not  g714 (n817, n343);
not  g715 (n1043, n217);
not  g716 (n733, n383);
not  g717 (n1026, n326);
not  g718 (n452, n301);
buf  g719 (n467, n346);
not  g720 (n688, n234);
not  g721 (n896, n260);
buf  g722 (n991, n325);
not  g723 (n854, n355);
not  g724 (n531, n322);
buf  g725 (n772, n205);
not  g726 (n820, n369);
not  g727 (n463, n309);
not  g728 (n978, n336);
not  g729 (n1047, n257);
not  g730 (n474, n269);
buf  g731 (n724, n341);
not  g732 (n420, n378);
not  g733 (n712, n374);
buf  g734 (n1008, n331);
not  g735 (n1055, n316);
not  g736 (n597, n345);
not  g737 (n668, n183);
not  g738 (n591, n261);
not  g739 (n572, n300);
not  g740 (n1017, n338);
buf  g741 (n540, n215);
buf  g742 (n822, n229);
buf  g743 (n477, n250);
buf  g744 (n979, n183);
not  g745 (n791, n196);
buf  g746 (n573, n393);
buf  g747 (n552, n383);
not  g748 (n653, n325);
not  g749 (n719, n291);
not  g750 (n682, n292);
buf  g751 (n754, n364);
buf  g752 (n904, n237);
not  g753 (n937, n194);
buf  g754 (n757, n370);
buf  g755 (n793, n198);
not  g756 (n1033, n246);
buf  g757 (n751, n208);
not  g758 (n644, n214);
not  g759 (n884, n270);
buf  g760 (n963, n291);
not  g761 (n530, n354);
not  g762 (n960, n187);
buf  g763 (n980, n296);
buf  g764 (n1048, n324);
not  g765 (n1004, n317);
not  g766 (n689, n206);
buf  g767 (n571, n196);
buf  g768 (n766, n366);
buf  g769 (n623, n361);
not  g770 (n739, n392);
not  g771 (n771, n256);
buf  g772 (n680, n299);
not  g773 (n652, n304);
buf  g774 (n600, n241);
buf  g775 (n1050, n321);
not  g776 (n430, n396);
buf  g777 (n549, n203);
buf  g778 (n986, n190);
buf  g779 (n580, n370);
buf  g780 (n880, n329);
not  g781 (n574, n353);
buf  g782 (n606, n337);
not  g783 (n641, n365);
not  g784 (n434, n233);
buf  g785 (n455, n376);
not  g786 (n1025, n202);
not  g787 (n734, n182);
buf  g788 (n737, n280);
buf  g789 (n441, n283);
not  g790 (n685, n239);
not  g791 (n556, n337);
buf  g792 (n691, n363);
not  g793 (n933, n268);
buf  g794 (n955, n385);
not  g795 (n818, n236);
not  g796 (n438, n293);
not  g797 (n876, n346);
not  g798 (n578, n188);
not  g799 (n604, n184);
not  g800 (n631, n394);
not  g801 (n1040, n209);
buf  g802 (n907, n333);
not  g803 (n825, n290);
not  g804 (n664, n202);
not  g805 (n996, n339);
not  g806 (n823, n276);
buf  g807 (n753, n238);
not  g808 (n872, n245);
not  g809 (n510, n365);
buf  g810 (n518, n245);
not  g811 (n683, n216);
not  g812 (n953, n362);
not  g813 (n1049, n358);
buf  g814 (n666, n198);
buf  g815 (n1032, n381);
buf  g816 (n404, n204);
buf  g817 (n588, n352);
not  g818 (n670, n210);
buf  g819 (n894, n222);
buf  g820 (n776, n213);
not  g821 (n493, n375);
not  g822 (n694, n254);
buf  g823 (n875, n363);
not  g824 (n905, n362);
buf  g825 (n931, n309);
not  g826 (n801, n348);
buf  g827 (n422, n298);
buf  g828 (n713, n312);
not  g829 (n469, n382);
buf  g830 (n827, n260);
not  g831 (n1018, n191);
not  g832 (n973, n196);
buf  g833 (n638, n258);
not  g834 (n399, n197);
buf  g835 (n437, n186);
buf  g836 (n761, n269);
not  g837 (n480, n322);
buf  g838 (n778, n184);
buf  g839 (n942, n265);
not  g840 (n952, n344);
buf  g841 (n1038, n226);
not  g842 (n989, n205);
buf  g843 (n487, n185);
not  g844 (n439, n278);
buf  g845 (n735, n216);
not  g846 (n545, n335);
buf  g847 (n866, n214);
not  g848 (n1039, n202);
buf  g849 (n741, n200);
not  g850 (n464, n375);
buf  g851 (n496, n200);
not  g852 (n1003, n242);
not  g853 (n537, n244);
buf  g854 (n515, n360);
buf  g855 (n492, n218);
buf  g856 (n886, n307);
not  g857 (n642, n287);
buf  g858 (n885, n321);
buf  g859 (n1024, n225);
buf  g860 (n497, n351);
not  g861 (n589, n227);
buf  g862 (n541, n391);
buf  g863 (n669, n284);
not  g864 (n488, n381);
buf  g865 (n985, n285);
buf  g866 (n975, n262);
not  g867 (n609, n242);
not  g868 (n654, n237);
buf  g869 (n871, n226);
not  g870 (n982, n258);
not  g871 (n788, n384);
not  g872 (n976, n254);
not  g873 (n1022, n381);
not  g874 (n410, n193);
buf  g875 (n684, n330);
not  g876 (n579, n296);
not  g877 (n607, n369);
not  g878 (n568, n274);
not  g879 (n471, n357);
not  g880 (n450, n188);
not  g881 (n672, n236);
not  g882 (n774, n360);
buf  g883 (n913, n385);
buf  g884 (n900, n397);
not  g885 (n522, n351);
not  g886 (n558, n211);
buf  g887 (n941, n286);
buf  g888 (n639, n190);
buf  g889 (n889, n187);
not  g890 (n466, n310);
buf  g891 (n999, n353);
not  g892 (n749, n297);
not  g893 (n821, n218);
not  g894 (n442, n374);
not  g895 (n957, n216);
not  g896 (n768, n236);
not  g897 (n695, n277);
buf  g898 (n645, n384);
not  g899 (n629, n201);
buf  g900 (n566, n207);
not  g901 (n829, n261);
not  g902 (n990, n287);
buf  g903 (n1030, n196);
buf  g904 (n1013, n223);
not  g905 (n601, n389);
buf  g906 (n1054, n268);
buf  g907 (n968, n180);
not  g908 (n456, n346);
buf  g909 (n998, n341);
not  g910 (n663, n333);
buf  g911 (n592, n325);
buf  g912 (n729, n218);
buf  g913 (n687, n214);
buf  g914 (n1031, n228);
not  g915 (n944, n377);
not  g916 (n732, n281);
buf  g917 (n764, n212);
buf  g918 (n503, n181);
not  g919 (n615, n374);
buf  g920 (n903, n187);
not  g921 (n775, n298);
buf  g922 (n655, n294);
not  g923 (n524, n327);
not  g924 (n1023, n272);
not  g925 (n535, n313);
not  g926 (n559, n344);
not  g927 (n850, n357);
not  g928 (n728, n324);
not  g929 (n618, n304);
not  g930 (n790, n281);
buf  g931 (n967, n351);
buf  g932 (n693, n261);
buf  g933 (n714, n207);
not  g934 (n419, n352);
buf  g935 (n485, n179);
not  g936 (n874, n242);
buf  g937 (n408, n354);
buf  g938 (n436, n380);
not  g939 (n1001, n387);
not  g940 (n815, n338);
buf  g941 (n1037, n257);
not  g942 (n650, n355);
buf  g943 (n924, n232);
not  g944 (n679, n297);
not  g945 (n831, n335);
xnor g946 (n860, n368, n397, n351, n339);
xor  g947 (n736, n290, n295, n373, n230);
nor  g948 (n560, n266, n305, n380, n289);
or   g949 (n665, n290, n226, n255, n302);
nor  g950 (n834, n318, n387, n207, n316);
and  g951 (n462, n198, n181, n209, n253);
nor  g952 (n458, n220, n291, n203, n363);
or   g953 (n690, n230, n244, n315, n251);
or   g954 (n716, n359, n345, n340, n194);
nor  g955 (n938, n241, n354, n210, n280);
xor  g956 (n505, n261, n368, n227, n293);
and  g957 (n811, n389, n285, n376, n314);
xnor g958 (n784, n326, n372, n192, n267);
or   g959 (n816, n220, n251, n350, n317);
nand g960 (n923, n225, n272, n183, n255);
xnor g961 (n630, n309, n381, n250, n268);
or   g962 (n1006, n229, n245, n348, n394);
or   g963 (n830, n394, n239, n344, n395);
or   g964 (n868, n333, n288, n247, n259);
nor  g965 (n1016, n283, n199, n281, n201);
xnor g966 (n479, n320, n221, n343, n380);
and  g967 (n468, n331, n340, n396, n364);
nor  g968 (n925, n235, n280, n329, n215);
or   g969 (n582, n181, n369, n313, n185);
or   g970 (n603, n279, n390, n327, n322);
nor  g971 (n892, n263, n194, n317, n299);
and  g972 (n806, n217, n329, n324, n267);
or   g973 (n867, n334, n188, n215, n201);
xnor g974 (n512, n232, n319, n249, n361);
xor  g975 (n974, n288, n359, n382, n297);
nor  g976 (n951, n266, n315, n300, n391);
xor  g977 (n760, n248, n270, n249, n318);
xor  g978 (n948, n276, n216, n294, n356);
nand g979 (n703, n265, n356, n392, n362);
nand g980 (n1057, n360, n311, n179, n332);
or   g981 (n532, n182, n291, n307, n231);
or   g982 (n759, n349, n189, n326, n289);
xor  g983 (n646, n288, n374, n274, n293);
nor  g984 (n490, n390, n344, n375, n189);
xor  g985 (n413, n276, n292, n190, n224);
nand g986 (n966, n312, n191, n355, n309);
nor  g987 (n756, n195, n223, n281, n316);
xor  g988 (n1051, n338, n186, n313, n249);
nand g989 (n851, n365, n252, n238, n277);
or   g990 (n425, n359, n253, n296, n367);
nor  g991 (n555, n219, n349, n386, n301);
xnor g992 (n451, n328, n189, n347, n248);
nor  g993 (n780, n387, n266, n271, n361);
nand g994 (n620, n258, n204, n368, n262);
xor  g995 (n814, n347, n240, n279, n236);
xor  g996 (n943, n373, n190, n377, n303);
and  g997 (n870, n299, n330, n347, n317);
xnor g998 (n499, n334, n350, n328, n305);
xnor g999 (n869, n284, n247, n327, n275);
or   g1000 (n730, n244, n375, n379, n249);
xor  g1001 (n507, n262, n379, n212, n308);
and  g1002 (n562, n323, n221, n201, n180);
or   g1003 (n845, n318, n287, n342, n266);
xor  g1004 (n661, n279, n395, n256, n330);
xor  g1005 (n453, n294, n234, n390, n282);
nand g1006 (n877, n339, n200, n231, n276);
xor  g1007 (n1029, n388, n343, n366, n385);
xnor g1008 (n443, n184, n294, n348, n345);
xnor g1009 (n423, n313, n334, n311, n382);
nor  g1010 (n705, n185, n308, n323, n210);
xnor g1011 (n770, n213, n225, n206, n303);
nand g1012 (n783, n331, n182, n210, n197);
and  g1013 (n536, n282, n373, n300, n371);
xor  g1014 (n465, n253, n227, n195, n272);
nand g1015 (n842, n213, n364, n286, n248);
xor  g1016 (n417, n329, n304, n343, n259);
xnor g1017 (n932, n318, n241, n192, n235);
xor  g1018 (n657, n361, n200, n187, n370);
or   g1019 (n1074, n551, n457, n789, n429);
xor  g1020 (n1085, n539, n683, n840, n553);
nand g1021 (n1121, n529, n795, n565, n451);
xnor g1022 (n1172, n721, n688, n643, n412);
xnor g1023 (n1160, n636, n908, n434, n816);
xor  g1024 (n1153, n727, n562, n824, n420);
nand g1025 (n1127, n768, n668, n557, n530);
nand g1026 (n1155, n836, n411, n606, n613);
or   g1027 (n1147, n733, n750, n794, n574);
xnor g1028 (n1132, n588, n525, n728, n575);
xor  g1029 (n1063, n459, n738, n492, n855);
xor  g1030 (n1099, n642, n475, n659, n616);
xnor g1031 (n1087, n674, n497, n503, n607);
xnor g1032 (n1165, n630, n481, n569, n909);
nor  g1033 (n1122, n517, n414, n788, n784);
xor  g1034 (n1175, n637, n640, n549, n535);
nor  g1035 (n1174, n604, n558, n469, n678);
and  g1036 (n1119, n744, n447, n591, n596);
nor  g1037 (n1113, n899, n473, n739, n778);
xnor g1038 (n1167, n566, n590, n536, n452);
xnor g1039 (n1126, n781, n725, n737, n699);
and  g1040 (n1186, n670, n743, n443, n520);
nor  g1041 (n1089, n560, n757, n495, n809);
or   g1042 (n1060, n792, n458, n564, n639);
xnor g1043 (n1073, n599, n779, n409, n417);
xor  g1044 (n1177, n680, n446, n839, n532);
or   g1045 (n1066, n405, n504, n499, n759);
xnor g1046 (n1136, n843, n402, n505, n802);
xnor g1047 (n1114, n877, n518, n437, n398);
xnor g1048 (n1168, n449, n807, n478, n825);
nor  g1049 (n1183, n863, n658, n489, n468);
nand g1050 (n1094, n881, n701, n498, n656);
nor  g1051 (n1143, n718, n764, n787, n598);
nand g1052 (n1170, n577, n521, n480, n772);
or   g1053 (n1117, n651, n780, n608, n901);
xnor g1054 (n1163, n769, n586, n887, n399);
xor  g1055 (n1148, n682, n485, n556, n488);
xor  g1056 (n1071, n482, n403, n477, n888);
xnor g1057 (n1091, n673, n775, n548, n799);
and  g1058 (n1161, n552, n430, n646, n878);
xnor g1059 (n1059, n634, n767, n490, n770);
nand g1060 (n1100, n442, n421, n664, n587);
and  g1061 (n1134, n626, n568, n828, n419);
and  g1062 (n1115, n487, n423, n837, n435);
nand g1063 (n1065, n691, n791, n461, n804);
or   g1064 (n1109, n713, n415, n818, n748);
nor  g1065 (n1144, n486, n508, n675, n669);
xnor g1066 (n1101, n885, n777, n582, n762);
nor  g1067 (n1173, n677, n693, n635, n666);
xor  g1068 (n1118, n621, n709, n690, n559);
or   g1069 (n1107, n844, n722, n614, n679);
nand g1070 (n1124, n870, n823, n662, n858);
nand g1071 (n1080, n796, n879, n522, n790);
xnor g1072 (n1083, n861, n523, n502, n612);
nor  g1073 (n1095, n627, n644, n515, n864);
xor  g1074 (n1072, n715, n745, n689, n652);
nand g1075 (n1108, n866, n584, n544, n433);
nor  g1076 (n1125, n625, n650, n705, n852);
xor  g1077 (n1096, n793, n413, n467, n841);
xnor g1078 (n1164, n883, n734, n810, n550);
xor  g1079 (n1162, n755, n814, n526, n519);
xnor g1080 (n1102, n661, n826, n890, n835);
and  g1081 (n1176, n660, n753, n605, n867);
or   g1082 (n1088, n479, n638, n424, n506);
xor  g1083 (n1110, n484, n404, n408, n501);
nand g1084 (n1152, n869, n692, n578, n554);
xnor g1085 (n1068, n425, n533, n774, n902);
nand g1086 (n1184, n717, n573, n712, n834);
or   g1087 (n1082, n815, n538, n724, n742);
xnor g1088 (n1070, n628, n454, n812, n471);
xor  g1089 (n1141, n831, n561, n821, n893);
or   g1090 (n1185, n440, n813, n543, n541);
and  g1091 (n1106, n580, n747, n401, n703);
nor  g1092 (n1157, n882, n589, n545, n464);
nor  g1093 (n1146, n798, n624, n555, n672);
nand g1094 (n1064, n513, n845, n862, n752);
nor  g1095 (n1061, n681, n671, n832, n460);
nor  g1096 (n1138, n874, n428, n441, n426);
nor  g1097 (n1062, n450, n884, n524, n579);
nand g1098 (n1097, n763, n886, n771, n811);
xor  g1099 (n1151, n455, n773, n494, n629);
and  g1100 (n1075, n406, n463, n873, n546);
xnor g1101 (n1137, n619, n740, n422, n849);
xnor g1102 (n1103, n857, n594, n694, n611);
or   g1103 (n1086, n853, n697, n581, n714);
nor  g1104 (n1181, n906, n766, n758, n645);
xor  g1105 (n1178, n685, n500, n765, n407);
or   g1106 (n1079, n601, n547, n410, n622);
xnor g1107 (n1179, n905, n817, n749, n875);
xnor g1108 (n1084, n527, n592, n702, n856);
and  g1109 (n1081, n648, n760, n491, n465);
and  g1110 (n1145, n438, n631, n496, n453);
or   g1111 (n1123, n400, n667, n512, n756);
and  g1112 (n1130, n829, n432, n830, n786);
xnor g1113 (n1182, n585, n716, n900, n860);
and  g1114 (n1166, n448, n700, n708, n754);
xnor g1115 (n1171, n761, n903, n620, n618);
xnor g1116 (n1158, n597, n805, n583, n880);
xnor g1117 (n1140, n706, n483, n842, n665);
nand g1118 (n1116, n704, n735, n595, n808);
nand g1119 (n1169, n603, n470, n695, n531);
and  g1120 (n1092, n570, n686, n609, n847);
and  g1121 (n1090, n801, n472, n820, n846);
or   g1122 (n1150, n466, n427, n436, n707);
nor  g1123 (n1111, n797, n871, n782, n510);
nor  g1124 (n1105, n563, n850, n439, n610);
xor  g1125 (n1098, n676, n741, n444, n723);
nor  g1126 (n1093, n615, n736, n868, n663);
nor  g1127 (n1069, n567, n537, n746, n833);
xnor g1128 (n1076, n730, n800, n896, n571);
or   g1129 (n1078, n848, n540, n516, n687);
nand g1130 (n1156, n593, n726, n456, n418);
xor  g1131 (n1135, n576, n633, n649, n783);
xor  g1132 (n1112, n719, n785, n416, n528);
xnor g1133 (n1159, n751, n872, n827, n865);
or   g1134 (n1077, n534, n819, n710, n892);
or   g1135 (n1142, n509, n895, n851, n776);
xor  g1136 (n1131, n854, n696, n632, n889);
or   g1137 (n1104, n898, n514, n654, n657);
or   g1138 (n1180, n476, n907, n729, n838);
or   g1139 (n1154, n623, n894, n431, n822);
nor  g1140 (n1133, n655, n507, n462, n684);
and  g1141 (n1129, n859, n653, n542, n641);
nor  g1142 (n1067, n897, n803, n731, n904);
or   g1143 (n1128, n602, n732, n600, n572);
nor  g1144 (n1139, n493, n891, n711, n698);
xnor g1145 (n1149, n876, n806, n617, n720);
and  g1146 (n1120, n511, n445, n474, n647);
buf  g1147 (n1197, n1080);
not  g1148 (n1205, n1081);
not  g1149 (n1213, n1090);
buf  g1150 (n1196, n1084);
buf  g1151 (n1190, n1089);
not  g1152 (n1218, n1066);
buf  g1153 (n1195, n1060);
buf  g1154 (n1212, n1078);
not  g1155 (n1191, n1088);
not  g1156 (n1192, n1075);
not  g1157 (n1204, n1087);
buf  g1158 (n1200, n1072);
not  g1159 (n1187, n1070);
buf  g1160 (n1211, n1077);
not  g1161 (n1215, n1067);
buf  g1162 (n1208, n1068);
not  g1163 (n1210, n1074);
buf  g1164 (n1203, n1061);
buf  g1165 (n1199, n1079);
buf  g1166 (n1189, n1083);
not  g1167 (n1198, n1062);
not  g1168 (n1206, n1064);
not  g1169 (n1217, n1085);
buf  g1170 (n1201, n1073);
buf  g1171 (n1207, n1069);
buf  g1172 (n1214, n1071);
buf  g1173 (n1216, n1082);
buf  g1174 (n1194, n1063);
not  g1175 (n1188, n1065);
buf  g1176 (n1193, n1076);
buf  g1177 (n1202, n1086);
buf  g1178 (n1209, n1059);
xor  g1179 (n1226, n1193, n1189);
nand g1180 (n1220, n1190, n1091);
nor  g1181 (n1222, n1199, n1198);
xnor g1182 (n1221, n1196, n1187);
xor  g1183 (n1219, n1197, n1194);
nand g1184 (n1225, n1195, n1188);
xnor g1185 (n1224, n1192, n1200);
and  g1186 (n1223, n1199, n1191);
xnor g1187 (n1235, n1221, n1225, n1226);
nand g1188 (n1234, n1204, n1206, n1226);
or   g1189 (n1227, n1201, n1202, n1220);
or   g1190 (n1231, n1204, n1225, n1203);
and  g1191 (n1230, n1205, n1203, n1222);
nor  g1192 (n1228, n1203, n1205, n1204);
xor  g1193 (n1233, n1204, n1202);
xnor g1194 (n1232, n1202, n1203, n1201);
or   g1195 (n1236, n1219, n1205, n1223);
xnor g1196 (n1229, n1200, n1201, n1224);
xnor g1197 (n1237, n943, n920, n1236, n933);
xnor g1198 (n1266, n991, n910, n1207);
xnor g1199 (n1272, n912, n1207, n930, n1229);
and  g1200 (n1276, n1209, n1228, n1006, n934);
xor  g1201 (n1273, n941, n927, n996, n1001);
or   g1202 (n1253, n1228, n940, n924, n1231);
xor  g1203 (n1249, n1231, n953, n952, n945);
xor  g1204 (n1267, n981, n1230, n979, n1231);
or   g1205 (n1268, n936, n970, n1003, n1227);
xor  g1206 (n1247, n959, n928, n1209, n938);
nand g1207 (n1254, n1100, n1000, n966, n913);
nor  g1208 (n1262, n963, n1207, n1098, n957);
nand g1209 (n1269, n990, n1229, n972, n977);
or   g1210 (n1263, n998, n914, n931, n1206);
or   g1211 (n1256, n1231, n932, n915, n971);
and  g1212 (n1274, n988, n976, n1232, n1235);
xnor g1213 (n1240, n1234, n1233, n965, n978);
or   g1214 (n1242, n1232, n1233, n958, n985);
nand g1215 (n1257, n946, n926, n1235, n984);
xnor g1216 (n1248, n1233, n989, n1235, n917);
or   g1217 (n1271, n937, n935, n1096, n1004);
or   g1218 (n1255, n918, n1206, n964);
or   g1219 (n1261, n1208, n942, n925, n992);
nor  g1220 (n1265, n929, n1228, n1002, n916);
xor  g1221 (n1264, n1228, n1232, n987, n919);
or   g1222 (n1260, n1233, n973, n962, n1230);
or   g1223 (n1239, n999, n983, n967, n961);
xnor g1224 (n1259, n1094, n1229, n993);
xnor g1225 (n1270, n950, n1234, n982);
or   g1226 (n1246, n923, n1230, n1093, n921);
and  g1227 (n1245, n1236, n948, n974, n949);
nor  g1228 (n1241, n1227, n975, n956, n944);
or   g1229 (n1258, n980, n1007, n951, n939);
nand g1230 (n1244, n969, n1232, n994, n1230);
or   g1231 (n1251, n1227, n955, n947, n1095);
nor  g1232 (n1243, n1208, n1235, n968, n1099);
or   g1233 (n1250, n1234, n1092, n1236, n1227);
or   g1234 (n1252, n986, n954, n1005, n1097);
xnor g1235 (n1275, n960, n1208, n911);
or   g1236 (n1238, n922, n995, n997, n1236);
or   g1237 (n1280, n1115, n1111, n1106, n1237);
nor  g1238 (n1282, n1104, n1114, n1112, n1238);
xor  g1239 (n1277, n1238, n1117, n1237, n1110);
xor  g1240 (n1279, n1237, n1101, n1113, n1109);
and  g1241 (n1278, n1102, n1103, n1237, n1108);
and  g1242 (n1281, n1116, n1105, n1118, n1107);
buf  g1243 (n1295, n1280);
not  g1244 (n1298, n1281);
not  g1245 (n1283, n1282);
not  g1246 (n1292, n1209);
buf  g1247 (n1296, n1282);
buf  g1248 (n1286, n1277);
buf  g1249 (n1284, n1282);
buf  g1250 (n1293, n1279);
not  g1251 (n1285, n1281);
not  g1252 (n1297, n1280);
not  g1253 (n1290, n1281);
buf  g1254 (n1289, n1280);
not  g1255 (n1287, n1211);
xor  g1256 (n1299, n1278, n1210);
xnor g1257 (n1291, n1279, n1210);
xor  g1258 (n1294, n1282, n1281, n1210);
xor  g1259 (n1288, n1209, n1278, n1280);
buf  g1260 (n1310, n1298);
buf  g1261 (n1343, n1294);
buf  g1262 (n1355, n1284);
not  g1263 (n1346, n1293);
buf  g1264 (n1302, n1286);
not  g1265 (n1321, n1213);
buf  g1266 (n1304, n1296);
buf  g1267 (n1354, n1297);
buf  g1268 (n1352, n1299);
not  g1269 (n1347, n1298);
not  g1270 (n1309, n1287);
buf  g1271 (n1327, n1286);
not  g1272 (n1357, n1292);
not  g1273 (n1341, n1286);
not  g1274 (n1315, n1214);
not  g1275 (n1349, n1285);
buf  g1276 (n1319, n1213);
not  g1277 (n1340, n1299);
not  g1278 (n1313, n1211);
buf  g1279 (n1350, n1295);
not  g1280 (n1331, n1285);
not  g1281 (n1308, n1287);
not  g1282 (n1336, n1285);
buf  g1283 (n1329, n1290);
buf  g1284 (n1328, n1288);
not  g1285 (n1306, n1212);
buf  g1286 (n1314, n1295);
not  g1287 (n1301, n1121);
not  g1288 (n1317, n1284);
not  g1289 (n1332, n1294);
not  g1290 (n1324, n1293);
not  g1291 (n1339, n1211);
buf  g1292 (n1345, n1290);
buf  g1293 (n1337, n1297);
not  g1294 (n1359, n1287);
not  g1295 (n1344, n1294);
not  g1296 (n1322, n1295);
not  g1297 (n1305, n1283);
buf  g1298 (n1351, n1283);
buf  g1299 (n1342, n1296);
not  g1300 (n1353, n1287);
buf  g1301 (n1318, n1296);
not  g1302 (n1356, n1288);
not  g1303 (n1333, n1285);
buf  g1304 (n1316, n1212);
not  g1305 (n1330, n1296);
not  g1306 (n1323, n1299);
buf  g1307 (n1307, n1214);
buf  g1308 (n1334, n1289);
buf  g1309 (n1325, n1293);
and  g1310 (n1326, n1299, n1298, n1288);
nor  g1311 (n1311, n1297, n1289, n1284);
nor  g1312 (n1320, n1215, n1120, n1293, n1291);
and  g1313 (n1338, n1286, n1291, n1290);
or   g1314 (n1335, n1212, n1283, n1122, n1294);
nor  g1315 (n1358, n1283, n1284, n1213, n1289);
and  g1316 (n1312, n1295, n1298, n1292, n1212);
or   g1317 (n1300, n1297, n1119, n1292);
xor  g1318 (n1303, n1213, n1291, n1289, n1288);
or   g1319 (n1348, n1211, n1290, n1214);
buf  g1320 (n1366, n1305);
buf  g1321 (n1379, n1308);
not  g1322 (n1370, n1307);
not  g1323 (n1369, n1309);
buf  g1324 (n1363, n1300);
buf  g1325 (n1372, n1304);
not  g1326 (n1362, n1313);
not  g1327 (n1377, n1302);
not  g1328 (n1375, n1314);
not  g1329 (n1368, n1319);
not  g1330 (n1371, n1318);
not  g1331 (n1365, n1303);
buf  g1332 (n1361, n1310);
buf  g1333 (n1376, n1317);
buf  g1334 (n1367, n1315);
not  g1335 (n1378, n1306);
not  g1336 (n1360, n1312);
buf  g1337 (n1364, n1301);
not  g1338 (n1373, n1316);
buf  g1339 (n1374, n1311);
buf  g1340 (n1408, n1243);
not  g1341 (n1418, n1257);
buf  g1342 (n1428, n1248);
buf  g1343 (n1425, n1215);
buf  g1344 (n1387, n1255);
not  g1345 (n1415, n1368);
not  g1346 (n1419, n1369);
not  g1347 (n1442, n1379);
not  g1348 (n1396, n1372);
not  g1349 (n1403, n1253);
buf  g1350 (n1447, n1371);
buf  g1351 (n1390, n1377);
not  g1352 (n1431, n1374);
not  g1353 (n1413, n1238);
buf  g1354 (n1407, n1368);
buf  g1355 (n1438, n1258);
buf  g1356 (n1411, n1260);
not  g1357 (n1454, n1365);
not  g1358 (n1426, n1261);
not  g1359 (n1414, n1271);
buf  g1360 (n1436, n1372);
not  g1361 (n1451, n1371);
buf  g1362 (n1433, n1240);
not  g1363 (n1424, n1366);
buf  g1364 (n1391, n1266);
buf  g1365 (n1420, n1369);
buf  g1366 (n1402, n1249);
buf  g1367 (n1455, n1262);
not  g1368 (n1439, n1270);
not  g1369 (n1380, n1264);
not  g1370 (n1430, n1262);
or   g1371 (n1384, n1364, n1251);
nand g1372 (n1457, n1260, n1245, n1370, n1374);
xnor g1373 (n1392, n1367, n1241, n1378, n1216);
xnor g1374 (n1445, n1374, n1245, n38, n1263);
xnor g1375 (n1459, n1253, n1242, n1240, n1269);
nor  g1376 (n1409, n1269, n1255, n1365);
or   g1377 (n1427, n1376, n1362, n1244, n1268);
and  g1378 (n1429, n1258, n1361, n1371, n1379);
and  g1379 (n1452, n37, n1266, n1257, n1375);
xor  g1380 (n1386, n1362, n1363, n1250, n1373);
xor  g1381 (n1444, n1372, n1268, n1244, n1260);
nor  g1382 (n1404, n1369, n1361, n1241, n1370);
nand g1383 (n1458, n1248, n1251, n1216, n1364);
and  g1384 (n1432, n1379, n1378, n1269, n1367);
xor  g1385 (n1388, n1361, n1238, n1263, n1265);
and  g1386 (n1441, n1370, n1270, n1264, n1261);
nand g1387 (n1406, n1360, n1366, n1255, n1249);
xnor g1388 (n1440, n1271, n1245, n1243, n1362);
and  g1389 (n1383, n1375, n1364, n1374, n1271);
nand g1390 (n1456, n1270, n1267, n1363, n1245);
nor  g1391 (n1382, n1253, n1259, n1250, n1264);
nand g1392 (n1412, n1241, n1363, n1378, n1377);
nand g1393 (n1422, n1259, n1247, n1377, n1373);
nand g1394 (n1434, n1251, n38, n1267, n1262);
nand g1395 (n1389, n1246, n1248, n1269, n1368);
nand g1396 (n1400, n1253, n1248, n1379, n1361);
nor  g1397 (n1405, n1262, n1246, n1265, n1368);
or   g1398 (n1453, n1267, n1244, n1360, n1367);
and  g1399 (n1401, n1216, n1256, n1251, n1254);
nor  g1400 (n1437, n1252, n1366, n1265, n1257);
and  g1401 (n1416, n38, n1249, n1242, n1252);
nor  g1402 (n1443, n1243, n1241, n1250, n1215);
nor  g1403 (n1450, n1258, n1242, n1246, n1362);
nand g1404 (n1423, n1216, n1247, n1242, n1377);
or   g1405 (n1410, n1260, n1256, n1378);
and  g1406 (n1381, n1259, n1239, n1365, n1375);
nor  g1407 (n1397, n1270, n1244, n1261, n1243);
xor  g1408 (n1394, n38, n1268, n1370, n1376);
or   g1409 (n1448, n1215, n1258, n1240, n1267);
or   g1410 (n1399, n1239, n1252, n1246);
or   g1411 (n1417, n1254, n1373, n1257, n1250);
or   g1412 (n1385, n1366, n1254, n1264);
xnor g1413 (n1449, n1255, n1239, n1360);
xnor g1414 (n1395, n1263, n1364, n1265, n1363);
nor  g1415 (n1398, n1240, n1268, n1261, n1263);
and  g1416 (n1446, n1376, n1376, n1369, n1247);
and  g1417 (n1421, n1249, n1367, n1266, n1373);
xnor g1418 (n1435, n1360, n1256, n1372, n1259);
nor  g1419 (n1393, n1371, n1247, n1266, n1375);
or   g1420 (n1462, n1387, n1413, n1447, n1431);
nand g1421 (n1463, n174, n1125, n1422, n1402);
xnor g1422 (n1471, n1400, n1380, n1396, n1453);
and  g1423 (n1481, n1448, n175, n1434, n1384);
xor  g1424 (n1467, n1451, n1127, n1425, n1391);
xnor g1425 (n1460, n1389, n174, n1420, n1430);
or   g1426 (n1466, n1459, n1429, n1406, n1446);
nor  g1427 (n1464, n1416, n1437, n1404, n1126);
or   g1428 (n1473, n1458, n1428, n1418, n1442);
nand g1429 (n1483, n1455, n1439, n176, n1454);
or   g1430 (n1475, n1441, n1426, n1397, n1394);
nor  g1431 (n1482, n175, n1452, n1124, n1385);
and  g1432 (n1469, n1438, n1412, n1427, n1392);
xor  g1433 (n1470, n1423, n1386, n1382, n1398);
xor  g1434 (n1465, n1433, n1410, n1393, n1432);
nor  g1435 (n1479, n1415, n1405, n1436, n1390);
and  g1436 (n1472, n1445, n1395, n1409, n1401);
or   g1437 (n1478, n1435, n175, n1388, n1450);
xor  g1438 (n1477, n1414, n1403, n1440, n1130);
nor  g1439 (n1480, n175, n1381, n1123, n174);
nor  g1440 (n1474, n1443, n1417, n1407, n1399);
and  g1441 (n1476, n1457, n1128, n1411, n1456);
xor  g1442 (n1461, n1444, n1129, n1408, n1383);
nor  g1443 (n1468, n1424, n1419, n1421, n1449);
not  g1444 (n1489, n1460);
not  g1445 (n1488, n1462);
buf  g1446 (n1485, n1463);
not  g1447 (n1487, n1467);
not  g1448 (n1491, n1465);
buf  g1449 (n1484, n1464);
buf  g1450 (n1486, n1461);
buf  g1451 (n1490, n1466);
and  g1452 (n1499, n1022, n1137, n1351, n1487);
xor  g1453 (n1520, n1343, n1032, n1323, n1042);
nand g1454 (n1497, n1016, n1320, n1348, n1009);
nand g1455 (n1517, n1485, n1031, n1324, n1133);
and  g1456 (n1495, n1035, n1048, n1484, n1029);
xor  g1457 (n1500, n1008, n1134, n1488, n1346);
xor  g1458 (n1513, n1484, n1036, n1488, n1034);
nand g1459 (n1507, n1025, n1038, n1027, n1056);
nand g1460 (n1501, n1039, n1030, n1028, n1023);
nor  g1461 (n1522, n1331, n1329, n1024, n1486);
xor  g1462 (n1511, n1490, n1043, n1349, n1013);
nand g1463 (n1508, n1340, n1347, n1350, n1490);
xor  g1464 (n1503, n1046, n1138, n1332, n1049);
xnor g1465 (n1521, n1469, n1484, n1033, n1132);
or   g1466 (n1510, n1487, n1055, n1490, n1135);
xor  g1467 (n1523, n1470, n1136, n1342, n1486);
xnor g1468 (n1519, n1019, n1328, n1485, n1344);
xor  g1469 (n1498, n1139, n1327, n1052, n1054);
xnor g1470 (n1516, n1336, n1491, n1489, n1050);
or   g1471 (n1504, n1040, n1321, n1322, n1217);
nor  g1472 (n1506, n1053, n1491, n1485);
xor  g1473 (n1493, n1045, n1487, n1140, n1334);
nor  g1474 (n1496, n1041, n1333, n1489, n1018);
xnor g1475 (n1518, n1012, n1486, n1491, n1341);
xnor g1476 (n1502, n1217, n1011, n1014, n1131);
nand g1477 (n1512, n1047, n1044, n1020, n1488);
or   g1478 (n1509, n1490, n1017, n1488, n1489);
xor  g1479 (n1505, n1345, n1026, n1335, n1010);
or   g1480 (n1515, n1491, n1484, n1021, n1337);
xnor g1481 (n1514, n1015, n1339, n1051, n1487);
xnor g1482 (n1494, n1325, n1037, n1468, n1338);
xor  g1483 (n1492, n1486, n1330, n1489, n1326);
buf  g1484 (n1524, n1492);
buf  g1485 (n1525, n1493);
xor  g1486 (n1526, n1142, n1525, n1143, n1141);
buf  g1487 (n1527, n1217);
xnor g1488 (n1528, n1217, n1526);
buf  g1489 (n1535, n1528);
buf  g1490 (n1529, n1527);
buf  g1491 (n1536, n1058);
buf  g1492 (n1534, n1528);
not  g1493 (n1530, n1527);
buf  g1494 (n1533, n1527);
xor  g1495 (n1532, n1057, n1527);
buf  g1496 (n1531, n1528);
buf  g1497 (n1537, n1146);
buf  g1498 (n1539, n1529);
or   g1499 (n1540, n1147, n1145);
or   g1500 (n1538, n1530, n1530, n1144, n1529);
nor  g1501 (n1541, n1540, n1148);
not  g1502 (n1543, n1541);
nor  g1503 (n1542, n1541, n1218);
not  g1504 (n1544, n1542);
buf  g1505 (n1545, n1150);
buf  g1506 (n1549, n1153);
buf  g1507 (n1547, n1152);
xnor g1508 (n1546, n1542, n1149, n1543, n1151);
nor  g1509 (n1548, n1154, n1543);
not  g1510 (n1557, n1354);
not  g1511 (n1559, n1536);
not  g1512 (n1568, n1531);
not  g1513 (n1567, n1549);
not  g1514 (n1561, n1352);
not  g1515 (n1556, n1534);
xnor g1516 (n1571, n1275, n1532);
xnor g1517 (n1566, n1534, n1536, n1545);
xnor g1518 (n1560, n1532, n1276, n1544);
and  g1519 (n1555, n1273, n1276, n1535, n1546);
nand g1520 (n1554, n1535, n1548, n1533);
nor  g1521 (n1551, n1533, n1534, n1272, n1549);
and  g1522 (n1563, n1534, n1530, n1531);
xor  g1523 (n1558, n1532, n1273, n1548, n1535);
xnor g1524 (n1553, n1533, n1273, n1531, n1218);
xor  g1525 (n1565, n1547, n1273, n1274, n1272);
or   g1526 (n1562, n1272, n1275, n1549, n1530);
xor  g1527 (n1564, n1353, n1547, n1546, n1545);
and  g1528 (n1570, n1544, n1274, n1545, n1549);
and  g1529 (n1572, n1272, n1276, n1274, n1548);
and  g1530 (n1550, n1546, n1536, n1545, n1275);
or   g1531 (n1552, n1275, n1547, n1544, n1274);
nand g1532 (n1573, n1218, n1533, n1544, n1546);
xnor g1533 (n1569, n1271, n1547, n1535, n1532);
not  g1534 (n1588, n1571);
buf  g1535 (n1592, n1564);
not  g1536 (n1593, n1562);
buf  g1537 (n1597, n1553);
not  g1538 (n1596, n1559);
buf  g1539 (n1582, n1554);
buf  g1540 (n1598, n1557);
buf  g1541 (n1594, n1550);
not  g1542 (n1605, n1561);
not  g1543 (n1583, n1568);
not  g1544 (n1578, n1558);
buf  g1545 (n1595, n1572);
not  g1546 (n1584, n1570);
buf  g1547 (n1587, n1565);
not  g1548 (n1579, n1571);
buf  g1549 (n1586, n1563);
not  g1550 (n1603, n1552);
not  g1551 (n1602, n1569);
not  g1552 (n1608, n1555);
buf  g1553 (n1607, n1566);
not  g1554 (n1604, n1551);
not  g1555 (n1590, n1571);
not  g1556 (n1577, n1560);
buf  g1557 (n1600, n1556);
buf  g1558 (n1609, n1570);
buf  g1559 (n1576, n1572);
buf  g1560 (n1581, n1570);
not  g1561 (n1585, n1573);
buf  g1562 (n1575, n1569);
not  g1563 (n1599, n1570);
buf  g1564 (n1591, n1567);
not  g1565 (n1606, n1572);
buf  g1566 (n1574, n1571);
buf  g1567 (n1601, n1572);
buf  g1568 (n1589, n1568);
buf  g1569 (n1580, n1573);
and  g1570 (n1613, n1594, n1574, n1605, n1606);
xor  g1571 (n1615, n1595, n1591, n1597, n1606);
nand g1572 (n1619, n1600, n1586, n1596, n1478);
nor  g1573 (n1621, n1593, n1583, n1576, n1473);
nand g1574 (n1620, n1580, n1604, n1480, n1592);
xor  g1575 (n1614, n1585, n1471, n1606, n1588);
nand g1576 (n1616, n1602, n1578, n1155, n1156);
nand g1577 (n1618, n1606, n1475, n1477, n1598);
and  g1578 (n1617, n1601, n1579, n1603, n1472);
xor  g1579 (n1612, n1575, n1587, n1599, n1476);
xnor g1580 (n1611, n1577, n1479, n1590, n1584);
xor  g1581 (n1610, n1582, n1474, n1589, n1581);
not  g1582 (n1622, n1617);
buf  g1583 (n1627, n1619);
buf  g1584 (n1626, n1620);
buf  g1585 (n1623, n1618);
not  g1586 (n1624, n1483);
xnor g1587 (n1625, n1616, n1482, n1481, n1621);
or   g1588 (n1633, n1498, n1357, n1497, n1521);
nand g1589 (n1641, n1496, n1625, n1626, n1506);
nor  g1590 (n1637, n1626, n1522, n1627, n39);
xor  g1591 (n1631, n1508, n1624, n39, n1503);
xor  g1592 (n1632, n1515, n1509, n1514, n1495);
xor  g1593 (n1638, n1520, n1523, n1519, n1627);
or   g1594 (n1628, n1358, n1505, n176, n1624);
xor  g1595 (n1640, n1626, n1623, n1511, n1507);
nor  g1596 (n1635, n1356, n1500, n1523, n177);
and  g1597 (n1643, n1513, n1359, n1517, n1494);
xor  g1598 (n1636, n176, n1627, n177);
or   g1599 (n1629, n1355, n1625, n1518, n39);
nor  g1600 (n1642, n1512, n176, n39, n1499);
nor  g1601 (n1634, n1622, n1501, n1523, n1625);
xnor g1602 (n1630, n1625, n1502, n1516, n1510);
nand g1603 (n1639, n177, n1504, n1626, n1523);
nor  g1604 (n1644, n177, n1573, n1643);
or   g1605 (n1645, n1644, n1609, n1607);
xnor g1606 (n1647, n1644, n1607, n1608);
or   g1607 (n1646, n1609, n1608, n1607);
and  g1608 (n1648, n1607, n1609, n1644);
nor  g1609 (n1657, n1157, n1184, n1648, n1159);
nand g1610 (n1656, n1158, n1174, n1163, n1173);
nor  g1611 (n1658, n1171, n1168, n1176, n1648);
and  g1612 (n1649, n1175, n1167, n1180, n1169);
or   g1613 (n1652, n1165, n1160, n1646, n1185);
nand g1614 (n1655, n1164, n1183, n1647, n1170);
xor  g1615 (n1653, n1181, n1166, n1647, n1161);
xor  g1616 (n1651, n1179, n1178, n1648, n1177);
or   g1617 (n1650, n1172, n1162, n1186, n1645);
nand g1618 (n1654, n1648, n1182, n1647);
endmodule
