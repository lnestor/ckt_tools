// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_687_1440 written by SynthGen on 2021/05/24 19:48:29
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_687_1440 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18,
 n660, n696, n694, n698, n686, n704, n699, n705,
 n695, n702, n693, n700, n691, n701, n688, n697,
 n687, n689, n692, n703, n690);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18;

output n660, n696, n694, n698, n686, n704, n699, n705,
 n695, n702, n693, n700, n691, n701, n688, n697,
 n687, n689, n692, n703, n690;

wire n19, n20, n21, n22, n23, n24, n25, n26,
 n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n487, n488, n489, n490,
 n491, n492, n493, n494, n495, n496, n497, n498,
 n499, n500, n501, n502, n503, n504, n505, n506,
 n507, n508, n509, n510, n511, n512, n513, n514,
 n515, n516, n517, n518, n519, n520, n521, n522,
 n523, n524, n525, n526, n527, n528, n529, n530,
 n531, n532, n533, n534, n535, n536, n537, n538,
 n539, n540, n541, n542, n543, n544, n545, n546,
 n547, n548, n549, n550, n551, n552, n553, n554,
 n555, n556, n557, n558, n559, n560, n561, n562,
 n563, n564, n565, n566, n567, n568, n569, n570,
 n571, n572, n573, n574, n575, n576, n577, n578,
 n579, n580, n581, n582, n583, n584, n585, n586,
 n587, n588, n589, n590, n591, n592, n593, n594,
 n595, n596, n597, n598, n599, n600, n601, n602,
 n603, n604, n605, n606, n607, n608, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685;

not  g0 (n71, n2);
not  g1 (n68, n15);
buf  g2 (n41, n1);
not  g3 (n73, n10);
buf  g4 (n43, n8);
not  g5 (n21, n3);
buf  g6 (n45, n6);
not  g7 (n26, n4);
not  g8 (n76, n14);
buf  g9 (n59, n7);
buf  g10 (n63, n1);
not  g11 (n72, n15);
not  g12 (n33, n13);
not  g13 (n64, n10);
buf  g14 (n35, n11);
buf  g15 (n52, n7);
not  g16 (n62, n5);
not  g17 (n28, n15);
not  g18 (n32, n8);
buf  g19 (n23, n3);
buf  g20 (n78, n12);
buf  g21 (n44, n6);
buf  g22 (n77, n5);
buf  g23 (n29, n10);
not  g24 (n51, n15);
buf  g25 (n46, n11);
buf  g26 (n67, n4);
buf  g27 (n30, n5);
not  g28 (n27, n14);
buf  g29 (n53, n5);
not  g30 (n20, n12);
not  g31 (n48, n11);
buf  g32 (n56, n7);
buf  g33 (n70, n4);
not  g34 (n75, n11);
not  g35 (n36, n3);
not  g36 (n69, n3);
not  g37 (n55, n12);
buf  g38 (n74, n1);
buf  g39 (n34, n10);
not  g40 (n49, n1);
not  g41 (n50, n13);
not  g42 (n40, n6);
buf  g43 (n58, n14);
not  g44 (n54, n9);
buf  g45 (n37, n9);
not  g46 (n57, n2);
not  g47 (n24, n12);
buf  g48 (n65, n2);
buf  g49 (n39, n14);
not  g50 (n31, n13);
buf  g51 (n60, n13);
not  g52 (n42, n2);
buf  g53 (n19, n9);
not  g54 (n66, n7);
buf  g55 (n61, n4);
not  g56 (n22, n9);
buf  g57 (n38, n8);
not  g58 (n25, n8);
not  g59 (n47, n6);
not  g60 (n126, n27);
buf  g61 (n121, n27);
buf  g62 (n122, n21);
not  g63 (n80, n22);
buf  g64 (n109, n28);
not  g65 (n128, n21);
not  g66 (n86, n24);
buf  g67 (n120, n25);
not  g68 (n84, n28);
buf  g69 (n102, n24);
buf  g70 (n110, n31);
not  g71 (n98, n23);
not  g72 (n115, n22);
not  g73 (n95, n20);
buf  g74 (n101, n26);
buf  g75 (n112, n22);
not  g76 (n124, n25);
buf  g77 (n114, n20);
buf  g78 (n103, n24);
buf  g79 (n85, n19);
not  g80 (n100, n23);
buf  g81 (n106, n25);
not  g82 (n107, n30);
not  g83 (n82, n27);
not  g84 (n90, n24);
buf  g85 (n81, n30);
not  g86 (n108, n29);
not  g87 (n104, n27);
buf  g88 (n117, n29);
not  g89 (n93, n25);
not  g90 (n105, n31);
not  g91 (n89, n28);
not  g92 (n127, n28);
not  g93 (n118, n21);
buf  g94 (n97, n29);
not  g95 (n96, n22);
not  g96 (n116, n20);
buf  g97 (n79, n20);
buf  g98 (n94, n19);
not  g99 (n99, n30);
buf  g100 (n119, n30);
not  g101 (n87, n19);
buf  g102 (n113, n23);
not  g103 (n88, n29);
not  g104 (n83, n19);
not  g105 (n91, n23);
not  g106 (n111, n26);
buf  g107 (n125, n21);
buf  g108 (n92, n26);
buf  g109 (n123, n26);
not  g110 (n315, n52);
buf  g111 (n149, n65);
not  g112 (n220, n98);
not  g113 (n179, n46);
buf  g114 (n163, n37);
not  g115 (n323, n90);
buf  g116 (n296, n126);
buf  g117 (n211, n107);
buf  g118 (n253, n51);
not  g119 (n131, n87);
buf  g120 (n203, n35);
buf  g121 (n311, n66);
buf  g122 (n153, n47);
buf  g123 (n286, n117);
not  g124 (n192, n84);
buf  g125 (n167, n110);
buf  g126 (n200, n114);
not  g127 (n252, n48);
not  g128 (n133, n45);
buf  g129 (n181, n107);
buf  g130 (n235, n43);
not  g131 (n303, n50);
not  g132 (n264, n94);
buf  g133 (n166, n68);
buf  g134 (n258, n35);
buf  g135 (n232, n69);
not  g136 (n278, n39);
not  g137 (n294, n34);
buf  g138 (n213, n101);
buf  g139 (n229, n32);
buf  g140 (n287, n104);
not  g141 (n322, n46);
not  g142 (n187, n88);
buf  g143 (n151, n70);
not  g144 (n234, n16);
not  g145 (n271, n86);
buf  g146 (n280, n71);
buf  g147 (n241, n16);
buf  g148 (n255, n120);
buf  g149 (n282, n49);
buf  g150 (n301, n103);
buf  g151 (n288, n102);
buf  g152 (n221, n113);
buf  g153 (n225, n89);
not  g154 (n162, n90);
buf  g155 (n186, n123);
not  g156 (n257, n73);
not  g157 (n157, n120);
buf  g158 (n169, n61);
not  g159 (n173, n125);
buf  g160 (n297, n37);
buf  g161 (n132, n38);
buf  g162 (n197, n119);
not  g163 (n214, n95);
not  g164 (n134, n76);
not  g165 (n231, n111);
buf  g166 (n292, n81);
buf  g167 (n269, n74);
not  g168 (n175, n87);
not  g169 (n219, n60);
not  g170 (n245, n109);
not  g171 (n277, n49);
not  g172 (n304, n41);
buf  g173 (n272, n127);
buf  g174 (n310, n42);
not  g175 (n250, n46);
buf  g176 (n161, n53);
buf  g177 (n152, n97);
not  g178 (n247, n104);
buf  g179 (n246, n119);
buf  g180 (n140, n84);
buf  g181 (n146, n50);
buf  g182 (n298, n71);
buf  g183 (n218, n17);
buf  g184 (n177, n35);
not  g185 (n198, n17);
not  g186 (n279, n91);
buf  g187 (n222, n44);
not  g188 (n307, n120);
buf  g189 (n138, n71);
not  g190 (n202, n96);
buf  g191 (n160, n96);
not  g192 (n281, n62);
not  g193 (n230, n17);
buf  g194 (n205, n31);
buf  g195 (n312, n95);
not  g196 (n195, n54);
buf  g197 (n191, n106);
not  g198 (n249, n99);
not  g199 (n150, n37);
buf  g200 (n159, n47);
not  g201 (n154, n60);
not  g202 (n236, n111);
not  g203 (n129, n36);
not  g204 (n156, n39);
not  g205 (n299, n55);
not  g206 (n130, n34);
buf  g207 (n283, n36);
not  g208 (n289, n125);
buf  g209 (n243, n108);
buf  g210 (n325, n51);
buf  g211 (n141, n111);
not  g212 (n240, n66);
not  g213 (n256, n40);
not  g214 (n212, n94);
buf  g215 (n204, n53);
buf  g216 (n270, n87);
not  g217 (n237, n113);
not  g218 (n254, n48);
not  g219 (n233, n83);
not  g220 (n188, n105);
not  g221 (n178, n63);
buf  g222 (n275, n80);
buf  g223 (n170, n121);
not  g224 (n300, n74);
not  g225 (n319, n79);
buf  g226 (n135, n124);
buf  g227 (n215, n41);
buf  g228 (n314, n108);
buf  g229 (n242, n72);
buf  g230 (n313, n38);
not  g231 (n321, n111);
not  g232 (n144, n18);
buf  g233 (n308, n44);
not  g234 (n266, n74);
buf  g235 (n185, n115);
buf  g236 (n155, n101);
not  g237 (n305, n118);
buf  g238 (n263, n54);
buf  g239 (n196, n32);
buf  g240 (n244, n96);
buf  g241 (n265, n64);
and  g242 (n317, n43, n55);
xnor g243 (n183, n53, n123, n109, n121);
nor  g244 (n201, n39, n117, n95, n88);
nor  g245 (n293, n128, n60, n118, n103);
and  g246 (n206, n83, n101, n79, n59);
xnor g247 (n268, n102, n52, n73, n97);
nand g248 (n223, n99, n128, n122, n72);
xnor g249 (n228, n114, n116, n124, n47);
nor  g250 (n290, n58, n44, n75, n72);
and  g251 (n309, n58, n68, n98, n75);
or   g252 (n172, n54, n110, n82, n123);
nand g253 (n306, n56, n112, n76, n59);
nand g254 (n262, n106, n98, n113, n89);
nand g255 (n217, n119, n70, n112, n58);
or   g256 (n226, n45, n95, n115, n89);
nand g257 (n143, n70, n100, n122, n18);
nor  g258 (n260, n58, n38, n112, n18);
xnor g259 (n291, n114, n105, n97, n102);
nand g260 (n158, n48, n124, n89);
xor  g261 (n137, n83, n128, n56, n80);
xnor g262 (n174, n81, n81, n127, n103);
and  g263 (n168, n92, n71, n128, n121);
and  g264 (n180, n31, n104, n91, n97);
nor  g265 (n251, n116, n112, n60, n92);
nand g266 (n176, n126, n36, n122, n73);
xnor g267 (n147, n78, n105, n67, n69);
xnor g268 (n238, n52, n107, n91, n57);
and  g269 (n318, n105, n110, n109, n59);
and  g270 (n139, n33, n118, n108, n82);
xnor g271 (n189, n127, n86, n125, n67);
nand g272 (n171, n33, n69, n63, n123);
or   g273 (n284, n56, n42, n57, n119);
or   g274 (n210, n117, n78, n110, n41);
or   g275 (n316, n109, n99, n43, n61);
nand g276 (n142, n43, n117, n93, n90);
or   g277 (n267, n79, n114, n88, n118);
xor  g278 (n302, n44, n108, n82, n78);
and  g279 (n276, n52, n73, n34, n45);
nor  g280 (n320, n93, n54, n49, n76);
nand g281 (n182, n57, n126, n127, n80);
nor  g282 (n224, n80, n40, n67, n61);
or   g283 (n136, n115, n92, n50, n65);
nand g284 (n248, n120, n36, n51, n90);
xnor g285 (n209, n96, n106, n81, n75);
or   g286 (n274, n84, n103, n94, n93);
nor  g287 (n199, n78, n65, n32, n77);
xnor g288 (n273, n18, n113, n40, n62);
or   g289 (n261, n75, n63, n64);
and  g290 (n326, n68, n107, n56, n53);
xor  g291 (n285, n100, n100, n86, n59);
nor  g292 (n165, n98, n99, n76, n74);
and  g293 (n259, n85, n64, n34, n101);
xnor g294 (n193, n122, n38, n116, n40);
nand g295 (n184, n51, n57, n55, n50);
nor  g296 (n194, n79, n82, n16, n126);
and  g297 (n324, n106, n32, n42, n83);
nand g298 (n145, n39, n33, n49, n69);
nand g299 (n295, n77, n87, n65, n41);
and  g300 (n207, n115, n33, n66, n100);
xor  g301 (n328, n72, n116, n92, n66);
or   g302 (n208, n46, n88, n64, n93);
xor  g303 (n190, n62, n125, n121, n86);
nor  g304 (n164, n48, n70, n62, n84);
and  g305 (n327, n91, n37, n68, n17);
xnor g306 (n216, n35, n85, n55, n42);
xnor g307 (n239, n94, n47, n45, n102);
or   g308 (n148, n77, n16, n85);
nand g309 (n227, n61, n67, n77, n104);
not  g310 (n331, n132);
not  g311 (n340, n130);
not  g312 (n330, n138);
buf  g313 (n339, n140);
buf  g314 (n333, n131);
not  g315 (n336, n129);
not  g316 (n332, n135);
not  g317 (n337, n139);
not  g318 (n335, n134);
not  g319 (n329, n136);
buf  g320 (n338, n137);
buf  g321 (n334, n133);
xor  g322 (n352, n172, n335, n161, n145);
nor  g323 (n355, n162, n329, n175, n169);
and  g324 (n347, n175, n174, n166, n331);
nor  g325 (n356, n144, n165, n172, n335);
nand g326 (n349, n157, n329, n149, n175);
and  g327 (n351, n154, n164, n174, n332);
and  g328 (n341, n169, n160, n155, n151);
and  g329 (n346, n174, n337, n172, n153);
nor  g330 (n353, n170, n173, n330, n333);
nor  g331 (n348, n332, n152, n167, n142);
and  g332 (n345, n156, n158, n336, n159);
nor  g333 (n350, n163, n146, n143, n334);
xor  g334 (n357, n171, n168, n148);
xnor g335 (n354, n170, n336, n172, n330);
or   g336 (n342, n334, n147, n171, n173);
nor  g337 (n343, n333, n141, n173, n150);
or   g338 (n344, n174, n173, n175, n331);
nand g339 (n375, n346, n186, n344, n196);
and  g340 (n382, n201, n184, n189, n177);
xor  g341 (n365, n197, n344, n187);
nand g342 (n366, n191, n349, n183, n195);
nand g343 (n376, n184, n201, n198, n200);
xnor g344 (n384, n189, n346, n181, n342);
nor  g345 (n391, n176, n348, n196, n184);
or   g346 (n358, n200, n179, n348);
nor  g347 (n385, n180, n180, n185, n199);
or   g348 (n364, n186, n192, n199, n188);
and  g349 (n371, n342, n197, n183, n345);
nor  g350 (n392, n183, n184, n195, n343);
or   g351 (n389, n341, n191, n343, n186);
nor  g352 (n360, n194, n349, n176, n193);
xor  g353 (n387, n341, n198, n191, n345);
xor  g354 (n381, n177, n187, n199);
or   g355 (n377, n178, n196, n189, n180);
xnor g356 (n372, n342, n347, n344);
and  g357 (n390, n177, n201, n190, n176);
xor  g358 (n383, n182, n198, n178, n343);
and  g359 (n368, n182, n194, n185, n345);
nand g360 (n361, n200, n190, n180, n185);
xor  g361 (n362, n346, n345, n344, n194);
xor  g362 (n359, n192, n200, n181);
xnor g363 (n367, n202, n183, n193, n177);
nand g364 (n370, n188, n342, n348, n185);
xor  g365 (n373, n197, n193);
nor  g366 (n374, n199, n194, n181, n176);
xor  g367 (n378, n186, n201, n349, n188);
xor  g368 (n386, n178, n341, n190, n195);
nand g369 (n379, n196, n343, n190, n195);
nand g370 (n369, n191, n192, n198, n188);
xor  g371 (n388, n178, n182, n347, n341);
xor  g372 (n380, n346, n192, n179, n348);
nand g373 (n363, n179, n182, n189, n347);
and  g374 (n429, n233, n210, n204, n236);
and  g375 (n399, n225, n205, n354);
xor  g376 (n411, n232, n236, n350, n235);
and  g377 (n421, n368, n211, n218, n228);
xor  g378 (n431, n241, n236, n207, n223);
xnor g379 (n410, n362, n211, n363, n219);
nand g380 (n393, n206, n240, n237, n239);
xnor g381 (n447, n203, n353, n242, n372);
or   g382 (n446, n209, n355, n238, n212);
and  g383 (n435, n213, n216, n352, n223);
and  g384 (n432, n230, n390, n224, n229);
and  g385 (n436, n237, n235, n208, n366);
or   g386 (n424, n376, n374, n240, n375);
nand g387 (n430, n210, n218, n212, n216);
xnor g388 (n404, n227, n350, n354, n228);
xor  g389 (n449, n364, n386, n219, n237);
and  g390 (n402, n243, n383, n222, n205);
xnor g391 (n456, n206, n229, n349, n204);
or   g392 (n438, n232, n383, n214, n213);
or   g393 (n420, n377, n212, n232, n373);
xnor g394 (n427, n354, n365, n207, n211);
nor  g395 (n414, n352, n242, n211, n369);
and  g396 (n397, n226, n234, n351, n222);
and  g397 (n451, n374, n226, n236, n230);
or   g398 (n422, n379, n352, n351, n227);
nor  g399 (n417, n240, n213, n203, n367);
xor  g400 (n407, n206, n205, n224, n212);
and  g401 (n398, n217, n226, n209, n204);
xor  g402 (n418, n225, n241, n219, n234);
xor  g403 (n439, n234, n238, n215, n242);
and  g404 (n415, n218, n372, n352, n240);
xnor g405 (n433, n215, n351, n387, n370);
nand g406 (n395, n392, n220, n359, n382);
or   g407 (n400, n234, n354, n203, n353);
nand g408 (n413, n221, n239, n218, n237);
xnor g409 (n406, n385, n350, n231, n235);
nand g410 (n448, n384, n214, n238, n228);
or   g411 (n441, n233, n221, n215);
xor  g412 (n425, n381, n207, n227, n391);
and  g413 (n416, n221, n239, n220, n360);
nand g414 (n419, n209, n382, n368, n230);
nor  g415 (n396, n216, n208, n377, n206);
and  g416 (n394, n369, n207, n209, n223);
nand g417 (n445, n231, n210, n239, n356);
nand g418 (n454, n353, n227, n225, n364);
nor  g419 (n401, n214, n365, n243, n389);
nor  g420 (n440, n229, n231, n355, n366);
and  g421 (n409, n356, n380, n386, n217);
nor  g422 (n452, n367, n204, n213, n216);
or   g423 (n403, n242, n203, n378, n224);
nand g424 (n437, n230, n241, n385, n210);
nor  g425 (n443, n355, n231, n225, n202);
or   g426 (n426, n370, n351, n379, n217);
nand g427 (n453, n228, n391, n388, n350);
xor  g428 (n412, n355, n233, n371, n375);
xnor g429 (n455, n381, n238, n389, n380);
nor  g430 (n444, n384, n232, n373, n388);
nand g431 (n423, n353, n208, n361, n235);
nand g432 (n442, n220, n226, n222, n241);
xor  g433 (n434, n222, n215, n390, n224);
and  g434 (n405, n214, n229, n202, n376);
xor  g435 (n450, n387, n233, n223, n219);
nand g436 (n428, n378, n392, n358, n208);
xor  g437 (n408, n202, n217, n371, n220);
not  g438 (n457, n393);
buf  g439 (n459, n244);
xor  g440 (n458, n244, n393);
or   g441 (n460, n393, n243);
xnor g442 (n475, n458, n402, n394, n398);
xor  g443 (n464, n402, n457, n244, n396);
and  g444 (n476, n399, n400, n460, n459);
xnor g445 (n469, n395, n459, n400);
xor  g446 (n463, n397, n398, n246);
or   g447 (n474, n396, n245, n246);
xor  g448 (n472, n397, n395, n458, n457);
xnor g449 (n467, n245, n247, n398, n399);
or   g450 (n468, n395, n402, n401, n458);
and  g451 (n466, n458, n394, n399, n401);
nand g452 (n473, n394, n244, n245, n247);
and  g453 (n465, n246, n459, n400, n399);
nand g454 (n461, n460, n457, n401, n395);
and  g455 (n470, n397, n460, n457, n394);
xnor g456 (n462, n396, n459, n398, n397);
nor  g457 (n471, n402, n401, n460, n396);
or   g458 (n484, n417, n461, n419, n471);
xor  g459 (n507, n411, n252, n423, n471);
nand g460 (n521, n425, n424, n472, n429);
xor  g461 (n527, n415, n472, n419, n255);
and  g462 (n525, n405, n475, n407, n251);
xnor g463 (n489, n254, n251, n337, n357);
and  g464 (n498, n474, n461, n417, n432);
nor  g465 (n535, n407, n416, n423, n418);
xor  g466 (n481, n429, n253, n468, n413);
nor  g467 (n485, n432, n408, n411, n256);
xor  g468 (n494, n464, n253, n433, n421);
and  g469 (n524, n423, n249, n253, n465);
and  g470 (n522, n256, n465, n469, n420);
nand g471 (n488, n407, n249, n252, n419);
nor  g472 (n534, n428, n474, n422, n466);
nand g473 (n490, n421, n430, n427, n473);
xor  g474 (n486, n412, n247, n462, n248);
or   g475 (n529, n255, n411, n413, n415);
nand g476 (n523, n409, n249, n467, n356);
or   g477 (n508, n422, n471, n249, n252);
nor  g478 (n510, n467, n339, n461, n429);
nor  g479 (n491, n338, n417, n426, n432);
or   g480 (n487, n357, n405, n426, n416);
xnor g481 (n482, n416, n431, n420, n408);
and  g482 (n477, n431, n409, n407, n404);
or   g483 (n518, n412, n433, n248, n414);
xor  g484 (n506, n431, n428, n463, n414);
xor  g485 (n499, n339, n357, n426, n412);
and  g486 (n517, n470, n250, n464, n254);
nor  g487 (n532, n468, n464, n417, n467);
and  g488 (n509, n466, n473, n250, n424);
nand g489 (n520, n422, n404, n425, n250);
or   g490 (n512, n405, n254, n465, n340);
or   g491 (n504, n423, n410, n474, n430);
nand g492 (n503, n252, n470, n422, n404);
nand g493 (n493, n413, n251, n404, n339);
and  g494 (n500, n462, n425, n428, n433);
xnor g495 (n492, n405, n414, n357, n465);
nor  g496 (n526, n428, n468, n403, n248);
or   g497 (n497, n464, n412, n247, n427);
and  g498 (n530, n418, n408, n340, n420);
xor  g499 (n515, n416, n466, n472, n255);
xnor g500 (n511, n429, n410, n473, n415);
nor  g501 (n501, n420, n475, n253, n421);
nor  g502 (n483, n410, n424, n425, n469);
nor  g503 (n480, n255, n406, n426, n431);
xor  g504 (n496, n462, n427, n474, n418);
nand g505 (n502, n472, n403, n406, n463);
nor  g506 (n513, n256, n410, n409, n254);
nor  g507 (n531, n470, n432, n403, n463);
or   g508 (n495, n248, n469, n411, n418);
xnor g509 (n528, n427, n406, n466);
xor  g510 (n478, n251, n433, n408, n338);
nor  g511 (n479, n461, n256, n424, n421);
xor  g512 (n505, n339, n356, n409, n413);
nor  g513 (n516, n470, n473, n430);
nand g514 (n514, n467, n403, n475, n419);
nor  g515 (n533, n415, n414, n250, n469);
and  g516 (n519, n463, n468, n462, n471);
xnor g517 (n626, n308, n321, n326, n318);
or   g518 (n594, n309, n270, n285, n326);
nand g519 (n627, n273, n300, n260, n272);
xnor g520 (n570, n312, n526, n279, n289);
and  g521 (n576, n531, n313, n269, n267);
or   g522 (n610, n286, n526, n499, n314);
nor  g523 (n631, n535, n317, n257, n314);
and  g524 (n538, n259, n280, n264, n283);
nand g525 (n581, n311, n265, n320, n281);
xor  g526 (n551, n526, n510, n305, n261);
xnor g527 (n608, n504, n267, n270, n525);
and  g528 (n539, n294, n313, n259, n501);
xor  g529 (n628, n263, n296, n322, n518);
xnor g530 (n564, n306, n528, n481, n305);
nand g531 (n543, n479, n317, n527, n295);
and  g532 (n625, n325, n320, n273, n291);
nand g533 (n550, n494, n529, n298, n286);
nor  g534 (n566, n276, n274, n523);
xnor g535 (n582, n306, n315, n507, n262);
and  g536 (n567, n261, n258, n516, n299);
xor  g537 (n606, n290, n505, n281, n316);
nand g538 (n609, n297, n305, n277, n274);
xnor g539 (n549, n266, n312, n315, n327);
nand g540 (n548, n324, n280, n292, n511);
xnor g541 (n630, n490, n301, n283, n296);
xnor g542 (n569, n284, n298, n485, n274);
xnor g543 (n590, n302, n325, n491, n508);
nand g544 (n547, n517, n326, n294, n291);
or   g545 (n574, n328, n488, n300, n258);
xnor g546 (n591, n279, n324, n320, n274);
nor  g547 (n589, n286, n278, n275, n291);
nand g548 (n577, n519, n306, n257, n293);
nor  g549 (n618, n275, n312, n531, n326);
and  g550 (n612, n321, n279, n317, n318);
xor  g551 (n586, n311, n281, n265, n324);
xnor g552 (n613, n288, n268, n531, n271);
or   g553 (n554, n500, n272, n284, n300);
or   g554 (n583, n328, n514, n529, n307);
and  g555 (n558, n520, n280, n524, n302);
nor  g556 (n565, n268, n308, n259, n293);
nand g557 (n545, n273, n275, n503, n282);
or   g558 (n603, n281, n309, n282, n528);
nand g559 (n593, n295, n272, n527, n484);
and  g560 (n573, n287, n306, n309, n323);
nand g561 (n561, n257, n284, n304, n289);
and  g562 (n621, n261, n278, n319, n285);
or   g563 (n588, n515, n299, n292, n316);
and  g564 (n542, n319, n323, n305, n269);
or   g565 (n596, n299, n497, n268, n328);
nor  g566 (n553, n272, n322, n276, n267);
xnor g567 (n552, n284, n301, n310, n277);
and  g568 (n602, n486, n294, n512, n527);
and  g569 (n604, n327, n276, n263, n311);
and  g570 (n623, n532, n533, n320, n283);
nand g571 (n629, n492, n321, n266, n264);
xor  g572 (n568, n482, n534, n297, n314);
and  g573 (n599, n312, n299, n288, n270);
xnor g574 (n597, n295, n322, n483, n524);
or   g575 (n617, n304, n315, n327, n289);
xor  g576 (n601, n285, n509, n524, n325);
nand g577 (n544, n308, n496, n521, n477);
nand g578 (n556, n265, n480, n313, n288);
xor  g579 (n616, n297, n262, n266, n528);
xnor g580 (n571, n260, n273, n294, n293);
or   g581 (n615, n535, n493, n303);
or   g582 (n611, n534, n530, n277, n292);
xor  g583 (n600, n321, n263, n259, n502);
or   g584 (n614, n291, n533, n287, n532);
nor  g585 (n585, n530, n275, n271, n513);
xor  g586 (n584, n525, n260, n530, n304);
or   g587 (n537, n263, n495, n307, n527);
nor  g588 (n592, n278, n269, n528, n271);
and  g589 (n540, n533, n290, n303, n277);
and  g590 (n559, n266, n296, n292, n307);
and  g591 (n580, n260, n287, n319, n262);
nand g592 (n536, n295, n535, n301, n533);
and  g593 (n624, n310, n532, n322, n293);
nor  g594 (n605, n268, n309, n258, n323);
xnor g595 (n557, n289, n279, n317, n302);
xnor g596 (n560, n308, n524, n298, n283);
xor  g597 (n555, n314, n531, n325, n526);
and  g598 (n563, n311, n328, n257, n304);
xnor g599 (n598, n535, n261, n318, n310);
nand g600 (n578, n282, n506, n276, n258);
nor  g601 (n622, n287, n286, n302, n324);
nand g602 (n619, n534, n290, n282, n318);
xor  g603 (n572, n522, n323, n525, n489);
xor  g604 (n607, n300, n265, n290, n303);
xnor g605 (n595, n280, n262, n316, n296);
xnor g606 (n620, n278, n316, n264, n285);
or   g607 (n579, n297, n271, n529, n525);
xor  g608 (n541, n530, n267, n532, n327);
nor  g609 (n546, n487, n307, n534, n310);
xor  g610 (n587, n478, n529, n264, n288);
and  g611 (n562, n313, n269, n298, n319);
nand g612 (n575, n315, n270, n301, n498);
nand g613 (n635, n562, n441, n442);
or   g614 (n653, n449, n561, n438, n559);
xnor g615 (n641, n536, n447, n455, n448);
and  g616 (n648, n434, n435, n456, n453);
xnor g617 (n642, n454, n450, n436, n446);
nor  g618 (n659, n439, n548, n543, n447);
nor  g619 (n647, n451, n443, n554, n452);
xnor g620 (n663, n555, n434, n446, n449);
xor  g621 (n639, n454, n558, n438, n537);
nor  g622 (n652, n435, n541, n440, n448);
and  g623 (n651, n449, n453, n437, n564);
or   g624 (n649, n456, n549, n538, n441);
and  g625 (n632, n445, n455, n438, n435);
or   g626 (n658, n452, n444, n539, n434);
nor  g627 (n637, n439, n442, n340, n552);
xnor g628 (n644, n447, n456, n448, n557);
nor  g629 (n640, n434, n446, n542, n476);
xnor g630 (n662, n455, n455, n565, n441);
or   g631 (n636, n566, n440, n476, n444);
nand g632 (n657, n441, n437, n452);
xor  g633 (n645, n560, n449, n439, n568);
xor  g634 (n643, n445, n547, n544, n553);
xor  g635 (n646, n435, n563, n451, n551);
and  g636 (n656, n445, n436, n437, n444);
or   g637 (n660, n456, n453, n447, n444);
and  g638 (n634, n451, n439, n450, n545);
xnor g639 (n664, n450, n445, n476, n443);
nor  g640 (n654, n438, n454, n550, n475);
nor  g641 (n650, n436, n442, n443, n440);
xnor g642 (n638, n540, n476, n453, n446);
nand g643 (n661, n450, n546, n451, n448);
or   g644 (n655, n567, n437, n436, n454);
xor  g645 (n633, n440, n340, n556, n443);
nor  g646 (n673, n649, n604, n599, n622);
xnor g647 (n678, n603, n614, n612, n628);
and  g648 (n667, n575, n592, n647, n636);
or   g649 (n684, n579, n572, n648, n610);
xnor g650 (n677, n620, n598, n606, n645);
nand g651 (n675, n624, n619, n613, n648);
and  g652 (n674, n641, n638, n630, n581);
and  g653 (n672, n618, n632, n626, n609);
nor  g654 (n671, n586, n621, n635, n596);
xnor g655 (n676, n607, n577, n580, n616);
xor  g656 (n685, n649, n644, n576, n639);
xor  g657 (n669, n569, n608, n578, n588);
xnor g658 (n668, n573, n602, n590, n623);
or   g659 (n666, n595, n633, n593, n584);
and  g660 (n680, n642, n570, n571, n617);
nand g661 (n682, n625, n594, n600, n587);
and  g662 (n681, n582, n574, n627, n650);
or   g663 (n683, n591, n643, n629, n601);
xnor g664 (n679, n583, n646, n611, n634);
and  g665 (n665, n631, n597, n585, n637);
or   g666 (n670, n589, n640, n605, n615);
nor  g667 (n695, n663, n653, n651, n684);
nor  g668 (n693, n680, n653, n662, n655);
xnor g669 (n687, n653, n650, n661, n685);
or   g670 (n698, n659, n651, n658, n682);
xor  g671 (n686, n652, n681, n675, n669);
and  g672 (n704, n656, n653, n662);
xor  g673 (n703, n663, n673, n655);
nor  g674 (n692, n651, n650, n658, n663);
xnor g675 (n699, n679, n664, n665, n656);
nor  g676 (n691, n677, n671, n652, n661);
and  g677 (n694, n656, n654, n664, n659);
xnor g678 (n701, n660, n672, n661, n656);
nor  g679 (n696, n658, n676, n655, n662);
xor  g680 (n688, n660, n663, n652, n654);
nor  g681 (n697, n654, n657, n664, n658);
or   g682 (n702, n667, n650, n674, n683);
xnor g683 (n700, n659, n657);
or   g684 (n689, n661, n651, n659, n652);
and  g685 (n705, n678, n660, n654);
xnor g686 (n690, n670, n666, n664, n668);
endmodule
