

module Stat_976_2713
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n968,
  n970,
  n975,
  n972,
  n986,
  n967,
  n980,
  n978,
  n966,
  n984,
  n985,
  n981,
  n974,
  n983,
  n976,
  n979,
  n969,
  n989,
  n971,
  n982,
  n988,
  n977,
  n991,
  n1001,
  n999,
  n1000,
  n1002,
  n998,
  n1003,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n968;
  output n970;
  output n975;
  output n972;
  output n986;
  output n967;
  output n980;
  output n978;
  output n966;
  output n984;
  output n985;
  output n981;
  output n974;
  output n983;
  output n976;
  output n979;
  output n969;
  output n989;
  output n971;
  output n982;
  output n988;
  output n977;
  output n991;
  output n1001;
  output n999;
  output n1000;
  output n1002;
  output n998;
  output n1003;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n973;
  wire n987;
  wire n990;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n42,
    n17
  );


  buf
  g1
  (
    n77,
    n13
  );


  buf
  g2
  (
    n53,
    n5
  );


  not
  g3
  (
    n37,
    n14
  );


  buf
  g4
  (
    n78,
    n9
  );


  not
  g5
  (
    n32,
    n13
  );


  not
  g6
  (
    n36,
    n9
  );


  buf
  g7
  (
    n55,
    n4
  );


  not
  g8
  (
    n79,
    n14
  );


  buf
  g9
  (
    n63,
    n7
  );


  not
  g10
  (
    n28,
    n7
  );


  not
  g11
  (
    n34,
    n17
  );


  not
  g12
  (
    n40,
    n10
  );


  buf
  g13
  (
    n31,
    n4
  );


  buf
  g14
  (
    n64,
    n12
  );


  not
  g15
  (
    n71,
    n12
  );


  not
  g16
  (
    n82,
    n12
  );


  not
  g17
  (
    n62,
    n11
  );


  buf
  g18
  (
    n66,
    n8
  );


  buf
  g19
  (
    n59,
    n18
  );


  not
  g20
  (
    n72,
    n14
  );


  not
  g21
  (
    n45,
    n3
  );


  not
  g22
  (
    n81,
    n11
  );


  not
  g23
  (
    n51,
    n12
  );


  not
  g24
  (
    n30,
    n13
  );


  buf
  g25
  (
    n33,
    n16
  );


  not
  g26
  (
    KeyWire_0_54,
    n10
  );


  not
  g27
  (
    n56,
    n2
  );


  not
  g28
  (
    n44,
    n19
  );


  buf
  g29
  (
    n69,
    n13
  );


  buf
  g30
  (
    n80,
    n18
  );


  not
  g31
  (
    n43,
    n19
  );


  buf
  g32
  (
    n41,
    n16
  );


  buf
  g33
  (
    n60,
    n6
  );


  buf
  g34
  (
    KeyWire_0_7,
    n15
  );


  not
  g35
  (
    n52,
    n3
  );


  not
  g36
  (
    n73,
    n1
  );


  not
  g37
  (
    n54,
    n8
  );


  not
  g38
  (
    n39,
    n17
  );


  not
  g39
  (
    n68,
    n5
  );


  not
  g40
  (
    n35,
    n16
  );


  buf
  g41
  (
    n29,
    n2
  );


  buf
  g42
  (
    n47,
    n11
  );


  not
  g43
  (
    n46,
    n10
  );


  not
  g44
  (
    n75,
    n15
  );


  buf
  g45
  (
    n65,
    n11
  );


  buf
  g46
  (
    n76,
    n18
  );


  buf
  g47
  (
    n70,
    n16
  );


  buf
  g48
  (
    n38,
    n14
  );


  not
  g49
  (
    n57,
    n18
  );


  buf
  g50
  (
    n50,
    n1
  );


  not
  g51
  (
    n61,
    n15
  );


  not
  g52
  (
    n49,
    n6
  );


  not
  g53
  (
    n74,
    n17
  );


  not
  g54
  (
    n83,
    n10
  );


  buf
  g55
  (
    n58,
    n15
  );


  buf
  g56
  (
    n165,
    n54
  );


  buf
  g57
  (
    n116,
    n48
  );


  not
  g58
  (
    n146,
    n51
  );


  buf
  g59
  (
    n163,
    n31
  );


  buf
  g60
  (
    n90,
    n29
  );


  buf
  g61
  (
    n153,
    n39
  );


  buf
  g62
  (
    n157,
    n47
  );


  buf
  g63
  (
    n161,
    n54
  );


  not
  g64
  (
    n105,
    n30
  );


  not
  g65
  (
    n143,
    n65
  );


  not
  g66
  (
    n117,
    n49
  );


  not
  g67
  (
    n131,
    n34
  );


  not
  g68
  (
    n127,
    n62
  );


  not
  g69
  (
    n132,
    n45
  );


  not
  g70
  (
    n122,
    n28
  );


  buf
  g71
  (
    n98,
    n28
  );


  buf
  g72
  (
    KeyWire_0_46,
    n37
  );


  buf
  g73
  (
    n151,
    n61
  );


  buf
  g74
  (
    n104,
    n68
  );


  buf
  g75
  (
    KeyWire_0_21,
    n46
  );


  buf
  g76
  (
    n112,
    n40
  );


  not
  g77
  (
    KeyWire_0_52,
    n50
  );


  buf
  g78
  (
    n110,
    n39
  );


  not
  g79
  (
    n92,
    n32
  );


  buf
  g80
  (
    n152,
    n43
  );


  buf
  g81
  (
    n135,
    n41
  );


  buf
  g82
  (
    n111,
    n33
  );


  buf
  g83
  (
    n102,
    n36
  );


  not
  g84
  (
    KeyWire_0_39,
    n48
  );


  not
  g85
  (
    n148,
    n49
  );


  not
  g86
  (
    n149,
    n37
  );


  not
  g87
  (
    n89,
    n56
  );


  buf
  g88
  (
    n100,
    n61
  );


  not
  g89
  (
    n106,
    n44
  );


  not
  g90
  (
    n164,
    n56
  );


  not
  g91
  (
    n147,
    n67
  );


  buf
  g92
  (
    n138,
    n58
  );


  buf
  g93
  (
    n109,
    n57
  );


  buf
  g94
  (
    n126,
    n57
  );


  buf
  g95
  (
    n97,
    n32
  );


  not
  g96
  (
    n136,
    n46
  );


  not
  g97
  (
    n154,
    n30
  );


  buf
  g98
  (
    n124,
    n58
  );


  not
  g99
  (
    n119,
    n50
  );


  buf
  g100
  (
    n128,
    n38
  );


  not
  g101
  (
    n120,
    n45
  );


  not
  g102
  (
    n145,
    n52
  );


  not
  g103
  (
    n107,
    n38
  );


  buf
  g104
  (
    n166,
    n62
  );


  not
  g105
  (
    n142,
    n51
  );


  not
  g106
  (
    n144,
    n42
  );


  not
  g107
  (
    n88,
    n47
  );


  buf
  g108
  (
    n101,
    n53
  );


  not
  g109
  (
    n113,
    n33
  );


  not
  g110
  (
    n133,
    n67
  );


  buf
  g111
  (
    n159,
    n66
  );


  buf
  g112
  (
    n94,
    n53
  );


  buf
  g113
  (
    n118,
    n60
  );


  buf
  g114
  (
    n91,
    n63
  );


  not
  g115
  (
    n125,
    n63
  );


  buf
  g116
  (
    n150,
    n55
  );


  buf
  g117
  (
    n129,
    n64
  );


  buf
  g118
  (
    n86,
    n41
  );


  not
  g119
  (
    n121,
    n65
  );


  buf
  g120
  (
    n160,
    n60
  );


  buf
  g121
  (
    n84,
    n44
  );


  not
  g122
  (
    n96,
    n42
  );


  not
  g123
  (
    n85,
    n35
  );


  buf
  g124
  (
    n162,
    n34
  );


  buf
  g125
  (
    n115,
    n59
  );


  buf
  g126
  (
    n99,
    n31
  );


  not
  g127
  (
    n95,
    n64
  );


  buf
  g128
  (
    n103,
    n36
  );


  buf
  g129
  (
    n156,
    n35
  );


  buf
  g130
  (
    n93,
    n68
  );


  buf
  g131
  (
    n139,
    n55
  );


  not
  g132
  (
    n155,
    n43
  );


  not
  g133
  (
    n123,
    n52
  );


  not
  g134
  (
    n158,
    n29
  );


  buf
  g135
  (
    n137,
    n66
  );


  not
  g136
  (
    n114,
    n40
  );


  buf
  g137
  (
    n141,
    n69
  );


  not
  g138
  (
    n87,
    n59
  );


  not
  g139
  (
    n226,
    n98
  );


  not
  g140
  (
    n237,
    n138
  );


  buf
  g141
  (
    n173,
    n161
  );


  not
  g142
  (
    n280,
    n127
  );


  buf
  g143
  (
    n246,
    n150
  );


  buf
  g144
  (
    n261,
    n144
  );


  buf
  g145
  (
    n214,
    n87
  );


  buf
  g146
  (
    n180,
    n120
  );


  not
  g147
  (
    n232,
    n155
  );


  not
  g148
  (
    n221,
    n140
  );


  not
  g149
  (
    n259,
    n114
  );


  not
  g150
  (
    n279,
    n99
  );


  not
  g151
  (
    n270,
    n143
  );


  not
  g152
  (
    n168,
    n90
  );


  buf
  g153
  (
    n216,
    n111
  );


  not
  g154
  (
    n217,
    n155
  );


  not
  g155
  (
    KeyWire_0_22,
    n147
  );


  not
  g156
  (
    n231,
    n138
  );


  buf
  g157
  (
    n182,
    n106
  );


  not
  g158
  (
    n169,
    n117
  );


  buf
  g159
  (
    n178,
    n151
  );


  not
  g160
  (
    n273,
    n131
  );


  buf
  g161
  (
    n204,
    n104
  );


  buf
  g162
  (
    n252,
    n133
  );


  buf
  g163
  (
    n256,
    n156
  );


  not
  g164
  (
    n170,
    n136
  );


  buf
  g165
  (
    n268,
    n153
  );


  buf
  g166
  (
    n251,
    n159
  );


  not
  g167
  (
    n236,
    n140
  );


  not
  g168
  (
    n206,
    n154
  );


  buf
  g169
  (
    n271,
    n148
  );


  buf
  g170
  (
    n265,
    n159
  );


  not
  g171
  (
    n275,
    n108
  );


  not
  g172
  (
    n201,
    n84
  );


  not
  g173
  (
    n192,
    n137
  );


  buf
  g174
  (
    n185,
    n88
  );


  not
  g175
  (
    n183,
    n96
  );


  not
  g176
  (
    n200,
    n93
  );


  not
  g177
  (
    n278,
    n103
  );


  not
  g178
  (
    n228,
    n110
  );


  not
  g179
  (
    n195,
    n142
  );


  not
  g180
  (
    n172,
    n148
  );


  not
  g181
  (
    n171,
    n163
  );


  buf
  g182
  (
    n235,
    n121
  );


  not
  g183
  (
    n197,
    n145
  );


  not
  g184
  (
    n238,
    n131
  );


  buf
  g185
  (
    n230,
    n154
  );


  buf
  g186
  (
    n225,
    n136
  );


  buf
  g187
  (
    n167,
    n134
  );


  not
  g188
  (
    n220,
    n129
  );


  buf
  g189
  (
    n277,
    n153
  );


  not
  g190
  (
    n208,
    n132
  );


  not
  g191
  (
    n244,
    n124
  );


  not
  g192
  (
    n202,
    n123
  );


  buf
  g193
  (
    n209,
    n145
  );


  not
  g194
  (
    n219,
    n139
  );


  buf
  g195
  (
    n207,
    n146
  );


  buf
  g196
  (
    KeyWire_0_47,
    n113
  );


  not
  g197
  (
    n260,
    n132
  );


  buf
  g198
  (
    n198,
    n150
  );


  not
  g199
  (
    n240,
    n101
  );


  not
  g200
  (
    n239,
    n107
  );


  buf
  g201
  (
    n247,
    n149
  );


  buf
  g202
  (
    n186,
    n160
  );


  buf
  g203
  (
    n262,
    n133
  );


  not
  g204
  (
    n263,
    n102
  );


  buf
  g205
  (
    n176,
    n141
  );


  not
  g206
  (
    n223,
    n152
  );


  not
  g207
  (
    n210,
    n92
  );


  not
  g208
  (
    n233,
    n128
  );


  buf
  g209
  (
    n184,
    n105
  );


  buf
  g210
  (
    n264,
    n85
  );


  not
  g211
  (
    n224,
    n157
  );


  buf
  g212
  (
    n242,
    n86
  );


  buf
  g213
  (
    n199,
    n162
  );


  buf
  g214
  (
    n211,
    n112
  );


  not
  g215
  (
    n253,
    n95
  );


  buf
  g216
  (
    n248,
    n158
  );


  buf
  g217
  (
    n258,
    n118
  );


  buf
  g218
  (
    n193,
    n100
  );


  not
  g219
  (
    n241,
    n139
  );


  buf
  g220
  (
    n205,
    n89
  );


  not
  g221
  (
    KeyWire_0_42,
    n97
  );


  not
  g222
  (
    n203,
    n147
  );


  buf
  g223
  (
    n255,
    n160
  );


  not
  g224
  (
    n257,
    n134
  );


  buf
  g225
  (
    n249,
    n149
  );


  buf
  g226
  (
    n250,
    n161
  );


  buf
  g227
  (
    n196,
    n130
  );


  buf
  g228
  (
    n269,
    n157
  );


  not
  g229
  (
    n266,
    n162
  );


  not
  g230
  (
    n272,
    n91
  );


  buf
  g231
  (
    KeyWire_0_59,
    n125
  );


  not
  g232
  (
    n175,
    n156
  );


  not
  g233
  (
    n229,
    n116
  );


  buf
  g234
  (
    n274,
    n122
  );


  not
  g235
  (
    n189,
    n152
  );


  buf
  g236
  (
    n190,
    n135
  );


  buf
  g237
  (
    KeyWire_0_40,
    n144
  );


  not
  g238
  (
    n267,
    n126
  );


  buf
  g239
  (
    KeyWire_0_30,
    n130
  );


  buf
  g240
  (
    n243,
    n151
  );


  buf
  g241
  (
    n227,
    n115
  );


  buf
  g242
  (
    n254,
    n119
  );


  buf
  g243
  (
    n213,
    n109
  );


  buf
  g244
  (
    n187,
    n135
  );


  buf
  g245
  (
    n215,
    n141
  );


  buf
  g246
  (
    n181,
    n143
  );


  not
  g247
  (
    KeyWire_0_33,
    n129
  );


  not
  g248
  (
    n212,
    n142
  );


  buf
  g249
  (
    n179,
    n146
  );


  not
  g250
  (
    n174,
    n94
  );


  not
  g251
  (
    n191,
    n158
  );


  buf
  g252
  (
    KeyWire_0_2,
    n137
  );


  buf
  g253
  (
    n300,
    n168
  );


  not
  g254
  (
    n289,
    n171
  );


  buf
  g255
  (
    n292,
    n177
  );


  not
  g256
  (
    n296,
    n176
  );


  not
  g257
  (
    n291,
    n174
  );


  not
  g258
  (
    n293,
    n169
  );


  not
  g259
  (
    n282,
    n176
  );


  not
  g260
  (
    n301,
    n175
  );


  buf
  g261
  (
    n283,
    n170
  );


  buf
  g262
  (
    n299,
    n171
  );


  buf
  g263
  (
    n288,
    n169
  );


  not
  g264
  (
    n298,
    n172
  );


  buf
  g265
  (
    n297,
    n174
  );


  not
  g266
  (
    n290,
    n168
  );


  buf
  g267
  (
    n287,
    n175
  );


  buf
  g268
  (
    n302,
    n167
  );


  not
  g269
  (
    n285,
    n170
  );


  buf
  g270
  (
    n294,
    n172
  );


  buf
  g271
  (
    n295,
    n173
  );


  buf
  g272
  (
    n286,
    n167
  );


  not
  g273
  (
    n284,
    n173
  );


  not
  g274
  (
    n281,
    n177
  );


  not
  g275
  (
    n309,
    n292
  );


  not
  g276
  (
    n315,
    n286
  );


  not
  g277
  (
    n307,
    n285
  );


  not
  g278
  (
    n311,
    n293
  );


  buf
  g279
  (
    n305,
    n287
  );


  not
  g280
  (
    n317,
    n291
  );


  buf
  g281
  (
    n312,
    n281
  );


  buf
  g282
  (
    n306,
    n296
  );


  not
  g283
  (
    n308,
    n178
  );


  buf
  g284
  (
    n304,
    n179
  );


  nor
  g285
  (
    n310,
    n180,
    n294
  );


  or
  g286
  (
    KeyWire_0_29,
    n295,
    n282
  );


  xnor
  g287
  (
    n313,
    n288,
    n180
  );


  xor
  g288
  (
    KeyWire_0_11,
    n178,
    n179
  );


  and
  g289
  (
    n303,
    n284,
    n283
  );


  xnor
  g290
  (
    n318,
    n290,
    n289
  );


  not
  g291
  (
    n357,
    n307
  );


  buf
  g292
  (
    n371,
    n318
  );


  buf
  g293
  (
    n346,
    n306
  );


  not
  g294
  (
    n339,
    n308
  );


  buf
  g295
  (
    n323,
    n311
  );


  buf
  g296
  (
    n364,
    n303
  );


  buf
  g297
  (
    n335,
    n310
  );


  buf
  g298
  (
    n324,
    n306
  );


  not
  g299
  (
    n347,
    n312
  );


  not
  g300
  (
    n329,
    n304
  );


  buf
  g301
  (
    n328,
    n311
  );


  buf
  g302
  (
    n320,
    n310
  );


  buf
  g303
  (
    n340,
    n305
  );


  not
  g304
  (
    n363,
    n314
  );


  not
  g305
  (
    KeyWire_0_53,
    n312
  );


  buf
  g306
  (
    n369,
    n315
  );


  not
  g307
  (
    n336,
    n307
  );


  not
  g308
  (
    n334,
    n318
  );


  buf
  g309
  (
    n337,
    n308
  );


  buf
  g310
  (
    n360,
    n315
  );


  buf
  g311
  (
    n368,
    n303
  );


  not
  g312
  (
    n319,
    n314
  );


  buf
  g313
  (
    n372,
    n303
  );


  not
  g314
  (
    n355,
    n317
  );


  buf
  g315
  (
    n365,
    n313
  );


  not
  g316
  (
    n381,
    n304
  );


  buf
  g317
  (
    n341,
    n313
  );


  not
  g318
  (
    n327,
    n304
  );


  buf
  g319
  (
    KeyWire_0_45,
    n316
  );


  buf
  g320
  (
    n366,
    n307
  );


  buf
  g321
  (
    n353,
    n311
  );


  not
  g322
  (
    n348,
    n305
  );


  buf
  g323
  (
    n351,
    n314
  );


  buf
  g324
  (
    n321,
    n313
  );


  not
  g325
  (
    n343,
    n305
  );


  buf
  g326
  (
    n332,
    n303
  );


  not
  g327
  (
    n370,
    n317
  );


  buf
  g328
  (
    n377,
    n316
  );


  not
  g329
  (
    n326,
    n305
  );


  buf
  g330
  (
    KeyWire_0_1,
    n317
  );


  not
  g331
  (
    n376,
    n306
  );


  not
  g332
  (
    n345,
    n315
  );


  buf
  g333
  (
    n359,
    n315
  );


  not
  g334
  (
    n361,
    n312
  );


  buf
  g335
  (
    n338,
    n308
  );


  buf
  g336
  (
    n379,
    n314
  );


  not
  g337
  (
    n367,
    n313
  );


  not
  g338
  (
    n333,
    n308
  );


  not
  g339
  (
    n322,
    n309
  );


  not
  g340
  (
    n358,
    n317
  );


  not
  g341
  (
    n352,
    n309
  );


  buf
  g342
  (
    n342,
    n304
  );


  not
  g343
  (
    n344,
    n307
  );


  not
  g344
  (
    n375,
    n311
  );


  not
  g345
  (
    n354,
    n312
  );


  not
  g346
  (
    n374,
    n318
  );


  buf
  g347
  (
    n380,
    n310
  );


  not
  g348
  (
    n331,
    n309
  );


  buf
  g349
  (
    n330,
    n310
  );


  not
  g350
  (
    n373,
    n316
  );


  buf
  g351
  (
    n325,
    n309
  );


  not
  g352
  (
    n356,
    n306
  );


  buf
  g353
  (
    n362,
    n316
  );


  not
  g354
  (
    KeyWire_0_5,
    n187
  );


  buf
  g355
  (
    n415,
    n339
  );


  not
  g356
  (
    n403,
    n344
  );


  not
  g357
  (
    n390,
    n337
  );


  buf
  g358
  (
    n417,
    n325
  );


  buf
  g359
  (
    n407,
    n346
  );


  buf
  g360
  (
    n401,
    n333
  );


  not
  g361
  (
    KeyWire_0_62,
    n331
  );


  not
  g362
  (
    n414,
    n182
  );


  not
  g363
  (
    n400,
    n193
  );


  not
  g364
  (
    n394,
    n181
  );


  buf
  g365
  (
    n416,
    n341
  );


  buf
  g366
  (
    n404,
    n322
  );


  buf
  g367
  (
    n385,
    n192
  );


  buf
  g368
  (
    n413,
    n334
  );


  not
  g369
  (
    n409,
    n335
  );


  buf
  g370
  (
    n388,
    n186
  );


  buf
  g371
  (
    n418,
    n352
  );


  buf
  g372
  (
    n402,
    n330
  );


  buf
  g373
  (
    n384,
    n345
  );


  buf
  g374
  (
    KeyWire_0_43,
    n338
  );


  buf
  g375
  (
    n391,
    n323
  );


  not
  g376
  (
    n386,
    n183
  );


  not
  g377
  (
    n412,
    n343
  );


  not
  g378
  (
    n383,
    n332
  );


  buf
  g379
  (
    n382,
    n328
  );


  buf
  g380
  (
    n408,
    n342
  );


  not
  g381
  (
    n406,
    n192
  );


  and
  g382
  (
    n395,
    n185,
    n326,
    n336
  );


  nor
  g383
  (
    n398,
    n190,
    n340,
    n188,
    n182
  );


  xnor
  g384
  (
    n399,
    n354,
    n181,
    n187,
    n347
  );


  xnor
  g385
  (
    n410,
    n324,
    n190,
    n321,
    n185
  );


  nor
  g386
  (
    n392,
    n355,
    n320,
    n191,
    n353
  );


  xnor
  g387
  (
    n389,
    n183,
    n184,
    n348,
    n188
  );


  or
  g388
  (
    n405,
    n350,
    n319,
    n184,
    n329
  );


  or
  g389
  (
    n387,
    n189,
    n191,
    n186,
    n327
  );


  nand
  g390
  (
    n396,
    n351,
    n189,
    n349,
    n193
  );


  nand
  g391
  (
    n429,
    n393,
    n24,
    n395,
    n394
  );


  and
  g392
  (
    n452,
    n383,
    n297,
    n20,
    n399
  );


  or
  g393
  (
    n444,
    n359,
    n378,
    n393,
    n398
  );


  and
  g394
  (
    KeyWire_0_19,
    n394,
    n22,
    n383
  );


  nor
  g395
  (
    n433,
    n298,
    n367,
    n383,
    n392
  );


  xnor
  g396
  (
    n460,
    n383,
    n24,
    n358,
    n22
  );


  xnor
  g397
  (
    n441,
    n370,
    n26,
    n378,
    n364
  );


  xor
  g398
  (
    n451,
    n26,
    n386,
    n362,
    n374
  );


  nor
  g399
  (
    n456,
    n20,
    n21,
    n375,
    n376
  );


  nor
  g400
  (
    n427,
    n363,
    n362,
    n396,
    n357
  );


  and
  g401
  (
    n436,
    n25,
    n400,
    n377,
    n356
  );


  or
  g402
  (
    n426,
    n392,
    n24,
    n373,
    n397
  );


  nand
  g403
  (
    n442,
    n21,
    n19,
    n360,
    n385
  );


  and
  g404
  (
    n453,
    n389,
    n365,
    n397,
    n381
  );


  xnor
  g405
  (
    n458,
    n373,
    n23,
    n361,
    n385
  );


  or
  g406
  (
    n421,
    n23,
    n398,
    n395,
    n25
  );


  nor
  g407
  (
    n446,
    n24,
    n374,
    n392,
    n388
  );


  and
  g408
  (
    n434,
    n388,
    n359,
    n20,
    n360
  );


  nand
  g409
  (
    n457,
    n391,
    n372,
    n198,
    n377
  );


  nor
  g410
  (
    n430,
    n21,
    n384,
    n386,
    n26
  );


  nor
  g411
  (
    KeyWire_0_44,
    n387,
    n300,
    n381,
    n197
  );


  xnor
  g412
  (
    n455,
    n392,
    n197,
    n380,
    n379
  );


  xnor
  g413
  (
    n459,
    n387,
    n382,
    n21,
    n388
  );


  xor
  g414
  (
    n439,
    n371,
    n389,
    n366,
    n368
  );


  xor
  g415
  (
    n425,
    n194,
    n386,
    n363,
    n391
  );


  xnor
  g416
  (
    n419,
    n380,
    n26,
    n395,
    n25
  );


  and
  g417
  (
    n447,
    n398,
    n399,
    n369,
    n384
  );


  xnor
  g418
  (
    n420,
    n23,
    n299,
    n391,
    n393
  );


  xnor
  g419
  (
    n454,
    n390,
    n364,
    n361,
    n393
  );


  xor
  g420
  (
    n448,
    n382,
    n385,
    n375,
    n379
  );


  and
  g421
  (
    n437,
    n23,
    n368,
    n196,
    n387
  );


  nor
  g422
  (
    n428,
    n398,
    n195,
    n382,
    n390
  );


  xor
  g423
  (
    n438,
    n365,
    n399,
    n386,
    n384
  );


  xor
  g424
  (
    n449,
    n372,
    n397,
    n396
  );


  nor
  g425
  (
    n440,
    n389,
    n196,
    n382,
    n390
  );


  or
  g426
  (
    n450,
    n25,
    n376,
    n396,
    n399
  );


  xor
  g427
  (
    n431,
    n389,
    n194,
    n367,
    n385
  );


  or
  g428
  (
    n424,
    n19,
    n371,
    n384,
    n20
  );


  xor
  g429
  (
    KeyWire_0_3,
    n387,
    n400,
    n395,
    n394
  );


  or
  g430
  (
    n422,
    n388,
    n369,
    n397,
    n22
  );


  nand
  g431
  (
    n445,
    n391,
    n366,
    n394,
    n370
  );


  or
  g432
  (
    KeyWire_0_51,
    n301,
    n390,
    n302,
    n195
  );


  xnor
  g433
  (
    n474,
    n412,
    n411,
    n437
  );


  and
  g434
  (
    n469,
    n404,
    n405,
    n428,
    n400
  );


  xnor
  g435
  (
    n478,
    n408,
    n425,
    n405,
    n414
  );


  nor
  g436
  (
    n483,
    n422,
    n405,
    n424,
    n403
  );


  xor
  g437
  (
    n462,
    n414,
    n433,
    n420,
    n409
  );


  nor
  g438
  (
    n475,
    n432,
    n411,
    n405,
    n409
  );


  nor
  g439
  (
    KeyWire_0_0,
    n401,
    n406,
    n418,
    n408
  );


  nand
  g440
  (
    n481,
    n409,
    n401,
    n418,
    n443
  );


  nand
  g441
  (
    n473,
    n415,
    n414,
    n416,
    n413
  );


  nor
  g442
  (
    n463,
    n418,
    n415,
    n426,
    n404
  );


  xor
  g443
  (
    n479,
    n403,
    n414,
    n415,
    n412
  );


  or
  g444
  (
    n471,
    n417,
    n408,
    n402
  );


  xor
  g445
  (
    n485,
    n407,
    n406,
    n401,
    n417
  );


  nand
  g446
  (
    n464,
    n439,
    n407,
    n431,
    n413
  );


  or
  g447
  (
    n465,
    n412,
    n430,
    n409,
    n436
  );


  nand
  g448
  (
    n468,
    n403,
    n406,
    n412,
    n416
  );


  xnor
  g449
  (
    n484,
    n413,
    n417,
    n402,
    n408
  );


  or
  g450
  (
    n470,
    n438,
    n442,
    n417,
    n418
  );


  and
  g451
  (
    n466,
    n401,
    n429,
    n406,
    n404
  );


  or
  g452
  (
    n480,
    n407,
    n403,
    n416,
    n421
  );


  and
  g453
  (
    n467,
    n435,
    n400,
    n427,
    n419
  );


  nor
  g454
  (
    n472,
    n434,
    n411,
    n407,
    n404
  );


  xor
  g455
  (
    n461,
    n415,
    n410,
    n441,
    n423
  );


  xnor
  g456
  (
    KeyWire_0_12,
    n410,
    n413,
    n440,
    n402
  );


  or
  g457
  (
    n482,
    n410,
    n410,
    n416,
    n318
  );


  buf
  g458
  (
    n507,
    n466
  );


  buf
  g459
  (
    n508,
    n470
  );


  not
  g460
  (
    n509,
    n468
  );


  buf
  g461
  (
    n511,
    n463
  );


  buf
  g462
  (
    n499,
    n470
  );


  not
  g463
  (
    n501,
    n465
  );


  buf
  g464
  (
    n498,
    n469
  );


  buf
  g465
  (
    n503,
    n467
  );


  not
  g466
  (
    n504,
    n466
  );


  not
  g467
  (
    n487,
    n462
  );


  buf
  g468
  (
    KeyWire_0_55,
    n469
  );


  not
  g469
  (
    n497,
    n461
  );


  buf
  g470
  (
    n494,
    n462
  );


  not
  g471
  (
    n505,
    n469
  );


  not
  g472
  (
    n502,
    n469
  );


  buf
  g473
  (
    n486,
    n464
  );


  buf
  g474
  (
    n492,
    n468
  );


  not
  g475
  (
    n496,
    n467
  );


  not
  g476
  (
    n491,
    n464
  );


  buf
  g477
  (
    n493,
    n463
  );


  not
  g478
  (
    n510,
    n470
  );


  not
  g479
  (
    n513,
    n468
  );


  buf
  g480
  (
    n489,
    n471
  );


  not
  g481
  (
    n495,
    n468
  );


  buf
  g482
  (
    n514,
    n461
  );


  buf
  g483
  (
    n490,
    n465
  );


  not
  g484
  (
    n512,
    n471
  );


  buf
  g485
  (
    n500,
    n470
  );


  not
  g486
  (
    n488,
    n467
  );


  not
  g487
  (
    n515,
    n486
  );


  not
  g488
  (
    n522,
    n487
  );


  buf
  g489
  (
    n518,
    n472
  );


  buf
  g490
  (
    n520,
    n472
  );


  buf
  g491
  (
    n526,
    n472
  );


  buf
  g492
  (
    n525,
    n488
  );


  buf
  g493
  (
    n516,
    n488
  );


  not
  g494
  (
    n524,
    n471
  );


  xor
  g495
  (
    n521,
    n487,
    n472,
    n473,
    n471
  );


  xor
  g496
  (
    n523,
    n488,
    n487,
    n474
  );


  xnor
  g497
  (
    KeyWire_0_58,
    n473,
    n486,
    n474
  );


  nor
  g498
  (
    n517,
    n486,
    n473,
    n488
  );


  not
  g499
  (
    n530,
    n496
  );


  not
  g500
  (
    n549,
    n453
  );


  not
  g501
  (
    n561,
    n496
  );


  buf
  g502
  (
    n543,
    n449
  );


  buf
  g503
  (
    n538,
    n448
  );


  buf
  g504
  (
    n551,
    n454
  );


  buf
  g505
  (
    n554,
    n494
  );


  buf
  g506
  (
    KeyWire_0_14,
    n444
  );


  buf
  g507
  (
    n529,
    n200
  );


  not
  g508
  (
    n536,
    n519
  );


  buf
  g509
  (
    n558,
    n494
  );


  xnor
  g510
  (
    n539,
    n494,
    n520,
    n491
  );


  xnor
  g511
  (
    n531,
    n525,
    n451,
    n490,
    n515
  );


  and
  g512
  (
    n528,
    n497,
    n498,
    n446,
    n526
  );


  xor
  g513
  (
    n559,
    n202,
    n523,
    n492,
    n445
  );


  nand
  g514
  (
    n552,
    n201,
    n521,
    n497,
    n493
  );


  or
  g515
  (
    n560,
    n492,
    n456,
    n491,
    n495
  );


  xor
  g516
  (
    n556,
    n457,
    n526,
    n497,
    n490
  );


  xnor
  g517
  (
    n557,
    n517,
    n489,
    n518,
    n495
  );


  or
  g518
  (
    KeyWire_0_27,
    n497,
    n498,
    n525,
    n526
  );


  nand
  g519
  (
    n553,
    n522,
    n494,
    n499,
    n492
  );


  nor
  g520
  (
    n555,
    n493,
    n496,
    n199,
    n489
  );


  nand
  g521
  (
    n542,
    n447,
    n490,
    n521,
    n523
  );


  xor
  g522
  (
    n532,
    n199,
    n499,
    n524
  );


  and
  g523
  (
    KeyWire_0_24,
    n499,
    n459,
    n460,
    n455
  );


  and
  g524
  (
    n535,
    n516,
    n452,
    n517,
    n492
  );


  xnor
  g525
  (
    n534,
    n493,
    n450,
    n521,
    n518
  );


  nand
  g526
  (
    n527,
    n496,
    n522,
    n198,
    n489
  );


  or
  g527
  (
    n547,
    n163,
    n525,
    n515,
    n200
  );


  xnor
  g528
  (
    n548,
    n519,
    n491,
    n495,
    n516
  );


  xnor
  g529
  (
    n550,
    n522,
    n526,
    n491,
    n490
  );


  and
  g530
  (
    n545,
    n498,
    n458,
    n164,
    n489
  );


  xor
  g531
  (
    n541,
    n493,
    n524,
    n201,
    n498
  );


  xor
  g532
  (
    n537,
    n495,
    n522,
    n523,
    n524
  );


  nand
  g533
  (
    n544,
    n523,
    n525,
    n520,
    n524
  );


  not
  g534
  (
    n616,
    n551
  );


  not
  g535
  (
    n585,
    n550
  );


  not
  g536
  (
    n659,
    n530
  );


  not
  g537
  (
    n603,
    n548
  );


  not
  g538
  (
    n581,
    n531
  );


  buf
  g539
  (
    n656,
    n550
  );


  buf
  g540
  (
    n649,
    n534
  );


  buf
  g541
  (
    n576,
    n529
  );


  not
  g542
  (
    KeyWire_0_56,
    n540
  );


  not
  g543
  (
    n583,
    n531
  );


  buf
  g544
  (
    n622,
    n547
  );


  not
  g545
  (
    n634,
    n538
  );


  buf
  g546
  (
    n580,
    n536
  );


  buf
  g547
  (
    KeyWire_0_4,
    n545
  );


  buf
  g548
  (
    n600,
    n546
  );


  not
  g549
  (
    n602,
    n551
  );


  not
  g550
  (
    n609,
    n538
  );


  not
  g551
  (
    KeyWire_0_16,
    n547
  );


  buf
  g552
  (
    n658,
    n538
  );


  not
  g553
  (
    KeyWire_0_28,
    n533
  );


  not
  g554
  (
    n618,
    n543
  );


  not
  g555
  (
    n575,
    n551
  );


  buf
  g556
  (
    n662,
    n532
  );


  not
  g557
  (
    n654,
    n534
  );


  not
  g558
  (
    n570,
    n529
  );


  buf
  g559
  (
    n626,
    n536
  );


  buf
  g560
  (
    n646,
    n538
  );


  buf
  g561
  (
    n571,
    n541
  );


  not
  g562
  (
    n615,
    n528
  );


  buf
  g563
  (
    n655,
    n550
  );


  buf
  g564
  (
    n577,
    n547
  );


  not
  g565
  (
    n630,
    n548
  );


  buf
  g566
  (
    n610,
    n534
  );


  buf
  g567
  (
    n617,
    n549
  );


  not
  g568
  (
    n613,
    n527
  );


  not
  g569
  (
    n606,
    n536
  );


  not
  g570
  (
    n599,
    n544
  );


  buf
  g571
  (
    n657,
    n530
  );


  not
  g572
  (
    KeyWire_0_9,
    n545
  );


  buf
  g573
  (
    n564,
    n536
  );


  buf
  g574
  (
    n627,
    n543
  );


  buf
  g575
  (
    n637,
    n550
  );


  buf
  g576
  (
    n601,
    n545
  );


  buf
  g577
  (
    n647,
    n532
  );


  not
  g578
  (
    n653,
    n544
  );


  buf
  g579
  (
    n623,
    n546
  );


  not
  g580
  (
    n628,
    n541
  );


  not
  g581
  (
    n621,
    n546
  );


  not
  g582
  (
    n652,
    n548
  );


  buf
  g583
  (
    n586,
    n529
  );


  buf
  g584
  (
    n639,
    n549
  );


  buf
  g585
  (
    n596,
    n540
  );


  not
  g586
  (
    n614,
    n537
  );


  not
  g587
  (
    n632,
    n531
  );


  buf
  g588
  (
    n578,
    n535
  );


  buf
  g589
  (
    n619,
    n541
  );


  buf
  g590
  (
    KeyWire_0_41,
    n532
  );


  buf
  g591
  (
    n604,
    n535
  );


  not
  g592
  (
    n608,
    n530
  );


  not
  g593
  (
    n591,
    n551
  );


  buf
  g594
  (
    n629,
    n533
  );


  buf
  g595
  (
    KeyWire_0_36,
    n544
  );


  buf
  g596
  (
    n611,
    n552
  );


  buf
  g597
  (
    n612,
    n552
  );


  buf
  g598
  (
    n638,
    n552
  );


  not
  g599
  (
    n589,
    n535
  );


  buf
  g600
  (
    n605,
    n549
  );


  buf
  g601
  (
    n572,
    n537
  );


  buf
  g602
  (
    n640,
    n534
  );


  not
  g603
  (
    n663,
    n532
  );


  not
  g604
  (
    n620,
    n528
  );


  not
  g605
  (
    n592,
    n527
  );


  buf
  g606
  (
    n562,
    n535
  );


  buf
  g607
  (
    n598,
    n530
  );


  buf
  g608
  (
    n666,
    n527
  );


  not
  g609
  (
    n590,
    n533
  );


  not
  g610
  (
    n587,
    n549
  );


  not
  g611
  (
    n633,
    n541
  );


  not
  g612
  (
    n642,
    n531
  );


  not
  g613
  (
    n563,
    n540
  );


  not
  g614
  (
    n569,
    n539
  );


  not
  g615
  (
    n643,
    n547
  );


  buf
  g616
  (
    n661,
    n542
  );


  not
  g617
  (
    n597,
    n544
  );


  not
  g618
  (
    KeyWire_0_61,
    n528
  );


  buf
  g619
  (
    n644,
    n529
  );


  buf
  g620
  (
    n645,
    n540
  );


  buf
  g621
  (
    n595,
    n537
  );


  not
  g622
  (
    n636,
    n543
  );


  not
  g623
  (
    n660,
    n539
  );


  not
  g624
  (
    n566,
    n533
  );


  buf
  g625
  (
    n573,
    n553
  );


  buf
  g626
  (
    n624,
    n543
  );


  not
  g627
  (
    n664,
    n537
  );


  buf
  g628
  (
    n651,
    n553
  );


  not
  g629
  (
    n568,
    n539
  );


  not
  g630
  (
    n582,
    n528
  );


  not
  g631
  (
    n625,
    n552
  );


  buf
  g632
  (
    n667,
    n548
  );


  buf
  g633
  (
    n607,
    n539
  );


  not
  g634
  (
    n665,
    n545
  );


  not
  g635
  (
    n588,
    n546
  );


  buf
  g636
  (
    n635,
    n542
  );


  buf
  g637
  (
    n579,
    n542
  );


  buf
  g638
  (
    n594,
    n542
  );


  buf
  g639
  (
    n584,
    n527
  );


  xor
  g640
  (
    n683,
    n506,
    n503,
    n567,
    n589
  );


  and
  g641
  (
    n677,
    n574,
    n507,
    n555,
    n483
  );


  xor
  g642
  (
    n713,
    n561,
    n590,
    n508,
    n481
  );


  or
  g643
  (
    n680,
    n556,
    n503,
    n513,
    n479
  );


  xnor
  g644
  (
    n711,
    n502,
    n511,
    n509,
    n481
  );


  nand
  g645
  (
    n679,
    n580,
    n594,
    n505,
    n586
  );


  xor
  g646
  (
    n706,
    n553,
    n555,
    n481,
    n587
  );


  nor
  g647
  (
    n712,
    n502,
    n582,
    n575,
    n506
  );


  or
  g648
  (
    n696,
    n476,
    n561,
    n514,
    n502
  );


  xor
  g649
  (
    n700,
    n563,
    n559,
    n478,
    n477
  );


  xor
  g650
  (
    KeyWire_0_8,
    n560,
    n484,
    n508,
    n581
  );


  or
  g651
  (
    n715,
    n500,
    n582,
    n506,
    n556
  );


  xnor
  g652
  (
    n695,
    n558,
    n594,
    n482,
    n500
  );


  xor
  g653
  (
    n716,
    n593,
    n511,
    n514,
    n508
  );


  and
  g654
  (
    n694,
    n568,
    n588,
    n579,
    n505
  );


  xor
  g655
  (
    n678,
    n554,
    n507,
    n592,
    n566
  );


  or
  g656
  (
    n681,
    n564,
    n554,
    n583,
    n476
  );


  and
  g657
  (
    n671,
    n480,
    n572,
    n514
  );


  xnor
  g658
  (
    n684,
    n513,
    n500,
    n571,
    n564
  );


  and
  g659
  (
    n718,
    n596,
    n503,
    n482,
    n559
  );


  and
  g660
  (
    n669,
    n595,
    n568,
    n475,
    n512
  );


  nand
  g661
  (
    n686,
    n569,
    n573,
    n559,
    n476
  );


  xnor
  g662
  (
    n688,
    n475,
    n567,
    n500,
    n509
  );


  nand
  g663
  (
    KeyWire_0_32,
    n587,
    n584,
    n554,
    n575
  );


  nand
  g664
  (
    n672,
    n586,
    n477,
    n596,
    n505
  );


  nor
  g665
  (
    KeyWire_0_26,
    n565,
    n562,
    n555,
    n502
  );


  nand
  g666
  (
    n685,
    n565,
    n585,
    n501
  );


  nor
  g667
  (
    n674,
    n510,
    n511,
    n479,
    n579
  );


  xor
  g668
  (
    n670,
    n480,
    n510,
    n591,
    n474
  );


  xor
  g669
  (
    n673,
    n513,
    n558,
    n504,
    n501
  );


  nand
  g670
  (
    n692,
    n503,
    n557,
    n569,
    n511
  );


  nor
  g671
  (
    n668,
    n556,
    n580,
    n509,
    n584
  );


  nand
  g672
  (
    n710,
    n509,
    n475,
    n557,
    n478
  );


  nand
  g673
  (
    n717,
    n483,
    n560,
    n482,
    n504
  );


  or
  g674
  (
    n702,
    n576,
    n570,
    n571,
    n513
  );


  xnor
  g675
  (
    n704,
    n572,
    n560,
    n581,
    n561
  );


  nand
  g676
  (
    n705,
    n480,
    n476,
    n478,
    n477
  );


  xnor
  g677
  (
    n693,
    n570,
    n501,
    n588,
    n477
  );


  xor
  g678
  (
    n689,
    n597,
    n583,
    n557,
    n593
  );


  nand
  g679
  (
    n714,
    n504,
    n510,
    n589,
    n559
  );


  or
  g680
  (
    n699,
    n563,
    n595,
    n482,
    n558
  );


  nand
  g681
  (
    KeyWire_0_31,
    n590,
    n573,
    n562,
    n592
  );


  and
  g682
  (
    n709,
    n507,
    n555,
    n557,
    n591
  );


  xor
  g683
  (
    n703,
    n553,
    n556,
    n576,
    n479
  );


  xnor
  g684
  (
    n682,
    n566,
    n501,
    n483,
    n505
  );


  xor
  g685
  (
    n687,
    n507,
    n474,
    n561,
    n578
  );


  xnor
  g686
  (
    n691,
    n574,
    n483,
    n554,
    n512
  );


  xor
  g687
  (
    n701,
    n560,
    n475,
    n504,
    n480
  );


  nor
  g688
  (
    n676,
    n479,
    n512,
    n577
  );


  or
  g689
  (
    n690,
    n478,
    n506,
    n481,
    n510
  );


  nor
  g690
  (
    n698,
    n578,
    n512,
    n508,
    n558
  );


  buf
  g691
  (
    n732,
    n614
  );


  buf
  g692
  (
    n722,
    n629
  );


  buf
  g693
  (
    n745,
    n603
  );


  buf
  g694
  (
    n749,
    n670
  );


  not
  g695
  (
    n739,
    n676
  );


  not
  g696
  (
    KeyWire_0_15,
    n608
  );


  nor
  g697
  (
    n741,
    n612,
    n679
  );


  nor
  g698
  (
    n742,
    n626,
    n673
  );


  xor
  g699
  (
    n748,
    n613,
    n598,
    n601,
    n612
  );


  or
  g700
  (
    n747,
    n627,
    n610,
    n607,
    n680
  );


  or
  g701
  (
    n736,
    n626,
    n621,
    n630,
    n676
  );


  xor
  g702
  (
    n743,
    n674,
    n608,
    n675,
    n680
  );


  or
  g703
  (
    n733,
    n633,
    n631,
    n617
  );


  nand
  g704
  (
    n738,
    n603,
    n670,
    n629,
    n617
  );


  or
  g705
  (
    n724,
    n610,
    n619,
    n607,
    n621
  );


  nor
  g706
  (
    n750,
    n683,
    n674,
    n679,
    n682
  );


  nand
  g707
  (
    n746,
    n598,
    n630,
    n616,
    n597
  );


  xor
  g708
  (
    n740,
    n609,
    n611,
    n619,
    n615
  );


  or
  g709
  (
    n731,
    n682,
    n620,
    n675,
    n611
  );


  and
  g710
  (
    n726,
    n614,
    n622,
    n618,
    n623
  );


  and
  g711
  (
    n728,
    n625,
    n681,
    n632,
    n620
  );


  nor
  g712
  (
    n720,
    n605,
    n600,
    n623,
    n602
  );


  xor
  g713
  (
    n729,
    n628,
    n599,
    n615,
    n678
  );


  xor
  g714
  (
    n735,
    n668,
    n605,
    n613,
    n600
  );


  or
  g715
  (
    n719,
    n632,
    n627,
    n672,
    n677
  );


  nor
  g716
  (
    n730,
    n618,
    n606,
    n677,
    n683
  );


  nand
  g717
  (
    n744,
    n668,
    n624,
    n633,
    n681
  );


  and
  g718
  (
    n727,
    n609,
    n602,
    n604
  );


  xor
  g719
  (
    n725,
    n606,
    n625,
    n628,
    n624
  );


  xnor
  g720
  (
    n723,
    n634,
    n669,
    n601
  );


  xor
  g721
  (
    n721,
    n672,
    n673,
    n671,
    n678
  );


  nand
  g722
  (
    n737,
    n622,
    n671,
    n616,
    n599
  );


  or
  g723
  (
    n761,
    n686,
    n166,
    n690,
    n689
  );


  nand
  g724
  (
    n770,
    n717,
    n69,
    n699,
    n165
  );


  xor
  g725
  (
    n778,
    n705,
    n734,
    n724,
    n728
  );


  or
  g726
  (
    KeyWire_0_20,
    n700,
    n73,
    n699,
    n712
  );


  xnor
  g727
  (
    n765,
    n705,
    n701,
    n725,
    n702
  );


  and
  g728
  (
    KeyWire_0_34,
    n695,
    n74,
    n720,
    n688
  );


  or
  g729
  (
    n773,
    n72,
    n697,
    n691,
    n706
  );


  and
  g730
  (
    n780,
    n716,
    n710,
    n687,
    n715
  );


  xnor
  g731
  (
    n753,
    n731,
    n693,
    n165,
    n716
  );


  or
  g732
  (
    n766,
    n702,
    n733,
    n730,
    n732
  );


  or
  g733
  (
    n759,
    n698,
    n719,
    n714,
    n703
  );


  and
  g734
  (
    n768,
    n697,
    n701,
    n709,
    n691
  );


  nand
  g735
  (
    n775,
    n717,
    n685,
    n716,
    n729
  );


  nand
  g736
  (
    n769,
    n728,
    n717,
    n709,
    n712
  );


  and
  g737
  (
    n777,
    n727,
    n726,
    n715,
    n692
  );


  xnor
  g738
  (
    n767,
    n733,
    n721,
    n723,
    n695
  );


  nand
  g739
  (
    n758,
    n70,
    n72,
    n696,
    n71
  );


  nand
  g740
  (
    KeyWire_0_60,
    n75,
    n700,
    n694,
    n704
  );


  xor
  g741
  (
    n757,
    n708,
    n715,
    n726,
    n75
  );


  nor
  g742
  (
    n776,
    n729,
    n76,
    n720,
    n164
  );


  nor
  g743
  (
    n755,
    n730,
    n71,
    n732,
    n684
  );


  xnor
  g744
  (
    n760,
    n722,
    n686,
    n711,
    n713
  );


  and
  g745
  (
    n764,
    n689,
    n707,
    n714
  );


  xnor
  g746
  (
    n754,
    n74,
    n708,
    n713,
    n727
  );


  nand
  g747
  (
    n779,
    n723,
    n703,
    n719,
    n73
  );


  xor
  g748
  (
    n771,
    n731,
    n684,
    n715,
    n724
  );


  and
  g749
  (
    n772,
    n706,
    n711,
    n693,
    n70
  );


  xnor
  g750
  (
    n781,
    n704,
    n690,
    n77,
    n721
  );


  and
  g751
  (
    n752,
    n687,
    n725,
    n698,
    n710
  );


  xnor
  g752
  (
    n751,
    n688,
    n76,
    n694,
    n716
  );


  and
  g753
  (
    n762,
    n722,
    n685,
    n692,
    n696
  );


  or
  g754
  (
    n786,
    n652,
    n646,
    n657,
    n662
  );


  and
  g755
  (
    n791,
    n758,
    n637,
    n767,
    n660
  );


  xor
  g756
  (
    n790,
    n635,
    n665,
    n765,
    n657
  );


  xor
  g757
  (
    n796,
    n640,
    n766,
    n639,
    n666
  );


  nand
  g758
  (
    n802,
    n761,
    n650,
    n753,
    n653
  );


  nand
  g759
  (
    n800,
    n667,
    n648,
    n637,
    n764
  );


  xnor
  g760
  (
    n804,
    n649,
    n659,
    n634,
    n772
  );


  xnor
  g761
  (
    n782,
    n762,
    n754,
    n643,
    n647
  );


  xnor
  g762
  (
    n799,
    n771,
    n770,
    n642,
    n769
  );


  nand
  g763
  (
    n784,
    n773,
    n651,
    n645
  );


  nand
  g764
  (
    n789,
    n640,
    n203,
    n760,
    n755
  );


  xnor
  g765
  (
    n794,
    n661,
    n658,
    n756,
    n638
  );


  xor
  g766
  (
    n787,
    n648,
    n636,
    n644,
    n752
  );


  or
  g767
  (
    n801,
    n642,
    n653,
    n664,
    n655
  );


  or
  g768
  (
    n785,
    n646,
    n661,
    n649,
    n757
  );


  xnor
  g769
  (
    n793,
    n656,
    n641,
    n659,
    n663
  );


  nand
  g770
  (
    n788,
    n638,
    n768,
    n654,
    n663
  );


  xor
  g771
  (
    n783,
    n644,
    n660,
    n667,
    n647
  );


  nand
  g772
  (
    n795,
    n651,
    n639,
    n666,
    n662
  );


  nand
  g773
  (
    n792,
    n641,
    n202,
    n759,
    n665
  );


  xnor
  g774
  (
    n798,
    n664,
    n650,
    n751,
    n643
  );


  nand
  g775
  (
    n797,
    n636,
    n654,
    n656,
    n655
  );


  and
  g776
  (
    n803,
    n635,
    n652,
    n763,
    n658
  );


  not
  g777
  (
    n806,
    n790
  );


  not
  g778
  (
    n811,
    n799
  );


  buf
  g779
  (
    n832,
    n206
  );


  buf
  g780
  (
    KeyWire_0_38,
    n796
  );


  buf
  g781
  (
    n808,
    n217
  );


  not
  g782
  (
    n830,
    n206
  );


  xor
  g783
  (
    n827,
    n782,
    n222,
    n212
  );


  xnor
  g784
  (
    n819,
    n799,
    n205,
    n220
  );


  nor
  g785
  (
    n820,
    n803,
    n718,
    n222
  );


  xor
  g786
  (
    n815,
    n792,
    n783,
    n785
  );


  nand
  g787
  (
    n833,
    n205,
    n804,
    n218
  );


  and
  g788
  (
    n824,
    n804,
    n203,
    n798
  );


  or
  g789
  (
    n821,
    n214,
    n204,
    n801
  );


  or
  g790
  (
    n805,
    n214,
    n717,
    n786
  );


  xor
  g791
  (
    n810,
    n212,
    n789,
    n718
  );


  xnor
  g792
  (
    n828,
    n224,
    n217,
    n207
  );


  nor
  g793
  (
    n826,
    n221,
    n802,
    n223
  );


  and
  g794
  (
    n813,
    n784,
    n213,
    n221
  );


  xor
  g795
  (
    n823,
    n788,
    n223,
    n216
  );


  xor
  g796
  (
    n829,
    n794,
    n215
  );


  xor
  g797
  (
    n809,
    n787,
    n219,
    n216
  );


  xnor
  g798
  (
    n818,
    n718,
    n207,
    n209
  );


  xor
  g799
  (
    n812,
    n213,
    n718,
    n219
  );


  nand
  g800
  (
    n817,
    n208,
    n802,
    n800
  );


  or
  g801
  (
    n814,
    n791,
    n224,
    n220
  );


  and
  g802
  (
    n807,
    n795,
    n793,
    n210
  );


  or
  g803
  (
    n822,
    n204,
    n208,
    n218
  );


  nand
  g804
  (
    n834,
    n209,
    n800,
    n803
  );


  nor
  g805
  (
    n816,
    n798,
    n797,
    n211
  );


  nor
  g806
  (
    n831,
    n211,
    n210,
    n801
  );


  xor
  g807
  (
    n837,
    n741,
    n747,
    n750,
    n746
  );


  nor
  g808
  (
    n842,
    n739,
    n485,
    n814
  );


  nor
  g809
  (
    n847,
    n747,
    n807,
    n739,
    n736
  );


  xor
  g810
  (
    n839,
    n737,
    n748,
    n741
  );


  xor
  g811
  (
    n835,
    n744,
    n740,
    n748,
    n742
  );


  nand
  g812
  (
    n852,
    n225,
    n806,
    n743,
    n739
  );


  and
  g813
  (
    n843,
    n750,
    n741,
    n813,
    n738
  );


  or
  g814
  (
    KeyWire_0_35,
    n749,
    n735,
    n736
  );


  nand
  g815
  (
    n845,
    n735,
    n816,
    n815,
    n806
  );


  nor
  g816
  (
    n841,
    n811,
    n748,
    n746
  );


  nand
  g817
  (
    n846,
    n737,
    n745,
    n750,
    n749
  );


  nor
  g818
  (
    KeyWire_0_23,
    n747,
    n742,
    n810,
    n485
  );


  and
  g819
  (
    n856,
    n809,
    n742,
    n807,
    n808
  );


  xnor
  g820
  (
    n853,
    n745,
    n745,
    n735,
    n741
  );


  nor
  g821
  (
    KeyWire_0_37,
    n484,
    n809,
    n744,
    n746
  );


  nor
  g822
  (
    n850,
    n739,
    n750,
    n747,
    n812
  );


  or
  g823
  (
    n854,
    n738,
    n743,
    n484
  );


  nand
  g824
  (
    n840,
    n812,
    n735,
    n749,
    n745
  );


  nor
  g825
  (
    n848,
    n808,
    n740,
    n737,
    n805
  );


  or
  g826
  (
    n836,
    n811,
    n805,
    n749,
    n740
  );


  nand
  g827
  (
    n858,
    n814,
    n737,
    n484,
    n738
  );


  xnor
  g828
  (
    n855,
    n743,
    n742,
    n740,
    n736
  );


  nand
  g829
  (
    n838,
    n813,
    n744,
    n810
  );


  xnor
  g830
  (
    n851,
    n734,
    n815,
    n816,
    n738
  );


  and
  g831
  (
    n927,
    n238,
    n826,
    n80,
    n835
  );


  nor
  g832
  (
    n867,
    n250,
    n27,
    n274,
    n857
  );


  or
  g833
  (
    n932,
    n270,
    n27,
    n278,
    n263
  );


  and
  g834
  (
    n887,
    n230,
    n829,
    n855,
    n841
  );


  nand
  g835
  (
    n897,
    n854,
    n849,
    n842,
    n853
  );


  or
  g836
  (
    n914,
    n853,
    n846,
    n280,
    n830
  );


  nand
  g837
  (
    n920,
    n832,
    n259,
    n827,
    n853
  );


  or
  g838
  (
    n921,
    n79,
    n269,
    n240
  );


  nand
  g839
  (
    n869,
    n774,
    n265,
    n273,
    n827
  );


  or
  g840
  (
    KeyWire_0_18,
    n828,
    n852,
    n256,
    n260
  );


  or
  g841
  (
    n879,
    n246,
    n276,
    n239,
    n258
  );


  xor
  g842
  (
    n865,
    n819,
    n228,
    n241,
    n858
  );


  nand
  g843
  (
    n868,
    n849,
    n262,
    n858,
    n259
  );


  xor
  g844
  (
    n931,
    n244,
    n279,
    n272,
    n858
  );


  or
  g845
  (
    n859,
    n279,
    n850,
    n280
  );


  nor
  g846
  (
    n878,
    n250,
    n280,
    n258,
    n271
  );


  nor
  g847
  (
    n898,
    n839,
    n828,
    n779,
    n276
  );


  and
  g848
  (
    n902,
    n232,
    n837,
    n236,
    n265
  );


  nand
  g849
  (
    n892,
    n261,
    n823,
    n852,
    n271
  );


  xor
  g850
  (
    n910,
    n778,
    n81,
    n226,
    n266
  );


  nor
  g851
  (
    n894,
    n855,
    n848,
    n825,
    n79
  );


  xnor
  g852
  (
    KeyWire_0_48,
    n838,
    n242,
    n274,
    n260
  );


  or
  g853
  (
    n901,
    n279,
    n264,
    n275,
    n278
  );


  nor
  g854
  (
    n886,
    n822,
    n851,
    n857,
    n846
  );


  nor
  g855
  (
    KeyWire_0_13,
    n843,
    n237,
    n829,
    n239
  );


  nor
  g856
  (
    n907,
    n848,
    n256,
    n244,
    n260
  );


  xor
  g857
  (
    n871,
    n234,
    n272,
    n260,
    n840
  );


  or
  g858
  (
    n875,
    n837,
    n280,
    n233,
    n817
  );


  and
  g859
  (
    n924,
    n781,
    n836,
    n858,
    n818
  );


  xnor
  g860
  (
    n863,
    n266,
    n272,
    n234,
    n851
  );


  xnor
  g861
  (
    n872,
    n241,
    n845,
    n228,
    n245
  );


  or
  g862
  (
    n870,
    n854,
    n255,
    n842,
    n833
  );


  or
  g863
  (
    n899,
    n847,
    n819,
    n841,
    n817
  );


  nand
  g864
  (
    n905,
    n81,
    n830,
    n855,
    n836
  );


  nor
  g865
  (
    n911,
    n261,
    n823,
    n263,
    n246
  );


  nor
  g866
  (
    KeyWire_0_17,
    n834,
    n275,
    n831
  );


  or
  g867
  (
    n926,
    n826,
    n857,
    n251,
    n847
  );


  xor
  g868
  (
    n888,
    n818,
    n277,
    n267,
    n851
  );


  xor
  g869
  (
    n884,
    n267,
    n78,
    n856,
    n831
  );


  or
  g870
  (
    n929,
    n236,
    n846,
    n258,
    n833
  );


  xnor
  g871
  (
    n873,
    n850,
    n852,
    n856,
    n263
  );


  nor
  g872
  (
    n860,
    n845,
    n226,
    n248,
    n259
  );


  and
  g873
  (
    n925,
    n242,
    n232,
    n265,
    n829
  );


  or
  g874
  (
    n861,
    n843,
    n857,
    n279,
    n827
  );


  xor
  g875
  (
    n866,
    n820,
    n251,
    n822,
    n845
  );


  nand
  g876
  (
    n885,
    n833,
    n776,
    n821,
    n249
  );


  xor
  g877
  (
    n916,
    n267,
    n831,
    n834,
    n252
  );


  nand
  g878
  (
    KeyWire_0_6,
    n854,
    n775,
    n832,
    n830
  );


  nand
  g879
  (
    n880,
    n276,
    n272,
    n267,
    n265
  );


  xnor
  g880
  (
    n919,
    n82,
    n273,
    n277,
    n485
  );


  xor
  g881
  (
    n904,
    n270,
    n840,
    n238,
    n849
  );


  xnor
  g882
  (
    n889,
    n269,
    n273,
    n276,
    n253
  );


  xor
  g883
  (
    n935,
    n832,
    n227,
    n835,
    n847
  );


  or
  g884
  (
    KeyWire_0_25,
    n247,
    n247,
    n263,
    n243
  );


  and
  g885
  (
    KeyWire_0_49,
    n231,
    n839,
    n824,
    n254
  );


  nand
  g886
  (
    n933,
    n821,
    n229,
    n853,
    n262
  );


  nand
  g887
  (
    n876,
    n845,
    n834,
    n233,
    n277
  );


  xor
  g888
  (
    n923,
    n847,
    n848,
    n254
  );


  xor
  g889
  (
    n893,
    n271,
    n257,
    n844,
    n824
  );


  nor
  g890
  (
    n862,
    n838,
    n249,
    n849,
    n830
  );


  and
  g891
  (
    n890,
    n844,
    n828,
    n237,
    n833
  );


  or
  g892
  (
    n896,
    n227,
    n78,
    n266,
    n856
  );


  nor
  g893
  (
    n903,
    n261,
    n245,
    n832,
    n225
  );


  or
  g894
  (
    n930,
    n275,
    n780,
    n278,
    n268
  );


  and
  g895
  (
    n909,
    n850,
    n264,
    n856,
    n844
  );


  and
  g896
  (
    n934,
    n274,
    n80,
    n278,
    n820
  );


  nand
  g897
  (
    n928,
    n231,
    n229,
    n27,
    n855
  );


  and
  g898
  (
    n891,
    n268,
    n262,
    n266,
    n827
  );


  or
  g899
  (
    n883,
    n270,
    n230,
    n243,
    n852
  );


  and
  g900
  (
    n881,
    n851,
    n264,
    n277,
    n252
  );


  or
  g901
  (
    n908,
    n77,
    n235,
    n248,
    n271
  );


  xnor
  g902
  (
    n864,
    n269,
    n834,
    n828,
    n273
  );


  and
  g903
  (
    n913,
    n846,
    n253,
    n264,
    n261
  );


  xnor
  g904
  (
    n918,
    n854,
    n262,
    n235,
    n829
  );


  nor
  g905
  (
    n917,
    n274,
    n777,
    n831,
    n268
  );


  or
  g906
  (
    n912,
    n825,
    n82,
    n268,
    n270
  );


  and
  g907
  (
    n906,
    n255,
    n240,
    n257,
    n259
  );


  not
  g908
  (
    n950,
    n869
  );


  not
  g909
  (
    n936,
    n870
  );


  buf
  g910
  (
    n961,
    n881
  );


  buf
  g911
  (
    n938,
    n882
  );


  buf
  g912
  (
    KeyWire_0_10,
    n867
  );


  buf
  g913
  (
    n941,
    n859
  );


  not
  g914
  (
    n955,
    n880
  );


  buf
  g915
  (
    n963,
    n885
  );


  not
  g916
  (
    n965,
    n876
  );


  buf
  g917
  (
    n943,
    n887
  );


  not
  g918
  (
    n953,
    n872
  );


  buf
  g919
  (
    n964,
    n886
  );


  buf
  g920
  (
    n959,
    n862
  );


  not
  g921
  (
    n962,
    n888
  );


  not
  g922
  (
    n954,
    n863
  );


  not
  g923
  (
    n958,
    n873
  );


  not
  g924
  (
    KeyWire_0_63,
    n884
  );


  not
  g925
  (
    n945,
    n879
  );


  buf
  g926
  (
    n957,
    n878
  );


  buf
  g927
  (
    n949,
    n877
  );


  not
  g928
  (
    n937,
    n860
  );


  not
  g929
  (
    n942,
    n875
  );


  buf
  g930
  (
    n951,
    n871
  );


  buf
  g931
  (
    n947,
    n864
  );


  buf
  g932
  (
    n960,
    n866
  );


  buf
  g933
  (
    KeyWire_0_57,
    n883
  );


  buf
  g934
  (
    n948,
    n868
  );


  buf
  g935
  (
    n952,
    n874
  );


  buf
  g936
  (
    n956,
    n861
  );


  not
  g937
  (
    n939,
    n865
  );


  xnor
  g938
  (
    n975,
    n936,
    n922,
    n895,
    n959
  );


  xnor
  g939
  (
    n987,
    n946,
    n907,
    n913,
    n957
  );


  nor
  g940
  (
    n979,
    n960,
    n941,
    n942,
    n954
  );


  xnor
  g941
  (
    n973,
    n904,
    n936,
    n940,
    n950
  );


  nor
  g942
  (
    n971,
    n940,
    n945,
    n960,
    n890
  );


  or
  g943
  (
    n969,
    n910,
    n897,
    n937,
    n956
  );


  and
  g944
  (
    n984,
    n908,
    n915,
    n921,
    n898
  );


  nand
  g945
  (
    n980,
    n949,
    n943,
    n942,
    n952
  );


  and
  g946
  (
    n989,
    n953,
    n949,
    n914,
    n939
  );


  xnor
  g947
  (
    n966,
    n950,
    n961,
    n891,
    n901
  );


  nand
  g948
  (
    n974,
    n948,
    n954,
    n937,
    n945
  );


  xor
  g949
  (
    n983,
    n951,
    n944,
    n946,
    n952
  );


  and
  g950
  (
    n972,
    n959,
    n951,
    n903,
    n902
  );


  and
  g951
  (
    n985,
    n938,
    n899,
    n959,
    n900
  );


  xor
  g952
  (
    n970,
    n906,
    n919,
    n912,
    n961
  );


  and
  g953
  (
    n967,
    n956,
    n959,
    n894,
    n917
  );


  xnor
  g954
  (
    n976,
    n916,
    n943,
    n960,
    n958
  );


  or
  g955
  (
    n981,
    n958,
    n947,
    n905,
    n961
  );


  and
  g956
  (
    n977,
    n939,
    n911,
    n918,
    n955
  );


  nor
  g957
  (
    KeyWire_0_50,
    n893,
    n892,
    n961,
    n944
  );


  nand
  g958
  (
    n982,
    n957,
    n889,
    n953,
    n941
  );


  or
  g959
  (
    n978,
    n962,
    n920,
    n938,
    n947
  );


  xnor
  g960
  (
    n986,
    n948,
    n962,
    n958,
    n960
  );


  and
  g961
  (
    n988,
    n955,
    n896,
    n958,
    n909
  );


  or
  g962
  (
    n990,
    n988,
    n962,
    n963
  );


  buf
  g963
  (
    n991,
    n990
  );


  not
  g964
  (
    n992,
    n990
  );


  xor
  g965
  (
    n993,
    n963,
    n992
  );


  xnor
  g966
  (
    n996,
    n964,
    n965,
    n963
  );


  xnor
  g967
  (
    n994,
    n965,
    n964
  );


  nor
  g968
  (
    n995,
    n965,
    n993
  );


  and
  g969
  (
    n997,
    n965,
    n964,
    n963,
    n993
  );


  and
  g970
  (
    n1001,
    n934,
    n926,
    n931,
    n924
  );


  nand
  g971
  (
    n1000,
    n933,
    n83,
    n994
  );


  or
  g972
  (
    n1003,
    n927,
    n995,
    n935,
    n27
  );


  xnor
  g973
  (
    n998,
    n923,
    n930,
    n997
  );


  xor
  g974
  (
    n1002,
    n932,
    n929,
    n928,
    n996
  );


  or
  g975
  (
    n999,
    n166,
    n996,
    n989,
    n925
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n476,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n349,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n188,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n423,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n567,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n393,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n882,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n67,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n707,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n574,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n946,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n316,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n477,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n900,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n533,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n734,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n648,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n874,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n915,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n435,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n756,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n130,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n222,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n857,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n540,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n922,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n708,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n546,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n593,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n314,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n194,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n675,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n697,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n276,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n763,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n849,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n565,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n844,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n825,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n134,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n234,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n631,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n177,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n411,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n432,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n378,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n108,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n218,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n895,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n877,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n968,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n443,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n140,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n350,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n48,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n506,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n650,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n944,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n519,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n245,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n774,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n641,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n397,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n940,
    KeyNOTWire_0_63
  );


endmodule

