

module Stat_3904_76_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n3042,
  n3044,
  n3032,
  n3049,
  n3353,
  n3348,
  n3345,
  n3351,
  n3338,
  n3352,
  n3339,
  n3350,
  n3341,
  n3344,
  n3349,
  n3340,
  n3346,
  n3491,
  n3526,
  n3529,
  n3524,
  n3530,
  n3521,
  n3522,
  n3531,
  n3923,
  n3921,
  n3922,
  n3924,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n3042;
  output n3044;
  output n3032;
  output n3049;
  output n3353;
  output n3348;
  output n3345;
  output n3351;
  output n3338;
  output n3352;
  output n3339;
  output n3350;
  output n3341;
  output n3344;
  output n3349;
  output n3340;
  output n3346;
  output n3491;
  output n3526;
  output n3529;
  output n3524;
  output n3530;
  output n3521;
  output n3522;
  output n3531;
  output n3923;
  output n3921;
  output n3922;
  output n3924;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire n3030;
  wire n3031;
  wire n3033;
  wire n3034;
  wire n3035;
  wire n3036;
  wire n3037;
  wire n3038;
  wire n3039;
  wire n3040;
  wire n3041;
  wire n3043;
  wire n3045;
  wire n3046;
  wire n3047;
  wire n3048;
  wire n3050;
  wire n3051;
  wire n3052;
  wire n3053;
  wire n3054;
  wire n3055;
  wire n3056;
  wire n3057;
  wire n3058;
  wire n3059;
  wire n3060;
  wire n3061;
  wire n3062;
  wire n3063;
  wire n3064;
  wire n3065;
  wire n3066;
  wire n3067;
  wire n3068;
  wire n3069;
  wire n3070;
  wire n3071;
  wire n3072;
  wire n3073;
  wire n3074;
  wire n3075;
  wire n3076;
  wire n3077;
  wire n3078;
  wire n3079;
  wire n3080;
  wire n3081;
  wire n3082;
  wire n3083;
  wire n3084;
  wire n3085;
  wire n3086;
  wire n3087;
  wire n3088;
  wire n3089;
  wire n3090;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire n3095;
  wire n3096;
  wire n3097;
  wire n3098;
  wire n3099;
  wire n3100;
  wire n3101;
  wire n3102;
  wire n3103;
  wire n3104;
  wire n3105;
  wire n3106;
  wire n3107;
  wire n3108;
  wire n3109;
  wire n3110;
  wire n3111;
  wire n3112;
  wire n3113;
  wire n3114;
  wire n3115;
  wire n3116;
  wire n3117;
  wire n3118;
  wire n3119;
  wire n3120;
  wire n3121;
  wire n3122;
  wire n3123;
  wire n3124;
  wire n3125;
  wire n3126;
  wire n3127;
  wire n3128;
  wire n3129;
  wire n3130;
  wire n3131;
  wire n3132;
  wire n3133;
  wire n3134;
  wire n3135;
  wire n3136;
  wire n3137;
  wire n3138;
  wire n3139;
  wire n3140;
  wire n3141;
  wire n3142;
  wire n3143;
  wire n3144;
  wire n3145;
  wire n3146;
  wire n3147;
  wire n3148;
  wire n3149;
  wire n3150;
  wire n3151;
  wire n3152;
  wire n3153;
  wire n3154;
  wire n3155;
  wire n3156;
  wire n3157;
  wire n3158;
  wire n3159;
  wire n3160;
  wire n3161;
  wire n3162;
  wire n3163;
  wire n3164;
  wire n3165;
  wire n3166;
  wire n3167;
  wire n3168;
  wire n3169;
  wire n3170;
  wire n3171;
  wire n3172;
  wire n3173;
  wire n3174;
  wire n3175;
  wire n3176;
  wire n3177;
  wire n3178;
  wire n3179;
  wire n3180;
  wire n3181;
  wire n3182;
  wire n3183;
  wire n3184;
  wire n3185;
  wire n3186;
  wire n3187;
  wire n3188;
  wire n3189;
  wire n3190;
  wire n3191;
  wire n3192;
  wire n3193;
  wire n3194;
  wire n3195;
  wire n3196;
  wire n3197;
  wire n3198;
  wire n3199;
  wire n3200;
  wire n3201;
  wire n3202;
  wire n3203;
  wire n3204;
  wire n3205;
  wire n3206;
  wire n3207;
  wire n3208;
  wire n3209;
  wire n3210;
  wire n3211;
  wire n3212;
  wire n3213;
  wire n3214;
  wire n3215;
  wire n3216;
  wire n3217;
  wire n3218;
  wire n3219;
  wire n3220;
  wire n3221;
  wire n3222;
  wire n3223;
  wire n3224;
  wire n3225;
  wire n3226;
  wire n3227;
  wire n3228;
  wire n3229;
  wire n3230;
  wire n3231;
  wire n3232;
  wire n3233;
  wire n3234;
  wire n3235;
  wire n3236;
  wire n3237;
  wire n3238;
  wire n3239;
  wire n3240;
  wire n3241;
  wire n3242;
  wire n3243;
  wire n3244;
  wire n3245;
  wire n3246;
  wire n3247;
  wire n3248;
  wire n3249;
  wire n3250;
  wire n3251;
  wire n3252;
  wire n3253;
  wire n3254;
  wire n3255;
  wire n3256;
  wire n3257;
  wire n3258;
  wire n3259;
  wire n3260;
  wire n3261;
  wire n3262;
  wire n3263;
  wire n3264;
  wire n3265;
  wire n3266;
  wire n3267;
  wire n3268;
  wire n3269;
  wire n3270;
  wire n3271;
  wire n3272;
  wire n3273;
  wire n3274;
  wire n3275;
  wire n3276;
  wire n3277;
  wire n3278;
  wire n3279;
  wire n3280;
  wire n3281;
  wire n3282;
  wire n3283;
  wire n3284;
  wire n3285;
  wire n3286;
  wire n3287;
  wire n3288;
  wire n3289;
  wire n3290;
  wire n3291;
  wire n3292;
  wire n3293;
  wire n3294;
  wire n3295;
  wire n3296;
  wire n3297;
  wire n3298;
  wire n3299;
  wire n3300;
  wire n3301;
  wire n3302;
  wire n3303;
  wire n3304;
  wire n3305;
  wire n3306;
  wire n3307;
  wire n3308;
  wire n3309;
  wire n3310;
  wire n3311;
  wire n3312;
  wire n3313;
  wire n3314;
  wire n3315;
  wire n3316;
  wire n3317;
  wire n3318;
  wire n3319;
  wire n3320;
  wire n3321;
  wire n3322;
  wire n3323;
  wire n3324;
  wire n3325;
  wire n3326;
  wire n3327;
  wire n3328;
  wire n3329;
  wire n3330;
  wire n3331;
  wire n3332;
  wire n3333;
  wire n3334;
  wire n3335;
  wire n3336;
  wire n3337;
  wire n3342;
  wire n3343;
  wire n3347;
  wire n3354;
  wire n3355;
  wire n3356;
  wire n3357;
  wire n3358;
  wire n3359;
  wire n3360;
  wire n3361;
  wire n3362;
  wire n3363;
  wire n3364;
  wire n3365;
  wire n3366;
  wire n3367;
  wire n3368;
  wire n3369;
  wire n3370;
  wire n3371;
  wire n3372;
  wire n3373;
  wire n3374;
  wire n3375;
  wire n3376;
  wire n3377;
  wire n3378;
  wire n3379;
  wire n3380;
  wire n3381;
  wire n3382;
  wire n3383;
  wire n3384;
  wire n3385;
  wire n3386;
  wire n3387;
  wire n3388;
  wire n3389;
  wire n3390;
  wire n3391;
  wire n3392;
  wire n3393;
  wire n3394;
  wire n3395;
  wire n3396;
  wire n3397;
  wire n3398;
  wire n3399;
  wire n3400;
  wire n3401;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3407;
  wire n3408;
  wire n3409;
  wire n3410;
  wire n3411;
  wire n3412;
  wire n3413;
  wire n3414;
  wire n3415;
  wire n3416;
  wire n3417;
  wire n3418;
  wire n3419;
  wire n3420;
  wire n3421;
  wire n3422;
  wire n3423;
  wire n3424;
  wire n3425;
  wire n3426;
  wire n3427;
  wire n3428;
  wire n3429;
  wire n3430;
  wire n3431;
  wire n3432;
  wire n3433;
  wire n3434;
  wire n3435;
  wire n3436;
  wire n3437;
  wire n3438;
  wire n3439;
  wire n3440;
  wire n3441;
  wire n3442;
  wire n3443;
  wire n3444;
  wire n3445;
  wire n3446;
  wire n3447;
  wire n3448;
  wire n3449;
  wire n3450;
  wire n3451;
  wire n3452;
  wire n3453;
  wire n3454;
  wire n3455;
  wire n3456;
  wire n3457;
  wire n3458;
  wire n3459;
  wire n3460;
  wire n3461;
  wire n3462;
  wire n3463;
  wire n3464;
  wire n3465;
  wire n3466;
  wire n3467;
  wire n3468;
  wire n3469;
  wire n3470;
  wire n3471;
  wire n3472;
  wire n3473;
  wire n3474;
  wire n3475;
  wire n3476;
  wire n3477;
  wire n3478;
  wire n3479;
  wire n3480;
  wire n3481;
  wire n3482;
  wire n3483;
  wire n3484;
  wire n3485;
  wire n3486;
  wire n3487;
  wire n3488;
  wire n3489;
  wire n3490;
  wire n3492;
  wire n3493;
  wire n3494;
  wire n3495;
  wire n3496;
  wire n3497;
  wire n3498;
  wire n3499;
  wire n3500;
  wire n3501;
  wire n3502;
  wire n3503;
  wire n3504;
  wire n3505;
  wire n3506;
  wire n3507;
  wire n3508;
  wire n3509;
  wire n3510;
  wire n3511;
  wire n3512;
  wire n3513;
  wire n3514;
  wire n3515;
  wire n3516;
  wire n3517;
  wire n3518;
  wire n3519;
  wire n3520;
  wire n3523;
  wire n3525;
  wire n3527;
  wire n3528;
  wire n3532;
  wire n3533;
  wire n3534;
  wire n3535;
  wire n3536;
  wire n3537;
  wire n3538;
  wire n3539;
  wire n3540;
  wire n3541;
  wire n3542;
  wire n3543;
  wire n3544;
  wire n3545;
  wire n3546;
  wire n3547;
  wire n3548;
  wire n3549;
  wire n3550;
  wire n3551;
  wire n3552;
  wire n3553;
  wire n3554;
  wire n3555;
  wire n3556;
  wire n3557;
  wire n3558;
  wire n3559;
  wire n3560;
  wire n3561;
  wire n3562;
  wire n3563;
  wire n3564;
  wire n3565;
  wire n3566;
  wire n3567;
  wire n3568;
  wire n3569;
  wire n3570;
  wire n3571;
  wire n3572;
  wire n3573;
  wire n3574;
  wire n3575;
  wire n3576;
  wire n3577;
  wire n3578;
  wire n3579;
  wire n3580;
  wire n3581;
  wire n3582;
  wire n3583;
  wire n3584;
  wire n3585;
  wire n3586;
  wire n3587;
  wire n3588;
  wire n3589;
  wire n3590;
  wire n3591;
  wire n3592;
  wire n3593;
  wire n3594;
  wire n3595;
  wire n3596;
  wire n3597;
  wire n3598;
  wire n3599;
  wire n3600;
  wire n3601;
  wire n3602;
  wire n3603;
  wire n3604;
  wire n3605;
  wire n3606;
  wire n3607;
  wire n3608;
  wire n3609;
  wire n3610;
  wire n3611;
  wire n3612;
  wire n3613;
  wire n3614;
  wire n3615;
  wire n3616;
  wire n3617;
  wire n3618;
  wire n3619;
  wire n3620;
  wire n3621;
  wire n3622;
  wire n3623;
  wire n3624;
  wire n3625;
  wire n3626;
  wire n3627;
  wire n3628;
  wire n3629;
  wire n3630;
  wire n3631;
  wire n3632;
  wire n3633;
  wire n3634;
  wire n3635;
  wire n3636;
  wire n3637;
  wire n3638;
  wire n3639;
  wire n3640;
  wire n3641;
  wire n3642;
  wire n3643;
  wire n3644;
  wire n3645;
  wire n3646;
  wire n3647;
  wire n3648;
  wire n3649;
  wire n3650;
  wire n3651;
  wire n3652;
  wire n3653;
  wire n3654;
  wire n3655;
  wire n3656;
  wire n3657;
  wire n3658;
  wire n3659;
  wire n3660;
  wire n3661;
  wire n3662;
  wire n3663;
  wire n3664;
  wire n3665;
  wire n3666;
  wire n3667;
  wire n3668;
  wire n3669;
  wire n3670;
  wire n3671;
  wire n3672;
  wire n3673;
  wire n3674;
  wire n3675;
  wire n3676;
  wire n3677;
  wire n3678;
  wire n3679;
  wire n3680;
  wire n3681;
  wire n3682;
  wire n3683;
  wire n3684;
  wire n3685;
  wire n3686;
  wire n3687;
  wire n3688;
  wire n3689;
  wire n3690;
  wire n3691;
  wire n3692;
  wire n3693;
  wire n3694;
  wire n3695;
  wire n3696;
  wire n3697;
  wire n3698;
  wire n3699;
  wire n3700;
  wire n3701;
  wire n3702;
  wire n3703;
  wire n3704;
  wire n3705;
  wire n3706;
  wire n3707;
  wire n3708;
  wire n3709;
  wire n3710;
  wire n3711;
  wire n3712;
  wire n3713;
  wire n3714;
  wire n3715;
  wire n3716;
  wire n3717;
  wire n3718;
  wire n3719;
  wire n3720;
  wire n3721;
  wire n3722;
  wire n3723;
  wire n3724;
  wire n3725;
  wire n3726;
  wire n3727;
  wire n3728;
  wire n3729;
  wire n3730;
  wire n3731;
  wire n3732;
  wire n3733;
  wire n3734;
  wire n3735;
  wire n3736;
  wire n3737;
  wire n3738;
  wire n3739;
  wire n3740;
  wire n3741;
  wire n3742;
  wire n3743;
  wire n3744;
  wire n3745;
  wire n3746;
  wire n3747;
  wire n3748;
  wire n3749;
  wire n3750;
  wire n3751;
  wire n3752;
  wire n3753;
  wire n3754;
  wire n3755;
  wire n3756;
  wire n3757;
  wire n3758;
  wire n3759;
  wire n3760;
  wire n3761;
  wire n3762;
  wire n3763;
  wire n3764;
  wire n3765;
  wire n3766;
  wire n3767;
  wire n3768;
  wire n3769;
  wire n3770;
  wire n3771;
  wire n3772;
  wire n3773;
  wire n3774;
  wire n3775;
  wire n3776;
  wire n3777;
  wire n3778;
  wire n3779;
  wire n3780;
  wire n3781;
  wire n3782;
  wire n3783;
  wire n3784;
  wire n3785;
  wire n3786;
  wire n3787;
  wire n3788;
  wire n3789;
  wire n3790;
  wire n3791;
  wire n3792;
  wire n3793;
  wire n3794;
  wire n3795;
  wire n3796;
  wire n3797;
  wire n3798;
  wire n3799;
  wire n3800;
  wire n3801;
  wire n3802;
  wire n3803;
  wire n3804;
  wire n3805;
  wire n3806;
  wire n3807;
  wire n3808;
  wire n3809;
  wire n3810;
  wire n3811;
  wire n3812;
  wire n3813;
  wire n3814;
  wire n3815;
  wire n3816;
  wire n3817;
  wire n3818;
  wire n3819;
  wire n3820;
  wire n3821;
  wire n3822;
  wire n3823;
  wire n3824;
  wire n3825;
  wire n3826;
  wire n3827;
  wire n3828;
  wire n3829;
  wire n3830;
  wire n3831;
  wire n3832;
  wire n3833;
  wire n3834;
  wire n3835;
  wire n3836;
  wire n3837;
  wire n3838;
  wire n3839;
  wire n3840;
  wire n3841;
  wire n3842;
  wire n3843;
  wire n3844;
  wire n3845;
  wire n3846;
  wire n3847;
  wire n3848;
  wire n3849;
  wire n3850;
  wire n3851;
  wire n3852;
  wire n3853;
  wire n3854;
  wire n3855;
  wire n3856;
  wire n3857;
  wire n3858;
  wire n3859;
  wire n3860;
  wire n3861;
  wire n3862;
  wire n3863;
  wire n3864;
  wire n3865;
  wire n3866;
  wire n3867;
  wire n3868;
  wire n3869;
  wire n3870;
  wire n3871;
  wire n3872;
  wire n3873;
  wire n3874;
  wire n3875;
  wire n3876;
  wire n3877;
  wire n3878;
  wire n3879;
  wire n3880;
  wire n3881;
  wire n3882;
  wire n3883;
  wire n3884;
  wire n3885;
  wire n3886;
  wire n3887;
  wire n3888;
  wire n3889;
  wire n3890;
  wire n3891;
  wire n3892;
  wire n3893;
  wire n3894;
  wire n3895;
  wire n3896;
  wire n3897;
  wire n3898;
  wire n3899;
  wire n3900;
  wire n3901;
  wire n3902;
  wire n3903;
  wire n3904;
  wire n3905;
  wire n3906;
  wire n3907;
  wire n3908;
  wire n3909;
  wire n3910;
  wire n3911;
  wire n3912;
  wire n3913;
  wire n3914;
  wire n3915;
  wire n3916;
  wire n3917;
  wire n3918;
  wire n3919;
  wire n3920;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n43,
    n12
  );


  buf
  g1
  (
    n28,
    n1
  );


  not
  g2
  (
    n69,
    n10
  );


  buf
  g3
  (
    n64,
    n4
  );


  not
  g4
  (
    n48,
    n1
  );


  not
  g5
  (
    n33,
    n7
  );


  buf
  g6
  (
    n67,
    n9
  );


  buf
  g7
  (
    n59,
    n10
  );


  not
  g8
  (
    n56,
    n2
  );


  not
  g9
  (
    n54,
    n3
  );


  not
  g10
  (
    n22,
    n4
  );


  buf
  g11
  (
    n44,
    n9
  );


  not
  g12
  (
    n68,
    n7
  );


  buf
  g13
  (
    n53,
    n5
  );


  not
  g14
  (
    n38,
    n1
  );


  not
  g15
  (
    n25,
    n9
  );


  buf
  g16
  (
    n51,
    n13
  );


  not
  g17
  (
    n31,
    n6
  );


  not
  g18
  (
    n50,
    n11
  );


  not
  g19
  (
    n65,
    n5
  );


  not
  g20
  (
    n35,
    n6
  );


  buf
  g21
  (
    n34,
    n5
  );


  buf
  g22
  (
    n66,
    n11
  );


  buf
  g23
  (
    n23,
    n7
  );


  buf
  g24
  (
    n29,
    n5
  );


  not
  g25
  (
    n46,
    n8
  );


  not
  g26
  (
    n37,
    n10
  );


  not
  g27
  (
    n55,
    n9
  );


  buf
  g28
  (
    KeyWire_0_15,
    n6
  );


  not
  g29
  (
    n62,
    n12
  );


  buf
  g30
  (
    n49,
    n4
  );


  buf
  g31
  (
    n60,
    n3
  );


  not
  g32
  (
    KeyWire_0_10,
    n2
  );


  buf
  g33
  (
    n40,
    n7
  );


  buf
  g34
  (
    n58,
    n2
  );


  buf
  g35
  (
    n45,
    n12
  );


  buf
  g36
  (
    n24,
    n3
  );


  buf
  g37
  (
    n47,
    n4
  );


  not
  g38
  (
    n30,
    n8
  );


  not
  g39
  (
    n61,
    n11
  );


  buf
  g40
  (
    n36,
    n1
  );


  buf
  g41
  (
    n26,
    n3
  );


  not
  g42
  (
    n63,
    n6
  );


  not
  g43
  (
    n42,
    n12
  );


  buf
  g44
  (
    n27,
    n11
  );


  buf
  g45
  (
    n52,
    n8
  );


  not
  g46
  (
    n39,
    n8
  );


  not
  g47
  (
    n32,
    n2
  );


  buf
  g48
  (
    n41,
    n10
  );


  not
  g49
  (
    n71,
    n21
  );


  buf
  g50
  (
    n70,
    n21
  );


  not
  g51
  (
    n77,
    n70
  );


  not
  g52
  (
    n79,
    n70
  );


  not
  g53
  (
    n74,
    n71
  );


  buf
  g54
  (
    n73,
    n70
  );


  buf
  g55
  (
    n72,
    n71
  );


  not
  g56
  (
    n75,
    n70
  );


  buf
  g57
  (
    n78,
    n71
  );


  buf
  g58
  (
    n76,
    n71
  );


  not
  g59
  (
    n88,
    n76
  );


  not
  g60
  (
    n95,
    n76
  );


  buf
  g61
  (
    n100,
    n74
  );


  not
  g62
  (
    n86,
    n73
  );


  not
  g63
  (
    n103,
    n75
  );


  not
  g64
  (
    n94,
    n77
  );


  buf
  g65
  (
    n104,
    n74
  );


  buf
  g66
  (
    n106,
    n77
  );


  not
  g67
  (
    n101,
    n72
  );


  buf
  g68
  (
    n92,
    n73
  );


  not
  g69
  (
    KeyWire_0_1,
    n78
  );


  buf
  g70
  (
    n96,
    n74
  );


  buf
  g71
  (
    n98,
    n76
  );


  not
  g72
  (
    n85,
    n72
  );


  not
  g73
  (
    n105,
    n79
  );


  buf
  g74
  (
    n84,
    n74
  );


  not
  g75
  (
    n108,
    n72
  );


  buf
  g76
  (
    n87,
    n73
  );


  not
  g77
  (
    n81,
    n72
  );


  not
  g78
  (
    n102,
    n75
  );


  not
  g79
  (
    n90,
    n78
  );


  buf
  g80
  (
    n82,
    n78
  );


  not
  g81
  (
    n91,
    n79
  );


  buf
  g82
  (
    n93,
    n75
  );


  not
  g83
  (
    n99,
    n76
  );


  not
  g84
  (
    n97,
    n77
  );


  buf
  g85
  (
    n83,
    n78
  );


  not
  g86
  (
    n107,
    n77
  );


  or
  g87
  (
    n89,
    n73,
    n75
  );


  buf
  g88
  (
    n207,
    n87
  );


  buf
  g89
  (
    n167,
    n83
  );


  buf
  g90
  (
    n121,
    n90
  );


  not
  g91
  (
    n196,
    n99
  );


  not
  g92
  (
    n211,
    n95
  );


  buf
  g93
  (
    n162,
    n105
  );


  not
  g94
  (
    n178,
    n97
  );


  buf
  g95
  (
    n143,
    n97
  );


  not
  g96
  (
    n135,
    n89
  );


  not
  g97
  (
    n132,
    n82
  );


  buf
  g98
  (
    n158,
    n95
  );


  not
  g99
  (
    n214,
    n103
  );


  not
  g100
  (
    n110,
    n107
  );


  buf
  g101
  (
    n113,
    n86
  );


  not
  g102
  (
    n131,
    n91
  );


  not
  g103
  (
    n138,
    n96
  );


  not
  g104
  (
    n198,
    n93
  );


  not
  g105
  (
    n197,
    n83
  );


  not
  g106
  (
    n177,
    n83
  );


  not
  g107
  (
    n193,
    n94
  );


  not
  g108
  (
    n115,
    n82
  );


  buf
  g109
  (
    n134,
    n100
  );


  not
  g110
  (
    n187,
    n92
  );


  buf
  g111
  (
    n163,
    n80
  );


  buf
  g112
  (
    n218,
    n87
  );


  buf
  g113
  (
    n149,
    n89
  );


  buf
  g114
  (
    n156,
    n81
  );


  not
  g115
  (
    n140,
    n100
  );


  not
  g116
  (
    n200,
    n88
  );


  buf
  g117
  (
    n148,
    n99
  );


  buf
  g118
  (
    n146,
    n102
  );


  not
  g119
  (
    n142,
    n80
  );


  buf
  g120
  (
    n125,
    n89
  );


  buf
  g121
  (
    n186,
    n81
  );


  not
  g122
  (
    n209,
    n104
  );


  not
  g123
  (
    n194,
    n85
  );


  not
  g124
  (
    n202,
    n93
  );


  not
  g125
  (
    n176,
    n88
  );


  not
  g126
  (
    n151,
    n105
  );


  buf
  g127
  (
    n179,
    n80
  );


  buf
  g128
  (
    n122,
    n100
  );


  buf
  g129
  (
    n206,
    n96
  );


  not
  g130
  (
    n170,
    n87
  );


  buf
  g131
  (
    n133,
    n91
  );


  not
  g132
  (
    n185,
    n94
  );


  not
  g133
  (
    n150,
    n80
  );


  not
  g134
  (
    n199,
    n106
  );


  buf
  g135
  (
    n137,
    n106
  );


  not
  g136
  (
    n109,
    n101
  );


  not
  g137
  (
    n171,
    n90
  );


  buf
  g138
  (
    n173,
    n86
  );


  buf
  g139
  (
    n161,
    n101
  );


  buf
  g140
  (
    n117,
    n91
  );


  buf
  g141
  (
    n154,
    n81
  );


  not
  g142
  (
    n180,
    n98
  );


  buf
  g143
  (
    n114,
    n98
  );


  not
  g144
  (
    n215,
    n106
  );


  not
  g145
  (
    n174,
    n81
  );


  buf
  g146
  (
    n191,
    n105
  );


  not
  g147
  (
    n160,
    n96
  );


  buf
  g148
  (
    n159,
    n94
  );


  buf
  g149
  (
    n175,
    n89
  );


  not
  g150
  (
    n128,
    n85
  );


  buf
  g151
  (
    n129,
    n85
  );


  buf
  g152
  (
    n145,
    n88
  );


  not
  g153
  (
    n111,
    n99
  );


  buf
  g154
  (
    n210,
    n104
  );


  not
  g155
  (
    n201,
    n82
  );


  buf
  g156
  (
    KeyWire_0_23,
    n98
  );


  buf
  g157
  (
    n144,
    n103
  );


  not
  g158
  (
    n130,
    n84
  );


  buf
  g159
  (
    n166,
    n104
  );


  buf
  g160
  (
    n165,
    n91
  );


  buf
  g161
  (
    n124,
    n93
  );


  not
  g162
  (
    n190,
    n87
  );


  buf
  g163
  (
    n184,
    n93
  );


  not
  g164
  (
    n152,
    n98
  );


  buf
  g165
  (
    n216,
    n90
  );


  not
  g166
  (
    n169,
    n106
  );


  buf
  g167
  (
    n172,
    n95
  );


  buf
  g168
  (
    n126,
    n107
  );


  buf
  g169
  (
    n127,
    n82
  );


  not
  g170
  (
    n212,
    n102
  );


  not
  g171
  (
    n213,
    n84
  );


  not
  g172
  (
    n157,
    n103
  );


  buf
  g173
  (
    n192,
    n86
  );


  not
  g174
  (
    n189,
    n101
  );


  not
  g175
  (
    n195,
    n100
  );


  buf
  g176
  (
    n183,
    n95
  );


  not
  g177
  (
    n204,
    n90
  );


  not
  g178
  (
    n168,
    n84
  );


  not
  g179
  (
    n208,
    n94
  );


  buf
  g180
  (
    n205,
    n104
  );


  buf
  g181
  (
    n123,
    n84
  );


  buf
  g182
  (
    n155,
    n102
  );


  buf
  g183
  (
    n181,
    n92
  );


  not
  g184
  (
    n147,
    n97
  );


  buf
  g185
  (
    n119,
    n88
  );


  not
  g186
  (
    n139,
    n86
  );


  not
  g187
  (
    n217,
    n101
  );


  not
  g188
  (
    n188,
    n92
  );


  not
  g189
  (
    n203,
    n102
  );


  not
  g190
  (
    n136,
    n97
  );


  not
  g191
  (
    n153,
    n96
  );


  buf
  g192
  (
    n141,
    n103
  );


  buf
  g193
  (
    n112,
    n99
  );


  not
  g194
  (
    n118,
    n92
  );


  not
  g195
  (
    n182,
    n105
  );


  buf
  g196
  (
    n164,
    n85
  );


  not
  g197
  (
    n120,
    n83
  );


  nor
  g198
  (
    n309,
    n152,
    n142,
    n146,
    n191
  );


  xor
  g199
  (
    n288,
    n194,
    n200,
    n137,
    n174
  );


  xor
  g200
  (
    n314,
    n165,
    n147,
    n125,
    n164
  );


  xor
  g201
  (
    n254,
    n183,
    n188,
    n173,
    n159
  );


  or
  g202
  (
    n235,
    n115,
    n182,
    n196,
    n166
  );


  and
  g203
  (
    n295,
    n170,
    n120,
    n163,
    n199
  );


  xor
  g204
  (
    n281,
    n167,
    n19,
    n116
  );


  xnor
  g205
  (
    n306,
    n17,
    n191,
    n109
  );


  and
  g206
  (
    n264,
    n153,
    n123,
    n192,
    n15
  );


  xor
  g207
  (
    n279,
    n111,
    n163,
    n144,
    n154
  );


  nor
  g208
  (
    n298,
    n143,
    n158,
    n18,
    n151
  );


  and
  g209
  (
    n313,
    n125,
    n172,
    n127,
    n117
  );


  or
  g210
  (
    n239,
    n171,
    n149,
    n166,
    n131
  );


  and
  g211
  (
    n251,
    n117,
    n181,
    n109,
    n165
  );


  and
  g212
  (
    n299,
    n19,
    n127,
    n157,
    n186
  );


  xnor
  g213
  (
    n317,
    n128,
    n119,
    n193,
    n156
  );


  and
  g214
  (
    n243,
    n160,
    n155,
    n195,
    n123
  );


  xnor
  g215
  (
    n252,
    n139,
    n13,
    n114,
    n149
  );


  nand
  g216
  (
    n260,
    n182,
    n112,
    n156,
    n148
  );


  nor
  g217
  (
    n236,
    n132,
    n161,
    n175,
    n138
  );


  nor
  g218
  (
    n228,
    n200,
    n156,
    n17,
    n196
  );


  and
  g219
  (
    n280,
    n119,
    n173,
    n157,
    n14
  );


  xor
  g220
  (
    n238,
    n151,
    n158,
    n201,
    n162
  );


  or
  g221
  (
    n305,
    n197,
    n188,
    n129,
    n174
  );


  and
  g222
  (
    n265,
    n133,
    n117,
    n14
  );


  or
  g223
  (
    n272,
    n137,
    n157,
    n15,
    n134
  );


  nand
  g224
  (
    n296,
    n110,
    n186,
    n159,
    n192
  );


  nor
  g225
  (
    n282,
    n142,
    n162,
    n169,
    n111
  );


  nor
  g226
  (
    KeyWire_0_26,
    n130,
    n135,
    n190,
    n199
  );


  or
  g227
  (
    n271,
    n198,
    n138,
    n121,
    n188
  );


  or
  g228
  (
    n245,
    n149,
    n195,
    n157,
    n200
  );


  xnor
  g229
  (
    n266,
    n111,
    n192,
    n174,
    n176
  );


  or
  g230
  (
    n229,
    n124,
    n148,
    n143,
    n140
  );


  xnor
  g231
  (
    n246,
    n159,
    n185,
    n144,
    n121
  );


  xor
  g232
  (
    n292,
    n131,
    n132,
    n198,
    n163
  );


  nand
  g233
  (
    n315,
    n129,
    n170,
    n126,
    n137
  );


  or
  g234
  (
    n230,
    n118,
    n134,
    n184
  );


  nand
  g235
  (
    n277,
    n16,
    n194,
    n130,
    n165
  );


  xor
  g236
  (
    n283,
    n193,
    n118,
    n133,
    n159
  );


  xor
  g237
  (
    n274,
    n189,
    n119,
    n152,
    n135
  );


  nand
  g238
  (
    n276,
    n120,
    n133,
    n114,
    n124
  );


  nor
  g239
  (
    n307,
    n181,
    n109,
    n139,
    n18
  );


  nand
  g240
  (
    n231,
    n138,
    n137,
    n178,
    n187
  );


  xnor
  g241
  (
    n316,
    n133,
    n194,
    n128,
    n144
  );


  and
  g242
  (
    n250,
    n154,
    n164,
    n160,
    n138
  );


  xor
  g243
  (
    n267,
    n191,
    n146,
    n13,
    n167
  );


  and
  g244
  (
    KeyWire_0_2,
    n186,
    n150,
    n166,
    n172
  );


  nand
  g245
  (
    n258,
    n169,
    n187,
    n155,
    n161
  );


  xor
  g246
  (
    n261,
    n190,
    n116,
    n158,
    n130
  );


  xnor
  g247
  (
    n249,
    n127,
    n116,
    n185,
    n177
  );


  xor
  g248
  (
    n294,
    n192,
    n180,
    n173,
    n153
  );


  or
  g249
  (
    n269,
    n173,
    n169,
    n16,
    n126
  );


  and
  g250
  (
    n284,
    n116,
    n152,
    n198,
    n202
  );


  nand
  g251
  (
    n227,
    n150,
    n190,
    n115,
    n136
  );


  or
  g252
  (
    n268,
    n147,
    n199,
    n196,
    n124
  );


  xor
  g253
  (
    n225,
    n125,
    n199,
    n146,
    n142
  );


  and
  g254
  (
    n275,
    n160,
    n125,
    n170,
    n171
  );


  nor
  g255
  (
    n262,
    n123,
    n149,
    n162,
    n175
  );


  and
  g256
  (
    n220,
    n130,
    n197,
    n134,
    n15
  );


  xor
  g257
  (
    n244,
    n182,
    n136,
    n118,
    n172
  );


  or
  g258
  (
    n237,
    n179,
    n115,
    n196,
    n144
  );


  xor
  g259
  (
    n248,
    n190,
    n164,
    n111,
    n168
  );


  and
  g260
  (
    n293,
    n146,
    n110,
    n14
  );


  or
  g261
  (
    n308,
    n172,
    n168,
    n153,
    n193
  );


  nor
  g262
  (
    n241,
    n126,
    n124,
    n119,
    n132
  );


  xor
  g263
  (
    n234,
    n161,
    n140,
    n174,
    n136
  );


  nor
  g264
  (
    n240,
    n18,
    n186,
    n183,
    n168
  );


  nand
  g265
  (
    n302,
    n153,
    n17,
    n148,
    n198
  );


  xnor
  g266
  (
    n300,
    n181,
    n178,
    n164,
    n131
  );


  nor
  g267
  (
    n233,
    n158,
    n194,
    n170,
    n163
  );


  xnor
  g268
  (
    n290,
    n177,
    n14,
    n201,
    n152
  );


  xor
  g269
  (
    n301,
    n179,
    n135,
    n110,
    n113
  );


  and
  g270
  (
    KeyWire_0_28,
    n185,
    n15,
    n17,
    n169
  );


  and
  g271
  (
    n318,
    n184,
    n145,
    n161,
    n155
  );


  and
  g272
  (
    n257,
    n114,
    n184,
    n195,
    n150
  );


  nand
  g273
  (
    n270,
    n202,
    n122,
    n143,
    n201
  );


  or
  g274
  (
    n297,
    n126,
    n175,
    n132,
    n121
  );


  nand
  g275
  (
    n247,
    n139,
    n147,
    n112,
    n154
  );


  or
  g276
  (
    n278,
    n166,
    n141,
    n151,
    n187
  );


  nand
  g277
  (
    n286,
    n16,
    n114,
    n180,
    n197
  );


  or
  g278
  (
    n259,
    n120,
    n187,
    n147,
    n171
  );


  and
  g279
  (
    n273,
    n188,
    n145,
    n179,
    n165
  );


  nand
  g280
  (
    n222,
    n135,
    n145,
    n193,
    n168
  );


  nor
  g281
  (
    n223,
    n131,
    n129,
    n182,
    n178
  );


  nand
  g282
  (
    n242,
    n191,
    n156,
    n183,
    n151
  );


  xnor
  g283
  (
    n263,
    n120,
    n167,
    n162,
    n128
  );


  and
  g284
  (
    n289,
    n189,
    n128,
    n143,
    n180
  );


  xor
  g285
  (
    n291,
    n175,
    n113,
    n201,
    n140
  );


  xnor
  g286
  (
    n310,
    n118,
    n112,
    n171,
    n181
  );


  xnor
  g287
  (
    n221,
    n123,
    n176,
    n180,
    n184
  );


  or
  g288
  (
    n232,
    n113,
    n200,
    n142,
    n112
  );


  nor
  g289
  (
    n256,
    n185,
    n195,
    n141
  );


  xnor
  g290
  (
    n287,
    n136,
    n183,
    n122,
    n189
  );


  nor
  g291
  (
    n219,
    n139,
    n177,
    n148,
    n154
  );


  nand
  g292
  (
    n255,
    n155,
    n129,
    n150,
    n141
  );


  nand
  g293
  (
    n303,
    n18,
    n178,
    n115,
    n122
  );


  xor
  g294
  (
    n224,
    n140,
    n13,
    n121,
    n122
  );


  xor
  g295
  (
    n304,
    n113,
    n189,
    n160,
    n176
  );


  xnor
  g296
  (
    n226,
    n197,
    n127,
    n16,
    n177
  );


  nand
  g297
  (
    n311,
    n179,
    n176,
    n145,
    n167
  );


  buf
  g298
  (
    n488,
    n305
  );


  not
  g299
  (
    n598,
    n303
  );


  buf
  g300
  (
    n602,
    n56
  );


  not
  g301
  (
    n464,
    n37
  );


  not
  g302
  (
    n478,
    n54
  );


  not
  g303
  (
    n630,
    n271
  );


  buf
  g304
  (
    n644,
    n299
  );


  not
  g305
  (
    n567,
    n50
  );


  not
  g306
  (
    n594,
    n236
  );


  not
  g307
  (
    n361,
    n249
  );


  not
  g308
  (
    n390,
    n309
  );


  buf
  g309
  (
    n638,
    n311
  );


  not
  g310
  (
    n486,
    n35
  );


  not
  g311
  (
    n398,
    n289
  );


  not
  g312
  (
    n528,
    n48
  );


  not
  g313
  (
    n495,
    n258
  );


  not
  g314
  (
    n351,
    n300
  );


  not
  g315
  (
    n492,
    n293
  );


  not
  g316
  (
    n608,
    n49
  );


  buf
  g317
  (
    n462,
    n286
  );


  buf
  g318
  (
    n424,
    n293
  );


  buf
  g319
  (
    n516,
    n248
  );


  buf
  g320
  (
    n575,
    n271
  );


  not
  g321
  (
    n490,
    n222
  );


  not
  g322
  (
    n384,
    n241
  );


  buf
  g323
  (
    n672,
    n31
  );


  not
  g324
  (
    n447,
    n305
  );


  buf
  g325
  (
    n694,
    n310
  );


  buf
  g326
  (
    KeyWire_0_18,
    n68
  );


  not
  g327
  (
    n596,
    n40
  );


  buf
  g328
  (
    n335,
    n60
  );


  not
  g329
  (
    n417,
    n308
  );


  not
  g330
  (
    n552,
    n240
  );


  not
  g331
  (
    n373,
    n292
  );


  buf
  g332
  (
    n499,
    n290
  );


  buf
  g333
  (
    n482,
    n27
  );


  buf
  g334
  (
    n321,
    n51
  );


  buf
  g335
  (
    n553,
    n233
  );


  buf
  g336
  (
    n660,
    n226
  );


  not
  g337
  (
    n584,
    n269
  );


  not
  g338
  (
    n662,
    n239
  );


  buf
  g339
  (
    n476,
    n228
  );


  not
  g340
  (
    n532,
    n247
  );


  not
  g341
  (
    n376,
    n220
  );


  buf
  g342
  (
    n381,
    n226
  );


  not
  g343
  (
    n623,
    n222
  );


  not
  g344
  (
    n481,
    n263
  );


  buf
  g345
  (
    n663,
    n256
  );


  not
  g346
  (
    n433,
    n61
  );


  buf
  g347
  (
    n400,
    n64
  );


  buf
  g348
  (
    n671,
    n223
  );


  not
  g349
  (
    n645,
    n299
  );


  buf
  g350
  (
    n382,
    n238
  );


  not
  g351
  (
    n619,
    n260
  );


  buf
  g352
  (
    n558,
    n63
  );


  not
  g353
  (
    n412,
    n59
  );


  buf
  g354
  (
    n467,
    n219
  );


  not
  g355
  (
    n333,
    n68
  );


  buf
  g356
  (
    n442,
    n39
  );


  buf
  g357
  (
    n425,
    n268
  );


  buf
  g358
  (
    n714,
    n234
  );


  not
  g359
  (
    n519,
    n247
  );


  buf
  g360
  (
    n523,
    n55
  );


  buf
  g361
  (
    n517,
    n258
  );


  not
  g362
  (
    n549,
    n242
  );


  buf
  g363
  (
    n325,
    n229
  );


  buf
  g364
  (
    n601,
    n312
  );


  buf
  g365
  (
    n401,
    n287
  );


  not
  g366
  (
    n568,
    n269
  );


  buf
  g367
  (
    n473,
    n63
  );


  not
  g368
  (
    n649,
    n49
  );


  buf
  g369
  (
    n665,
    n295
  );


  buf
  g370
  (
    n697,
    n244
  );


  buf
  g371
  (
    n520,
    n22
  );


  not
  g372
  (
    n359,
    n269
  );


  not
  g373
  (
    n421,
    n247
  );


  not
  g374
  (
    n348,
    n306
  );


  buf
  g375
  (
    n378,
    n66
  );


  buf
  g376
  (
    n624,
    n309
  );


  not
  g377
  (
    n484,
    n239
  );


  not
  g378
  (
    n542,
    n253
  );


  buf
  g379
  (
    n439,
    n240
  );


  buf
  g380
  (
    n580,
    n55
  );


  buf
  g381
  (
    n324,
    n273
  );


  not
  g382
  (
    n657,
    n267
  );


  not
  g383
  (
    n380,
    n234
  );


  not
  g384
  (
    n597,
    n312
  );


  not
  g385
  (
    n673,
    n245
  );


  buf
  g386
  (
    n328,
    n230
  );


  buf
  g387
  (
    n675,
    n232
  );


  not
  g388
  (
    n605,
    n243
  );


  not
  g389
  (
    n428,
    n257
  );


  not
  g390
  (
    n345,
    n228
  );


  not
  g391
  (
    n544,
    n255
  );


  not
  g392
  (
    n561,
    n317
  );


  buf
  g393
  (
    n537,
    n284
  );


  buf
  g394
  (
    n559,
    n45
  );


  not
  g395
  (
    n522,
    n292
  );


  buf
  g396
  (
    n620,
    n62
  );


  not
  g397
  (
    n684,
    n69
  );


  buf
  g398
  (
    n468,
    n250
  );


  buf
  g399
  (
    n547,
    n27
  );


  not
  g400
  (
    n666,
    n300
  );


  buf
  g401
  (
    n546,
    n264
  );


  not
  g402
  (
    n536,
    n289
  );


  not
  g403
  (
    n459,
    n294
  );


  not
  g404
  (
    n329,
    n24
  );


  buf
  g405
  (
    n677,
    n288
  );


  not
  g406
  (
    n573,
    n262
  );


  buf
  g407
  (
    n422,
    n274
  );


  buf
  g408
  (
    n338,
    n270
  );


  not
  g409
  (
    n385,
    n270
  );


  not
  g410
  (
    n477,
    n39
  );


  not
  g411
  (
    n450,
    n241
  );


  buf
  g412
  (
    n642,
    n291
  );


  not
  g413
  (
    n661,
    n52
  );


  buf
  g414
  (
    n524,
    n308
  );


  buf
  g415
  (
    n341,
    n301
  );


  not
  g416
  (
    n676,
    n227
  );


  not
  g417
  (
    n713,
    n233
  );


  not
  g418
  (
    n527,
    n25
  );


  buf
  g419
  (
    n610,
    n63
  );


  buf
  g420
  (
    n670,
    n285
  );


  not
  g421
  (
    n545,
    n239
  );


  buf
  g422
  (
    n703,
    n236
  );


  not
  g423
  (
    n399,
    n314
  );


  buf
  g424
  (
    n578,
    n231
  );


  buf
  g425
  (
    n678,
    n234
  );


  buf
  g426
  (
    n353,
    n25
  );


  not
  g427
  (
    n540,
    n41
  );


  buf
  g428
  (
    n629,
    n34
  );


  buf
  g429
  (
    n648,
    n278
  );


  buf
  g430
  (
    n514,
    n299
  );


  buf
  g431
  (
    n331,
    n25
  );


  buf
  g432
  (
    n330,
    n288
  );


  buf
  g433
  (
    n538,
    n268
  );


  buf
  g434
  (
    n408,
    n245
  );


  buf
  g435
  (
    n655,
    n291
  );


  buf
  g436
  (
    n680,
    n43
  );


  buf
  g437
  (
    n403,
    n38
  );


  not
  g438
  (
    n530,
    n65
  );


  not
  g439
  (
    n501,
    n36
  );


  not
  g440
  (
    n455,
    n279
  );


  buf
  g441
  (
    n705,
    n41
  );


  not
  g442
  (
    n413,
    n249
  );


  buf
  g443
  (
    n414,
    n259
  );


  buf
  g444
  (
    n491,
    n316
  );


  not
  g445
  (
    n591,
    n254
  );


  buf
  g446
  (
    n562,
    n36
  );


  not
  g447
  (
    n589,
    n303
  );


  not
  g448
  (
    n364,
    n255
  );


  not
  g449
  (
    n504,
    n296
  );


  not
  g450
  (
    n535,
    n53
  );


  not
  g451
  (
    n571,
    n243
  );


  buf
  g452
  (
    n487,
    n38
  );


  buf
  g453
  (
    n592,
    n314
  );


  buf
  g454
  (
    n430,
    n300
  );


  buf
  g455
  (
    n692,
    n29
  );


  buf
  g456
  (
    n458,
    n288
  );


  buf
  g457
  (
    n386,
    n248
  );


  buf
  g458
  (
    n465,
    n253
  );


  buf
  g459
  (
    n693,
    n266
  );


  not
  g460
  (
    n685,
    n290
  );


  buf
  g461
  (
    n687,
    n28
  );


  buf
  g462
  (
    KeyWire_0_20,
    n301
  );


  buf
  g463
  (
    n632,
    n33
  );


  buf
  g464
  (
    n449,
    n37
  );


  buf
  g465
  (
    n460,
    n264
  );


  not
  g466
  (
    n709,
    n24
  );


  not
  g467
  (
    n440,
    n313
  );


  not
  g468
  (
    n456,
    n298
  );


  not
  g469
  (
    n388,
    n259
  );


  not
  g470
  (
    n698,
    n225
  );


  buf
  g471
  (
    n457,
    n219
  );


  buf
  g472
  (
    n689,
    n302
  );


  buf
  g473
  (
    n706,
    n225
  );


  not
  g474
  (
    n643,
    n236
  );


  not
  g475
  (
    n690,
    n23
  );


  buf
  g476
  (
    n667,
    n33
  );


  buf
  g477
  (
    n548,
    n247
  );


  buf
  g478
  (
    n656,
    n265
  );


  not
  g479
  (
    n391,
    n244
  );


  buf
  g480
  (
    n659,
    n29
  );


  not
  g481
  (
    n498,
    n307
  );


  not
  g482
  (
    n534,
    n289
  );


  buf
  g483
  (
    n708,
    n226
  );


  buf
  g484
  (
    n368,
    n307
  );


  buf
  g485
  (
    n323,
    n246
  );


  not
  g486
  (
    KeyWire_0_19,
    n272
  );


  not
  g487
  (
    n543,
    n250
  );


  not
  g488
  (
    n654,
    n54
  );


  buf
  g489
  (
    n647,
    n273
  );


  not
  g490
  (
    n363,
    n296
  );


  not
  g491
  (
    n525,
    n263
  );


  not
  g492
  (
    n337,
    n302
  );


  buf
  g493
  (
    n683,
    n315
  );


  buf
  g494
  (
    n340,
    n292
  );


  not
  g495
  (
    n510,
    n297
  );


  not
  g496
  (
    n479,
    n299
  );


  not
  g497
  (
    n612,
    n67
  );


  not
  g498
  (
    n357,
    n44
  );


  not
  g499
  (
    n650,
    n47
  );


  buf
  g500
  (
    n393,
    n44
  );


  not
  g501
  (
    n441,
    n50
  );


  buf
  g502
  (
    n480,
    n271
  );


  not
  g503
  (
    n365,
    n249
  );


  buf
  g504
  (
    n370,
    n32
  );


  not
  g505
  (
    n434,
    n51
  );


  buf
  g506
  (
    n453,
    n231
  );


  not
  g507
  (
    n529,
    n30
  );


  not
  g508
  (
    n541,
    n242
  );


  not
  g509
  (
    n358,
    n315
  );


  not
  g510
  (
    n415,
    n28
  );


  not
  g511
  (
    n507,
    n223
  );


  not
  g512
  (
    n626,
    n304
  );


  buf
  g513
  (
    n349,
    n284
  );


  not
  g514
  (
    n668,
    n283
  );


  buf
  g515
  (
    n572,
    n260
  );


  buf
  g516
  (
    n585,
    n22
  );


  buf
  g517
  (
    n410,
    n230
  );


  not
  g518
  (
    n595,
    n221
  );


  not
  g519
  (
    n712,
    n316
  );


  not
  g520
  (
    n423,
    n69
  );


  not
  g521
  (
    n445,
    n221
  );


  not
  g522
  (
    n515,
    n276
  );


  buf
  g523
  (
    n371,
    n23
  );


  buf
  g524
  (
    n395,
    n49
  );


  buf
  g525
  (
    n429,
    n43
  );


  not
  g526
  (
    n627,
    n311
  );


  not
  g527
  (
    n352,
    n47
  );


  buf
  g528
  (
    n511,
    n254
  );


  not
  g529
  (
    n640,
    n264
  );


  not
  g530
  (
    n344,
    n224
  );


  buf
  g531
  (
    n702,
    n61
  );


  buf
  g532
  (
    n463,
    n274
  );


  buf
  g533
  (
    n446,
    n265
  );


  buf
  g534
  (
    n531,
    n219
  );


  buf
  g535
  (
    n471,
    n22
  );


  not
  g536
  (
    n669,
    n305
  );


  buf
  g537
  (
    n356,
    n60
  );


  not
  g538
  (
    n617,
    n258
  );


  not
  g539
  (
    n416,
    n58
  );


  not
  g540
  (
    n494,
    n56
  );


  buf
  g541
  (
    n607,
    n252
  );


  buf
  g542
  (
    n696,
    n228
  );


  buf
  g543
  (
    n618,
    n63
  );


  buf
  g544
  (
    n682,
    n219
  );


  buf
  g545
  (
    n686,
    n266
  );


  not
  g546
  (
    n664,
    n25
  );


  buf
  g547
  (
    n564,
    n260
  );


  buf
  g548
  (
    n461,
    n261
  );


  buf
  g549
  (
    n658,
    n50
  );


  not
  g550
  (
    n563,
    n291
  );


  buf
  g551
  (
    n320,
    n251
  );


  buf
  g552
  (
    n419,
    n295
  );


  buf
  g553
  (
    n653,
    n42
  );


  not
  g554
  (
    n707,
    n42
  );


  not
  g555
  (
    n437,
    n42
  );


  not
  g556
  (
    n389,
    n281
  );


  buf
  g557
  (
    n366,
    n220
  );


  not
  g558
  (
    n505,
    n37
  );


  not
  g559
  (
    n583,
    n275
  );


  buf
  g560
  (
    n674,
    n220
  );


  buf
  g561
  (
    n616,
    n308
  );


  not
  g562
  (
    n646,
    n32
  );


  not
  g563
  (
    n533,
    n48
  );


  not
  g564
  (
    n360,
    n232
  );


  not
  g565
  (
    n588,
    n265
  );


  not
  g566
  (
    n496,
    n317
  );


  buf
  g567
  (
    n443,
    n23
  );


  buf
  g568
  (
    n319,
    n30
  );


  not
  g569
  (
    n409,
    n286
  );


  not
  g570
  (
    n334,
    n279
  );


  not
  g571
  (
    n394,
    n225
  );


  not
  g572
  (
    n469,
    n248
  );


  not
  g573
  (
    n604,
    n296
  );


  buf
  g574
  (
    n715,
    n306
  );


  buf
  g575
  (
    n557,
    n235
  );


  not
  g576
  (
    n362,
    n286
  );


  not
  g577
  (
    n379,
    n272
  );


  not
  g578
  (
    n420,
    n240
  );


  not
  g579
  (
    n448,
    n227
  );


  buf
  g580
  (
    n350,
    n289
  );


  buf
  g581
  (
    n550,
    n43
  );


  buf
  g582
  (
    n509,
    n285
  );


  not
  g583
  (
    n586,
    n66
  );


  not
  g584
  (
    n322,
    n256
  );


  buf
  g585
  (
    n603,
    n257
  );


  not
  g586
  (
    n451,
    n291
  );


  buf
  g587
  (
    n405,
    n45
  );


  not
  g588
  (
    n699,
    n33
  );


  not
  g589
  (
    n502,
    n252
  );


  not
  g590
  (
    n474,
    n62
  );


  buf
  g591
  (
    n374,
    n27
  );


  not
  g592
  (
    n711,
    n250
  );


  buf
  g593
  (
    n569,
    n67
  );


  buf
  g594
  (
    n342,
    n243
  );


  buf
  g595
  (
    n375,
    n281
  );


  buf
  g596
  (
    n652,
    n257
  );


  buf
  g597
  (
    n570,
    n267
  );


  not
  g598
  (
    n622,
    n228
  );


  buf
  g599
  (
    n621,
    n248
  );


  buf
  g600
  (
    n639,
    n37
  );


  not
  g601
  (
    n611,
    n244
  );


  not
  g602
  (
    n444,
    n65
  );


  not
  g603
  (
    n427,
    n249
  );


  buf
  g604
  (
    n339,
    n302
  );


  not
  g605
  (
    n614,
    n67
  );


  buf
  g606
  (
    n633,
    n304
  );


  buf
  g607
  (
    n631,
    n245
  );


  not
  g608
  (
    n581,
    n274
  );


  not
  g609
  (
    n634,
    n26
  );


  buf
  g610
  (
    n369,
    n253
  );


  not
  g611
  (
    n336,
    n53
  );


  not
  g612
  (
    n565,
    n300
  );


  not
  g613
  (
    n377,
    n29
  );


  not
  g614
  (
    n392,
    n243
  );


  buf
  g615
  (
    n681,
    n285
  );


  buf
  g616
  (
    n452,
    n231
  );


  buf
  g617
  (
    n636,
    n306
  );


  buf
  g618
  (
    n411,
    n278
  );


  buf
  g619
  (
    n688,
    n309
  );


  buf
  g620
  (
    n466,
    n235
  );


  buf
  g621
  (
    n489,
    n311
  );


  not
  g622
  (
    n651,
    n258
  );


  not
  g623
  (
    n483,
    n290
  );


  buf
  g624
  (
    n518,
    n46
  );


  buf
  g625
  (
    n355,
    n23
  );


  buf
  g626
  (
    n574,
    n231
  );


  buf
  g627
  (
    n628,
    n303
  );


  buf
  g628
  (
    n396,
    n246
  );


  not
  g629
  (
    n539,
    n224
  );


  nand
  g630
  (
    n435,
    n286,
    n235,
    n34,
    n272
  );


  nor
  g631
  (
    n404,
    n277,
    n314,
    n230,
    n242
  );


  and
  g632
  (
    n346,
    n298,
    n40,
    n68,
    n285
  );


  nand
  g633
  (
    n526,
    n57,
    n262,
    n282,
    n292
  );


  nand
  g634
  (
    n710,
    n275,
    n287,
    n54,
    n44
  );


  nand
  g635
  (
    n576,
    n52,
    n274,
    n39,
    n287
  );


  and
  g636
  (
    n582,
    n242,
    n223,
    n251,
    n259
  );


  or
  g637
  (
    n577,
    n47,
    n50,
    n46,
    n317
  );


  nor
  g638
  (
    n566,
    n277,
    n58,
    n237,
    n253
  );


  xor
  g639
  (
    n347,
    n271,
    n69,
    n283,
    n312
  );


  xor
  g640
  (
    n609,
    n312,
    n36,
    n256,
    n267
  );


  xnor
  g641
  (
    n432,
    n284,
    n280,
    n252,
    n279
  );


  nor
  g642
  (
    n397,
    n281,
    n35,
    n52,
    n273
  );


  and
  g643
  (
    n637,
    n245,
    n240,
    n238,
    n280
  );


  xor
  g644
  (
    n704,
    n266,
    n237,
    n224,
    n280
  );


  xor
  g645
  (
    n695,
    n318,
    n57,
    n277,
    n273
  );


  and
  g646
  (
    n436,
    n21,
    n301,
    n282,
    n238
  );


  nor
  g647
  (
    n512,
    n256,
    n56,
    n281,
    n279
  );


  xnor
  g648
  (
    n470,
    n250,
    n310,
    n59,
    n298
  );


  and
  g649
  (
    n485,
    n48,
    n27,
    n278,
    n238
  );


  and
  g650
  (
    n508,
    n227,
    n257,
    n45,
    n241
  );


  and
  g651
  (
    n438,
    n28,
    n36,
    n268,
    n239
  );


  nand
  g652
  (
    n426,
    n35,
    n52,
    n306,
    n229
  );


  and
  g653
  (
    n606,
    n53,
    n254,
    n310
  );


  xor
  g654
  (
    n701,
    n278,
    n41,
    n24,
    n66
  );


  nand
  g655
  (
    n475,
    n293,
    n69,
    n47,
    n59
  );


  and
  g656
  (
    n554,
    n61,
    n267,
    n284,
    n270
  );


  nor
  g657
  (
    n590,
    n237,
    n40,
    n304,
    n269
  );


  or
  g658
  (
    n326,
    n313,
    n233,
    n57,
    n272
  );


  or
  g659
  (
    n497,
    n290,
    n264,
    n24,
    n311
  );


  nor
  g660
  (
    n383,
    n255,
    n40,
    n57,
    n32
  );


  xor
  g661
  (
    n613,
    n252,
    n230,
    n234,
    n295
  );


  nand
  g662
  (
    n579,
    n33,
    n262,
    n223,
    n61
  );


  xor
  g663
  (
    n343,
    n303,
    n255,
    n53,
    n260
  );


  nand
  g664
  (
    n372,
    n315,
    n55,
    n301,
    n49
  );


  xnor
  g665
  (
    n700,
    n54,
    n280,
    n224,
    n22
  );


  xnor
  g666
  (
    n418,
    n315,
    n39,
    n227,
    n275
  );


  or
  g667
  (
    n431,
    n283,
    n296,
    n60,
    n59
  );


  nor
  g668
  (
    n500,
    n236,
    n259,
    n65,
    n262
  );


  or
  g669
  (
    n691,
    n287,
    n232,
    n64
  );


  nand
  g670
  (
    n354,
    n276,
    n44,
    n65,
    n294
  );


  nor
  g671
  (
    n599,
    n45,
    n261,
    n307,
    n30
  );


  nand
  g672
  (
    n615,
    n38,
    n246,
    n51,
    n28
  );


  xor
  g673
  (
    n503,
    n294,
    n26,
    n275,
    n220
  );


  and
  g674
  (
    n332,
    n221,
    n316,
    n34,
    n29
  );


  nand
  g675
  (
    n587,
    n261,
    n288,
    n304,
    n282
  );


  or
  g676
  (
    n641,
    n241,
    n251,
    n222,
    n229
  );


  xnor
  g677
  (
    n367,
    n48,
    n265,
    n38,
    n222
  );


  xor
  g678
  (
    n555,
    n31,
    n56,
    n41,
    n51
  );


  xor
  g679
  (
    n406,
    n251,
    n68,
    n276,
    n46
  );


  xor
  g680
  (
    n556,
    n55,
    n26,
    n229,
    n67
  );


  nand
  g681
  (
    n454,
    n297,
    n298,
    n276,
    n307
  );


  and
  g682
  (
    n513,
    n270,
    n107,
    n244,
    n32
  );


  xor
  g683
  (
    n600,
    n31,
    n64,
    n42,
    n66
  );


  nor
  g684
  (
    n521,
    n266,
    n233,
    n297,
    n316
  );


  nand
  g685
  (
    n472,
    n34,
    n263,
    n282,
    n221
  );


  nand
  g686
  (
    n625,
    n21,
    n246,
    n58,
    n237
  );


  xor
  g687
  (
    n407,
    n317,
    n308,
    n31,
    n313
  );


  and
  g688
  (
    n493,
    n297,
    n43,
    n283,
    n46
  );


  or
  g689
  (
    n506,
    n277,
    n64,
    n26,
    n30
  );


  nor
  g690
  (
    n402,
    n58,
    n60,
    n268,
    n35
  );


  xnor
  g691
  (
    n551,
    n313,
    n226,
    n235,
    n225
  );


  and
  g692
  (
    n593,
    n254,
    n293,
    n309,
    n62
  );


  and
  g693
  (
    n560,
    n302,
    n305,
    n294,
    n314
  );


  nor
  g694
  (
    n635,
    n62,
    n261,
    n263,
    n295
  );


  buf
  g695
  (
    n1442,
    n422
  );


  not
  g696
  (
    n1700,
    n362
  );


  buf
  g697
  (
    n1791,
    n698
  );


  buf
  g698
  (
    n2190,
    n376
  );


  not
  g699
  (
    n1105,
    n379
  );


  not
  g700
  (
    n1802,
    n655
  );


  buf
  g701
  (
    n830,
    n666
  );


  not
  g702
  (
    n1670,
    n634
  );


  buf
  g703
  (
    n741,
    n442
  );


  not
  g704
  (
    n905,
    n510
  );


  buf
  g705
  (
    n1531,
    n596
  );


  buf
  g706
  (
    n1808,
    n568
  );


  not
  g707
  (
    n2086,
    n461
  );


  buf
  g708
  (
    n2047,
    n596
  );


  buf
  g709
  (
    n2161,
    n647
  );


  not
  g710
  (
    n2288,
    n714
  );


  buf
  g711
  (
    n1045,
    n340
  );


  buf
  g712
  (
    n2171,
    n617
  );


  not
  g713
  (
    n2076,
    n328
  );


  buf
  g714
  (
    n1667,
    n654
  );


  buf
  g715
  (
    n746,
    n673
  );


  not
  g716
  (
    n1939,
    n498
  );


  buf
  g717
  (
    n1421,
    n574
  );


  not
  g718
  (
    n1782,
    n568
  );


  not
  g719
  (
    n2023,
    n206
  );


  buf
  g720
  (
    n1735,
    n207
  );


  not
  g721
  (
    n976,
    n489
  );


  not
  g722
  (
    n1694,
    n388
  );


  not
  g723
  (
    n1770,
    n699
  );


  not
  g724
  (
    n1224,
    n340
  );


  not
  g725
  (
    n1773,
    n414
  );


  buf
  g726
  (
    n964,
    n695
  );


  not
  g727
  (
    n1816,
    n204
  );


  buf
  g728
  (
    n975,
    n586
  );


  not
  g729
  (
    n2182,
    n484
  );


  not
  g730
  (
    n2010,
    n530
  );


  not
  g731
  (
    n2138,
    n697
  );


  not
  g732
  (
    n1339,
    n550
  );


  not
  g733
  (
    n961,
    n418
  );


  buf
  g734
  (
    n2252,
    n397
  );


  not
  g735
  (
    n1737,
    n544
  );


  buf
  g736
  (
    n1261,
    n591
  );


  buf
  g737
  (
    n2088,
    n373
  );


  not
  g738
  (
    n1292,
    n403
  );


  not
  g739
  (
    n1824,
    n324
  );


  not
  g740
  (
    n2264,
    n605
  );


  not
  g741
  (
    n1803,
    n553
  );


  not
  g742
  (
    n1961,
    n692
  );


  not
  g743
  (
    n1249,
    n645
  );


  not
  g744
  (
    n1908,
    n352
  );


  not
  g745
  (
    n1898,
    n383
  );


  not
  g746
  (
    n799,
    n552
  );


  buf
  g747
  (
    n1477,
    n426
  );


  buf
  g748
  (
    n738,
    n666
  );


  buf
  g749
  (
    n1083,
    n398
  );


  not
  g750
  (
    n1362,
    n411
  );


  not
  g751
  (
    n1327,
    n427
  );


  buf
  g752
  (
    n2041,
    n627
  );


  buf
  g753
  (
    n1619,
    n326
  );


  buf
  g754
  (
    n1147,
    n593
  );


  not
  g755
  (
    n1853,
    n354
  );


  not
  g756
  (
    n1934,
    n364
  );


  not
  g757
  (
    n2224,
    n490
  );


  buf
  g758
  (
    n1199,
    n320
  );


  not
  g759
  (
    n1801,
    n325
  );


  not
  g760
  (
    n2119,
    n555
  );


  buf
  g761
  (
    n1676,
    n583
  );


  not
  g762
  (
    n1946,
    n684
  );


  buf
  g763
  (
    n1376,
    n589
  );


  not
  g764
  (
    n803,
    n429
  );


  buf
  g765
  (
    n995,
    n674
  );


  not
  g766
  (
    n2122,
    n350
  );


  not
  g767
  (
    n1532,
    n404
  );


  not
  g768
  (
    n2147,
    n644
  );


  buf
  g769
  (
    n1457,
    n592
  );


  buf
  g770
  (
    n2060,
    n370
  );


  buf
  g771
  (
    n1574,
    n494
  );


  not
  g772
  (
    n1515,
    n206
  );


  buf
  g773
  (
    n1091,
    n608
  );


  buf
  g774
  (
    n856,
    n501
  );


  buf
  g775
  (
    n2294,
    n542
  );


  buf
  g776
  (
    n1564,
    n580
  );


  not
  g777
  (
    n939,
    n331
  );


  buf
  g778
  (
    n2039,
    n703
  );


  buf
  g779
  (
    n1309,
    n489
  );


  buf
  g780
  (
    n980,
    n628
  );


  not
  g781
  (
    n1765,
    n393
  );


  not
  g782
  (
    n2095,
    n567
  );


  not
  g783
  (
    n1566,
    n367
  );


  not
  g784
  (
    n2205,
    n386
  );


  buf
  g785
  (
    n842,
    n436
  );


  buf
  g786
  (
    n1825,
    n567
  );


  buf
  g787
  (
    n1223,
    n634
  );


  buf
  g788
  (
    n1089,
    n445
  );


  buf
  g789
  (
    n900,
    n679
  );


  buf
  g790
  (
    n1271,
    n406
  );


  buf
  g791
  (
    n1377,
    n625
  );


  buf
  g792
  (
    n1208,
    n477
  );


  buf
  g793
  (
    n1635,
    n427
  );


  buf
  g794
  (
    n2134,
    n557
  );


  not
  g795
  (
    n2097,
    n508
  );


  not
  g796
  (
    n1634,
    n603
  );


  not
  g797
  (
    n1538,
    n574
  );


  not
  g798
  (
    n1661,
    n627
  );


  buf
  g799
  (
    n1864,
    n693
  );


  buf
  g800
  (
    n1328,
    n687
  );


  not
  g801
  (
    n1245,
    n529
  );


  buf
  g802
  (
    n2136,
    n468
  );


  not
  g803
  (
    n904,
    n349
  );


  not
  g804
  (
    n732,
    n344
  );


  buf
  g805
  (
    n2280,
    n488
  );


  not
  g806
  (
    n1962,
    n424
  );


  not
  g807
  (
    n1805,
    n497
  );


  buf
  g808
  (
    n824,
    n321
  );


  buf
  g809
  (
    n1390,
    n699
  );


  buf
  g810
  (
    n1965,
    n449
  );


  buf
  g811
  (
    n997,
    n479
  );


  not
  g812
  (
    n1892,
    n640
  );


  not
  g813
  (
    n1493,
    n634
  );


  not
  g814
  (
    n1783,
    n546
  );


  buf
  g815
  (
    n1313,
    n319
  );


  buf
  g816
  (
    n1907,
    n454
  );


  buf
  g817
  (
    n1144,
    n379
  );


  buf
  g818
  (
    n1970,
    n546
  );


  buf
  g819
  (
    n1752,
    n436
  );


  buf
  g820
  (
    n909,
    n621
  );


  not
  g821
  (
    n1507,
    n569
  );


  buf
  g822
  (
    n1828,
    n208
  );


  not
  g823
  (
    n1932,
    n613
  );


  buf
  g824
  (
    n1929,
    n334
  );


  not
  g825
  (
    n1657,
    n390
  );


  buf
  g826
  (
    n1546,
    n630
  );


  buf
  g827
  (
    n1052,
    n514
  );


  not
  g828
  (
    n1641,
    n564
  );


  not
  g829
  (
    n1451,
    n524
  );


  not
  g830
  (
    n1433,
    n500
  );


  buf
  g831
  (
    n1145,
    n533
  );


  buf
  g832
  (
    n935,
    n611
  );


  buf
  g833
  (
    n1659,
    n361
  );


  not
  g834
  (
    n1734,
    n629
  );


  not
  g835
  (
    n1882,
    n693
  );


  not
  g836
  (
    n2152,
    n535
  );


  not
  g837
  (
    n2167,
    n438
  );


  buf
  g838
  (
    n2258,
    n607
  );


  buf
  g839
  (
    n1523,
    n460
  );


  not
  g840
  (
    n1076,
    n217
  );


  not
  g841
  (
    n1902,
    n446
  );


  not
  g842
  (
    n1088,
    n451
  );


  not
  g843
  (
    KeyWire_0_25,
    n217
  );


  not
  g844
  (
    n1236,
    n527
  );


  not
  g845
  (
    n1118,
    n582
  );


  not
  g846
  (
    n1890,
    n577
  );


  not
  g847
  (
    n2087,
    n615
  );


  not
  g848
  (
    n1745,
    n475
  );


  not
  g849
  (
    n990,
    n559
  );


  buf
  g850
  (
    n2070,
    n516
  );


  not
  g851
  (
    n1494,
    n439
  );


  not
  g852
  (
    n1479,
    n682
  );


  buf
  g853
  (
    n866,
    n543
  );


  buf
  g854
  (
    n731,
    n649
  );


  buf
  g855
  (
    n1601,
    n358
  );


  buf
  g856
  (
    n1446,
    n342
  );


  not
  g857
  (
    n1235,
    n474
  );


  buf
  g858
  (
    n2213,
    n649
  );


  buf
  g859
  (
    n1817,
    n212
  );


  not
  g860
  (
    n1547,
    n582
  );


  buf
  g861
  (
    n1498,
    n709
  );


  buf
  g862
  (
    n2094,
    n492
  );


  buf
  g863
  (
    n1696,
    n686
  );


  not
  g864
  (
    n1420,
    n689
  );


  buf
  g865
  (
    n1660,
    n595
  );


  buf
  g866
  (
    n1002,
    n606
  );


  buf
  g867
  (
    n1300,
    n365
  );


  not
  g868
  (
    n1813,
    n353
  );


  buf
  g869
  (
    n1107,
    n656
  );


  buf
  g870
  (
    n1852,
    n359
  );


  buf
  g871
  (
    n901,
    n576
  );


  buf
  g872
  (
    n2265,
    n642
  );


  buf
  g873
  (
    n820,
    n434
  );


  not
  g874
  (
    n1146,
    n507
  );


  buf
  g875
  (
    n772,
    n348
  );


  buf
  g876
  (
    n844,
    n587
  );


  not
  g877
  (
    n1578,
    n354
  );


  not
  g878
  (
    n1520,
    n493
  );


  buf
  g879
  (
    n1203,
    n494
  );


  not
  g880
  (
    n1015,
    n652
  );


  not
  g881
  (
    n2042,
    n452
  );


  buf
  g882
  (
    n1681,
    n601
  );


  not
  g883
  (
    n1533,
    n585
  );


  buf
  g884
  (
    n1198,
    n618
  );


  buf
  g885
  (
    n1140,
    n554
  );


  not
  g886
  (
    n1407,
    n705
  );


  not
  g887
  (
    n1410,
    n369
  );


  not
  g888
  (
    n1304,
    n408
  );


  buf
  g889
  (
    n1256,
    n710
  );


  buf
  g890
  (
    n1098,
    n679
  );


  buf
  g891
  (
    n2084,
    n596
  );


  not
  g892
  (
    n1607,
    n375
  );


  not
  g893
  (
    n1597,
    n472
  );


  not
  g894
  (
    n1826,
    n693
  );


  buf
  g895
  (
    n1586,
    n576
  );


  not
  g896
  (
    n849,
    n713
  );


  not
  g897
  (
    n1218,
    n324
  );


  buf
  g898
  (
    n1286,
    n409
  );


  buf
  g899
  (
    n1190,
    n360
  );


  not
  g900
  (
    n1951,
    n79
  );


  buf
  g901
  (
    n1980,
    n531
  );


  not
  g902
  (
    n1189,
    n666
  );


  buf
  g903
  (
    n1373,
    n432
  );


  buf
  g904
  (
    n840,
    n581
  );


  buf
  g905
  (
    n1733,
    n493
  );


  not
  g906
  (
    n1889,
    n486
  );


  buf
  g907
  (
    n1363,
    n499
  );


  not
  g908
  (
    n1192,
    n627
  );


  buf
  g909
  (
    n1947,
    n359
  );


  buf
  g910
  (
    n1881,
    n594
  );


  not
  g911
  (
    n1220,
    n559
  );


  buf
  g912
  (
    n954,
    n499
  );


  buf
  g913
  (
    n1480,
    n469
  );


  buf
  g914
  (
    n1637,
    n413
  );


  not
  g915
  (
    n2002,
    n366
  );


  not
  g916
  (
    n1003,
    n520
  );


  buf
  g917
  (
    n1374,
    n470
  );


  not
  g918
  (
    n1150,
    n475
  );


  not
  g919
  (
    n984,
    n345
  );


  buf
  g920
  (
    n1713,
    n541
  );


  not
  g921
  (
    n940,
    n499
  );


  not
  g922
  (
    n1758,
    n683
  );


  buf
  g923
  (
    n1943,
    n603
  );


  buf
  g924
  (
    n2110,
    n552
  );


  buf
  g925
  (
    n1093,
    n534
  );


  not
  g926
  (
    n925,
    n460
  );


  not
  g927
  (
    n874,
    n491
  );


  not
  g928
  (
    n761,
    n504
  );


  not
  g929
  (
    n2072,
    n480
  );


  not
  g930
  (
    n1857,
    n457
  );


  buf
  g931
  (
    n1127,
    n615
  );


  not
  g932
  (
    n1900,
    n688
  );


  not
  g933
  (
    n1799,
    n425
  );


  buf
  g934
  (
    n2046,
    n214
  );


  not
  g935
  (
    n1682,
    n534
  );


  not
  g936
  (
    n2292,
    n597
  );


  buf
  g937
  (
    n1345,
    n514
  );


  buf
  g938
  (
    n1811,
    n466
  );


  buf
  g939
  (
    n2185,
    n449
  );


  buf
  g940
  (
    n1280,
    n367
  );


  buf
  g941
  (
    n2090,
    n690
  );


  buf
  g942
  (
    n1307,
    n401
  );


  not
  g943
  (
    n1720,
    n203
  );


  buf
  g944
  (
    n1398,
    n675
  );


  buf
  g945
  (
    n721,
    n335
  );


  buf
  g946
  (
    n1312,
    n418
  );


  buf
  g947
  (
    n2052,
    n561
  );


  buf
  g948
  (
    n771,
    n575
  );


  not
  g949
  (
    n2186,
    n538
  );


  not
  g950
  (
    n1129,
    n366
  );


  not
  g951
  (
    n1549,
    n444
  );


  buf
  g952
  (
    n1899,
    n620
  );


  not
  g953
  (
    n2108,
    n674
  );


  buf
  g954
  (
    n739,
    n624
  );


  not
  g955
  (
    n1982,
    n412
  );


  buf
  g956
  (
    n2151,
    n629
  );


  buf
  g957
  (
    n807,
    n678
  );


  buf
  g958
  (
    n1094,
    n683
  );


  not
  g959
  (
    n1579,
    n463
  );


  not
  g960
  (
    n949,
    n454
  );


  buf
  g961
  (
    n972,
    n472
  );


  buf
  g962
  (
    n1971,
    n620
  );


  buf
  g963
  (
    n1877,
    n697
  );


  buf
  g964
  (
    n1695,
    n608
  );


  not
  g965
  (
    n1596,
    n337
  );


  not
  g966
  (
    n850,
    n697
  );


  not
  g967
  (
    n1840,
    n480
  );


  buf
  g968
  (
    n1592,
    n488
  );


  buf
  g969
  (
    n1253,
    n518
  );


  not
  g970
  (
    n2170,
    n553
  );


  buf
  g971
  (
    n2049,
    n345
  );


  not
  g972
  (
    n854,
    n496
  );


  not
  g973
  (
    n1671,
    n695
  );


  not
  g974
  (
    n2035,
    n447
  );


  not
  g975
  (
    n1101,
    n537
  );


  buf
  g976
  (
    n1958,
    n512
  );


  buf
  g977
  (
    n718,
    n339
  );


  buf
  g978
  (
    n2123,
    n502
  );


  not
  g979
  (
    n1933,
    n506
  );


  buf
  g980
  (
    n1722,
    n503
  );


  not
  g981
  (
    n1460,
    n428
  );


  buf
  g982
  (
    n2121,
    n672
  );


  not
  g983
  (
    n784,
    n450
  );


  buf
  g984
  (
    n1148,
    n507
  );


  buf
  g985
  (
    n915,
    n520
  );


  not
  g986
  (
    n1501,
    n636
  );


  not
  g987
  (
    n1171,
    n423
  );


  not
  g988
  (
    n1035,
    n588
  );


  not
  g989
  (
    n2053,
    n529
  );


  buf
  g990
  (
    n1402,
    n451
  );


  not
  g991
  (
    n1760,
    n483
  );


  not
  g992
  (
    n1909,
    n632
  );


  buf
  g993
  (
    n2263,
    n582
  );


  buf
  g994
  (
    n1204,
    n594
  );


  not
  g995
  (
    n2293,
    n436
  );


  buf
  g996
  (
    n717,
    n617
  );


  buf
  g997
  (
    n1378,
    n625
  );


  buf
  g998
  (
    n1509,
    n544
  );


  not
  g999
  (
    n1931,
    n361
  );


  not
  g1000
  (
    n1797,
    n573
  );


  buf
  g1001
  (
    n1184,
    n506
  );


  buf
  g1002
  (
    n1417,
    n554
  );


  buf
  g1003
  (
    n1866,
    n419
  );


  buf
  g1004
  (
    n2183,
    n481
  );


  not
  g1005
  (
    n1250,
    n698
  );


  not
  g1006
  (
    n1488,
    n670
  );


  not
  g1007
  (
    n1196,
    n667
  );


  buf
  g1008
  (
    n1954,
    n391
  );


  not
  g1009
  (
    n1551,
    n698
  );


  not
  g1010
  (
    n2191,
    n538
  );


  buf
  g1011
  (
    n1880,
    n427
  );


  buf
  g1012
  (
    n2256,
    n659
  );


  not
  g1013
  (
    n1413,
    n337
  );


  not
  g1014
  (
    n1483,
    n412
  );


  buf
  g1015
  (
    n1205,
    n350
  );


  buf
  g1016
  (
    n2003,
    n323
  );


  buf
  g1017
  (
    n1941,
    n639
  );


  not
  g1018
  (
    n920,
    n413
  );


  buf
  g1019
  (
    n876,
    n496
  );


  not
  g1020
  (
    n1335,
    n336
  );


  not
  g1021
  (
    n1258,
    n638
  );


  buf
  g1022
  (
    n2162,
    n688
  );


  not
  g1023
  (
    n2251,
    n637
  );


  not
  g1024
  (
    n1461,
    n587
  );


  buf
  g1025
  (
    n1589,
    n557
  );


  buf
  g1026
  (
    n1133,
    n657
  );


  buf
  g1027
  (
    n791,
    n525
  );


  not
  g1028
  (
    n2139,
    n623
  );


  buf
  g1029
  (
    n769,
    n213
  );


  not
  g1030
  (
    n911,
    n608
  );


  buf
  g1031
  (
    n1357,
    n602
  );


  not
  g1032
  (
    n1974,
    n439
  );


  buf
  g1033
  (
    n1879,
    n573
  );


  buf
  g1034
  (
    n1210,
    n215
  );


  not
  g1035
  (
    n2021,
    n654
  );


  buf
  g1036
  (
    n835,
    n679
  );


  buf
  g1037
  (
    n983,
    n532
  );


  buf
  g1038
  (
    n765,
    n385
  );


  buf
  g1039
  (
    n1775,
    n646
  );


  buf
  g1040
  (
    n916,
    n455
  );


  not
  g1041
  (
    n1439,
    n407
  );


  buf
  g1042
  (
    n1216,
    n538
  );


  buf
  g1043
  (
    n1059,
    n371
  );


  not
  g1044
  (
    n730,
    n456
  );


  buf
  g1045
  (
    n1244,
    n707
  );


  buf
  g1046
  (
    n1215,
    n563
  );


  not
  g1047
  (
    n1856,
    n399
  );


  not
  g1048
  (
    n1058,
    n371
  );


  buf
  g1049
  (
    n838,
    n482
  );


  not
  g1050
  (
    n1871,
    n663
  );


  not
  g1051
  (
    n882,
    n513
  );


  buf
  g1052
  (
    n970,
    n547
  );


  buf
  g1053
  (
    n2019,
    n207
  );


  not
  g1054
  (
    n1382,
    n424
  );


  not
  g1055
  (
    n1301,
    n476
  );


  not
  g1056
  (
    n1703,
    n656
  );


  buf
  g1057
  (
    n1161,
    n692
  );


  not
  g1058
  (
    n1126,
    n696
  );


  not
  g1059
  (
    n1438,
    n418
  );


  buf
  g1060
  (
    n1102,
    n329
  );


  not
  g1061
  (
    n1379,
    n581
  );


  buf
  g1062
  (
    n1525,
    n535
  );


  buf
  g1063
  (
    n1495,
    n423
  );


  buf
  g1064
  (
    n1553,
    n374
  );


  buf
  g1065
  (
    n2159,
    n212
  );


  buf
  g1066
  (
    n960,
    n468
  );


  buf
  g1067
  (
    n1257,
    n485
  );


  not
  g1068
  (
    n1834,
    n557
  );


  not
  g1069
  (
    n1863,
    n652
  );


  buf
  g1070
  (
    n1921,
    n619
  );


  not
  g1071
  (
    n1677,
    n711
  );


  buf
  g1072
  (
    n2279,
    n341
  );


  buf
  g1073
  (
    n1023,
    n337
  );


  not
  g1074
  (
    n1251,
    n409
  );


  not
  g1075
  (
    n2005,
    n366
  );


  buf
  g1076
  (
    n1977,
    n456
  );


  not
  g1077
  (
    n2176,
    n565
  );


  buf
  g1078
  (
    n1743,
    n331
  );


  not
  g1079
  (
    n1370,
    n692
  );


  buf
  g1080
  (
    n1473,
    n341
  );


  not
  g1081
  (
    n1613,
    n691
  );


  not
  g1082
  (
    n852,
    n444
  );


  buf
  g1083
  (
    n1702,
    n339
  );


  not
  g1084
  (
    n1492,
    n509
  );


  not
  g1085
  (
    n1066,
    n423
  );


  buf
  g1086
  (
    n989,
    n432
  );


  buf
  g1087
  (
    n749,
    n704
  );


  buf
  g1088
  (
    n1367,
    n415
  );


  buf
  g1089
  (
    n1875,
    n500
  );


  buf
  g1090
  (
    n2179,
    n669
  );


  not
  g1091
  (
    n1818,
    n604
  );


  buf
  g1092
  (
    n1359,
    n346
  );


  not
  g1093
  (
    n1424,
    n381
  );


  not
  g1094
  (
    n1600,
    n688
  );


  buf
  g1095
  (
    n1202,
    n356
  );


  buf
  g1096
  (
    n1057,
    n410
  );


  buf
  g1097
  (
    n2209,
    n467
  );


  buf
  g1098
  (
    n1618,
    n671
  );


  buf
  g1099
  (
    n1310,
    n213
  );


  buf
  g1100
  (
    n1375,
    n370
  );


  not
  g1101
  (
    n1807,
    n411
  );


  not
  g1102
  (
    n2045,
    n555
  );


  buf
  g1103
  (
    n958,
    n578
  );


  buf
  g1104
  (
    n1711,
    n642
  );


  buf
  g1105
  (
    n2063,
    n463
  );


  buf
  g1106
  (
    n1165,
    n550
  );


  not
  g1107
  (
    n1777,
    n377
  );


  buf
  g1108
  (
    n2101,
    n468
  );


  buf
  g1109
  (
    n1873,
    n410
  );


  buf
  g1110
  (
    n1609,
    n395
  );


  buf
  g1111
  (
    n2141,
    n611
  );


  buf
  g1112
  (
    n1690,
    n585
  );


  not
  g1113
  (
    n1688,
    n475
  );


  buf
  g1114
  (
    n888,
    n484
  );


  buf
  g1115
  (
    n2201,
    n516
  );


  buf
  g1116
  (
    n1673,
    n215
  );


  not
  g1117
  (
    n1764,
    n502
  );


  buf
  g1118
  (
    n1496,
    n669
  );


  not
  g1119
  (
    n2056,
    n609
  );


  not
  g1120
  (
    n1726,
    n551
  );


  buf
  g1121
  (
    n2301,
    n537
  );


  not
  g1122
  (
    n1542,
    n570
  );


  buf
  g1123
  (
    n1883,
    n214
  );


  buf
  g1124
  (
    n998,
    n408
  );


  not
  g1125
  (
    n1463,
    n668
  );


  buf
  g1126
  (
    n832,
    n576
  );


  buf
  g1127
  (
    n804,
    n325
  );


  buf
  g1128
  (
    n1746,
    n528
  );


  not
  g1129
  (
    n1099,
    n496
  );


  not
  g1130
  (
    n2143,
    n512
  );


  not
  g1131
  (
    n843,
    n382
  );


  not
  g1132
  (
    n2081,
    n661
  );


  buf
  g1133
  (
    n2000,
    n585
  );


  buf
  g1134
  (
    n1638,
    n613
  );


  buf
  g1135
  (
    n2098,
    n696
  );


  not
  g1136
  (
    n2275,
    n320
  );


  not
  g1137
  (
    n2073,
    n393
  );


  not
  g1138
  (
    n1815,
    n210
  );


  not
  g1139
  (
    n1543,
    n465
  );


  buf
  g1140
  (
    n1485,
    n519
  );


  buf
  g1141
  (
    n1662,
    n524
  );


  not
  g1142
  (
    n973,
    n384
  );


  not
  g1143
  (
    n1399,
    n508
  );


  not
  g1144
  (
    n2018,
    n454
  );


  buf
  g1145
  (
    n1512,
    n511
  );


  not
  g1146
  (
    n1437,
    n355
  );


  buf
  g1147
  (
    n2120,
    n415
  );


  buf
  g1148
  (
    n1135,
    n592
  );


  buf
  g1149
  (
    n1858,
    n607
  );


  not
  g1150
  (
    n1298,
    n678
  );


  not
  g1151
  (
    n740,
    n337
  );


  not
  g1152
  (
    n1394,
    n641
  );


  buf
  g1153
  (
    n2029,
    n387
  );


  not
  g1154
  (
    n1436,
    n665
  );


  buf
  g1155
  (
    n1503,
    n672
  );


  not
  g1156
  (
    n1404,
    n564
  );


  not
  g1157
  (
    n716,
    n483
  );


  buf
  g1158
  (
    n2077,
    n395
  );


  buf
  g1159
  (
    n1558,
    n354
  );


  not
  g1160
  (
    n1964,
    n504
  );


  buf
  g1161
  (
    n1295,
    n541
  );


  not
  g1162
  (
    n1915,
    n566
  );


  not
  g1163
  (
    n1391,
    n488
  );


  not
  g1164
  (
    n1632,
    n652
  );


  buf
  g1165
  (
    n1927,
    n569
  );


  buf
  g1166
  (
    n944,
    n510
  );


  buf
  g1167
  (
    n720,
    n583
  );


  buf
  g1168
  (
    n2061,
    n643
  );


  buf
  g1169
  (
    n1790,
    n345
  );


  buf
  g1170
  (
    n1839,
    n442
  );


  buf
  g1171
  (
    n2164,
    n342
  );


  buf
  g1172
  (
    n1319,
    n457
  );


  not
  g1173
  (
    n1903,
    n533
  );


  buf
  g1174
  (
    n1901,
    n513
  );


  buf
  g1175
  (
    n1936,
    n358
  );


  not
  g1176
  (
    n1472,
    n482
  );


  not
  g1177
  (
    n1047,
    n639
  );


  buf
  g1178
  (
    n747,
    n365
  );


  buf
  g1179
  (
    n1426,
    n321
  );


  not
  g1180
  (
    n1655,
    n549
  );


  not
  g1181
  (
    n1530,
    n368
  );


  not
  g1182
  (
    n1372,
    n631
  );


  buf
  g1183
  (
    n1022,
    n397
  );


  buf
  g1184
  (
    n1459,
    n630
  );


  buf
  g1185
  (
    n1835,
    n218
  );


  not
  g1186
  (
    n1810,
    n429
  );


  not
  g1187
  (
    n2196,
    n333
  );


  not
  g1188
  (
    n2055,
    n79
  );


  buf
  g1189
  (
    n1996,
    n518
  );


  not
  g1190
  (
    n1565,
    n658
  );


  buf
  g1191
  (
    n1195,
    n437
  );


  not
  g1192
  (
    n987,
    n543
  );


  buf
  g1193
  (
    n2034,
    n501
  );


  not
  g1194
  (
    n1036,
    n332
  );


  not
  g1195
  (
    n1675,
    n382
  );


  buf
  g1196
  (
    n1679,
    n357
  );


  buf
  g1197
  (
    n884,
    n502
  );


  not
  g1198
  (
    n1614,
    n494
  );


  buf
  g1199
  (
    n1874,
    n349
  );


  buf
  g1200
  (
    n966,
    n598
  );


  not
  g1201
  (
    n1110,
    n508
  );


  buf
  g1202
  (
    n1038,
    n371
  );


  not
  g1203
  (
    n1314,
    n602
  );


  not
  g1204
  (
    n1935,
    n359
  );


  buf
  g1205
  (
    n1185,
    n517
  );


  buf
  g1206
  (
    n834,
    n349
  );


  buf
  g1207
  (
    n1175,
    n625
  );


  not
  g1208
  (
    n1337,
    n676
  );


  buf
  g1209
  (
    n2216,
    n539
  );


  buf
  g1210
  (
    n1590,
    n673
  );


  buf
  g1211
  (
    n1944,
    n610
  );


  buf
  g1212
  (
    n1355,
    n429
  );


  buf
  g1213
  (
    n1913,
    n335
  );


  not
  g1214
  (
    n2237,
    n638
  );


  buf
  g1215
  (
    n2040,
    n580
  );


  buf
  g1216
  (
    n1612,
    n208
  );


  buf
  g1217
  (
    n1685,
    n525
  );


  buf
  g1218
  (
    n1653,
    n517
  );


  buf
  g1219
  (
    n1833,
    n706
  );


  not
  g1220
  (
    n1067,
    n351
  );


  buf
  g1221
  (
    n848,
    n616
  );


  not
  g1222
  (
    n932,
    n490
  );


  buf
  g1223
  (
    n1225,
    n401
  );


  not
  g1224
  (
    n902,
    n677
  );


  buf
  g1225
  (
    n2103,
    n207
  );


  not
  g1226
  (
    n2030,
    n548
  );


  buf
  g1227
  (
    n887,
    n539
  );


  not
  g1228
  (
    n1490,
    n363
  );


  buf
  g1229
  (
    n1604,
    n609
  );


  not
  g1230
  (
    n2239,
    n479
  );


  buf
  g1231
  (
    n1405,
    n656
  );


  not
  g1232
  (
    n2277,
    n633
  );


  buf
  g1233
  (
    n750,
    n426
  );


  buf
  g1234
  (
    n2217,
    n584
  );


  buf
  g1235
  (
    n1017,
    n526
  );


  buf
  g1236
  (
    n2100,
    n644
  );


  buf
  g1237
  (
    n1997,
    n416
  );


  not
  g1238
  (
    n1705,
    n606
  );


  buf
  g1239
  (
    n1534,
    n478
  );


  buf
  g1240
  (
    n1651,
    n344
  );


  buf
  g1241
  (
    n1724,
    n646
  );


  buf
  g1242
  (
    n1453,
    n419
  );


  buf
  g1243
  (
    n1278,
    n653
  );


  buf
  g1244
  (
    n1004,
    n691
  );


  buf
  g1245
  (
    n1134,
    n515
  );


  not
  g1246
  (
    n2220,
    n613
  );


  not
  g1247
  (
    n1322,
    n360
  );


  not
  g1248
  (
    n1645,
    n386
  );


  buf
  g1249
  (
    n2195,
    n657
  );


  not
  g1250
  (
    n1385,
    n323
  );


  buf
  g1251
  (
    n1241,
    n334
  );


  buf
  g1252
  (
    n1188,
    n439
  );


  buf
  g1253
  (
    n1289,
    n528
  );


  not
  g1254
  (
    n1595,
    n395
  );


  buf
  g1255
  (
    n778,
    n617
  );


  buf
  g1256
  (
    n1484,
    n458
  );


  buf
  g1257
  (
    n1238,
    n421
  );


  not
  g1258
  (
    n1621,
    n696
  );


  not
  g1259
  (
    n2017,
    n620
  );


  not
  g1260
  (
    n2012,
    n519
  );


  buf
  g1261
  (
    n1386,
    n479
  );


  buf
  g1262
  (
    n1894,
    n496
  );


  buf
  g1263
  (
    KeyWire_0_14,
    n552
  );


  not
  g1264
  (
    n1598,
    n681
  );


  not
  g1265
  (
    n1331,
    n487
  );


  not
  g1266
  (
    n1291,
    n340
  );


  not
  g1267
  (
    n1299,
    n689
  );


  not
  g1268
  (
    n1591,
    n602
  );


  not
  g1269
  (
    n827,
    n562
  );


  buf
  g1270
  (
    n1693,
    n509
  );


  not
  g1271
  (
    n1804,
    n396
  );


  buf
  g1272
  (
    n1212,
    n511
  );


  buf
  g1273
  (
    n1522,
    n381
  );


  not
  g1274
  (
    n1296,
    n341
  );


  buf
  g1275
  (
    n1469,
    n459
  );


  not
  g1276
  (
    n826,
    n687
  );


  buf
  g1277
  (
    n1193,
    n658
  );


  not
  g1278
  (
    n1684,
    n375
  );


  not
  g1279
  (
    n796,
    n530
  );


  buf
  g1280
  (
    n1786,
    n330
  );


  not
  g1281
  (
    n1876,
    n390
  );


  not
  g1282
  (
    n2145,
    n638
  );


  buf
  g1283
  (
    n948,
    n570
  );


  not
  g1284
  (
    n785,
    n462
  );


  not
  g1285
  (
    n1341,
    n708
  );


  buf
  g1286
  (
    n1610,
    n569
  );


  buf
  g1287
  (
    n1843,
    n632
  );


  not
  g1288
  (
    n1248,
    n622
  );


  not
  g1289
  (
    n1650,
    n649
  );


  not
  g1290
  (
    n1548,
    n711
  );


  buf
  g1291
  (
    n1738,
    n603
  );


  not
  g1292
  (
    n1822,
    n378
  );


  not
  g1293
  (
    n1077,
    n676
  );


  buf
  g1294
  (
    n2247,
    n368
  );


  buf
  g1295
  (
    n2272,
    n405
  );


  not
  g1296
  (
    n831,
    n210
  );


  buf
  g1297
  (
    n1854,
    n684
  );


  buf
  g1298
  (
    n894,
    n443
  );


  not
  g1299
  (
    n1832,
    n440
  );


  buf
  g1300
  (
    n1369,
    n445
  );


  buf
  g1301
  (
    n1294,
    n485
  );


  buf
  g1302
  (
    n1100,
    n703
  );


  buf
  g1303
  (
    n1065,
    n504
  );


  buf
  g1304
  (
    n1984,
    n590
  );


  not
  g1305
  (
    n1583,
    n209
  );


  buf
  g1306
  (
    n2178,
    n568
  );


  not
  g1307
  (
    n1279,
    n491
  );


  buf
  g1308
  (
    n1043,
    n545
  );


  not
  g1309
  (
    n1499,
    n715
  );


  not
  g1310
  (
    n1841,
    n675
  );


  not
  g1311
  (
    n1109,
    n451
  );


  not
  g1312
  (
    n2013,
    n455
  );


  not
  g1313
  (
    n2133,
    n518
  );


  not
  g1314
  (
    n1508,
    n565
  );


  not
  g1315
  (
    n1311,
    n414
  );


  buf
  g1316
  (
    n1012,
    n343
  );


  buf
  g1317
  (
    n723,
    n352
  );


  not
  g1318
  (
    n2004,
    n350
  );


  not
  g1319
  (
    n1097,
    n521
  );


  buf
  g1320
  (
    n2106,
    n628
  );


  not
  g1321
  (
    n1274,
    n565
  );


  buf
  g1322
  (
    n1584,
    n549
  );


  not
  g1323
  (
    n1986,
    n713
  );


  buf
  g1324
  (
    n777,
    n469
  );


  buf
  g1325
  (
    n1293,
    n378
  );


  not
  g1326
  (
    n1878,
    n399
  );


  not
  g1327
  (
    n1697,
    n497
  );


  buf
  g1328
  (
    n1981,
    n216
  );


  not
  g1329
  (
    n1518,
    n405
  );


  buf
  g1330
  (
    n1371,
    n212
  );


  buf
  g1331
  (
    n2112,
    n517
  );


  buf
  g1332
  (
    n783,
    n413
  );


  not
  g1333
  (
    n923,
    n662
  );


  buf
  g1334
  (
    n1648,
    n639
  );


  buf
  g1335
  (
    n2107,
    n338
  );


  not
  g1336
  (
    n1559,
    n319
  );


  buf
  g1337
  (
    n1080,
    n614
  );


  buf
  g1338
  (
    n1968,
    n667
  );


  not
  g1339
  (
    n1334,
    n445
  );


  not
  g1340
  (
    n1252,
    n338
  );


  not
  g1341
  (
    n2001,
    n206
  );


  buf
  g1342
  (
    n1297,
    n584
  );


  not
  g1343
  (
    n1170,
    n364
  );


  not
  g1344
  (
    n855,
    n480
  );


  buf
  g1345
  (
    n2129,
    n614
  );


  not
  g1346
  (
    n2093,
    n348
  );


  not
  g1347
  (
    n1476,
    n376
  );


  buf
  g1348
  (
    n1240,
    n478
  );


  not
  g1349
  (
    n2249,
    n401
  );


  not
  g1350
  (
    n2024,
    n407
  );


  buf
  g1351
  (
    n1418,
    n416
  );


  not
  g1352
  (
    n1287,
    n356
  );


  buf
  g1353
  (
    n1321,
    n593
  );


  buf
  g1354
  (
    n1957,
    n524
  );


  buf
  g1355
  (
    n1926,
    n458
  );


  not
  g1356
  (
    n1000,
    n415
  );


  not
  g1357
  (
    n2043,
    n694
  );


  buf
  g1358
  (
    n2269,
    n322
  );


  buf
  g1359
  (
    n1486,
    n636
  );


  not
  g1360
  (
    n1969,
    n655
  );


  not
  g1361
  (
    n845,
    n659
  );


  not
  g1362
  (
    n1422,
    n689
  );


  buf
  g1363
  (
    n1795,
    n419
  );


  buf
  g1364
  (
    n2131,
    n647
  );


  not
  g1365
  (
    n1288,
    n689
  );


  buf
  g1366
  (
    n937,
    n465
  );


  not
  g1367
  (
    n2109,
    n443
  );


  buf
  g1368
  (
    n2296,
    n435
  );


  not
  g1369
  (
    n1051,
    n386
  );


  not
  g1370
  (
    n1502,
    n434
  );


  not
  g1371
  (
    n860,
    n591
  );


  not
  g1372
  (
    n2207,
    n560
  );


  not
  g1373
  (
    n1654,
    n704
  );


  not
  g1374
  (
    n1112,
    n391
  );


  buf
  g1375
  (
    n1617,
    n467
  );


  buf
  g1376
  (
    n1615,
    n450
  );


  buf
  g1377
  (
    n991,
    n348
  );


  buf
  g1378
  (
    n1095,
    n659
  );


  not
  g1379
  (
    n2188,
    n672
  );


  not
  g1380
  (
    n756,
    n450
  );


  not
  g1381
  (
    n2080,
    n531
  );


  not
  g1382
  (
    n2211,
    n631
  );


  buf
  g1383
  (
    n2007,
    n573
  );


  not
  g1384
  (
    n1435,
    n461
  );


  buf
  g1385
  (
    n1988,
    n656
  );


  buf
  g1386
  (
    n1912,
    n478
  );


  buf
  g1387
  (
    n2243,
    n402
  );


  not
  g1388
  (
    n1013,
    n606
  );


  buf
  g1389
  (
    n1131,
    n391
  );


  buf
  g1390
  (
    n802,
    n487
  );


  buf
  g1391
  (
    n1178,
    n687
  );


  not
  g1392
  (
    n1847,
    n560
  );


  not
  g1393
  (
    n1169,
    n595
  );


  not
  g1394
  (
    n2192,
    n662
  );


  not
  g1395
  (
    n1571,
    n536
  );


  not
  g1396
  (
    n2174,
    n425
  );


  not
  g1397
  (
    n926,
    n462
  );


  buf
  g1398
  (
    n2238,
    n519
  );


  buf
  g1399
  (
    n1430,
    n711
  );


  not
  g1400
  (
    n1640,
    n604
  );


  not
  g1401
  (
    n1572,
    n332
  );


  not
  g1402
  (
    n2261,
    n209
  );


  buf
  g1403
  (
    n1924,
    n643
  );


  not
  g1404
  (
    n955,
    n578
  );


  buf
  g1405
  (
    n945,
    n529
  );


  not
  g1406
  (
    n1317,
    n682
  );


  not
  g1407
  (
    n2132,
    n355
  );


  not
  g1408
  (
    n1911,
    n704
  );


  buf
  g1409
  (
    n2082,
    n420
  );


  not
  g1410
  (
    n1963,
    n531
  );


  not
  g1411
  (
    n767,
    n559
  );


  not
  g1412
  (
    n1005,
    n668
  );


  not
  g1413
  (
    n1992,
    n550
  );


  not
  g1414
  (
    n2172,
    n428
  );


  buf
  g1415
  (
    n867,
    n449
  );


  buf
  g1416
  (
    n1104,
    n464
  );


  not
  g1417
  (
    n1930,
    n448
  );


  buf
  g1418
  (
    n1633,
    n507
  );


  not
  g1419
  (
    n1432,
    n328
  );


  not
  g1420
  (
    n1213,
    n665
  );


  not
  g1421
  (
    n1230,
    n471
  );


  buf
  g1422
  (
    n1096,
    n389
  );


  buf
  g1423
  (
    n1361,
    n532
  );


  buf
  g1424
  (
    n1068,
    n650
  );


  buf
  g1425
  (
    n1956,
    n410
  );


  not
  g1426
  (
    n1537,
    n587
  );


  buf
  g1427
  (
    n1276,
    n553
  );


  not
  g1428
  (
    n2038,
    n489
  );


  buf
  g1429
  (
    n1560,
    n599
  );


  buf
  g1430
  (
    n864,
    n645
  );


  buf
  g1431
  (
    n814,
    n649
  );


  not
  g1432
  (
    n1028,
    n409
  );


  not
  g1433
  (
    n1163,
    n713
  );


  not
  g1434
  (
    n1916,
    n335
  );


  buf
  g1435
  (
    n726,
    n336
  );


  buf
  g1436
  (
    n1744,
    n463
  );


  not
  g1437
  (
    n1728,
    n564
  );


  buf
  g1438
  (
    n2240,
    n611
  );


  buf
  g1439
  (
    n1789,
    n377
  );


  buf
  g1440
  (
    n1972,
    n690
  );


  buf
  g1441
  (
    n1060,
    n537
  );


  buf
  g1442
  (
    n2189,
    n527
  );


  buf
  g1443
  (
    n1979,
    n641
  );


  buf
  g1444
  (
    n1194,
    n700
  );


  not
  g1445
  (
    n2096,
    n657
  );


  not
  g1446
  (
    n2048,
    n574
  );


  not
  g1447
  (
    n2234,
    n554
  );


  not
  g1448
  (
    n1983,
    n605
  );


  buf
  g1449
  (
    n818,
    n416
  );


  buf
  g1450
  (
    n754,
    n712
  );


  not
  g1451
  (
    n752,
    n630
  );


  buf
  g1452
  (
    n1116,
    n700
  );


  not
  g1453
  (
    n2287,
    n449
  );


  buf
  g1454
  (
    n919,
    n630
  );


  not
  g1455
  (
    n2281,
    n492
  );


  not
  g1456
  (
    n1893,
    n392
  );


  not
  g1457
  (
    n2078,
    n349
  );


  not
  g1458
  (
    n1906,
    n409
  );


  not
  g1459
  (
    n1757,
    n577
  );


  buf
  g1460
  (
    n1324,
    n624
  );


  not
  g1461
  (
    n841,
    n366
  );


  not
  g1462
  (
    n1788,
    n211
  );


  not
  g1463
  (
    n956,
    n685
  );


  not
  g1464
  (
    n1255,
    n419
  );


  not
  g1465
  (
    n2067,
    n353
  );


  not
  g1466
  (
    n2253,
    n650
  );


  buf
  g1467
  (
    n2054,
    n211
  );


  buf
  g1468
  (
    n1425,
    n658
  );


  buf
  g1469
  (
    n781,
    n695
  );


  buf
  g1470
  (
    n1562,
    n389
  );


  buf
  g1471
  (
    n770,
    n618
  );


  not
  g1472
  (
    n1070,
    n659
  );


  not
  g1473
  (
    n1960,
    n386
  );


  buf
  g1474
  (
    KeyWire_0_3,
    n709
  );


  not
  g1475
  (
    n892,
    n661
  );


  not
  g1476
  (
    n2273,
    n325
  );


  not
  g1477
  (
    n971,
    n701
  );


  not
  g1478
  (
    n1955,
    n558
  );


  buf
  g1479
  (
    n811,
    n715
  );


  buf
  g1480
  (
    n1191,
    n620
  );


  not
  g1481
  (
    n1306,
    n345
  );


  not
  g1482
  (
    n1392,
    n521
  );


  not
  g1483
  (
    n978,
    n346
  );


  buf
  g1484
  (
    n1552,
    n334
  );


  not
  g1485
  (
    n1465,
    n436
  );


  buf
  g1486
  (
    n779,
    n396
  );


  buf
  g1487
  (
    n979,
    n329
  );


  buf
  g1488
  (
    n1452,
    n655
  );


  buf
  g1489
  (
    n1647,
    n482
  );


  not
  g1490
  (
    n1759,
    n431
  );


  buf
  g1491
  (
    n1505,
    n566
  );


  buf
  g1492
  (
    n797,
    n710
  );


  not
  g1493
  (
    n1725,
    n535
  );


  buf
  g1494
  (
    n969,
    n388
  );


  buf
  g1495
  (
    n1269,
    n647
  );


  buf
  g1496
  (
    n735,
    n709
  );


  not
  g1497
  (
    n2008,
    n637
  );


  not
  g1498
  (
    n1021,
    n464
  );


  not
  g1499
  (
    n967,
    n543
  );


  not
  g1500
  (
    n1061,
    n558
  );


  not
  g1501
  (
    n891,
    n601
  );


  buf
  g1502
  (
    n2218,
    n536
  );


  not
  g1503
  (
    n2246,
    n710
  );


  buf
  g1504
  (
    n938,
    n657
  );


  buf
  g1505
  (
    n1466,
    n575
  );


  buf
  g1506
  (
    n1732,
    n680
  );


  buf
  g1507
  (
    n933,
    n583
  );


  buf
  g1508
  (
    n1281,
    n378
  );


  buf
  g1509
  (
    n1689,
    n562
  );


  not
  g1510
  (
    n1141,
    n480
  );


  not
  g1511
  (
    n2219,
    n392
  );


  not
  g1512
  (
    n851,
    n361
  );


  not
  g1513
  (
    n2290,
    n713
  );


  not
  g1514
  (
    n1487,
    n416
  );


  not
  g1515
  (
    n1108,
    n378
  );


  not
  g1516
  (
    n1087,
    n481
  );


  buf
  g1517
  (
    n1042,
    n560
  );


  not
  g1518
  (
    n828,
    n653
  );


  buf
  g1519
  (
    n1784,
    n533
  );


  not
  g1520
  (
    n1468,
    n464
  );


  buf
  g1521
  (
    n1347,
    n583
  );


  buf
  g1522
  (
    n883,
    n358
  );


  not
  g1523
  (
    n875,
    n475
  );


  not
  g1524
  (
    n1998,
    n456
  );


  not
  g1525
  (
    n1152,
    n618
  );


  not
  g1526
  (
    n1991,
    n339
  );


  not
  g1527
  (
    n1217,
    n332
  );


  buf
  g1528
  (
    n813,
    n355
  );


  buf
  g1529
  (
    n1262,
    n708
  );


  buf
  g1530
  (
    n2026,
    n450
  );


  not
  g1531
  (
    n1401,
    n437
  );


  buf
  g1532
  (
    n1478,
    n204
  );


  buf
  g1533
  (
    n2267,
    n631
  );


  not
  g1534
  (
    n1073,
    n455
  );


  buf
  g1535
  (
    n1233,
    n566
  );


  buf
  g1536
  (
    n1138,
    n654
  );


  buf
  g1537
  (
    n1206,
    n561
  );


  buf
  g1538
  (
    n1664,
    n458
  );


  not
  g1539
  (
    n1605,
    n406
  );


  buf
  g1540
  (
    n1569,
    n684
  );


  not
  g1541
  (
    n1862,
    n610
  );


  not
  g1542
  (
    n1030,
    n705
  );


  not
  g1543
  (
    n1519,
    n638
  );


  buf
  g1544
  (
    n1277,
    n344
  );


  not
  g1545
  (
    n1162,
    n579
  );


  buf
  g1546
  (
    n1227,
    n382
  );


  not
  g1547
  (
    n1351,
    n537
  );


  not
  g1548
  (
    n1284,
    n487
  );


  buf
  g1549
  (
    n2228,
    n495
  );


  not
  g1550
  (
    n913,
    n522
  );


  not
  g1551
  (
    n1740,
    n644
  );


  not
  g1552
  (
    n1837,
    n333
  );


  buf
  g1553
  (
    n1514,
    n333
  );


  not
  g1554
  (
    n1285,
    n503
  );


  buf
  g1555
  (
    n930,
    n369
  );


  not
  g1556
  (
    n1920,
    n595
  );


  buf
  g1557
  (
    n1115,
    n622
  );


  not
  g1558
  (
    n1450,
    n453
  );


  not
  g1559
  (
    n2198,
    n612
  );


  not
  g1560
  (
    n1125,
    n321
  );


  not
  g1561
  (
    n1302,
    n609
  );


  buf
  g1562
  (
    n1754,
    n421
  );


  buf
  g1563
  (
    n2230,
    n367
  );


  buf
  g1564
  (
    n1447,
    n417
  );


  buf
  g1565
  (
    n2015,
    n462
  );


  not
  g1566
  (
    n2064,
    n391
  );


  not
  g1567
  (
    n806,
    n633
  );


  not
  g1568
  (
    n1056,
    n385
  );


  buf
  g1569
  (
    n1626,
    n205
  );


  buf
  g1570
  (
    n1290,
    n522
  );


  buf
  g1571
  (
    n2051,
    n706
  );


  buf
  g1572
  (
    n1475,
    n582
  );


  buf
  g1573
  (
    n2016,
    n438
  );


  buf
  g1574
  (
    n2229,
    n393
  );


  not
  g1575
  (
    n950,
    n671
  );


  not
  g1576
  (
    n1755,
    n654
  );


  not
  g1577
  (
    n1624,
    n682
  );


  not
  g1578
  (
    n1904,
    n488
  );


  buf
  g1579
  (
    n1727,
    n664
  );


  not
  g1580
  (
    n1575,
    n357
  );


  buf
  g1581
  (
    n1246,
    n677
  );


  buf
  g1582
  (
    n1938,
    n526
  );


  buf
  g1583
  (
    n1411,
    n600
  );


  buf
  g1584
  (
    n1868,
    n351
  );


  not
  g1585
  (
    n1174,
    n332
  );


  buf
  g1586
  (
    n1708,
    n590
  );


  buf
  g1587
  (
    n1157,
    n686
  );


  not
  g1588
  (
    n1639,
    n481
  );


  buf
  g1589
  (
    n825,
    n369
  );


  not
  g1590
  (
    n992,
    n448
  );


  not
  g1591
  (
    n1388,
    n705
  );


  buf
  g1592
  (
    n1316,
    n513
  );


  buf
  g1593
  (
    n2028,
    n396
  );


  not
  g1594
  (
    n1454,
    n443
  );


  not
  g1595
  (
    n1540,
    n363
  );


  buf
  g1596
  (
    n1646,
    n590
  );


  not
  g1597
  (
    n1809,
    n347
  );


  buf
  g1598
  (
    n1414,
    n340
  );


  buf
  g1599
  (
    n1850,
    n675
  );


  not
  g1600
  (
    n1187,
    n707
  );


  buf
  g1601
  (
    n1470,
    n621
  );


  buf
  g1602
  (
    n1137,
    n606
  );


  not
  g1603
  (
    n1456,
    n509
  );


  not
  g1604
  (
    n1075,
    n453
  );


  not
  g1605
  (
    n1016,
    n203
  );


  buf
  g1606
  (
    n2068,
    n331
  );


  buf
  g1607
  (
    n914,
    n351
  );


  not
  g1608
  (
    n898,
    n483
  );


  not
  g1609
  (
    n1766,
    n392
  );


  not
  g1610
  (
    n1283,
    n205
  );


  buf
  g1611
  (
    n871,
    n433
  );


  buf
  g1612
  (
    n745,
    n608
  );


  buf
  g1613
  (
    n865,
    n408
  );


  buf
  g1614
  (
    n1556,
    n399
  );


  not
  g1615
  (
    n2163,
    n368
  );


  buf
  g1616
  (
    n1209,
    n597
  );


  buf
  g1617
  (
    n1323,
    n501
  );


  not
  g1618
  (
    n1587,
    n500
  );


  buf
  g1619
  (
    n896,
    n613
  );


  not
  g1620
  (
    n1631,
    n523
  );


  not
  g1621
  (
    n2069,
    n331
  );


  not
  g1622
  (
    n1668,
    n216
  );


  not
  g1623
  (
    n1445,
    n211
  );


  buf
  g1624
  (
    n921,
    n632
  );


  buf
  g1625
  (
    n2278,
    n407
  );


  buf
  g1626
  (
    n1471,
    n401
  );


  not
  g1627
  (
    n729,
    n635
  );


  not
  g1628
  (
    n1872,
    n589
  );


  not
  g1629
  (
    n1905,
    n361
  );


  buf
  g1630
  (
    n1239,
    n333
  );


  buf
  g1631
  (
    n2025,
    n383
  );


  not
  g1632
  (
    n927,
    n440
  );


  buf
  g1633
  (
    n2126,
    n326
  );


  not
  g1634
  (
    n959,
    n213
  );


  not
  g1635
  (
    n1039,
    n369
  );


  not
  g1636
  (
    n792,
    n204
  );


  not
  g1637
  (
    n2271,
    n402
  );


  buf
  g1638
  (
    n1606,
    n641
  );


  buf
  g1639
  (
    n1781,
    n403
  );


  buf
  g1640
  (
    n1719,
    n440
  );


  not
  g1641
  (
    n1008,
    n470
  );


  buf
  g1642
  (
    n1937,
    n382
  );


  not
  g1643
  (
    n1416,
    n579
  );


  not
  g1644
  (
    n2020,
    n476
  );


  buf
  g1645
  (
    n1360,
    n380
  );


  buf
  g1646
  (
    n1181,
    n588
  );


  buf
  g1647
  (
    n1033,
    n658
  );


  not
  g1648
  (
    n1352,
    n463
  );


  buf
  g1649
  (
    n1967,
    n545
  );


  buf
  g1650
  (
    n1406,
    n503
  );


  not
  g1651
  (
    n1573,
    n400
  );


  not
  g1652
  (
    n2208,
    n510
  );


  buf
  g1653
  (
    n1320,
    n437
  );


  not
  g1654
  (
    n760,
    n319
  );


  not
  g1655
  (
    n1330,
    n520
  );


  not
  g1656
  (
    n2226,
    n661
  );


  buf
  g1657
  (
    n2286,
    n365
  );


  not
  g1658
  (
    n1053,
    n702
  );


  buf
  g1659
  (
    n1536,
    n468
  );


  not
  g1660
  (
    n2260,
    n592
  );


  not
  g1661
  (
    n727,
    n704
  );


  buf
  g1662
  (
    n1340,
    n377
  );


  not
  g1663
  (
    n1069,
    n504
  );


  buf
  g1664
  (
    n2115,
    n629
  );


  not
  g1665
  (
    n1497,
    n379
  );


  not
  g1666
  (
    n1567,
    n615
  );


  not
  g1667
  (
    n722,
    n712
  );


  buf
  g1668
  (
    n1687,
    n660
  );


  not
  g1669
  (
    n816,
    n698
  );


  not
  g1670
  (
    n1706,
    n584
  );


  not
  g1671
  (
    n766,
    n577
  );


  not
  g1672
  (
    n2036,
    n671
  );


  not
  g1673
  (
    n2248,
    n446
  );


  not
  g1674
  (
    n1007,
    n668
  );


  buf
  g1675
  (
    n2284,
    n445
  );


  buf
  g1676
  (
    n1403,
    n581
  );


  buf
  g1677
  (
    n1851,
    n459
  );


  not
  g1678
  (
    n2116,
    n343
  );


  not
  g1679
  (
    n947,
    n439
  );


  buf
  g1680
  (
    n1354,
    n383
  );


  not
  g1681
  (
    n1050,
    n662
  );


  buf
  g1682
  (
    n2099,
    n327
  );


  buf
  g1683
  (
    n1026,
    n623
  );


  buf
  g1684
  (
    n2236,
    n487
  );


  buf
  g1685
  (
    n1966,
    n395
  );


  buf
  g1686
  (
    n1329,
    n693
  );


  buf
  g1687
  (
    n789,
    n336
  );


  not
  g1688
  (
    n1010,
    n612
  );


  not
  g1689
  (
    n2146,
    n712
  );


  buf
  g1690
  (
    n751,
    n375
  );


  buf
  g1691
  (
    n2197,
    n650
  );


  buf
  g1692
  (
    n1482,
    n446
  );


  buf
  g1693
  (
    n1254,
    n526
  );


  not
  g1694
  (
    n877,
    n505
  );


  not
  g1695
  (
    n1855,
    n209
  );


  not
  g1696
  (
    n2245,
    n327
  );


  buf
  g1697
  (
    n1778,
    n549
  );


  not
  g1698
  (
    n1644,
    n561
  );


  not
  g1699
  (
    n801,
    n695
  );


  buf
  g1700
  (
    n1541,
    n525
  );


  buf
  g1701
  (
    n2105,
    n428
  );


  buf
  g1702
  (
    n1243,
    n545
  );


  buf
  g1703
  (
    n1709,
    n673
  );


  buf
  g1704
  (
    n1715,
    n663
  );


  not
  g1705
  (
    n1349,
    n586
  );


  not
  g1706
  (
    n794,
    n319
  );


  not
  g1707
  (
    n836,
    n568
  );


  buf
  g1708
  (
    n2268,
    n533
  );


  not
  g1709
  (
    n1780,
    n635
  );


  not
  g1710
  (
    n1124,
    n430
  );


  buf
  g1711
  (
    n872,
    n701
  );


  buf
  g1712
  (
    n1686,
    n544
  );


  not
  g1713
  (
    n1914,
    n643
  );


  buf
  g1714
  (
    n1861,
    n604
  );


  not
  g1715
  (
    n1177,
    n584
  );


  buf
  g1716
  (
    n2244,
    n660
  );


  buf
  g1717
  (
    n2276,
    n593
  );


  not
  g1718
  (
    n847,
    n433
  );


  not
  g1719
  (
    n837,
    n471
  );


  not
  g1720
  (
    n1785,
    n605
  );


  buf
  g1721
  (
    n1623,
    n204
  );


  not
  g1722
  (
    n1247,
    n632
  );


  not
  g1723
  (
    n1674,
    n572
  );


  buf
  g1724
  (
    n2033,
    n524
  );


  buf
  g1725
  (
    n1064,
    n618
  );


  buf
  g1726
  (
    n1895,
    n708
  );


  buf
  g1727
  (
    n1762,
    n474
  );


  buf
  g1728
  (
    n1019,
    n328
  );


  not
  g1729
  (
    n774,
    n471
  );


  buf
  g1730
  (
    n2075,
    n481
  );


  buf
  g1731
  (
    n858,
    n645
  );


  not
  g1732
  (
    n1229,
    n576
  );


  buf
  g1733
  (
    n1018,
    n681
  );


  buf
  g1734
  (
    n1267,
    n479
  );


  buf
  g1735
  (
    n2298,
    n477
  );


  buf
  g1736
  (
    n1120,
    n516
  );


  not
  g1737
  (
    n2202,
    n513
  );


  not
  g1738
  (
    n899,
    n535
  );


  buf
  g1739
  (
    n1761,
    n518
  );


  not
  g1740
  (
    n1897,
    n541
  );


  not
  g1741
  (
    n2297,
    n324
  );


  not
  g1742
  (
    n2124,
    n469
  );


  not
  g1743
  (
    n1029,
    n394
  );


  buf
  g1744
  (
    n782,
    n636
  );


  not
  g1745
  (
    n1774,
    n627
  );


  not
  g1746
  (
    n1827,
    n674
  );


  buf
  g1747
  (
    n1237,
    n397
  );


  buf
  g1748
  (
    n1630,
    n610
  );


  not
  g1749
  (
    n965,
    n375
  );


  not
  g1750
  (
    n2203,
    n326
  );


  buf
  g1751
  (
    n1683,
    n389
  );


  not
  g1752
  (
    n1353,
    n694
  );


  not
  g1753
  (
    n1344,
    n586
  );


  buf
  g1754
  (
    n985,
    n367
  );


  buf
  g1755
  (
    n1836,
    n365
  );


  not
  g1756
  (
    n951,
    n532
  );


  buf
  g1757
  (
    n790,
    n575
  );


  not
  g1758
  (
    n1049,
    n458
  );


  not
  g1759
  (
    n1511,
    n637
  );


  not
  g1760
  (
    n1994,
    n414
  );


  buf
  g1761
  (
    n2127,
    n422
  );


  not
  g1762
  (
    n1180,
    n338
  );


  buf
  g1763
  (
    n1136,
    n547
  );


  not
  g1764
  (
    n1232,
    n598
  );


  not
  g1765
  (
    n1747,
    n406
  );


  buf
  g1766
  (
    n742,
    n546
  );


  buf
  g1767
  (
    n1823,
    n353
  );


  buf
  g1768
  (
    n1806,
    n548
  );


  not
  g1769
  (
    n1186,
    n594
  );


  buf
  g1770
  (
    n897,
    n664
  );


  buf
  g1771
  (
    n1625,
    n380
  );


  not
  g1772
  (
    n1024,
    n558
  );


  not
  g1773
  (
    n1044,
    n385
  );


  buf
  g1774
  (
    n2160,
    n376
  );


  buf
  g1775
  (
    n2187,
    n203
  );


  not
  g1776
  (
    n1040,
    n685
  );


  buf
  g1777
  (
    n1628,
    n530
  );


  not
  g1778
  (
    n2232,
    n527
  );


  buf
  g1779
  (
    n1887,
    n360
  );


  buf
  g1780
  (
    n2091,
    n662
  );


  not
  g1781
  (
    n1973,
    n522
  );


  buf
  g1782
  (
    n1158,
    n478
  );


  not
  g1783
  (
    n1945,
    n536
  );


  not
  g1784
  (
    n2283,
    n538
  );


  not
  g1785
  (
    n1273,
    n476
  );


  not
  g1786
  (
    n795,
    n398
  );


  not
  g1787
  (
    n823,
    n668
  );


  not
  g1788
  (
    n981,
    n218
  );


  not
  g1789
  (
    n1009,
    n567
  );


  not
  g1790
  (
    n1739,
    n667
  );


  not
  g1791
  (
    n1649,
    n548
  );


  buf
  g1792
  (
    n2092,
    n370
  );


  not
  g1793
  (
    n1122,
    n604
  );


  not
  g1794
  (
    n931,
    n356
  );


  not
  g1795
  (
    n2193,
    n405
  );


  buf
  g1796
  (
    n2168,
    n544
  );


  buf
  g1797
  (
    n753,
    n216
  );


  not
  g1798
  (
    n1517,
    n339
  );


  not
  g1799
  (
    n1183,
    n357
  );


  not
  g1800
  (
    n2142,
    n647
  );


  buf
  g1801
  (
    n2177,
    n678
  );


  buf
  g1802
  (
    n1350,
    n563
  );


  buf
  g1803
  (
    n1348,
    n384
  );


  not
  g1804
  (
    n873,
    n680
  );


  buf
  g1805
  (
    KeyWire_0_13,
    n539
  );


  not
  g1806
  (
    n922,
    n371
  );


  buf
  g1807
  (
    n1959,
    n525
  );


  buf
  g1808
  (
    n2011,
    n421
  );


  buf
  g1809
  (
    n2031,
    n413
  );


  buf
  g1810
  (
    n988,
    n214
  );


  buf
  g1811
  (
    n1528,
    n712
  );


  buf
  g1812
  (
    n1942,
    n586
  );


  buf
  g1813
  (
    n1656,
    n347
  );


  not
  g1814
  (
    n1859,
    n205
  );


  not
  g1815
  (
    n1611,
    n402
  );


  not
  g1816
  (
    n977,
    n493
  );


  not
  g1817
  (
    n1387,
    n577
  );


  not
  g1818
  (
    n878,
    n636
  );


  not
  g1819
  (
    n2153,
    n601
  );


  buf
  g1820
  (
    n1308,
    n602
  );


  not
  g1821
  (
    n1041,
    n714
  );


  buf
  g1822
  (
    n908,
    n384
  );


  not
  g1823
  (
    n2117,
    n485
  );


  buf
  g1824
  (
    n2299,
    n444
  );


  not
  g1825
  (
    n1557,
    n705
  );


  not
  g1826
  (
    n993,
    n561
  );


  not
  g1827
  (
    n1282,
    n682
  );


  not
  g1828
  (
    n974,
    n217
  );


  buf
  g1829
  (
    n1415,
    n628
  );


  buf
  g1830
  (
    n1792,
    n671
  );


  buf
  g1831
  (
    n2130,
    n398
  );


  buf
  g1832
  (
    n1114,
    n437
  );


  not
  g1833
  (
    n1730,
    n626
  );


  not
  g1834
  (
    n1563,
    n448
  );


  buf
  g1835
  (
    n2200,
    n362
  );


  not
  g1836
  (
    n1489,
    n451
  );


  not
  g1837
  (
    n2014,
    n514
  );


  buf
  g1838
  (
    n2227,
    n715
  );


  buf
  g1839
  (
    n1149,
    n625
  );


  buf
  g1840
  (
    n1848,
    n617
  );


  buf
  g1841
  (
    n1113,
    n373
  );


  buf
  g1842
  (
    n744,
    n342
  );


  not
  g1843
  (
    n1153,
    n677
  );


  not
  g1844
  (
    n1062,
    n626
  );


  buf
  g1845
  (
    n1365,
    n453
  );


  not
  g1846
  (
    n1756,
    n403
  );


  not
  g1847
  (
    n1444,
    n597
  );


  buf
  g1848
  (
    KeyWire_0_29,
    n320
  );


  buf
  g1849
  (
    n1409,
    n679
  );


  buf
  g1850
  (
    n1953,
    n473
  );


  buf
  g1851
  (
    n1820,
    n515
  );


  buf
  g1852
  (
    n1260,
    n542
  );


  not
  g1853
  (
    n822,
    n473
  );


  not
  g1854
  (
    n1159,
    n587
  );


  buf
  g1855
  (
    n1698,
    n502
  );


  not
  g1856
  (
    n1526,
    n706
  );


  not
  g1857
  (
    n1568,
    n692
  );


  buf
  g1858
  (
    n1993,
    n540
  );


  buf
  g1859
  (
    n2165,
    n353
  );


  buf
  g1860
  (
    n1544,
    n670
  );


  buf
  g1861
  (
    n1772,
    n578
  );


  not
  g1862
  (
    n857,
    n517
  );


  not
  g1863
  (
    n2079,
    n347
  );


  buf
  g1864
  (
    n1714,
    n663
  );


  not
  g1865
  (
    n1397,
    n428
  );


  buf
  g1866
  (
    n1111,
    n635
  );


  not
  g1867
  (
    n2050,
    n601
  );


  buf
  g1868
  (
    n1691,
    n348
  );


  not
  g1869
  (
    n1336,
    n417
  );


  buf
  g1870
  (
    n1717,
    n626
  );


  not
  g1871
  (
    n2118,
    n208
  );


  buf
  g1872
  (
    n1776,
    n433
  );


  buf
  g1873
  (
    n1084,
    n534
  );


  buf
  g1874
  (
    n821,
    n358
  );


  not
  g1875
  (
    n1168,
    n441
  );


  buf
  g1876
  (
    n1048,
    n387
  );


  buf
  g1877
  (
    n2071,
    n599
  );


  not
  g1878
  (
    n1989,
    n648
  );


  not
  g1879
  (
    n1748,
    n660
  );


  buf
  g1880
  (
    n1491,
    n614
  );


  not
  g1881
  (
    n1588,
    n714
  );


  not
  g1882
  (
    n918,
    n585
  );


  buf
  g1883
  (
    n2111,
    n555
  );


  not
  g1884
  (
    n1860,
    n448
  );


  not
  g1885
  (
    n1464,
    n681
  );


  buf
  g1886
  (
    n755,
    n370
  );


  not
  g1887
  (
    n748,
    n207
  );


  buf
  g1888
  (
    n1867,
    n596
  );


  buf
  g1889
  (
    n1458,
    n476
  );


  not
  g1890
  (
    n1207,
    n547
  );


  not
  g1891
  (
    n1819,
    n425
  );


  buf
  g1892
  (
    n952,
    n350
  );


  not
  g1893
  (
    n1046,
    n206
  );


  buf
  g1894
  (
    n2300,
    n494
  );


  buf
  g1895
  (
    n1678,
    n655
  );


  not
  g1896
  (
    n1086,
    n540
  );


  not
  g1897
  (
    n1555,
    n336
  );


  buf
  g1898
  (
    n1001,
    n660
  );


  not
  g1899
  (
    n1831,
    n490
  );


  not
  g1900
  (
    n1710,
    n347
  );


  not
  g1901
  (
    n1629,
    n452
  );


  not
  g1902
  (
    n1085,
    n648
  );


  buf
  g1903
  (
    n734,
    n389
  );


  buf
  g1904
  (
    n1034,
    n322
  );


  buf
  g1905
  (
    n903,
    n600
  );


  buf
  g1906
  (
    n2155,
    n498
  );


  not
  g1907
  (
    n2173,
    n506
  );


  not
  g1908
  (
    n1940,
    n390
  );


  buf
  g1909
  (
    n1167,
    n593
  );


  not
  g1910
  (
    n968,
    n505
  );


  not
  g1911
  (
    n2266,
    n503
  );


  not
  g1912
  (
    n2166,
    n431
  );


  buf
  g1913
  (
    n793,
    n323
  );


  buf
  g1914
  (
    n1919,
    n697
  );


  buf
  g1915
  (
    n2057,
    n423
  );


  not
  g1916
  (
    n910,
    n211
  );


  buf
  g1917
  (
    n1692,
    n486
  );


  buf
  g1918
  (
    n1264,
    n528
  );


  buf
  g1919
  (
    n1793,
    n477
  );


  buf
  g1920
  (
    n895,
    n621
  );


  buf
  g1921
  (
    n1844,
    n562
  );


  buf
  g1922
  (
    n1665,
    n670
  );


  buf
  g1923
  (
    n1151,
    n364
  );


  not
  g1924
  (
    n890,
    n619
  );


  buf
  g1925
  (
    n1419,
    n522
  );


  buf
  g1926
  (
    n1381,
    n218
  );


  not
  g1927
  (
    n810,
    n536
  );


  not
  g1928
  (
    n1481,
    n432
  );


  not
  g1929
  (
    n1731,
    n699
  );


  buf
  g1930
  (
    n2255,
    n351
  );


  not
  g1931
  (
    n2241,
    n446
  );


  buf
  g1932
  (
    n2157,
    n610
  );


  not
  g1933
  (
    n2225,
    n557
  );


  buf
  g1934
  (
    n1272,
    n624
  );


  not
  g1935
  (
    n1771,
    n459
  );


  not
  g1936
  (
    n1032,
    n209
  );


  not
  g1937
  (
    n1949,
    n363
  );


  not
  g1938
  (
    n2291,
    n648
  );


  not
  g1939
  (
    n1123,
    n457
  );


  not
  g1940
  (
    n1749,
    n352
  );


  buf
  g1941
  (
    n1333,
    n614
  );


  not
  g1942
  (
    n2285,
    n420
  );


  not
  g1943
  (
    n2212,
    n352
  );


  buf
  g1944
  (
    n1037,
    n486
  );


  not
  g1945
  (
    n1164,
    n424
  );


  buf
  g1946
  (
    n1922,
    n683
  );


  buf
  g1947
  (
    n1121,
    n711
  );


  not
  g1948
  (
    n2022,
    n509
  );


  buf
  g1949
  (
    n2223,
    n588
  );


  not
  g1950
  (
    n1798,
    n399
  );


  not
  g1951
  (
    n1431,
    n438
  );


  buf
  g1952
  (
    n1622,
    n364
  );


  buf
  g1953
  (
    n1582,
    n642
  );


  buf
  g1954
  (
    n1396,
    n521
  );


  not
  g1955
  (
    n2044,
    n637
  );


  buf
  g1956
  (
    n1561,
    n570
  );


  not
  g1957
  (
    n2214,
    n663
  );


  buf
  g1958
  (
    n859,
    n581
  );


  not
  g1959
  (
    n880,
    n495
  );


  not
  g1960
  (
    n2074,
    n407
  );


  buf
  g1961
  (
    n893,
    n539
  );


  buf
  g1962
  (
    n1383,
    n676
  );


  not
  g1963
  (
    n1680,
    n688
  );


  buf
  g1964
  (
    n2184,
    n707
  );


  buf
  g1965
  (
    n1434,
    n691
  );


  buf
  g1966
  (
    n1594,
    n709
  );


  buf
  g1967
  (
    n1166,
    n394
  );


  not
  g1968
  (
    n758,
    n338
  );


  not
  g1969
  (
    n2085,
    n474
  );


  buf
  g1970
  (
    n1270,
    n329
  );


  not
  g1971
  (
    n1443,
    n498
  );


  not
  g1972
  (
    n2140,
    n510
  );


  not
  g1973
  (
    n862,
    n542
  );


  not
  g1974
  (
    n1132,
    n380
  );


  buf
  g1975
  (
    n1620,
    n472
  );


  buf
  g1976
  (
    n736,
    n385
  );


  not
  g1977
  (
    n1990,
    n422
  );


  buf
  g1978
  (
    n1128,
    n217
  );


  buf
  g1979
  (
    n2065,
    n591
  );


  not
  g1980
  (
    n868,
    n430
  );


  not
  g1981
  (
    n1576,
    n483
  );


  not
  g1982
  (
    n941,
    n615
  );


  buf
  g1983
  (
    n1616,
    n327
  );


  not
  g1984
  (
    n1130,
    n392
  );


  not
  g1985
  (
    n743,
    n506
  );


  buf
  g1986
  (
    n805,
    n464
  );


  buf
  g1987
  (
    n1265,
    n515
  );


  buf
  g1988
  (
    n1231,
    n572
  );


  not
  g1989
  (
    n1721,
    n387
  );


  not
  g1990
  (
    n1652,
    n453
  );


  not
  g1991
  (
    n1176,
    n373
  );


  buf
  g1992
  (
    n1356,
    n619
  );


  buf
  g1993
  (
    n2235,
    n629
  );


  not
  g1994
  (
    n763,
    n547
  );


  not
  g1995
  (
    n907,
    n482
  );


  not
  g1996
  (
    n1539,
    n427
  );


  buf
  g1997
  (
    n1985,
    n457
  );


  buf
  g1998
  (
    n2089,
    n397
  );


  not
  g1999
  (
    n986,
    n511
  );


  not
  g2000
  (
    n1242,
    n326
  );


  not
  g2001
  (
    n889,
    n675
  );


  buf
  g2002
  (
    n2114,
    n346
  );


  buf
  g2003
  (
    n1326,
    n600
  );


  not
  g2004
  (
    n846,
    n430
  );


  not
  g2005
  (
    n1663,
    n556
  );


  buf
  g2006
  (
    n2289,
    n329
  );


  buf
  g2007
  (
    n1408,
    n343
  );


  buf
  g2008
  (
    n2204,
    n376
  );


  not
  g2009
  (
    n1763,
    n466
  );


  buf
  g2010
  (
    n1535,
    n493
  );


  not
  g2011
  (
    n1570,
    n210
  );


  not
  g2012
  (
    n1787,
    n360
  );


  buf
  g2013
  (
    n2274,
    n651
  );


  not
  g2014
  (
    n815,
    n355
  );


  buf
  g2015
  (
    n1753,
    n664
  );


  buf
  g2016
  (
    n1580,
    n411
  );


  buf
  g2017
  (
    n2242,
    n565
  );


  buf
  g2018
  (
    n1449,
    n694
  );


  not
  g2019
  (
    n1928,
    n359
  );


  not
  g2020
  (
    n1506,
    n700
  );


  buf
  g2021
  (
    n1139,
    n426
  );


  buf
  g2022
  (
    n1885,
    n354
  );


  buf
  g2023
  (
    n2180,
    n330
  );


  not
  g2024
  (
    n2270,
    n344
  );


  not
  g2025
  (
    n787,
    n540
  );


  buf
  g2026
  (
    n1918,
    n640
  );


  buf
  g2027
  (
    n885,
    n665
  );


  not
  g2028
  (
    n957,
    n210
  );


  not
  g2029
  (
    n1886,
    n633
  );


  buf
  g2030
  (
    n819,
    n545
  );


  buf
  g2031
  (
    KeyWire_0_16,
    n495
  );


  buf
  g2032
  (
    n780,
    n681
  );


  buf
  g2033
  (
    n1342,
    n640
  );


  not
  g2034
  (
    n1769,
    n404
  );


  not
  g2035
  (
    n1751,
    n456
  );


  buf
  g2036
  (
    n800,
    n532
  );


  not
  g2037
  (
    n1627,
    n498
  );


  buf
  g2038
  (
    n924,
    n651
  );


  not
  g2039
  (
    n788,
    n580
  );


  buf
  g2040
  (
    n2144,
    n374
  );


  not
  g2041
  (
    n1513,
    n469
  );


  not
  g2042
  (
    n1516,
    n491
  );


  buf
  g2043
  (
    n1554,
    n466
  );


  buf
  g2044
  (
    n1441,
    n684
  );


  not
  g2045
  (
    n2194,
    n683
  );


  buf
  g2046
  (
    n2175,
    n635
  );


  not
  g2047
  (
    n1581,
    n325
  );


  buf
  g2048
  (
    KeyWire_0_17,
    n685
  );


  not
  g2049
  (
    n764,
    n641
  );


  not
  g2050
  (
    n1729,
    n708
  );


  buf
  g2051
  (
    n1577,
    n569
  );


  buf
  g2052
  (
    n1440,
    n633
  );


  buf
  g2053
  (
    n982,
    n341
  );


  buf
  g2054
  (
    n2181,
    n431
  );


  buf
  g2055
  (
    n1154,
    n579
  );


  not
  g2056
  (
    n869,
    n549
  );


  buf
  g2057
  (
    n2062,
    n612
  );


  not
  g2058
  (
    n1427,
    n612
  );


  buf
  g2059
  (
    n2250,
    n694
  );


  not
  g2060
  (
    n1768,
    n415
  );


  not
  g2061
  (
    n943,
    n406
  );


  not
  g2062
  (
    n1303,
    n334
  );


  not
  g2063
  (
    n1259,
    n665
  );


  not
  g2064
  (
    n1234,
    n202
  );


  buf
  g2065
  (
    n1474,
    n696
  );


  not
  g2066
  (
    n1545,
    n404
  );


  buf
  g2067
  (
    n1156,
    n590
  );


  buf
  g2068
  (
    n881,
    n429
  );


  not
  g2069
  (
    n2083,
    n208
  );


  not
  g2070
  (
    n1521,
    n216
  );


  buf
  g2071
  (
    n928,
    n472
  );


  buf
  g2072
  (
    n1830,
    n362
  );


  not
  g2073
  (
    n2262,
    n634
  );


  not
  g2074
  (
    n1999,
    n447
  );


  not
  g2075
  (
    n1455,
    n403
  );


  not
  g2076
  (
    n1380,
    n495
  );


  buf
  g2077
  (
    n2254,
    n639
  );


  buf
  g2078
  (
    n1510,
    n400
  );


  buf
  g2079
  (
    n1741,
    n421
  );


  not
  g2080
  (
    n817,
    n690
  );


  not
  g2081
  (
    n1779,
    n484
  );


  not
  g2082
  (
    n2113,
    n431
  );


  not
  g2083
  (
    n1884,
    n512
  );


  not
  g2084
  (
    n1142,
    n368
  );


  buf
  g2085
  (
    n1869,
    n393
  );


  not
  g2086
  (
    n1119,
    n543
  );


  not
  g2087
  (
    n1117,
    n443
  );


  buf
  g2088
  (
    n1699,
    n212
  );


  buf
  g2089
  (
    n1055,
    n372
  );


  not
  g2090
  (
    n1636,
    n454
  );


  buf
  g2091
  (
    n1978,
    n651
  );


  buf
  g2092
  (
    n2233,
    n214
  );


  not
  g2093
  (
    n2032,
    n542
  );


  buf
  g2094
  (
    n879,
    n372
  );


  not
  g2095
  (
    n1201,
    n589
  );


  not
  g2096
  (
    n1845,
    n677
  );


  not
  g2097
  (
    n2104,
    n616
  );


  not
  g2098
  (
    n1593,
    n442
  );


  buf
  g2099
  (
    n2009,
    n562
  );


  not
  g2100
  (
    n1222,
    n706
  );


  not
  g2101
  (
    n912,
    n374
  );


  buf
  g2102
  (
    n1891,
    n707
  );


  buf
  g2103
  (
    n737,
    n600
  );


  not
  g2104
  (
    n2148,
    n372
  );


  buf
  g2105
  (
    n757,
    n500
  );


  not
  g2106
  (
    n1228,
    n616
  );


  not
  g2107
  (
    n1143,
    n548
  );


  not
  g2108
  (
    n1389,
    n412
  );


  buf
  g2109
  (
    n1173,
    n566
  );


  buf
  g2110
  (
    n2206,
    n690
  );


  buf
  g2111
  (
    n953,
    n505
  );


  buf
  g2112
  (
    n724,
    n619
  );


  buf
  g2113
  (
    n1952,
    n402
  );


  buf
  g2114
  (
    n1838,
    n626
  );


  not
  g2115
  (
    n962,
    n203
  );


  not
  g2116
  (
    n2149,
    n710
  );


  buf
  g2117
  (
    n886,
    n465
  );


  buf
  g2118
  (
    n1020,
    n499
  );


  not
  g2119
  (
    n1063,
    n648
  );


  not
  g2120
  (
    n833,
    n330
  );


  buf
  g2121
  (
    n2221,
    n432
  );


  buf
  g2122
  (
    n1071,
    n678
  );


  not
  g2123
  (
    n1429,
    n571
  );


  buf
  g2124
  (
    n1550,
    n363
  );


  not
  g2125
  (
    n2128,
    n492
  );


  not
  g2126
  (
    n946,
    n465
  );


  buf
  g2127
  (
    n1865,
    n551
  );


  not
  g2128
  (
    n2295,
    n362
  );


  not
  g2129
  (
    n1800,
    n400
  );


  not
  g2130
  (
    n2027,
    n555
  );


  not
  g2131
  (
    n2037,
    n595
  );


  not
  g2132
  (
    n1467,
    n414
  );


  not
  g2133
  (
    n1412,
    n422
  );


  buf
  g2134
  (
    n1742,
    n523
  );


  buf
  g2135
  (
    n1006,
    n411
  );


  buf
  g2136
  (
    n1796,
    n215
  );


  buf
  g2137
  (
    n1750,
    n575
  );


  not
  g2138
  (
    n1896,
    n580
  );


  not
  g2139
  (
    n2154,
    n343
  );


  not
  g2140
  (
    n994,
    n669
  );


  buf
  g2141
  (
    n1462,
    n356
  );


  not
  g2142
  (
    n1829,
    n442
  );


  buf
  g2143
  (
    n1716,
    n519
  );


  buf
  g2144
  (
    n1332,
    n394
  );


  buf
  g2145
  (
    n1400,
    n473
  );


  buf
  g2146
  (
    KeyWire_0_0,
    n703
  );


  buf
  g2147
  (
    n861,
    n508
  );


  buf
  g2148
  (
    n1172,
    n563
  );


  not
  g2149
  (
    n1602,
    n651
  );


  not
  g2150
  (
    n936,
    n669
  );


  not
  g2151
  (
    n1090,
    n623
  );


  not
  g2152
  (
    n934,
    n540
  );


  not
  g2153
  (
    n1364,
    n484
  );


  not
  g2154
  (
    n725,
    n381
  );


  not
  g2155
  (
    n1346,
    n438
  );


  not
  g2156
  (
    n1917,
    n579
  );


  buf
  g2157
  (
    n762,
    n322
  );


  buf
  g2158
  (
    n2066,
    n327
  );


  not
  g2159
  (
    n1925,
    n687
  );


  not
  g2160
  (
    n1975,
    n515
  );


  not
  g2161
  (
    n1888,
    n388
  );


  not
  g2162
  (
    n906,
    n387
  );


  buf
  g2163
  (
    n2137,
    n512
  );


  buf
  g2164
  (
    n1214,
    n560
  );


  buf
  g2165
  (
    n1669,
    n440
  );


  not
  g2166
  (
    n2222,
    n572
  );


  buf
  g2167
  (
    KeyWire_0_4,
    n573
  );


  not
  g2168
  (
    n1976,
    n452
  );


  not
  g2169
  (
    n2259,
    n405
  );


  buf
  g2170
  (
    n2006,
    n321
  );


  not
  g2171
  (
    n2102,
    n390
  );


  not
  g2172
  (
    n1923,
    n384
  );


  buf
  g2173
  (
    n1358,
    n426
  );


  buf
  g2174
  (
    n1870,
    n396
  );


  buf
  g2175
  (
    n1266,
    n551
  );


  buf
  g2176
  (
    n1338,
    n507
  );


  not
  g2177
  (
    n1842,
    n516
  );


  not
  g2178
  (
    n1092,
    n571
  );


  not
  g2179
  (
    n1393,
    n408
  );


  buf
  g2180
  (
    n1448,
    n571
  );


  buf
  g2181
  (
    n1736,
    n425
  );


  not
  g2182
  (
    n2215,
    n441
  );


  not
  g2183
  (
    n1011,
    n624
  );


  buf
  g2184
  (
    n1767,
    n530
  );


  not
  g2185
  (
    n1179,
    n435
  );


  not
  g2186
  (
    n1325,
    n528
  );


  not
  g2187
  (
    n728,
    n400
  );


  not
  g2188
  (
    n1315,
    n441
  );


  buf
  g2189
  (
    n1910,
    n459
  );


  buf
  g2190
  (
    n1305,
    n607
  );


  buf
  g2191
  (
    n759,
    n646
  );


  buf
  g2192
  (
    n1072,
    n701
  );


  not
  g2193
  (
    n2282,
    n685
  );


  buf
  g2194
  (
    n853,
    n497
  );


  not
  g2195
  (
    n1527,
    n215
  );


  not
  g2196
  (
    n2169,
    n434
  );


  not
  g2197
  (
    n1103,
    n571
  );


  buf
  g2198
  (
    KeyWire_0_9,
    n410
  );


  buf
  g2199
  (
    n1712,
    n567
  );


  buf
  g2200
  (
    n1707,
    n460
  );


  buf
  g2201
  (
    n942,
    n564
  );


  buf
  g2202
  (
    n1504,
    n218
  );


  not
  g2203
  (
    n1987,
    n323
  );


  buf
  g2204
  (
    n719,
    n380
  );


  buf
  g2205
  (
    n929,
    n622
  );


  buf
  g2206
  (
    n1368,
    n546
  );


  not
  g2207
  (
    n1718,
    n623
  );


  buf
  g2208
  (
    n1642,
    n594
  );


  buf
  g2209
  (
    n1599,
    n474
  );


  not
  g2210
  (
    n2150,
    n574
  );


  buf
  g2211
  (
    n1666,
    n466
  );


  not
  g2212
  (
    n839,
    n379
  );


  not
  g2213
  (
    n963,
    n398
  );


  buf
  g2214
  (
    n1524,
    n550
  );


  not
  g2215
  (
    n808,
    n435
  );


  buf
  g2216
  (
    n1106,
    n640
  );


  not
  g2217
  (
    n1366,
    n424
  );


  not
  g2218
  (
    KeyWire_0_21,
    n556
  );


  not
  g2219
  (
    n2210,
    n552
  );


  buf
  g2220
  (
    n809,
    n605
  );


  not
  g2221
  (
    n2059,
    n455
  );


  not
  g2222
  (
    n2125,
    n597
  );


  not
  g2223
  (
    n1500,
    n420
  );


  not
  g2224
  (
    n1219,
    n461
  );


  buf
  g2225
  (
    n2231,
    n430
  );


  buf
  g2226
  (
    n829,
    n644
  );


  buf
  g2227
  (
    n1014,
    n383
  );


  not
  g2228
  (
    n1603,
    n650
  );


  buf
  g2229
  (
    n1197,
    n622
  );


  buf
  g2230
  (
    n1395,
    n700
  );


  not
  g2231
  (
    n1200,
    n452
  );


  not
  g2232
  (
    n1082,
    n628
  );


  not
  g2233
  (
    n2135,
    n570
  );


  buf
  g2234
  (
    n1268,
    n621
  );


  not
  g2235
  (
    n1074,
    n673
  );


  not
  g2236
  (
    n1078,
    n563
  );


  not
  g2237
  (
    n1025,
    n473
  );


  not
  g2238
  (
    n2156,
    n497
  );


  not
  g2239
  (
    n1275,
    n322
  );


  buf
  g2240
  (
    n1849,
    n491
  );


  not
  g2241
  (
    n1031,
    n607
  );


  buf
  g2242
  (
    n1027,
    n703
  );


  buf
  g2243
  (
    n1529,
    n373
  );


  buf
  g2244
  (
    n1343,
    n529
  );


  not
  g2245
  (
    KeyWire_0_8,
    n652
  );


  not
  g2246
  (
    n1428,
    n591
  );


  not
  g2247
  (
    n1081,
    n664
  );


  buf
  g2248
  (
    n798,
    n460
  );


  buf
  g2249
  (
    n776,
    n394
  );


  buf
  g2250
  (
    n2302,
    n556
  );


  buf
  g2251
  (
    n1318,
    n388
  );


  not
  g2252
  (
    n2158,
    n342
  );


  buf
  g2253
  (
    n1263,
    n330
  );


  not
  g2254
  (
    n1585,
    n715
  );


  not
  g2255
  (
    n1658,
    n702
  );


  not
  g2256
  (
    n1794,
    n433
  );


  buf
  g2257
  (
    n1226,
    n702
  );


  buf
  g2258
  (
    n812,
    n541
  );


  xnor
  g2259
  (
    n1643,
    n417,
    n412,
    n467,
    n346
  );


  nor
  g2260
  (
    n1182,
    n631,
    n680,
    n534,
    n357
  );


  nand
  g2261
  (
    n1995,
    n599,
    n520,
    n553,
    n420
  );


  nor
  g2262
  (
    n768,
    n572,
    n558,
    n435,
    n680
  );


  xor
  g2263
  (
    n1821,
    n444,
    n462,
    n676,
    n492
  );


  and
  g2264
  (
    n1079,
    n441,
    n471,
    n645,
    n523
  );


  or
  g2265
  (
    n1948,
    n611,
    n523,
    n589,
    n646
  );


  xnor
  g2266
  (
    n733,
    n372,
    n527,
    n470,
    n714
  );


  and
  g2267
  (
    n1054,
    n642,
    n699,
    n505,
    n554
  );


  and
  g2268
  (
    n773,
    n556,
    n447,
    n701,
    n691
  );


  and
  g2269
  (
    n999,
    n661,
    n417,
    n653,
    n559
  );


  or
  g2270
  (
    n1155,
    n461,
    n511,
    n592,
    n686
  );


  nor
  g2271
  (
    n996,
    n477,
    n588,
    n603,
    n531
  );


  nor
  g2272
  (
    n1950,
    n672,
    n418,
    n486,
    n616
  );


  xnor
  g2273
  (
    n863,
    n324,
    n609,
    n328,
    n467
  );


  and
  g2274
  (
    n1812,
    n598,
    n666,
    n374,
    n670
  );


  xnor
  g2275
  (
    n1723,
    n702,
    n578,
    n643,
    n526
  );


  xor
  g2276
  (
    n1608,
    n551,
    n202,
    n434,
    n470
  );


  nor
  g2277
  (
    n1846,
    n485,
    n490,
    n674,
    n598
  );


  and
  g2278
  (
    n1384,
    n686,
    n489,
    n320,
    n653
  );


  nor
  g2279
  (
    n775,
    n381,
    n377,
    n404,
    n667
  );


  nand
  g2280
  (
    n917,
    n447,
    n335,
    n213,
    n599
  );


  xor
  g2281
  (
    n1704,
    n521,
    n501,
    n514,
    n205
  );


  xor
  g2282
  (
    n2500,
    n1186,
    n1059,
    n1727,
    n1325
  );


  xor
  g2283
  (
    n2486,
    n1697,
    n1615,
    n1847,
    n745
  );


  nand
  g2284
  (
    n2738,
    n845,
    n1276,
    n1435,
    n1654
  );


  nand
  g2285
  (
    n2460,
    n1650,
    n1770,
    n848,
    n1529
  );


  nor
  g2286
  (
    n2863,
    n1341,
    n1103,
    n1418,
    n1528
  );


  and
  g2287
  (
    n2640,
    n1413,
    n1140,
    n1440,
    n906
  );


  nor
  g2288
  (
    n2347,
    n1442,
    n1677,
    n955,
    n1120
  );


  xnor
  g2289
  (
    n2860,
    n819,
    n1885,
    n1274,
    n1729
  );


  xnor
  g2290
  (
    n2340,
    n1176,
    n783,
    n914,
    n1797
  );


  nand
  g2291
  (
    n2703,
    n1870,
    n1421,
    n1858,
    n1662
  );


  xnor
  g2292
  (
    n2890,
    n1694,
    n1508,
    n822,
    n1646
  );


  or
  g2293
  (
    n2346,
    n1740,
    n1741,
    n1272,
    n1189
  );


  or
  g2294
  (
    n2492,
    n1641,
    n1487,
    n1486,
    n1506
  );


  and
  g2295
  (
    n2698,
    n1402,
    n996,
    n1166,
    n1404
  );


  xnor
  g2296
  (
    n2634,
    n951,
    n1559,
    n1003,
    n1118
  );


  nand
  g2297
  (
    n2385,
    n763,
    n1104,
    n1663,
    n868
  );


  xnor
  g2298
  (
    n2620,
    n1430,
    n1469,
    n1053,
    n1312
  );


  nor
  g2299
  (
    n2373,
    n832,
    n1377,
    n869,
    n859
  );


  nor
  g2300
  (
    n2454,
    n885,
    n1266,
    n1219,
    n1092
  );


  nand
  g2301
  (
    n2542,
    n1142,
    n1826,
    n1478,
    n1350
  );


  xor
  g2302
  (
    n2521,
    n1715,
    n1813,
    n1119,
    n989
  );


  and
  g2303
  (
    n2522,
    n1881,
    n1374,
    n1292,
    n1563
  );


  xor
  g2304
  (
    n2797,
    n1856,
    n1260,
    n1874,
    n837
  );


  nand
  g2305
  (
    n2651,
    n1682,
    n1810,
    n1545,
    n1033
  );


  xor
  g2306
  (
    n2538,
    n904,
    n1722,
    n1176,
    n1135
  );


  xor
  g2307
  (
    n2540,
    n1229,
    n1418,
    n1626,
    n1598
  );


  and
  g2308
  (
    n2880,
    n963,
    n1087,
    n970,
    n1824
  );


  xor
  g2309
  (
    n2719,
    n1345,
    n1288,
    n1053,
    n1524
  );


  nand
  g2310
  (
    n2390,
    n1607,
    n1297,
    n1405,
    n1266
  );


  nor
  g2311
  (
    n2881,
    n1831,
    n1799,
    n1602,
    n1130
  );


  nand
  g2312
  (
    n2425,
    n1264,
    n1728,
    n1191,
    n959
  );


  or
  g2313
  (
    n2856,
    n1754,
    n1634,
    n1393,
    n1587
  );


  nand
  g2314
  (
    n2585,
    n1805,
    n1041,
    n1342,
    n1798
  );


  or
  g2315
  (
    KeyWire_0_22,
    n1824,
    n1811,
    n1407,
    n832
  );


  or
  g2316
  (
    n2495,
    n1845,
    n1436,
    n1839,
    n1647
  );


  xnor
  g2317
  (
    n2883,
    n823,
    n1268,
    n1403,
    n1733
  );


  and
  g2318
  (
    n2770,
    n1740,
    n1550,
    n1873,
    n1530
  );


  and
  g2319
  (
    n2613,
    n1518,
    n808,
    n1008,
    n1524
  );


  and
  g2320
  (
    n2550,
    n1094,
    n763,
    n744,
    n854
  );


  and
  g2321
  (
    KeyWire_0_11,
    n1064,
    n995,
    n852,
    n1711
  );


  xor
  g2322
  (
    n2497,
    n1781,
    n721,
    n1160,
    n1569
  );


  nand
  g2323
  (
    n2740,
    n1328,
    n1531,
    n1179,
    n1734
  );


  nand
  g2324
  (
    n2333,
    n1385,
    n1383,
    n1443,
    n888
  );


  xor
  g2325
  (
    n2871,
    n733,
    n1891,
    n1086,
    n1143
  );


  or
  g2326
  (
    n2840,
    n1588,
    n774,
    n1761,
    n1696
  );


  or
  g2327
  (
    n2469,
    n1015,
    n1325,
    n1201,
    n1011
  );


  xnor
  g2328
  (
    n2851,
    n896,
    n739,
    n1566,
    n1127
  );


  nor
  g2329
  (
    n2687,
    n724,
    n1685,
    n1446,
    n1034
  );


  nand
  g2330
  (
    n2877,
    n1052,
    n1837,
    n1766,
    n1047
  );


  or
  g2331
  (
    n2337,
    n1302,
    n1073,
    n1381,
    n882
  );


  xor
  g2332
  (
    n2539,
    n1877,
    n1379,
    n1102,
    n1131
  );


  nand
  g2333
  (
    n2637,
    n896,
    n1141,
    n749,
    n1459
  );


  and
  g2334
  (
    n2598,
    n1735,
    n732,
    n1309,
    n1644
  );


  nand
  g2335
  (
    n2511,
    n974,
    n1593,
    n1242,
    n1269
  );


  nand
  g2336
  (
    n2426,
    n1429,
    n1031,
    n1572,
    n1183
  );


  or
  g2337
  (
    n2725,
    n1121,
    n1263,
    n1460,
    n1450
  );


  or
  g2338
  (
    n2749,
    n1071,
    n1779,
    n917,
    n1017
  );


  nand
  g2339
  (
    n2841,
    n1312,
    n1794,
    n1590,
    n1737
  );


  and
  g2340
  (
    n2536,
    n1700,
    n1704,
    n1523,
    n944
  );


  nor
  g2341
  (
    n2334,
    n1040,
    n1184,
    n1032,
    n1582
  );


  nor
  g2342
  (
    n2867,
    n1796,
    n1797,
    n1134,
    n939
  );


  xor
  g2343
  (
    n2517,
    n1580,
    n1474,
    n1160,
    n1083
  );


  xor
  g2344
  (
    n2577,
    n799,
    n779,
    n1493,
    n1025
  );


  xor
  g2345
  (
    n2862,
    n1539,
    n1619,
    n1002,
    n1074
  );


  nand
  g2346
  (
    n2361,
    n908,
    n1803,
    n1889,
    n1565
  );


  and
  g2347
  (
    n2695,
    n749,
    n1104,
    n1692,
    n1671
  );


  and
  g2348
  (
    n2354,
    n1452,
    n942,
    n1648,
    n1188
  );


  xnor
  g2349
  (
    n2506,
    n1753,
    n912,
    n998,
    n1764
  );


  and
  g2350
  (
    n2716,
    n1336,
    n1445,
    n1618,
    n1568
  );


  or
  g2351
  (
    n2836,
    n1809,
    n1512,
    n862,
    n785
  );


  nor
  g2352
  (
    n2670,
    n1843,
    n1393,
    n1523,
    n1291
  );


  or
  g2353
  (
    n2713,
    n947,
    n1806,
    n1631,
    n850
  );


  and
  g2354
  (
    n2413,
    n1417,
    n991,
    n1261,
    n778
  );


  xor
  g2355
  (
    n2665,
    n1363,
    n1706,
    n1079,
    n1662
  );


  xor
  g2356
  (
    n2400,
    n1807,
    n931,
    n844,
    n1619
  );


  xnor
  g2357
  (
    n2518,
    n1807,
    n1042,
    n1279,
    n759
  );


  or
  g2358
  (
    n2528,
    n911,
    n1528,
    n826,
    n1127
  );


  and
  g2359
  (
    n2818,
    n796,
    n1504,
    n1281,
    n1813
  );


  nand
  g2360
  (
    n2433,
    n1326,
    n1894,
    n1020,
    n1007
  );


  nand
  g2361
  (
    n2533,
    n879,
    n1300,
    n1583,
    n1782
  );


  nand
  g2362
  (
    n2833,
    n1749,
    n1380,
    n1377,
    n1189
  );


  nor
  g2363
  (
    n2855,
    n1367,
    n1246,
    n1334,
    n1673
  );


  or
  g2364
  (
    n2420,
    n1578,
    n913,
    n1039,
    n1303
  );


  and
  g2365
  (
    n2717,
    n1321,
    n1793,
    n973,
    n1223
  );


  or
  g2366
  (
    n2527,
    n1145,
    n849,
    n1526,
    n1162
  );


  and
  g2367
  (
    n2571,
    n1729,
    n1096,
    n1785,
    n1744
  );


  nor
  g2368
  (
    n2614,
    n1539,
    n1521,
    n1675,
    n1560
  );


  xor
  g2369
  (
    n2532,
    n1070,
    n1247,
    n991,
    n1365
  );


  or
  g2370
  (
    n2844,
    n791,
    n806,
    n1094,
    n1175
  );


  nor
  g2371
  (
    n2564,
    n1751,
    n1605,
    n1161,
    n1034
  );


  or
  g2372
  (
    n2364,
    n1128,
    n1136,
    n1204,
    n1802
  );


  xnor
  g2373
  (
    n2745,
    n871,
    n1779,
    n792,
    n1553
  );


  xnor
  g2374
  (
    n2336,
    n1466,
    n719,
    n1248,
    n823
  );


  and
  g2375
  (
    n2783,
    n934,
    n1861,
    n1791,
    n1555
  );


  and
  g2376
  (
    n2362,
    n795,
    n1121,
    n1395,
    n1875
  );


  xnor
  g2377
  (
    n2803,
    n1502,
    n1010,
    n1725,
    n1252
  );


  nand
  g2378
  (
    n2573,
    n1352,
    n1585,
    n976,
    n817
  );


  or
  g2379
  (
    n2475,
    n1275,
    n1742,
    n1448,
    n929
  );


  xnor
  g2380
  (
    n2671,
    n802,
    n1036,
    n1615,
    n837
  );


  or
  g2381
  (
    n2393,
    n1443,
    n1463,
    n1473,
    n1129
  );


  nor
  g2382
  (
    n2636,
    n1581,
    n1343,
    n1115,
    n935
  );


  xor
  g2383
  (
    n2647,
    n1125,
    n1638,
    n1544,
    n1244
  );


  nor
  g2384
  (
    n2878,
    n1492,
    n1542,
    n858,
    n910
  );


  xor
  g2385
  (
    n2315,
    n1013,
    n1185,
    n1256,
    n1525
  );


  xor
  g2386
  (
    n2342,
    n921,
    n926,
    n1462,
    n1207
  );


  xnor
  g2387
  (
    n2388,
    n1000,
    n1072,
    n1340,
    n898
  );


  and
  g2388
  (
    n2480,
    n1412,
    n1101,
    n1114,
    n937
  );


  and
  g2389
  (
    n2864,
    n1561,
    n1654,
    n856,
    n830
  );


  nor
  g2390
  (
    n2320,
    n1487,
    n843,
    n1635,
    n1335
  );


  and
  g2391
  (
    n2399,
    n922,
    n936,
    n1603,
    n1633
  );


  nor
  g2392
  (
    n2371,
    n716,
    n1803,
    n718,
    n870
  );


  nor
  g2393
  (
    n2391,
    n1808,
    n940,
    n1099,
    n1219
  );


  nor
  g2394
  (
    n2449,
    n962,
    n1859,
    n1849,
    n1828
  );


  xnor
  g2395
  (
    n2732,
    n1710,
    n1251,
    n747,
    n1431
  );


  xor
  g2396
  (
    n2859,
    n1427,
    n948,
    n1271,
    n1239
  );


  nand
  g2397
  (
    n2588,
    n1221,
    n1336,
    n861,
    n884
  );


  nand
  g2398
  (
    n2645,
    n1371,
    n1830,
    n1660,
    n1360
  );


  xor
  g2399
  (
    n2801,
    n760,
    n1171,
    n903,
    n1378
  );


  and
  g2400
  (
    n2847,
    n892,
    n1498,
    n1889,
    n748
  );


  xnor
  g2401
  (
    n2365,
    n1815,
    n1237,
    n1590,
    n1378
  );


  and
  g2402
  (
    n2567,
    n1113,
    n1403,
    n738,
    n1223
  );


  xnor
  g2403
  (
    n2872,
    n1571,
    n1576,
    n1199,
    n1161
  );


  or
  g2404
  (
    n2706,
    n1853,
    n1556,
    n755,
    n959
  );


  xor
  g2405
  (
    n2802,
    n866,
    n1259,
    n1847,
    n1702
  );


  xor
  g2406
  (
    n2826,
    n1431,
    n1220,
    n825,
    n1144
  );


  or
  g2407
  (
    n2611,
    n1774,
    n1607,
    n1156,
    n831
  );


  or
  g2408
  (
    n2547,
    n857,
    n1871,
    n811,
    n1839
  );


  nand
  g2409
  (
    n2555,
    n1096,
    n1328,
    n1309,
    n1091
  );


  nor
  g2410
  (
    n2606,
    n1134,
    n754,
    n734,
    n1280
  );


  and
  g2411
  (
    n2653,
    n1202,
    n1155,
    n1709,
    n1567
  );


  and
  g2412
  (
    n2601,
    n1082,
    n1222,
    n1769,
    n914
  );


  xnor
  g2413
  (
    n2383,
    n1119,
    n907,
    n736,
    n982
  );


  and
  g2414
  (
    n2657,
    n1339,
    n985,
    n1231,
    n1829
  );


  xnor
  g2415
  (
    n2845,
    n1835,
    n1126,
    n1492,
    n1214
  );


  and
  g2416
  (
    n2510,
    n953,
    n1210,
    n941,
    n1886
  );


  xnor
  g2417
  (
    n2531,
    n934,
    n1320,
    n1686,
    n1545
  );


  nand
  g2418
  (
    n2710,
    n1073,
    n1023,
    n947,
    n1594
  );


  nor
  g2419
  (
    n2356,
    n1569,
    n1738,
    n1676,
    n996
  );


  and
  g2420
  (
    n2696,
    n815,
    n1550,
    n1639,
    n1688
  );


  xor
  g2421
  (
    n2759,
    n887,
    n950,
    n1203,
    n1537
  );


  and
  g2422
  (
    n2694,
    n1605,
    n772,
    n805,
    n1814
  );


  nor
  g2423
  (
    n2473,
    n738,
    n1004,
    n1427,
    n1317
  );


  xor
  g2424
  (
    n2376,
    n1067,
    n1147,
    n1149,
    n1424
  );


  nand
  g2425
  (
    n2760,
    n1627,
    n1468,
    n1659,
    n860
  );


  or
  g2426
  (
    n2625,
    n1845,
    n969,
    n938,
    n807
  );


  or
  g2427
  (
    n2837,
    n866,
    n1761,
    n773,
    n1447
  );


  and
  g2428
  (
    n2854,
    n1316,
    n800,
    n1604,
    n1468
  );


  xnor
  g2429
  (
    n2584,
    n812,
    n1236,
    n1510,
    n1653
  );


  xnor
  g2430
  (
    n2496,
    n1481,
    n1760,
    n1186,
    n1897
  );


  and
  g2431
  (
    n2873,
    n1705,
    n1747,
    n810,
    n1552
  );


  xor
  g2432
  (
    n2525,
    n1456,
    n1515,
    n1785,
    n1520
  );


  and
  g2433
  (
    n2750,
    n1855,
    n891,
    n1494,
    n860
  );


  xor
  g2434
  (
    n2785,
    n1475,
    n1212,
    n1216,
    n816
  );


  or
  g2435
  (
    n2498,
    n1600,
    n1703,
    n1672,
    n1623
  );


  and
  g2436
  (
    n2341,
    n919,
    n1894,
    n1509,
    n1102
  );


  xor
  g2437
  (
    n2616,
    n1850,
    n1472,
    n1521,
    n1722
  );


  or
  g2438
  (
    n2396,
    n1584,
    n957,
    n1810,
    n921
  );


  xor
  g2439
  (
    n2705,
    n1137,
    n1399,
    n1337,
    n1748
  );


  nor
  g2440
  (
    n2462,
    n1355,
    n1527,
    n1448,
    n767
  );


  or
  g2441
  (
    n2644,
    n1876,
    n915,
    n723,
    n890
  );


  or
  g2442
  (
    n2368,
    n1795,
    n878,
    n1398,
    n803
  );


  nor
  g2443
  (
    n2779,
    n1331,
    n796,
    n1187,
    n946
  );


  xor
  g2444
  (
    n2664,
    n1516,
    n977,
    n825,
    n1419
  );


  nand
  g2445
  (
    n2378,
    n1089,
    n1267,
    n1311,
    n1452
  );


  nand
  g2446
  (
    n2551,
    n1314,
    n1333,
    n1525,
    n1068
  );


  nor
  g2447
  (
    n2592,
    n1045,
    n1572,
    n918,
    n863
  );


  and
  g2448
  (
    n2422,
    n1836,
    n1169,
    n813,
    n1600
  );


  nor
  g2449
  (
    n2596,
    n1450,
    n773,
    n1188,
    n1241
  );


  and
  g2450
  (
    n2316,
    n1098,
    n1230,
    n849,
    n1593
  );


  xor
  g2451
  (
    n2652,
    n1567,
    n735,
    n1513,
    n1493
  );


  nand
  g2452
  (
    n2810,
    n1652,
    n1306,
    n1438,
    n1684
  );


  nor
  g2453
  (
    n2467,
    n1357,
    n990,
    n830,
    n737
  );


  nor
  g2454
  (
    n2578,
    n913,
    n1351,
    n1884,
    n927
  );


  nor
  g2455
  (
    n2494,
    n1246,
    n1007,
    n1571,
    n841
  );


  xnor
  g2456
  (
    n2700,
    n1742,
    n1625,
    n839,
    n1025
  );


  xnor
  g2457
  (
    n2764,
    n989,
    n1295,
    n889,
    n1746
  );


  or
  g2458
  (
    n2363,
    n1038,
    n1834,
    n1099,
    n1500
  );


  nor
  g2459
  (
    n2787,
    n1484,
    n1105,
    n1757,
    n790
  );


  nor
  g2460
  (
    n2515,
    n789,
    n1433,
    n781,
    n730
  );


  xnor
  g2461
  (
    n2329,
    n1013,
    n980,
    n1088,
    n1519
  );


  xor
  g2462
  (
    n2884,
    n1806,
    n1390,
    n883,
    n1559
  );


  xnor
  g2463
  (
    n2782,
    n1586,
    n928,
    n988,
    n798
  );


  xnor
  g2464
  (
    n2650,
    n1163,
    n965,
    n1062,
    n1801
  );


  xor
  g2465
  (
    n2672,
    n1061,
    n867,
    n1721,
    n1300
  );


  nor
  g2466
  (
    n2463,
    n1274,
    n1085,
    n1825,
    n1848
  );


  and
  g2467
  (
    n2607,
    n772,
    n846,
    n1610,
    n818
  );


  nand
  g2468
  (
    n2404,
    n1152,
    n1736,
    n1812,
    n1868
  );


  nor
  g2469
  (
    n2846,
    n1384,
    n1663,
    n1495,
    n1712
  );


  and
  g2470
  (
    n2568,
    n1344,
    n781,
    n1522,
    n1371
  );


  nand
  g2471
  (
    n2470,
    n1631,
    n746,
    n960,
    n1086
  );


  xor
  g2472
  (
    n2436,
    n1863,
    n1110,
    n1277,
    n1558
  );


  nor
  g2473
  (
    n2471,
    n1364,
    n1774,
    n1780,
    n1636
  );


  and
  g2474
  (
    n2781,
    n790,
    n1556,
    n1517,
    n1887
  );


  xor
  g2475
  (
    n2520,
    n1072,
    n1895,
    n1707,
    n1899
  );


  nand
  g2476
  (
    n2673,
    n1145,
    n912,
    n1148,
    n1315
  );


  nor
  g2477
  (
    n2746,
    n1049,
    n1208,
    n1659,
    n1181
  );


  xor
  g2478
  (
    n2431,
    n1510,
    n1732,
    n1865,
    n1630
  );


  and
  g2479
  (
    n2344,
    n1190,
    n1898,
    n935,
    n808
  );


  and
  g2480
  (
    n2659,
    n1685,
    n1864,
    n1529,
    n853
  );


  and
  g2481
  (
    n2523,
    n752,
    n1177,
    n1503,
    n1180
  );


  nor
  g2482
  (
    n2784,
    n1772,
    n836,
    n1743,
    n1834
  );


  or
  g2483
  (
    n2441,
    n1308,
    n1240,
    n1110,
    n971
  );


  nor
  g2484
  (
    n2641,
    n1805,
    n1395,
    n1464,
    n1574
  );


  xnor
  g2485
  (
    n2805,
    n1388,
    n1527,
    n1899,
    n1065
  );


  xnor
  g2486
  (
    n2563,
    n1075,
    n1687,
    n1778,
    n762
  );


  nor
  g2487
  (
    n2627,
    n1036,
    n1628,
    n1143,
    n1250
  );


  xor
  g2488
  (
    n2649,
    n1775,
    n1809,
    n1819,
    n1876
  );


  nor
  g2489
  (
    n2546,
    n1767,
    n1690,
    n1477,
    n764
  );


  and
  g2490
  (
    n2505,
    n745,
    n1669,
    n1018,
    n1304
  );


  xor
  g2491
  (
    n2428,
    n1698,
    n1323,
    n1513,
    n740
  );


  xnor
  g2492
  (
    n2809,
    n1033,
    n757,
    n1726,
    n1151
  );


  nand
  g2493
  (
    n2587,
    n1892,
    n1723,
    n1612,
    n1670
  );


  xor
  g2494
  (
    n2381,
    n1784,
    n980,
    n1501,
    n791
  );


  or
  g2495
  (
    n2330,
    n1710,
    n816,
    n1865,
    n1831
  );


  and
  g2496
  (
    n2815,
    n1282,
    n1852,
    n1638,
    n1070
  );


  xnor
  g2497
  (
    n2452,
    n1185,
    n1137,
    n1595,
    n1838
  );


  xor
  g2498
  (
    n2786,
    n1614,
    n1879,
    n1258,
    n1875
  );


  nand
  g2499
  (
    n2739,
    n1833,
    n967,
    n1084,
    n1795
  );


  xnor
  g2500
  (
    n2351,
    n1522,
    n1217,
    n1195,
    n1122
  );


  nor
  g2501
  (
    n2767,
    n741,
    n1718,
    n1604,
    n1714
  );


  xnor
  g2502
  (
    n2526,
    n1392,
    n1286,
    n1887,
    n809
  );


  nor
  g2503
  (
    n2619,
    n1187,
    n1736,
    n1434,
    n1582
  );


  and
  g2504
  (
    n2434,
    n882,
    n1318,
    n771,
    n1399
  );


  nand
  g2505
  (
    n2604,
    n1478,
    n809,
    n1543,
    n1049
  );


  and
  g2506
  (
    n2524,
    n901,
    n875,
    n815,
    n1597
  );


  nand
  g2507
  (
    n2817,
    n1243,
    n1641,
    n805,
    n793
  );


  xor
  g2508
  (
    n2712,
    n1012,
    n1239,
    n1108,
    n1480
  );


  and
  g2509
  (
    n2885,
    n1850,
    n1410,
    n1629,
    n840
  );


  xnor
  g2510
  (
    n2655,
    n1275,
    n746,
    n1629,
    n1538
  );


  and
  g2511
  (
    n2658,
    n1409,
    n1630,
    n1128,
    n930
  );


  nand
  g2512
  (
    n2615,
    n964,
    n1664,
    n774,
    n1307
  );


  and
  g2513
  (
    n2502,
    n840,
    n1209,
    n1520,
    n1156
  );


  xnor
  g2514
  (
    n2309,
    n1133,
    n1307,
    n1408,
    n1728
  );


  nand
  g2515
  (
    n2446,
    n775,
    n1338,
    n1606,
    n820
  );


  nor
  g2516
  (
    n2850,
    n1048,
    n1057,
    n1091,
    n1112
  );


  nor
  g2517
  (
    n2317,
    n1158,
    n1592,
    n1692,
    n1090
  );


  xnor
  g2518
  (
    n2692,
    n1170,
    n1719,
    n1500,
    n865
  );


  nor
  g2519
  (
    n2887,
    n869,
    n1512,
    n999,
    n1471
  );


  or
  g2520
  (
    n2623,
    n1220,
    n1168,
    n1391,
    n1098
  );


  xnor
  g2521
  (
    n2734,
    n993,
    n857,
    n1506,
    n1201
  );


  or
  g2522
  (
    n2423,
    n1376,
    n1428,
    n1191,
    n726
  );


  xor
  g2523
  (
    n2387,
    n1037,
    n1397,
    n1077,
    n1413
  );


  xor
  g2524
  (
    n2453,
    n943,
    n895,
    n1709,
    n1179
  );


  xnor
  g2525
  (
    n2691,
    n1653,
    n1617,
    n1730,
    n1637
  );


  nor
  g2526
  (
    n2656,
    n891,
    n1819,
    n1577,
    n744
  );


  xor
  g2527
  (
    n2876,
    n1242,
    n1173,
    n1446,
    n983
  );


  xnor
  g2528
  (
    n2679,
    n1815,
    n1132,
    n1341,
    n1563
  );


  nor
  g2529
  (
    n2823,
    n1412,
    n1745,
    n1765,
    n1693
  );


  xnor
  g2530
  (
    n2729,
    n1755,
    n1611,
    n1716,
    n1555
  );


  nand
  g2531
  (
    n2326,
    n1290,
    n1147,
    n1319,
    n1758
  );


  and
  g2532
  (
    n2842,
    n986,
    n1451,
    n767,
    n1483
  );


  or
  g2533
  (
    n2458,
    n1821,
    n1861,
    n1460,
    n1200
  );


  xor
  g2534
  (
    n2835,
    n894,
    n1456,
    n1704,
    n1759
  );


  xor
  g2535
  (
    n2580,
    n1159,
    n1844,
    n1701,
    n1675
  );


  xnor
  g2536
  (
    n2704,
    n969,
    n1323,
    n1580,
    n1666
  );


  xor
  g2537
  (
    n2535,
    n1703,
    n1234,
    n1235,
    n1491
  );


  and
  g2538
  (
    n2776,
    n937,
    n1008,
    n1349,
    n821
  );


  xnor
  g2539
  (
    n2674,
    n1291,
    n1316,
    n1071,
    n1599
  );


  nand
  g2540
  (
    n2780,
    n894,
    n1449,
    n1869,
    n1843
  );


  and
  g2541
  (
    n2748,
    n862,
    n1532,
    n917,
    n1547
  );


  xor
  g2542
  (
    n2432,
    n911,
    n756,
    n1758,
    n1765
  );


  nor
  g2543
  (
    n2418,
    n1713,
    n1748,
    n1612,
    n1222
  );


  nand
  g2544
  (
    n2405,
    n1800,
    n1231,
    n1489,
    n797
  );


  xnor
  g2545
  (
    n2556,
    n1203,
    n1060,
    n1536,
    n1422
  );


  xor
  g2546
  (
    n2472,
    n768,
    n1714,
    n1090,
    n1793
  );


  xnor
  g2547
  (
    n2407,
    n954,
    n1241,
    n1050,
    n1282
  );


  and
  g2548
  (
    n2447,
    n988,
    n1453,
    n1024,
    n1283
  );


  or
  g2549
  (
    n2680,
    n1623,
    n1372,
    n1396,
    n1883
  );


  and
  g2550
  (
    n2882,
    n1198,
    n1217,
    n1480,
    n1470
  );


  or
  g2551
  (
    n2800,
    n1124,
    n1636,
    n1733,
    n752
  );


  xnor
  g2552
  (
    n2416,
    n1212,
    n902,
    n1125,
    n1647
  );


  nand
  g2553
  (
    n2490,
    n1666,
    n1365,
    n743,
    n1278
  );


  xor
  g2554
  (
    n2771,
    n1637,
    n1111,
    n1076,
    n872
  );


  xnor
  g2555
  (
    n2869,
    n1472,
    n804,
    n1329,
    n1488
  );


  xor
  g2556
  (
    n2411,
    n1088,
    n1514,
    n1296,
    n812
  );


  xor
  g2557
  (
    n2324,
    n1124,
    n1064,
    n1407,
    n1708
  );


  nor
  g2558
  (
    n2461,
    n1397,
    n1644,
    n1570,
    n1294
  );


  nand
  g2559
  (
    n2758,
    n787,
    n1419,
    n1240,
    n786
  );


  nand
  g2560
  (
    n2444,
    n1425,
    n968,
    n1101,
    n986
  );


  nor
  g2561
  (
    n2558,
    n925,
    n944,
    n1453,
    n1796
  );


  nand
  g2562
  (
    n2677,
    n1581,
    n1324,
    n1426,
    n1897
  );


  or
  g2563
  (
    n2667,
    n1327,
    n739,
    n1423,
    n1193
  );


  nor
  g2564
  (
    n2812,
    n1368,
    n848,
    n1857,
    n1056
  );


  or
  g2565
  (
    n2448,
    n1006,
    n803,
    n1215,
    n1640
  );


  or
  g2566
  (
    n2631,
    n1109,
    n1700,
    n1486,
    n916
  );


  and
  g2567
  (
    n2682,
    n1192,
    n1491,
    n794,
    n1485
  );


  nand
  g2568
  (
    n2618,
    n1695,
    n1444,
    n766,
    n789
  );


  xor
  g2569
  (
    n2360,
    n1100,
    n903,
    n1747,
    n1093
  );


  nand
  g2570
  (
    n2628,
    n1669,
    n1829,
    n1422,
    n1165
  );


  or
  g2571
  (
    n2791,
    n1599,
    n957,
    n1108,
    n1170
  );


  or
  g2572
  (
    n2825,
    n1055,
    n1689,
    n770,
    n1749
  );


  nand
  g2573
  (
    n2622,
    n1872,
    n883,
    n1602,
    n864
  );


  nor
  g2574
  (
    n2332,
    n754,
    n1777,
    n1757,
    n1210
  );


  xnor
  g2575
  (
    n2489,
    n893,
    n1461,
    n1674,
    n1224
  );


  xnor
  g2576
  (
    n2813,
    n1394,
    n1672,
    n999,
    n1253
  );


  xnor
  g2577
  (
    n2417,
    n963,
    n1154,
    n1310,
    n1206
  );


  xor
  g2578
  (
    n2874,
    n1330,
    n1068,
    n1549,
    n1376
  );


  and
  g2579
  (
    n2313,
    n979,
    n923,
    n833,
    n951
  );


  xor
  g2580
  (
    n2638,
    n1254,
    n1164,
    n1205,
    n1270
  );


  nor
  g2581
  (
    n2794,
    n1632,
    n993,
    n1624,
    n1211
  );


  and
  g2582
  (
    n2635,
    n1227,
    n1677,
    n1658,
    n1105
  );


  nand
  g2583
  (
    n2807,
    n1233,
    n835,
    n1040,
    n1711
  );


  xor
  g2584
  (
    n2777,
    n1541,
    n780,
    n1479,
    n1303
  );


  xor
  g2585
  (
    n2684,
    n1573,
    n1152,
    n977,
    n750
  );


  xor
  g2586
  (
    n2481,
    n1180,
    n1461,
    n757,
    n1651
  );


  nand
  g2587
  (
    n2372,
    n1353,
    n936,
    n750,
    n941
  );


  and
  g2588
  (
    n2733,
    n802,
    n1652,
    n1643,
    n800
  );


  nor
  g2589
  (
    n2709,
    n1400,
    n1515,
    n1862,
    n1665
  );


  xor
  g2590
  (
    n2654,
    n1597,
    n1601,
    n933,
    n1295
  );


  nor
  g2591
  (
    n2661,
    n1021,
    n1163,
    n854,
    n1032
  );


  nor
  g2592
  (
    n2646,
    n1726,
    n1469,
    n1664,
    n962
  );


  nor
  g2593
  (
    n2305,
    n1896,
    n1416,
    n1004,
    n1364
  );


  nand
  g2594
  (
    n2582,
    n1698,
    n1473,
    n1322,
    n1421
  );


  or
  g2595
  (
    n2370,
    n1535,
    n717,
    n1540,
    n952
  );


  and
  g2596
  (
    n2643,
    n1546,
    n954,
    n1755,
    n1626
  );


  or
  g2597
  (
    n2747,
    n1043,
    n1621,
    n1738,
    n1177
  );


  xnor
  g2598
  (
    n2579,
    n1691,
    n1357,
    n1621,
    n979
  );


  nor
  g2599
  (
    n2353,
    n1798,
    n1485,
    n1285,
    n1337
  );


  or
  g2600
  (
    n2429,
    n1289,
    n888,
    n1010,
    n1287
  );


  xor
  g2601
  (
    n2508,
    n1557,
    n753,
    n886,
    n1296
  );


  xor
  g2602
  (
    n2544,
    n1442,
    n1837,
    n1617,
    n1439
  );


  xnor
  g2603
  (
    n2485,
    n1583,
    n1029,
    n990,
    n1348
  );


  or
  g2604
  (
    n2566,
    n1657,
    n946,
    n1001,
    n1804
  );


  nor
  g2605
  (
    n2773,
    n1799,
    n1482,
    n1235,
    n1622
  );


  and
  g2606
  (
    n2830,
    n1057,
    n1087,
    n1115,
    n792
  );


  xnor
  g2607
  (
    n2414,
    n1683,
    n1823,
    n881,
    n974
  );


  or
  g2608
  (
    n2476,
    n1890,
    n747,
    n1721,
    n1117
  );


  or
  g2609
  (
    n2612,
    n1353,
    n1878,
    n1503,
    n846
  );


  nand
  g2610
  (
    n2788,
    n967,
    n1020,
    n1384,
    n1768
  );


  xor
  g2611
  (
    n2477,
    n842,
    n1297,
    n1731,
    n1574
  );


  or
  g2612
  (
    n2699,
    n1248,
    n1668,
    n1667,
    n1568
  );


  or
  g2613
  (
    n2468,
    n1014,
    n1379,
    n755,
    n1429
  );


  xor
  g2614
  (
    n2605,
    n1047,
    n1249,
    n932,
    n1402
  );


  and
  g2615
  (
    n2367,
    n1536,
    n1359,
    n1299,
    n1030
  );


  xor
  g2616
  (
    n2384,
    n1017,
    n1499,
    n1289,
    n1178
  );


  xor
  g2617
  (
    n2597,
    n1135,
    n1827,
    n1505,
    n811
  );


  nand
  g2618
  (
    n2852,
    n1244,
    n1406,
    n1359,
    n1867
  );


  nor
  g2619
  (
    n2728,
    n1081,
    n1530,
    n1823,
    n1465
  );


  nand
  g2620
  (
    n2406,
    n1394,
    n1355,
    n1770,
    n1247
  );


  xor
  g2621
  (
    n2335,
    n1226,
    n1885,
    n1752,
    n1730
  );


  and
  g2622
  (
    n2466,
    n1410,
    n1132,
    n1832,
    n1259
  );


  and
  g2623
  (
    n2402,
    n1154,
    n1006,
    n1463,
    n856
  );


  xnor
  g2624
  (
    n2427,
    n1228,
    n1541,
    n1716,
    n1131
  );


  nor
  g2625
  (
    n2735,
    n864,
    n859,
    n798,
    n1097
  );


  xnor
  g2626
  (
    n2727,
    n1059,
    n870,
    n1324,
    n1100
  );


  nor
  g2627
  (
    n2375,
    n1585,
    n1649,
    n1873,
    n1298
  );


  xor
  g2628
  (
    n2401,
    n1370,
    n972,
    n1734,
    n1846
  );


  or
  g2629
  (
    n2648,
    n1868,
    n948,
    n964,
    n827
  );


  xor
  g2630
  (
    n2744,
    n885,
    n1841,
    n1029,
    n1735
  );


  nand
  g2631
  (
    n2753,
    n1846,
    n1657,
    n1475,
    n1319
  );


  xor
  g2632
  (
    n2306,
    n1551,
    n1388,
    n1281,
    n1553
  );


  xor
  g2633
  (
    n2503,
    n1166,
    n1577,
    n961,
    n1820
  );


  and
  g2634
  (
    n2575,
    n978,
    n1095,
    n1867,
    n1182
  );


  nor
  g2635
  (
    n2723,
    n1565,
    n742,
    n1390,
    n1642
  );


  xor
  g2636
  (
    n2366,
    n1042,
    n997,
    n741,
    n1893
  );


  xor
  g2637
  (
    n2875,
    n1814,
    n1345,
    n1676,
    n1294
  );


  nand
  g2638
  (
    n2369,
    n1146,
    n1420,
    n765,
    n1633
  );


  xnor
  g2639
  (
    n2374,
    n794,
    n1476,
    n1649,
    n992
  );


  and
  g2640
  (
    n2772,
    n1794,
    n1821,
    n1543,
    n1343
  );


  nor
  g2641
  (
    n2701,
    n965,
    n1387,
    n1204,
    n1888
  );


  xor
  g2642
  (
    n2683,
    n1558,
    n1880,
    n782,
    n1725
  );


  nor
  g2643
  (
    n2724,
    n928,
    n1356,
    n1686,
    n1078
  );


  or
  g2644
  (
    n2829,
    n961,
    n1881,
    n768,
    n1562
  );


  xor
  g2645
  (
    n2557,
    n1272,
    n874,
    n1862,
    n1447
  );


  and
  g2646
  (
    n2543,
    n820,
    n1213,
    n1077,
    n1424
  );


  xnor
  g2647
  (
    n2819,
    n1404,
    n1374,
    n1080,
    n833
  );


  or
  g2648
  (
    n2410,
    n1474,
    n1157,
    n1773,
    n1680
  );


  nand
  g2649
  (
    n2730,
    n1699,
    n1783,
    n1306,
    n910
  );


  and
  g2650
  (
    n2565,
    n1830,
    n1406,
    n1750,
    n1027
  );


  nand
  g2651
  (
    n2311,
    n1380,
    n1046,
    n1339,
    n1656
  );


  and
  g2652
  (
    n2756,
    n817,
    n1441,
    n901,
    n1023
  );


  nand
  g2653
  (
    n2339,
    n1284,
    n892,
    n770,
    n1764
  );


  nor
  g2654
  (
    n2435,
    n1258,
    n1417,
    n1778,
    n978
  );


  or
  g2655
  (
    n2603,
    n1494,
    n932,
    n1237,
    n1792
  );


  nor
  g2656
  (
    n2459,
    n1715,
    n1081,
    n1002,
    n998
  );


  nor
  g2657
  (
    n2307,
    n1301,
    n838,
    n1773,
    n1437
  );


  or
  g2658
  (
    n2591,
    n1012,
    n898,
    n1717,
    n1026
  );


  and
  g2659
  (
    n2457,
    n1400,
    n976,
    n1882,
    n1759
  );


  nor
  g2660
  (
    n2857,
    n1298,
    n1083,
    n1750,
    n1858
  );


  xor
  g2661
  (
    n2888,
    n1708,
    n1268,
    n992,
    n1069
  );


  nand
  g2662
  (
    n2593,
    n760,
    n1234,
    n1892,
    n1532
  );


  xor
  g2663
  (
    n2827,
    n1816,
    n1476,
    n873,
    n1279
  );


  xor
  g2664
  (
    n2554,
    n1005,
    n1044,
    n1144,
    n907
  );


  and
  g2665
  (
    n2545,
    n1454,
    n1864,
    n1157,
    n1879
  );


  and
  g2666
  (
    n2594,
    n867,
    n1822,
    n1211,
    n1511
  );


  nor
  g2667
  (
    n2482,
    n939,
    n897,
    n1534,
    n966
  );


  and
  g2668
  (
    n2811,
    n1573,
    n1225,
    n942,
    n1009
  );


  or
  g2669
  (
    n2493,
    n1270,
    n1167,
    n1228,
    n1537
  );


  nor
  g2670
  (
    n2450,
    n1445,
    n1030,
    n975,
    n900
  );


  xnor
  g2671
  (
    n2352,
    n1299,
    n720,
    n1622,
    n1771
  );


  xor
  g2672
  (
    n2438,
    n1856,
    n1681,
    n761,
    n1458
  );


  nor
  g2673
  (
    n2408,
    n1392,
    n1489,
    n1173,
    n899
  );


  nand
  g2674
  (
    n2602,
    n1459,
    n1818,
    n940,
    n1435
  );


  or
  g2675
  (
    n2430,
    n1866,
    n884,
    n1058,
    n1790
  );


  xnor
  g2676
  (
    n2552,
    n1603,
    n1516,
    n1174,
    n1428
  );


  and
  g2677
  (
    n2678,
    n1028,
    n1383,
    n1634,
    n1035
  );


  nand
  g2678
  (
    n2806,
    n1366,
    n1332,
    n1465,
    n1643
  );


  nor
  g2679
  (
    n2504,
    n1123,
    n1505,
    n1542,
    n1595
  );


  and
  g2680
  (
    n2509,
    n886,
    n1369,
    n1167,
    n1504
  );


  xor
  g2681
  (
    n2715,
    n994,
    n797,
    n924,
    n1016
  );


  xnor
  g2682
  (
    n2792,
    n1254,
    n759,
    n933,
    n1356
  );


  or
  g2683
  (
    n2804,
    n1719,
    n1775,
    n1680,
    n1739
  );


  nor
  g2684
  (
    n2338,
    n1586,
    n1860,
    n1141,
    n895
  );


  xnor
  g2685
  (
    n2639,
    n1762,
    n1218,
    n1389,
    n1679
  );


  nand
  g2686
  (
    n2514,
    n1455,
    n1149,
    n881,
    n1069
  );


  xor
  g2687
  (
    n2559,
    n1287,
    n1391,
    n897,
    n1611
  );


  nand
  g2688
  (
    n2816,
    n1584,
    n987,
    n1398,
    n972
  );


  xnor
  g2689
  (
    n2762,
    n1112,
    n1625,
    n966,
    n1832
  );


  xor
  g2690
  (
    n2519,
    n893,
    n953,
    n1405,
    n1146
  );


  nor
  g2691
  (
    n2358,
    n1414,
    n1041,
    n1168,
    n1678
  );


  xnor
  g2692
  (
    n2456,
    n1679,
    n1882,
    n1346,
    n1158
  );


  nand
  g2693
  (
    n2693,
    n1278,
    n1826,
    n804,
    n756
  );


  xor
  g2694
  (
    n2778,
    n1628,
    n872,
    n1788,
    n1438
  );


  nand
  g2695
  (
    n2722,
    n1060,
    n1869,
    n1305,
    n1646
  );


  nor
  g2696
  (
    n2303,
    n1028,
    n1517,
    n1256,
    n1233
  );


  and
  g2697
  (
    n2737,
    n1076,
    n1578,
    n1660,
    n1015
  );


  xnor
  g2698
  (
    n2421,
    n1488,
    n1215,
    n1554,
    n1092
  );


  or
  g2699
  (
    n2357,
    n1713,
    n1264,
    n1330,
    n1457
  );


  or
  g2700
  (
    n2834,
    n793,
    n769,
    n1169,
    n1107
  );


  xnor
  g2701
  (
    n2688,
    n1196,
    n1575,
    n1432,
    n1800
  );


  nor
  g2702
  (
    n2866,
    n956,
    n1737,
    n1792,
    n1344
  );


  nor
  g2703
  (
    n2697,
    n1153,
    n1288,
    n1139,
    n1514
  );


  xnor
  g2704
  (
    n2843,
    n1227,
    n1787,
    n762,
    n1693
  );


  nand
  g2705
  (
    n2630,
    n1609,
    n1182,
    n1608,
    n1682
  );


  or
  g2706
  (
    n2529,
    n1361,
    n1003,
    n1411,
    n1816
  );


  nor
  g2707
  (
    n2848,
    n1827,
    n1065,
    n1320,
    n1695
  );


  or
  g2708
  (
    n2798,
    n1560,
    n1197,
    n1687,
    n1739
  );


  nor
  g2709
  (
    n2304,
    n1277,
    n871,
    n1712,
    n766
  );


  nor
  g2710
  (
    n2562,
    n1691,
    n727,
    n1745,
    n784
  );


  nand
  g2711
  (
    n2726,
    n1635,
    n1019,
    n1609,
    n1113
  );


  nor
  g2712
  (
    n2586,
    n847,
    n788,
    n1401,
    n1354
  );


  or
  g2713
  (
    n2849,
    n814,
    n1613,
    n1554,
    n1346
  );


  and
  g2714
  (
    n2395,
    n1817,
    n984,
    n1051,
    n1498
  );


  and
  g2715
  (
    n2455,
    n975,
    n1655,
    n1467,
    n1776
  );


  or
  g2716
  (
    n2419,
    n1490,
    n1482,
    n1606,
    n1301
  );


  or
  g2717
  (
    n2660,
    n1226,
    n1142,
    n1181,
    n1640
  );


  xor
  g2718
  (
    n2569,
    n1362,
    n1396,
    n831,
    n1754
  );


  and
  g2719
  (
    n2308,
    n960,
    n851,
    n1723,
    n1195
  );


  xnor
  g2720
  (
    n2488,
    n930,
    n834,
    n1895,
    n1123
  );


  xnor
  g2721
  (
    n2633,
    n1150,
    n1349,
    n1273,
    n877
  );


  and
  g2722
  (
    n2397,
    n1308,
    n1338,
    n1197,
    n729
  );


  nor
  g2723
  (
    n2743,
    n973,
    n742,
    n1564,
    n1037
  );


  nand
  g2724
  (
    n2808,
    n1706,
    n1771,
    n1720,
    n1872
  );


  or
  g2725
  (
    n2599,
    n1253,
    n1812,
    n889,
    n1608
  );


  xor
  g2726
  (
    n2707,
    n1420,
    n1844,
    n1432,
    n1063
  );


  and
  g2727
  (
    n2769,
    n1575,
    n821,
    n949,
    n1425
  );


  nor
  g2728
  (
    n2394,
    n1044,
    n1533,
    n1557,
    n777
  );


  nor
  g2729
  (
    n2870,
    n1627,
    n1232,
    n1546,
    n1502
  );


  or
  g2730
  (
    n2718,
    n1763,
    n1645,
    n1218,
    n853
  );


  xor
  g2731
  (
    n2814,
    n1054,
    n1511,
    n1038,
    n880
  );


  nand
  g2732
  (
    n2583,
    n1208,
    n1589,
    n1138,
    n1313
  );


  nor
  g2733
  (
    n2865,
    n1153,
    n1358,
    n1898,
    n1437
  );


  and
  g2734
  (
    n2530,
    n1171,
    n1024,
    n1842,
    n880
  );


  and
  g2735
  (
    n2721,
    n1386,
    n1851,
    n958,
    n876
  );


  or
  g2736
  (
    n2479,
    n1276,
    n1589,
    n971,
    n737
  );


  nand
  g2737
  (
    n2581,
    n843,
    n1852,
    n1019,
    n1111
  );


  and
  g2738
  (
    n2822,
    n1116,
    n1285,
    n807,
    n1026
  );


  nor
  g2739
  (
    n2765,
    n1103,
    n1194,
    n1109,
    n1587
  );


  or
  g2740
  (
    n2799,
    n806,
    n1079,
    n1690,
    n731
  );


  nor
  g2741
  (
    n2858,
    n1292,
    n1035,
    n1250,
    n1229
  );


  xnor
  g2742
  (
    n2676,
    n1078,
    n1462,
    n1842,
    n1368
  );


  nor
  g2743
  (
    n2310,
    n1251,
    n1048,
    n1097,
    n1031
  );


  and
  g2744
  (
    n2442,
    n1273,
    n1011,
    n1552,
    n1252
  );


  xnor
  g2745
  (
    n2589,
    n994,
    n1497,
    n1802,
    n1172
  );


  or
  g2746
  (
    n2853,
    n1269,
    n1075,
    n728,
    n828
  );


  xor
  g2747
  (
    n2755,
    n1697,
    n1054,
    n1592,
    n1507
  );


  xor
  g2748
  (
    n2513,
    n1454,
    n1620,
    n1681,
    n1804
  );


  nor
  g2749
  (
    n2534,
    n1871,
    n733,
    n1880,
    n1801
  );


  nand
  g2750
  (
    n2570,
    n943,
    n1519,
    n788,
    n1780
  );


  or
  g2751
  (
    n2832,
    n1089,
    n1789,
    n1414,
    n1678
  );


  and
  g2752
  (
    n2443,
    n1674,
    n1120,
    n1753,
    n877
  );


  xor
  g2753
  (
    n2626,
    n945,
    n1192,
    n1436,
    n949
  );


  and
  g2754
  (
    n2766,
    n1369,
    n1415,
    n1576,
    n1347
  );


  and
  g2755
  (
    n2886,
    n1164,
    n1763,
    n1661,
    n1642
  );


  and
  g2756
  (
    n2831,
    n1624,
    n1548,
    n1022,
    n1509
  );


  nand
  g2757
  (
    n2512,
    n1408,
    n1479,
    n1838,
    n1133
  );


  and
  g2758
  (
    n2720,
    n916,
    n863,
    n1183,
    n1386
  );


  and
  g2759
  (
    n2501,
    n779,
    n1245,
    n1415,
    n1720
  );


  nand
  g2760
  (
    n2318,
    n1214,
    n822,
    n819,
    n1001
  );


  xnor
  g2761
  (
    n2754,
    n1172,
    n929,
    n850,
    n1387
  );


  and
  g2762
  (
    n2379,
    n1080,
    n1411,
    n926,
    n1760
  );


  xor
  g2763
  (
    n2314,
    n1790,
    n1743,
    n1854,
    n905
  );


  xnor
  g2764
  (
    n2322,
    n758,
    n1650,
    n1833,
    n1350
  );


  nand
  g2765
  (
    n2328,
    n1471,
    n1786,
    n1818,
    n861
  );


  or
  g2766
  (
    n2415,
    n1051,
    n1689,
    n1082,
    n952
  );


  xor
  g2767
  (
    n2572,
    n983,
    n1302,
    n1477,
    n1039
  );


  nor
  g2768
  (
    n2624,
    n1534,
    n1317,
    n938,
    n1342
  );


  nor
  g2769
  (
    n2768,
    n1588,
    n1213,
    n799,
    n1334
  );


  nor
  g2770
  (
    n2828,
    n1267,
    n1262,
    n987,
    n1000
  );


  nor
  g2771
  (
    n2348,
    n801,
    n915,
    n955,
    n786
  );


  xor
  g2772
  (
    n2331,
    n1490,
    n1840,
    n1835,
    n722
  );


  and
  g2773
  (
    n2685,
    n1705,
    n801,
    n908,
    n1085
  );


  nand
  g2774
  (
    n2345,
    n1249,
    n1564,
    n1744,
    n1890
  );


  nand
  g2775
  (
    n2752,
    n879,
    n1430,
    n1434,
    n920
  );


  and
  g2776
  (
    KeyWire_0_30,
    n725,
    n1741,
    n858,
    n1198
  );


  nand
  g2777
  (
    n2821,
    n1271,
    n1768,
    n1548,
    n1061
  );


  and
  g2778
  (
    n2609,
    n1347,
    n1457,
    n1014,
    n1518
  );


  xnor
  g2779
  (
    n2507,
    n751,
    n1313,
    n1367,
    n1290
  );


  nand
  g2780
  (
    n2610,
    n1444,
    n1483,
    n1699,
    n925
  );


  xor
  g2781
  (
    n2763,
    n758,
    n1050,
    n1822,
    n1332
  );


  and
  g2782
  (
    KeyWire_0_24,
    n1225,
    n1165,
    n1526,
    n985
  );


  xnor
  g2783
  (
    n2669,
    n1209,
    n1499,
    n1891,
    n1150
  );


  and
  g2784
  (
    n2553,
    n1781,
    n1651,
    n1202,
    n1257
  );


  nand
  g2785
  (
    n2774,
    n924,
    n1598,
    n777,
    n1859
  );


  and
  g2786
  (
    n2478,
    n1366,
    n1074,
    n931,
    n826
  );


  and
  g2787
  (
    n2663,
    n1389,
    n783,
    n1114,
    n1808
  );


  xor
  g2788
  (
    n2403,
    n1286,
    n818,
    n838,
    n1016
  );


  or
  g2789
  (
    n2412,
    n1766,
    n1702,
    n834,
    n1360
  );


  and
  g2790
  (
    n2742,
    n1293,
    n1717,
    n1255,
    n1863
  );


  and
  g2791
  (
    n2343,
    n1373,
    n785,
    n1118,
    n875
  );


  xor
  g2792
  (
    n2675,
    n1052,
    n1857,
    n769,
    n1840
  );


  nand
  g2793
  (
    n2516,
    n1688,
    n1329,
    n905,
    n1314
  );


  nor
  g2794
  (
    n2838,
    n1451,
    n1540,
    n1694,
    n1614
  );


  xnor
  g2795
  (
    n2327,
    n1751,
    n1138,
    n1084,
    n1579
  );


  and
  g2796
  (
    n2736,
    n1238,
    n900,
    n1789,
    n778
  );


  nand
  g2797
  (
    n2689,
    n1549,
    n1596,
    n865,
    n1648
  );


  xor
  g2798
  (
    n2590,
    n1449,
    n927,
    n1860,
    n734
  );


  nor
  g2799
  (
    n2608,
    n1632,
    n1841,
    n845,
    n1481
  );


  xnor
  g2800
  (
    n2751,
    n1893,
    n1439,
    n1409,
    n918
  );


  xnor
  g2801
  (
    n2349,
    n1601,
    n1255,
    n1055,
    n1538
  );


  xor
  g2802
  (
    n2464,
    n1373,
    n1772,
    n775,
    n1507
  );


  nor
  g2803
  (
    n2775,
    n844,
    n982,
    n776,
    n1727
  );


  nand
  g2804
  (
    n2820,
    n1009,
    n1372,
    n1354,
    n1200
  );


  nor
  g2805
  (
    n2561,
    n1596,
    n876,
    n1877,
    n839
  );


  xnor
  g2806
  (
    n2386,
    n1058,
    n984,
    n945,
    n751
  );


  or
  g2807
  (
    n2839,
    n1174,
    n1535,
    n1262,
    n1791
  );


  xnor
  g2808
  (
    n2321,
    n1335,
    n855,
    n1351,
    n1455
  );


  nor
  g2809
  (
    n2380,
    n1616,
    n1732,
    n1645,
    n841
  );


  and
  g2810
  (
    n2824,
    n873,
    n795,
    n1224,
    n1005
  );


  nor
  g2811
  (
    n2789,
    n735,
    n1811,
    n827,
    n1495
  );


  xnor
  g2812
  (
    n2323,
    n1283,
    n1151,
    n956,
    n1665
  );


  and
  g2813
  (
    n2355,
    n1620,
    n1673,
    n1333,
    n1470
  );


  xnor
  g2814
  (
    n2741,
    n1361,
    n1066,
    n824,
    n1820
  );


  xor
  g2815
  (
    n2861,
    n1140,
    n784,
    n878,
    n1579
  );


  nand
  g2816
  (
    n2325,
    n1731,
    n1497,
    n1130,
    n1243
  );


  nor
  g2817
  (
    n2382,
    n1321,
    n1375,
    n1496,
    n1756
  );


  xor
  g2818
  (
    n2711,
    n1126,
    n1746,
    n981,
    n1221
  );


  or
  g2819
  (
    n2549,
    n1358,
    n1362,
    n1284,
    n1315
  );


  or
  g2820
  (
    n2465,
    n1756,
    n1854,
    n1305,
    n1257
  );


  nand
  g2821
  (
    n2484,
    n1878,
    n1027,
    n1591,
    n1618
  );


  nand
  g2822
  (
    n2487,
    n1159,
    n1056,
    n1331,
    n1466
  );


  xor
  g2823
  (
    n2621,
    n902,
    n743,
    n1707,
    n1236
  );


  xor
  g2824
  (
    n2440,
    n1232,
    n1423,
    n836,
    n981
  );


  xnor
  g2825
  (
    n2632,
    n1696,
    n906,
    n1382,
    n1265
  );


  and
  g2826
  (
    n2319,
    n1207,
    n1639,
    n923,
    n1853
  );


  and
  g2827
  (
    n2574,
    n1531,
    n1322,
    n776,
    n1769
  );


  and
  g2828
  (
    n2666,
    n1684,
    n1416,
    n1467,
    n1667
  );


  and
  g2829
  (
    n2681,
    n1190,
    n890,
    n1066,
    n1326
  );


  xnor
  g2830
  (
    n2377,
    n1129,
    n813,
    n1718,
    n1724
  );


  nor
  g2831
  (
    n2537,
    n1886,
    n1501,
    n1776,
    n1836
  );


  nor
  g2832
  (
    n2576,
    n1613,
    n1293,
    n887,
    n842
  );


  and
  g2833
  (
    n2793,
    n1043,
    n787,
    n1205,
    n1045
  );


  nor
  g2834
  (
    n2668,
    n1777,
    n1884,
    n1656,
    n1022
  );


  or
  g2835
  (
    n2389,
    n1245,
    n829,
    n764,
    n736
  );


  nor
  g2836
  (
    n2889,
    n1260,
    n1683,
    n1162,
    n1561
  );


  and
  g2837
  (
    n2617,
    n868,
    n1116,
    n1562,
    n852
  );


  nand
  g2838
  (
    n2879,
    n851,
    n1484,
    n1310,
    n1175
  );


  xor
  g2839
  (
    n2359,
    n1883,
    n1155,
    n1304,
    n1340
  );


  xnor
  g2840
  (
    n2541,
    n1817,
    n904,
    n1752,
    n1401
  );


  or
  g2841
  (
    n2600,
    n920,
    n1566,
    n1216,
    n1594
  );


  or
  g2842
  (
    n2690,
    n950,
    n1724,
    n1370,
    n1263
  );


  xnor
  g2843
  (
    n2714,
    n922,
    n1018,
    n1193,
    n1551
  );


  nor
  g2844
  (
    n2595,
    n1440,
    n1063,
    n753,
    n1095
  );


  nor
  g2845
  (
    n2409,
    n1363,
    n1441,
    n1767,
    n1670
  );


  and
  g2846
  (
    n2629,
    n1496,
    n970,
    n1784,
    n1280
  );


  and
  g2847
  (
    n2398,
    n1311,
    n1701,
    n1866,
    n1855
  );


  and
  g2848
  (
    n2761,
    n1616,
    n814,
    n1661,
    n919
  );


  xor
  g2849
  (
    n2445,
    n1851,
    n782,
    n1874,
    n780
  );


  nor
  g2850
  (
    n2731,
    n1385,
    n1117,
    n1782,
    n909
  );


  nand
  g2851
  (
    n2483,
    n1106,
    n1786,
    n909,
    n771
  );


  and
  g2852
  (
    n2451,
    n1426,
    n1093,
    n1896,
    n1381
  );


  nor
  g2853
  (
    n2437,
    n765,
    n828,
    n1178,
    n1348
  );


  nor
  g2854
  (
    n2392,
    n874,
    n1021,
    n1825,
    n732
  );


  and
  g2855
  (
    n2312,
    n1464,
    n829,
    n1327,
    n995
  );


  or
  g2856
  (
    n2439,
    n1067,
    n1433,
    n997,
    n1375
  );


  or
  g2857
  (
    n2702,
    n899,
    n1184,
    n968,
    n1671
  );


  or
  g2858
  (
    n2795,
    n824,
    n1136,
    n1199,
    n1265
  );


  xor
  g2859
  (
    n2662,
    n1658,
    n748,
    n1788,
    n847
  );


  xnor
  g2860
  (
    n2560,
    n810,
    n1533,
    n1888,
    n1194
  );


  nor
  g2861
  (
    n2548,
    n1783,
    n1230,
    n855,
    n1352
  );


  xor
  g2862
  (
    n2868,
    n835,
    n1547,
    n1318,
    n740
  );


  and
  g2863
  (
    n2708,
    n1238,
    n1139,
    n1046,
    n1591
  );


  nand
  g2864
  (
    n2491,
    n1762,
    n1655,
    n1828,
    n1848
  );


  xnor
  g2865
  (
    n2757,
    n958,
    n1508,
    n1668,
    n1122
  );


  xnor
  g2866
  (
    n2796,
    n1610,
    n1382,
    n1870,
    n1849
  );


  nand
  g2867
  (
    n2499,
    n1206,
    n1062,
    n1106,
    n1148
  );


  nor
  g2868
  (
    n2424,
    n1544,
    n1570,
    n1458,
    n1787
  );


  nor
  g2869
  (
    n2642,
    n1107,
    n761,
    n1196,
    n1261
  );


  nand
  g2870
  (
    n2902,
    n1900,
    n2366,
    n2482,
    n2307
  );


  xor
  g2871
  (
    n2906,
    n2467,
    n2327,
    n2312,
    n2425
  );


  and
  g2872
  (
    n2893,
    n2481,
    n2470,
    n2458,
    n2486
  );


  xor
  g2873
  (
    n2901,
    n2305,
    n2500,
    n2499,
    n2440
  );


  or
  g2874
  (
    n2899,
    n2415,
    n2455,
    n2402,
    n2419
  );


  or
  g2875
  (
    n2895,
    n2480,
    n1909,
    n2464,
    n2420
  );


  xnor
  g2876
  (
    n2919,
    n2447,
    n2308,
    n2475,
    n2370
  );


  or
  g2877
  (
    n2930,
    n1905,
    n2429,
    n2381,
    n2463
  );


  xnor
  g2878
  (
    n2941,
    n1907,
    n1906,
    n2477,
    n1901
  );


  nand
  g2879
  (
    n2896,
    n2501,
    n2365,
    n2414,
    n2445
  );


  nor
  g2880
  (
    n2937,
    n1908,
    n2433,
    n2483,
    n2442
  );


  nor
  g2881
  (
    n2942,
    n2472,
    n2399,
    n2401,
    n2346
  );


  nor
  g2882
  (
    n2926,
    n2311,
    n1900,
    n2310,
    n2319
  );


  and
  g2883
  (
    n2921,
    n2394,
    n2434,
    n1903,
    n2372
  );


  or
  g2884
  (
    n2891,
    n2352,
    n2484,
    n2396,
    n2323
  );


  and
  g2885
  (
    n2903,
    n2378,
    n2485,
    n2334,
    n2417
  );


  nor
  g2886
  (
    n2925,
    n2450,
    n2367,
    n2495,
    n2453
  );


  xnor
  g2887
  (
    n2911,
    n2331,
    n2329,
    n2479,
    n2322
  );


  nand
  g2888
  (
    n2908,
    n2416,
    n2471,
    n2386,
    n2318
  );


  xor
  g2889
  (
    n2892,
    n2324,
    n1901,
    n2466,
    n2326
  );


  xnor
  g2890
  (
    n2917,
    n2493,
    n2462,
    n2314,
    n2391
  );


  or
  g2891
  (
    n2936,
    n2379,
    n2474,
    n2451,
    n2347
  );


  nor
  g2892
  (
    n2933,
    n2380,
    n1905,
    n2338,
    n2337
  );


  nor
  g2893
  (
    n2943,
    n2444,
    n2358,
    n2357,
    n2342
  );


  or
  g2894
  (
    n2929,
    n1910,
    n1902,
    n2349,
    n2339
  );


  nor
  g2895
  (
    n2939,
    n2397,
    n2344,
    n2321,
    n2393
  );


  and
  g2896
  (
    n2907,
    n1904,
    n2497,
    n2385,
    n2377
  );


  and
  g2897
  (
    n2904,
    n2387,
    n2454,
    n2388,
    n2461
  );


  nor
  g2898
  (
    n2900,
    n1911,
    n2333,
    n2498,
    n2427
  );


  xor
  g2899
  (
    n2946,
    n2423,
    n2439,
    n1909,
    n2418
  );


  or
  g2900
  (
    n2912,
    n2361,
    n2487,
    n2309,
    n2428
  );


  xnor
  g2901
  (
    n2916,
    n2383,
    n2476,
    n2316,
    n2489
  );


  and
  g2902
  (
    n2910,
    n2448,
    n2407,
    n2375,
    n1910
  );


  nor
  g2903
  (
    n2918,
    n1907,
    n2435,
    n2494,
    n2356
  );


  xor
  g2904
  (
    n2932,
    n2320,
    n2465,
    n2496,
    n2469
  );


  nand
  g2905
  (
    n2898,
    n2354,
    n2313,
    n1902,
    n2353
  );


  or
  g2906
  (
    n2905,
    n2436,
    n2408,
    n2376,
    n2390
  );


  xnor
  g2907
  (
    n2914,
    n2413,
    n2371,
    n2317,
    n2395
  );


  and
  g2908
  (
    n2897,
    n2410,
    n2431,
    n2369,
    n2332
  );


  or
  g2909
  (
    n2924,
    n2340,
    n2335,
    n2432,
    n2409
  );


  xnor
  g2910
  (
    n2913,
    n2345,
    n2382,
    n2325,
    n2443
  );


  xor
  g2911
  (
    n2931,
    n2426,
    n2304,
    n2430,
    n2459
  );


  nand
  g2912
  (
    n2945,
    n2421,
    n2441,
    n2360,
    n2460
  );


  and
  g2913
  (
    n2909,
    n2384,
    n2392,
    n2336,
    n1903
  );


  xor
  g2914
  (
    n2938,
    n2412,
    n2303,
    n2364,
    n2449
  );


  xnor
  g2915
  (
    n2922,
    n2424,
    n2438,
    n2457,
    n2363
  );


  nor
  g2916
  (
    n2923,
    n2355,
    n2328,
    n2473,
    n2343
  );


  xor
  g2917
  (
    n2934,
    n2350,
    n2374,
    n2348,
    n2406
  );


  xnor
  g2918
  (
    n2920,
    n2403,
    n2411,
    n2405,
    n1904
  );


  xnor
  g2919
  (
    n2894,
    n2488,
    n2478,
    n2490,
    n2330
  );


  or
  g2920
  (
    n2944,
    n2492,
    n2351,
    n2468,
    n2373
  );


  xor
  g2921
  (
    n2928,
    n2368,
    n2359,
    n2456,
    n2502
  );


  nor
  g2922
  (
    n2915,
    n2437,
    n2398,
    n2452,
    n2389
  );


  nor
  g2923
  (
    n2940,
    n2400,
    n2422,
    n2315,
    n1908
  );


  nand
  g2924
  (
    n2935,
    n2404,
    n1906,
    n2341,
    n2503
  );


  or
  g2925
  (
    n2927,
    n2306,
    n2446,
    n2491,
    n2362
  );


  nor
  g2926
  (
    n2948,
    n1971,
    n1948,
    n1942,
    n2545
  );


  and
  g2927
  (
    n3016,
    n1978,
    n1940,
    n1957,
    n1980
  );


  xnor
  g2928
  (
    n3009,
    n1953,
    n1916,
    n1969,
    n1936
  );


  or
  g2929
  (
    n3024,
    n1930,
    n1973,
    n1917,
    n1947
  );


  nor
  g2930
  (
    n3029,
    n1953,
    n2932,
    n2581,
    n1984
  );


  xnor
  g2931
  (
    n3015,
    n1946,
    n2548,
    n2557,
    n2574
  );


  or
  g2932
  (
    n2951,
    n2938,
    n1948,
    n1952,
    n1951
  );


  xor
  g2933
  (
    n2989,
    n1960,
    n1997,
    n2906,
    n2556
  );


  nor
  g2934
  (
    n3007,
    n2939,
    n2570,
    n1987,
    n2534
  );


  or
  g2935
  (
    n2968,
    n1940,
    n1918,
    n1966,
    n1949
  );


  or
  g2936
  (
    n3008,
    n2918,
    n2579,
    n2546,
    n1994
  );


  nor
  g2937
  (
    n2964,
    n1960,
    n2922,
    n1921,
    n2555
  );


  nor
  g2938
  (
    n2973,
    n1970,
    n2945,
    n2544,
    n2930
  );


  nor
  g2939
  (
    n2993,
    n2908,
    n1968,
    n1958,
    n1974
  );


  nor
  g2940
  (
    n2960,
    n1954,
    n2580,
    n1975,
    n1945
  );


  xor
  g2941
  (
    n3013,
    n2899,
    n2519,
    n1930,
    n1922
  );


  xnor
  g2942
  (
    n2967,
    n2900,
    n2559,
    n1997,
    n2933
  );


  nand
  g2943
  (
    n2959,
    n1936,
    n2530,
    n2915,
    n1972
  );


  xor
  g2944
  (
    n2980,
    n1973,
    n1938,
    n2937,
    n1962
  );


  nor
  g2945
  (
    n3010,
    n1933,
    n1915,
    n2933,
    n1938
  );


  nand
  g2946
  (
    n3025,
    n2894,
    n1945,
    n1923,
    n2543
  );


  or
  g2947
  (
    n2995,
    n1987,
    n1931,
    n2940,
    n2567
  );


  nand
  g2948
  (
    n2956,
    n1959,
    n1982,
    n1935,
    n2525
  );


  nor
  g2949
  (
    n2953,
    n1957,
    n1941,
    n2898,
    n2936
  );


  or
  g2950
  (
    n2971,
    n2577,
    n1929,
    n2514,
    n1914
  );


  nand
  g2951
  (
    n2977,
    n2515,
    n1961,
    n1989,
    n2554
  );


  xnor
  g2952
  (
    n2974,
    n1932,
    n2944,
    n2902,
    n2578
  );


  nor
  g2953
  (
    n3011,
    n1992,
    n1962,
    n1966,
    n1956
  );


  xnor
  g2954
  (
    n2999,
    n2513,
    n2934,
    n2538,
    n1970
  );


  nand
  g2955
  (
    n2972,
    n2910,
    n1975,
    n2517,
    n2917
  );


  nor
  g2956
  (
    n2970,
    n1933,
    n1993,
    n1986,
    n1996
  );


  xor
  g2957
  (
    KeyWire_0_31,
    n2524,
    n1928,
    n1912,
    n2914
  );


  and
  g2958
  (
    n2952,
    n2893,
    n2528,
    n1937,
    n2518
  );


  nand
  g2959
  (
    n2978,
    n2568,
    n1935,
    n2533,
    n2912
  );


  or
  g2960
  (
    n2979,
    n2507,
    n1920,
    n1963,
    n1926
  );


  or
  g2961
  (
    n2954,
    n1984,
    n2941,
    n1959
  );


  nor
  g2962
  (
    n3018,
    n2521,
    n1969,
    n2535,
    n2541
  );


  xnor
  g2963
  (
    n2982,
    n2921,
    n2509,
    n1950,
    n2923
  );


  or
  g2964
  (
    n3028,
    n2916,
    n1982,
    n2566,
    n2897
  );


  nand
  g2965
  (
    n2998,
    n2508,
    n1980,
    n2549,
    n2942
  );


  nor
  g2966
  (
    n2950,
    n2935,
    n2553,
    n2919,
    n1919
  );


  or
  g2967
  (
    n2994,
    n1925,
    n2511,
    n1979,
    n1947
  );


  nand
  g2968
  (
    n3022,
    n2576,
    n2920,
    n1961,
    n1990
  );


  and
  g2969
  (
    n3004,
    n1920,
    n1964,
    n1952,
    n1985
  );


  xor
  g2970
  (
    n2947,
    n2942,
    n1916,
    n1934,
    n2933
  );


  xnor
  g2971
  (
    n2962,
    n1954,
    n1942,
    n1989,
    n2896
  );


  xor
  g2972
  (
    n2990,
    n1925,
    n2940,
    n1977,
    n1941
  );


  xor
  g2973
  (
    n2957,
    n2526,
    n2523,
    n1955,
    n1944
  );


  and
  g2974
  (
    n2961,
    n2512,
    n2936,
    n2561,
    n2505
  );


  nor
  g2975
  (
    n3026,
    n2901,
    n2529,
    n1939,
    n2931
  );


  nand
  g2976
  (
    n3006,
    n2909,
    n2940,
    n1988,
    n2536
  );


  or
  g2977
  (
    n2976,
    n1996,
    n1924,
    n2931,
    n2504
  );


  or
  g2978
  (
    n2969,
    n2938,
    n2506,
    n1972,
    n1914
  );


  xnor
  g2979
  (
    n3014,
    n2562,
    n2941,
    n1992,
    n1990
  );


  and
  g2980
  (
    n3027,
    n1913,
    n1911,
    n2935,
    n2904
  );


  nor
  g2981
  (
    n2966,
    n2895,
    n2542,
    n2934,
    n1927
  );


  and
  g2982
  (
    n2988,
    n2937,
    n2891,
    n2532,
    n1924
  );


  or
  g2983
  (
    n2991,
    n1976,
    n1919,
    n1983,
    n2552
  );


  nand
  g2984
  (
    n3019,
    n1977,
    n2522,
    n1926,
    n1991
  );


  xor
  g2985
  (
    n2955,
    n1918,
    n1951,
    n1978,
    n1964
  );


  nand
  g2986
  (
    n2963,
    n2563,
    n1923,
    n1946,
    n2926
  );


  xnor
  g2987
  (
    n3000,
    n1949,
    n1956,
    n2943,
    n1967
  );


  xor
  g2988
  (
    n2986,
    n1922,
    n1995,
    n1915,
    n2937
  );


  nor
  g2989
  (
    n2965,
    n1912,
    n2930,
    n2551,
    n2565
  );


  nor
  g2990
  (
    n2984,
    n2928,
    n1927,
    n2943,
    n2560
  );


  nor
  g2991
  (
    n3017,
    n2571,
    n2934,
    n1976,
    n2913
  );


  nor
  g2992
  (
    n3002,
    n1994,
    n2944,
    n2945,
    n2943
  );


  and
  g2993
  (
    n3020,
    n1958,
    n2945,
    n2925,
    n1944
  );


  nand
  g2994
  (
    n2981,
    n2539,
    n2938,
    n2939,
    n2942
  );


  xor
  g2995
  (
    n3003,
    n1913,
    n1981,
    n1993,
    n1955
  );


  nand
  g2996
  (
    n2996,
    n2905,
    n2510,
    n2527,
    n1986
  );


  xor
  g2997
  (
    n2997,
    n1928,
    n2573,
    n1967,
    n1937
  );


  and
  g2998
  (
    n3021,
    n2537,
    n1939,
    n2929,
    n2575
  );


  nor
  g2999
  (
    n3001,
    n2935,
    n2944,
    n1929,
    n1983
  );


  nand
  g3000
  (
    n2992,
    n2903,
    n1932,
    n1921,
    n1968
  );


  nand
  g3001
  (
    n2975,
    n2569,
    n2572,
    n1981,
    n2550
  );


  nor
  g3002
  (
    n3012,
    n1943,
    n1965,
    n1979,
    n1991
  );


  and
  g3003
  (
    n3030,
    n1985,
    n2564,
    n1934,
    n1974
  );


  nand
  g3004
  (
    n2949,
    n2924,
    n1931,
    n1917,
    n2907
  );


  or
  g3005
  (
    n2987,
    n1971,
    n1963,
    n2927,
    n2939
  );


  nor
  g3006
  (
    n2983,
    n1943,
    n1965,
    n2936,
    n2932
  );


  or
  g3007
  (
    n2985,
    n2558,
    n2531,
    n2516,
    n1950
  );


  xor
  g3008
  (
    n3005,
    n1995,
    n2520,
    n2540,
    n1988
  );


  xor
  g3009
  (
    n3023,
    n2547,
    n1998,
    n2911,
    n2892
  );


  and
  g3010
  (
    n3032,
    n2957,
    n2986,
    n2947,
    n2985
  );


  or
  g3011
  (
    n3045,
    n2970,
    n2985,
    n2954,
    n2983
  );


  xor
  g3012
  (
    n3049,
    n2958,
    n2984,
    n2974,
    n2965
  );


  nand
  g3013
  (
    n3031,
    n2985,
    n2982,
    n2966,
    n2979
  );


  xnor
  g3014
  (
    n3050,
    n2950,
    n2981,
    n2963,
    n2990
  );


  nand
  g3015
  (
    n3039,
    n2978,
    n2980,
    n2953,
    n2955
  );


  nand
  g3016
  (
    n3041,
    n2977,
    n2987,
    n2949,
    n2989
  );


  xor
  g3017
  (
    n3036,
    n1999,
    n2977,
    n2986,
    n2983
  );


  xnor
  g3018
  (
    n3046,
    n2989,
    n2979,
    n2976,
    n2973
  );


  or
  g3019
  (
    n3047,
    n2982,
    n2984,
    n2969,
    n2948
  );


  or
  g3020
  (
    n3034,
    n2991,
    n2000,
    n2978,
    n2976
  );


  or
  g3021
  (
    n3042,
    n2980,
    n2968,
    n1998,
    n2972
  );


  and
  g3022
  (
    n3038,
    n2989,
    n2975,
    n2977,
    n2000
  );


  xnor
  g3023
  (
    n3033,
    n2971,
    n2980,
    n2976,
    n2961
  );


  nor
  g3024
  (
    n3044,
    n2967,
    n2984,
    n2986,
    n2982
  );


  and
  g3025
  (
    n3037,
    n2960,
    n2952,
    n2964,
    n2962
  );


  xor
  g3026
  (
    n3035,
    n2988,
    n2990,
    n2979,
    n2956
  );


  xnor
  g3027
  (
    n3040,
    n2951,
    n2988,
    n2981,
    n1999
  );


  xor
  g3028
  (
    n3043,
    n2988,
    n2959,
    n2990,
    n2981
  );


  xnor
  g3029
  (
    n3048,
    n2978,
    n2983,
    n2987
  );


  nand
  g3030
  (
    n3058,
    n3043,
    n2002,
    n2007
  );


  nor
  g3031
  (
    n3062,
    n2009,
    n3047,
    n2012,
    n2013
  );


  xnor
  g3032
  (
    n3051,
    n2019,
    n2001,
    n2008,
    n2003
  );


  or
  g3033
  (
    n3061,
    n2011,
    n2003,
    n2002,
    n3038
  );


  xnor
  g3034
  (
    n3052,
    n2011,
    n2015,
    n2017,
    n2008
  );


  nand
  g3035
  (
    n3060,
    n3045,
    n2013,
    n2010,
    n3037
  );


  or
  g3036
  (
    n3057,
    n2004,
    n3044,
    n2009,
    n2001
  );


  nand
  g3037
  (
    n3059,
    n2015,
    n2017,
    n3040,
    n3036
  );


  nor
  g3038
  (
    n3063,
    n2016,
    n3041,
    n2014,
    n2010
  );


  nor
  g3039
  (
    n3055,
    n2014,
    n3046,
    n3035,
    n3042
  );


  xor
  g3040
  (
    n3056,
    n2006,
    n2006,
    n2019,
    n2012
  );


  xor
  g3041
  (
    n3053,
    n2007,
    n2005,
    n2018,
    n2004
  );


  nor
  g3042
  (
    n3054,
    n2005,
    n2018,
    n3039,
    n2016
  );


  xnor
  g3043
  (
    n3073,
    n2038,
    n2021,
    n3054,
    n2042
  );


  and
  g3044
  (
    n3069,
    n3057,
    n2033,
    n2025,
    n2021
  );


  xor
  g3045
  (
    n3072,
    n2036,
    n2035,
    n3052,
    n2034
  );


  nor
  g3046
  (
    n3068,
    n2039,
    n2032,
    n2020,
    n2027
  );


  nand
  g3047
  (
    n3064,
    n2022,
    n3060,
    n2023,
    n2030
  );


  nand
  g3048
  (
    n3078,
    n3062,
    n2035,
    n2037,
    n3063
  );


  xnor
  g3049
  (
    n3076,
    n2030,
    n3062,
    n3059,
    n2031
  );


  nand
  g3050
  (
    n3075,
    n3063,
    n2038,
    n2028,
    n2040
  );


  or
  g3051
  (
    n3070,
    n2031,
    n2025,
    n2020,
    n2041
  );


  or
  g3052
  (
    n3065,
    n2033,
    n2028,
    n2022,
    n2039
  );


  or
  g3053
  (
    n3067,
    n2027,
    n2029,
    n2036,
    n3061
  );


  nor
  g3054
  (
    n3066,
    n2026,
    n3056,
    n2041,
    n2024
  );


  nor
  g3055
  (
    n3071,
    n2023,
    n3051,
    n2024,
    n2040
  );


  xnor
  g3056
  (
    n3074,
    n2026,
    n2032,
    n3053,
    n3055
  );


  and
  g3057
  (
    n3077,
    n2029,
    n3058,
    n2037,
    n2034
  );


  or
  g3058
  (
    n3082,
    n2586,
    n2600,
    n2599,
    n3069
  );


  nand
  g3059
  (
    n3087,
    n2612,
    n3067,
    n2603,
    n2616
  );


  nand
  g3060
  (
    n3091,
    n2589,
    n2596,
    n2593,
    n2582
  );


  xnor
  g3061
  (
    n3092,
    n2615,
    n2606,
    n2584,
    n3070
  );


  nand
  g3062
  (
    n3085,
    n2614,
    n2622,
    n2618,
    n3070
  );


  xor
  g3063
  (
    n3084,
    n3065,
    n2617,
    n2583,
    n3068
  );


  and
  g3064
  (
    n3081,
    n2613,
    n2605,
    n3071,
    n2594
  );


  nor
  g3065
  (
    n3090,
    n3066,
    n2611,
    n3067,
    n3072
  );


  nand
  g3066
  (
    n3089,
    n3064,
    n2609,
    n2621,
    n3071
  );


  xnor
  g3067
  (
    n3080,
    n2595,
    n2620,
    n2601,
    n2623
  );


  xor
  g3068
  (
    n3086,
    n2597,
    n2585,
    n2602,
    n2607
  );


  or
  g3069
  (
    n3088,
    n3069,
    n3068,
    n2598,
    n2588
  );


  xor
  g3070
  (
    n3083,
    n2587,
    n2608,
    n2610,
    n2604
  );


  xor
  g3071
  (
    n3079,
    n2591,
    n2590,
    n2592,
    n2619
  );


  xor
  g3072
  (
    n3093,
    n3081,
    n3005,
    n3006,
    n3085
  );


  and
  g3073
  (
    n3116,
    n3003,
    n2999,
    n2994,
    n3080
  );


  or
  g3074
  (
    n3096,
    n3085,
    n3005,
    n3073,
    n2994
  );


  or
  g3075
  (
    n3105,
    n3074,
    n3000,
    n3081,
    n2998
  );


  nand
  g3076
  (
    n3102,
    n2998,
    n3088,
    n2995,
    n2045
  );


  nand
  g3077
  (
    n3110,
    n3001,
    n2044,
    n3086,
    n3088
  );


  nor
  g3078
  (
    n3107,
    n3084,
    n3074,
    n2993,
    n3082
  );


  nor
  g3079
  (
    n3095,
    n2993,
    n2998,
    n2997,
    n3087
  );


  and
  g3080
  (
    n3098,
    n2049,
    n3003,
    n2043,
    n3000
  );


  xnor
  g3081
  (
    n3103,
    n3079,
    n2991,
    n3088,
    n3084
  );


  xnor
  g3082
  (
    n3097,
    n3001,
    n2047,
    n2049,
    n3087
  );


  xnor
  g3083
  (
    n3101,
    n3082,
    n2994,
    n2999,
    n2992
  );


  or
  g3084
  (
    n3106,
    n2997,
    n2996,
    n2995,
    n2045
  );


  xnor
  g3085
  (
    n3104,
    n2991,
    n2992,
    n2999,
    n3079
  );


  xnor
  g3086
  (
    n3108,
    n2048,
    n3004,
    n3002
  );


  xnor
  g3087
  (
    n3115,
    n3083,
    n2997,
    n3003,
    n2042
  );


  and
  g3088
  (
    n3111,
    n2048,
    n2050,
    n107,
    n3081
  );


  nor
  g3089
  (
    n3100,
    n2992,
    n3083,
    n3004
  );


  and
  g3090
  (
    n3114,
    n3072,
    n2044,
    n3005,
    n2996
  );


  or
  g3091
  (
    n3099,
    n2996,
    n3087,
    n3084,
    n3086
  );


  xnor
  g3092
  (
    n3109,
    n3001,
    n3073,
    n3082,
    n2995
  );


  or
  g3093
  (
    n3112,
    n2043,
    n2046,
    n2624
  );


  nor
  g3094
  (
    n3113,
    n3085,
    n3000,
    n3086,
    n3002
  );


  nand
  g3095
  (
    n3094,
    n2047,
    n2993,
    n3004,
    n3080
  );


  buf
  g3096
  (
    n3129,
    n3094
  );


  buf
  g3097
  (
    n3117,
    n3007
  );


  not
  g3098
  (
    n3127,
    n3008
  );


  not
  g3099
  (
    n3128,
    n3097
  );


  buf
  g3100
  (
    n3125,
    n3009
  );


  not
  g3101
  (
    n3130,
    n3010
  );


  not
  g3102
  (
    n3120,
    n3101
  );


  not
  g3103
  (
    n3131,
    n3106
  );


  not
  g3104
  (
    n3118,
    n3108
  );


  buf
  g3105
  (
    n3124,
    n3009
  );


  not
  g3106
  (
    n3121,
    n3009
  );


  buf
  g3107
  (
    n3132,
    n3007
  );


  xor
  g3108
  (
    n3119,
    n3006,
    n3008,
    n3100,
    n3099
  );


  or
  g3109
  (
    n3122,
    n3107,
    n3008,
    n3006,
    n3096
  );


  or
  g3110
  (
    n3126,
    n3105,
    n3102,
    n3095,
    n3007
  );


  nand
  g3111
  (
    n3123,
    n3103,
    n3104,
    n3093,
    n3098
  );


  buf
  g3112
  (
    n3153,
    n3124
  );


  not
  g3113
  (
    n3150,
    n3122
  );


  not
  g3114
  (
    n3134,
    n3118
  );


  not
  g3115
  (
    n3135,
    n3119
  );


  buf
  g3116
  (
    n3151,
    n3120
  );


  not
  g3117
  (
    n3136,
    n3124
  );


  buf
  g3118
  (
    n3147,
    n3130
  );


  not
  g3119
  (
    n3133,
    n3127
  );


  buf
  g3120
  (
    n3154,
    n3129
  );


  not
  g3121
  (
    n3148,
    n3123
  );


  not
  g3122
  (
    n3139,
    n3129
  );


  not
  g3123
  (
    n3152,
    n3049
  );


  buf
  g3124
  (
    n3146,
    n3125
  );


  not
  g3125
  (
    n3142,
    n3128
  );


  buf
  g3126
  (
    n3156,
    n3123
  );


  buf
  g3127
  (
    n3138,
    n3125
  );


  nand
  g3128
  (
    n3157,
    n3130,
    n3132,
    n3010,
    n3048
  );


  nand
  g3129
  (
    n3144,
    n3126,
    n3118,
    n3122,
    n3119
  );


  nor
  g3130
  (
    n3149,
    n3128,
    n3123,
    n3121,
    n3127
  );


  xnor
  g3131
  (
    n3140,
    n3132,
    n3131,
    n3126,
    n3125
  );


  xnor
  g3132
  (
    n3137,
    n3131,
    n3129,
    n3118,
    n3120
  );


  xor
  g3133
  (
    n3145,
    n3010,
    n3117,
    n3121
  );


  and
  g3134
  (
    n3141,
    n3122,
    n3011,
    n3130,
    n3126
  );


  or
  g3135
  (
    n3143,
    n3128,
    n3050,
    n3132,
    n3119
  );


  xor
  g3136
  (
    n3155,
    n3131,
    n3124,
    n3120,
    n3127
  );


  xnor
  g3137
  (
    n3166,
    n3150,
    n3149,
    n3133,
    n3137
  );


  and
  g3138
  (
    n3163,
    n3142,
    n3136,
    n3139,
    n3146
  );


  and
  g3139
  (
    n3159,
    n3150,
    n3134,
    n2050
  );


  and
  g3140
  (
    n3158,
    n3147,
    n3145,
    n3150,
    n3137
  );


  nand
  g3141
  (
    n3169,
    n3148,
    n3135,
    n3138,
    n3145
  );


  xor
  g3142
  (
    n3165,
    n3135,
    n3138,
    n3141
  );


  nand
  g3143
  (
    n3170,
    n3136,
    n3143,
    n3133
  );


  nand
  g3144
  (
    n3161,
    n3139,
    n3149,
    n3134,
    n3138
  );


  or
  g3145
  (
    n3171,
    n3147,
    n3149,
    n3148,
    n3144
  );


  xnor
  g3146
  (
    n3167,
    n3145,
    n3140,
    n3133,
    n3146
  );


  xor
  g3147
  (
    n3164,
    n3151,
    n3140,
    n3144,
    n3135
  );


  xor
  g3148
  (
    n3162,
    n3137,
    n3150,
    n3143,
    n3147
  );


  nor
  g3149
  (
    n3172,
    n3148,
    n3141,
    n3140,
    n3136
  );


  xor
  g3150
  (
    n3168,
    n3148,
    n3142,
    n3144,
    n3146
  );


  nand
  g3151
  (
    n3160,
    n3151,
    n3139,
    n3149,
    n3142
  );


  and
  g3152
  (
    n3175,
    n2066,
    n2072,
    n2080,
    n2053
  );


  and
  g3153
  (
    n3206,
    n3171,
    n2063,
    n2080,
    n3172
  );


  and
  g3154
  (
    n3183,
    n2061,
    n2097,
    n2068,
    n2054
  );


  xnor
  g3155
  (
    n3205,
    n2093,
    n3161,
    n2092,
    n2100
  );


  and
  g3156
  (
    n3202,
    n3162,
    n2077,
    n2070,
    n3168
  );


  or
  g3157
  (
    n3177,
    n3170,
    n2087,
    n2095,
    n2062
  );


  and
  g3158
  (
    n3185,
    n2094,
    n2091,
    n2084,
    n2069
  );


  or
  g3159
  (
    n3201,
    n3172,
    n2096,
    n2069,
    n2095
  );


  or
  g3160
  (
    n3204,
    n2085,
    n2083,
    n3170,
    n2067
  );


  and
  g3161
  (
    n3180,
    n2051,
    n2065,
    n2091,
    n2085
  );


  xor
  g3162
  (
    n3188,
    n2075,
    n3163,
    n2097,
    n3171
  );


  xor
  g3163
  (
    n3179,
    n3168,
    n2067,
    n2074,
    n3166
  );


  nor
  g3164
  (
    n3173,
    n2088,
    n2096,
    n3161,
    n3158
  );


  xnor
  g3165
  (
    n3196,
    n2068,
    n3159,
    n2087,
    n2070
  );


  nand
  g3166
  (
    n3191,
    n2051,
    n3172,
    n2056,
    n2057
  );


  nor
  g3167
  (
    n3174,
    n2089,
    n2100,
    n3160,
    n3169
  );


  or
  g3168
  (
    n3203,
    n2065,
    n2078,
    n2090,
    n2074
  );


  nor
  g3169
  (
    n3197,
    n2076,
    n2071,
    n2082,
    n2073
  );


  nand
  g3170
  (
    n3186,
    n2098,
    n2063,
    n3167,
    n3162
  );


  nor
  g3171
  (
    n3199,
    n2084,
    n2066,
    n2058,
    n2064
  );


  nor
  g3172
  (
    n3194,
    n2099,
    n2072,
    n2078,
    n3165
  );


  nor
  g3173
  (
    n3195,
    n3165,
    n2081,
    n3158,
    n2090
  );


  or
  g3174
  (
    n3192,
    n2099,
    n2076,
    n2055,
    n3160
  );


  nor
  g3175
  (
    n3187,
    n3159,
    n2082,
    n2054,
    n3163
  );


  xor
  g3176
  (
    n3178,
    n2055,
    n2052,
    n2058,
    n2062
  );


  and
  g3177
  (
    n3176,
    n2094,
    n2086,
    n3164,
    n2101
  );


  nor
  g3178
  (
    n3181,
    n2079,
    n2071,
    n3167,
    n3166
  );


  or
  g3179
  (
    n3182,
    n2057,
    n2101,
    n2061,
    n2052
  );


  xor
  g3180
  (
    n3193,
    n2075,
    n3170,
    n3169,
    n2098
  );


  xor
  g3181
  (
    n3200,
    n2089,
    n2056,
    n2093,
    n3171
  );


  nor
  g3182
  (
    n3190,
    n2064,
    n2059,
    n2088,
    n3169
  );


  or
  g3183
  (
    n3184,
    n2081,
    n2059,
    n2073,
    n3164
  );


  and
  g3184
  (
    n3198,
    n2083,
    n2077,
    n2079,
    n2092
  );


  nand
  g3185
  (
    n3189,
    n2053,
    n2060,
    n2086
  );


  not
  g3186
  (
    n3209,
    n3180
  );


  not
  g3187
  (
    n3215,
    n3173
  );


  not
  g3188
  (
    n3208,
    n3184
  );


  buf
  g3189
  (
    n3219,
    n3177
  );


  not
  g3190
  (
    n3210,
    n3178
  );


  not
  g3191
  (
    n3218,
    n3185
  );


  not
  g3192
  (
    n3216,
    n3181
  );


  not
  g3193
  (
    n3213,
    n3179
  );


  buf
  g3194
  (
    n3214,
    n3183
  );


  buf
  g3195
  (
    n3207,
    n3175
  );


  not
  g3196
  (
    n3220,
    n3187
  );


  not
  g3197
  (
    n3212,
    n3174
  );


  not
  g3198
  (
    n3211,
    n3186
  );


  buf
  g3199
  (
    n3221,
    n3176
  );


  not
  g3200
  (
    n3217,
    n3182
  );


  and
  g3201
  (
    n3236,
    n3156,
    n3215,
    n3157,
    n3207
  );


  or
  g3202
  (
    n3229,
    n3116,
    n2946,
    n3011,
    n3153
  );


  xnor
  g3203
  (
    n3223,
    n3213,
    n3211,
    n3155,
    n3214
  );


  xnor
  g3204
  (
    n3234,
    n3218,
    n3219,
    n3221,
    n3151
  );


  xnor
  g3205
  (
    n3237,
    n3115,
    n3221,
    n3153,
    n2946
  );


  xnor
  g3206
  (
    n3230,
    n3152,
    n3154,
    n3155
  );


  nand
  g3207
  (
    n3222,
    n3153,
    n3115,
    n3157,
    n3219
  );


  and
  g3208
  (
    n3233,
    n2946,
    n3151,
    n3216,
    n3154
  );


  nor
  g3209
  (
    n3228,
    n3110,
    n3116,
    n3112,
    n3111
  );


  xor
  g3210
  (
    n3224,
    n3157,
    n3208,
    n3152
  );


  xor
  g3211
  (
    n3231,
    n3112,
    n3114,
    n3109,
    n3212
  );


  xnor
  g3212
  (
    n3232,
    n3217,
    n3156,
    n3154,
    n3155
  );


  nor
  g3213
  (
    n3226,
    n3114,
    n3218,
    n3153,
    n3157
  );


  xor
  g3214
  (
    n3225,
    n3217,
    n3216,
    n3113,
    n3152
  );


  and
  g3215
  (
    n3235,
    n3156,
    n3220,
    n3209
  );


  nor
  g3216
  (
    n3227,
    n3155,
    n3113,
    n3156,
    n3210
  );


  nor
  g3217
  (
    n3238,
    n2112,
    n2102,
    n2104,
    n2113
  );


  or
  g3218
  (
    n3244,
    n3225,
    n3228,
    n2124,
    n2115
  );


  xnor
  g3219
  (
    n3256,
    n3228,
    n2111,
    n2105,
    n2109
  );


  or
  g3220
  (
    n3254,
    n2116,
    n2125,
    n2105,
    n2123
  );


  xor
  g3221
  (
    n3243,
    n2128,
    n2104,
    n3225,
    n2126
  );


  xnor
  g3222
  (
    n3246,
    n2117,
    n3222,
    n2121,
    n2126
  );


  nor
  g3223
  (
    n3251,
    n2123,
    n2106,
    n2111,
    n3231
  );


  and
  g3224
  (
    n3245,
    n2122,
    n3229,
    n2110,
    n3224
  );


  and
  g3225
  (
    n3255,
    n2108,
    n2124,
    n2127,
    n3230
  );


  xor
  g3226
  (
    n3241,
    n2125,
    n2127,
    n2117,
    n3227
  );


  xor
  g3227
  (
    n3247,
    n2103,
    n2128,
    n2114,
    n2121
  );


  nand
  g3228
  (
    n3248,
    n2120,
    n3230,
    n3223,
    n2118
  );


  nand
  g3229
  (
    n3249,
    n2118,
    n3222,
    n2106,
    n3229
  );


  nor
  g3230
  (
    n3253,
    n2107,
    n2102,
    n2113,
    n3227
  );


  or
  g3231
  (
    n3242,
    n2129,
    n2109,
    n3223,
    n2119
  );


  and
  g3232
  (
    n3250,
    n2103,
    n2108,
    n2110,
    n2116
  );


  or
  g3233
  (
    n3252,
    n2112,
    n3226,
    n2115,
    n2129
  );


  xnor
  g3234
  (
    n3240,
    n2107,
    n2120,
    n2114,
    n2130
  );


  or
  g3235
  (
    n3239,
    n2122,
    n3226,
    n2119,
    n3224
  );


  and
  g3236
  (
    n3265,
    n2625,
    n2658,
    n3239,
    n3241
  );


  xnor
  g3237
  (
    n3269,
    n2629,
    n2639,
    n2627,
    n3241
  );


  xnor
  g3238
  (
    n3260,
    n3240,
    n3242,
    n2643,
    n2632
  );


  or
  g3239
  (
    n3271,
    n2664,
    n2665,
    n2631,
    n2635
  );


  and
  g3240
  (
    n3257,
    n2634,
    n2637,
    n3241,
    n2638
  );


  and
  g3241
  (
    n3264,
    n3243,
    n2668,
    n2660,
    n2667
  );


  nand
  g3242
  (
    n3262,
    n2654,
    n2647,
    n2651,
    n2630
  );


  or
  g3243
  (
    n3263,
    n2663,
    n2656,
    n2653,
    n2662
  );


  xor
  g3244
  (
    n3261,
    n2655,
    n3238,
    n3239,
    n3240
  );


  nor
  g3245
  (
    n3259,
    n2646,
    n3242,
    n2626,
    n2640
  );


  or
  g3246
  (
    n3272,
    n2644,
    n2670,
    n2652,
    n2649
  );


  and
  g3247
  (
    n3267,
    n2641,
    n2648,
    n2636,
    n2645
  );


  xor
  g3248
  (
    n3258,
    n2130,
    n3238,
    n2657,
    n2650
  );


  or
  g3249
  (
    n3268,
    n2671,
    n2669,
    n3238,
    n2642
  );


  and
  g3250
  (
    n3266,
    n2628,
    n2659,
    n3240,
    n3239
  );


  xnor
  g3251
  (
    n3270,
    n2633,
    n2661,
    n2666,
    n3242
  );


  nand
  g3252
  (
    n3273,
    n3257,
    n3258
  );


  not
  g3253
  (
    n3277,
    n3273
  );


  not
  g3254
  (
    n3274,
    n3189
  );


  nor
  g3255
  (
    n3275,
    n3259,
    n3273
  );


  nand
  g3256
  (
    n3276,
    n3190,
    n3273,
    n3188
  );


  and
  g3257
  (
    n3284,
    n3269,
    n3092,
    n3275,
    n3267
  );


  nand
  g3258
  (
    n3280,
    n3267,
    n3091,
    n3266,
    n3265
  );


  and
  g3259
  (
    n3286,
    n3089,
    n3274,
    n3276
  );


  and
  g3260
  (
    n3287,
    n3276,
    n2131,
    n3091,
    n3275
  );


  nand
  g3261
  (
    n3288,
    n3276,
    n3090,
    n3092
  );


  nand
  g3262
  (
    n3285,
    n3264,
    n3263,
    n3090,
    n3092
  );


  xnor
  g3263
  (
    n3281,
    n3265,
    n3262,
    n3089,
    n3091
  );


  xor
  g3264
  (
    n3282,
    n3275,
    n2672,
    n3269
  );


  and
  g3265
  (
    n3278,
    n3089,
    n3268,
    n3261
  );


  xnor
  g3266
  (
    n3279,
    n3275,
    n3262,
    n3266,
    n3274
  );


  and
  g3267
  (
    n3289,
    n3274,
    n3263,
    n3261,
    n3260
  );


  nor
  g3268
  (
    n3283,
    n3260,
    n3274,
    n3259,
    n3264
  );


  or
  g3269
  (
    n3297,
    n2147,
    n2133,
    n2149,
    n2135
  );


  xnor
  g3270
  (
    n3308,
    n2139,
    n2159,
    n3284,
    n2148
  );


  and
  g3271
  (
    n3295,
    n3287,
    n2157,
    n2154,
    n2142
  );


  xor
  g3272
  (
    n3292,
    n2159,
    n2158,
    n2161,
    n2134
  );


  xnor
  g3273
  (
    n3296,
    n3279,
    n2132,
    n3280,
    n2161
  );


  and
  g3274
  (
    n3305,
    n3286,
    n2135,
    n2162,
    n2140
  );


  and
  g3275
  (
    n3301,
    n3284,
    n2131,
    n2154,
    n2139
  );


  and
  g3276
  (
    n3309,
    n3285,
    n2137,
    n2152,
    n2138
  );


  nand
  g3277
  (
    n3306,
    n2141,
    n2134,
    n2136,
    n2153
  );


  nand
  g3278
  (
    n3298,
    n3282,
    n2155,
    n2136,
    n3288
  );


  xnor
  g3279
  (
    n3294,
    n2137,
    n3281,
    n2160,
    n2155
  );


  nand
  g3280
  (
    n3310,
    n2142,
    n3283,
    n2151,
    n2150
  );


  xnor
  g3281
  (
    n3300,
    n2147,
    n2141,
    n3278,
    n2145
  );


  nand
  g3282
  (
    n3304,
    n2149,
    n2152,
    n2158,
    n2156
  );


  nor
  g3283
  (
    n3293,
    n2151,
    n2140,
    n2146,
    n3278
  );


  or
  g3284
  (
    n3303,
    n3279,
    n2144,
    n3286,
    n3283
  );


  nand
  g3285
  (
    n3290,
    n2143,
    n2133,
    n2145,
    n2138
  );


  or
  g3286
  (
    n3302,
    n3285,
    n2144,
    n2148,
    n2162
  );


  nand
  g3287
  (
    n3291,
    n2160,
    n2150,
    n2157,
    n3287
  );


  nor
  g3288
  (
    n3307,
    n3281,
    n3282,
    n2156,
    n2153
  );


  and
  g3289
  (
    n3299,
    n2132,
    n3280,
    n2146,
    n2143
  );


  or
  g3290
  (
    n3314,
    n3246,
    n3290,
    n3250
  );


  xnor
  g3291
  (
    n3320,
    n3249,
    n3295,
    n3293,
    n3252
  );


  xnor
  g3292
  (
    n3318,
    n3255,
    n2678,
    n3250,
    n3247
  );


  nand
  g3293
  (
    n3323,
    n3253,
    n3292,
    n3255,
    n3254
  );


  and
  g3294
  (
    n3326,
    n3256,
    n3292,
    n3252,
    n3294
  );


  and
  g3295
  (
    n3312,
    n2680,
    n3244,
    n3253,
    n3243
  );


  xnor
  g3296
  (
    n3319,
    n3251,
    n3253,
    n3255,
    n3293
  );


  or
  g3297
  (
    n3327,
    n3248,
    n2677,
    n3245,
    n3291
  );


  xnor
  g3298
  (
    n3328,
    n3251,
    n3246,
    n3290,
    n3255
  );


  nand
  g3299
  (
    n3324,
    n3248,
    n3246,
    n3252,
    n3249
  );


  xor
  g3300
  (
    n3325,
    n3254,
    n3245,
    n2676,
    n3248
  );


  nor
  g3301
  (
    n3329,
    n3291,
    n3249,
    n3256
  );


  nor
  g3302
  (
    n3313,
    n3251,
    n3244,
    n3256,
    n2674
  );


  xor
  g3303
  (
    n3321,
    n3256,
    n3291,
    n3244,
    n3292
  );


  or
  g3304
  (
    n3322,
    n3251,
    n3295,
    n2675,
    n3294
  );


  and
  g3305
  (
    n3316,
    n3250,
    n3247,
    n3245,
    n3254
  );


  xor
  g3306
  (
    n3315,
    n3294,
    n3295,
    n2679,
    n3253
  );


  or
  g3307
  (
    n3311,
    n3243,
    n3247,
    n3254,
    n3293
  );


  nor
  g3308
  (
    n3317,
    n3296,
    n3252,
    n3290,
    n2673
  );


  buf
  g3309
  (
    n3330,
    n3311
  );


  not
  g3310
  (
    n3331,
    n3311
  );


  buf
  g3311
  (
    n3332,
    n3312
  );


  buf
  g3312
  (
    KeyWire_0_27,
    n3311
  );


  xnor
  g3313
  (
    n3334,
    n3013,
    n3014,
    n3330,
    n3012
  );


  or
  g3314
  (
    n3336,
    n3013,
    n3330,
    n3014,
    n3011
  );


  and
  g3315
  (
    n3335,
    n3015,
    n3012,
    n3331,
    n3330
  );


  nor
  g3316
  (
    n3337,
    n3013,
    n3014,
    n3015,
    n3012
  );


  or
  g3317
  (
    n3346,
    n3296,
    n3204,
    n3337,
    n3016
  );


  xnor
  g3318
  (
    n3350,
    n3337,
    n3336,
    n3297,
    n3203
  );


  xor
  g3319
  (
    n3352,
    n3298,
    n3198,
    n2681,
    n3334
  );


  or
  g3320
  (
    n3338,
    n3195,
    n3017,
    n3334,
    n2682
  );


  and
  g3321
  (
    n3351,
    n3335,
    n3199,
    n3191,
    n3337
  );


  xor
  g3322
  (
    n3345,
    n3206,
    n3277,
    n3017,
    n3205
  );


  nand
  g3323
  (
    n3342,
    n3337,
    n3296,
    n3298,
    n3299
  );


  nand
  g3324
  (
    n3353,
    n3300,
    n3298,
    n3200,
    n3336
  );


  xor
  g3325
  (
    n3341,
    n3203,
    n3206,
    n3297,
    n2163
  );


  xor
  g3326
  (
    n3349,
    n3192,
    n3277,
    n3017,
    n3202
  );


  nor
  g3327
  (
    n3348,
    n3196,
    n3197,
    n3334,
    n3016
  );


  xor
  g3328
  (
    n3344,
    n3205,
    n3015,
    n3201,
    n3204
  );


  nor
  g3329
  (
    n3343,
    n3016,
    n3202,
    n3335,
    n3194
  );


  xnor
  g3330
  (
    n3339,
    n3193,
    n3277,
    n3335,
    n3334
  );


  xnor
  g3331
  (
    n3347,
    n3277,
    n3299,
    n3201
  );


  nand
  g3332
  (
    n3340,
    n3335,
    n3297,
    n3336
  );


  or
  g3333
  (
    n3354,
    n3351,
    n3288,
    n3352
  );


  nand
  g3334
  (
    n3355,
    n3353,
    n3289
  );


  xnor
  g3335
  (
    n3360,
    n3355,
    n3300,
    n3354,
    n3304
  );


  nand
  g3336
  (
    n3356,
    n3303,
    n3305,
    n3301
  );


  nand
  g3337
  (
    n3359,
    n3304,
    n3303,
    n3302
  );


  or
  g3338
  (
    n3358,
    n3302,
    n3355,
    n3354,
    n3303
  );


  xnor
  g3339
  (
    n3357,
    n3300,
    n3355,
    n3304,
    n3301
  );


  nand
  g3340
  (
    n3361,
    n3313,
    n3356
  );


  or
  g3341
  (
    n3362,
    n3356,
    n3312,
    n3313
  );


  xor
  g3342
  (
    n3363,
    n3361,
    n3270
  );


  buf
  g3343
  (
    n3364,
    n3363
  );


  xnor
  g3344
  (
    n3366,
    n2165,
    n2163,
    n3364
  );


  xor
  g3345
  (
    n3365,
    n2165,
    n2166,
    n2164
  );


  buf
  g3346
  (
    n3370,
    n3365
  );


  not
  g3347
  (
    n3371,
    n3366
  );


  buf
  g3348
  (
    n3368,
    n3365
  );


  buf
  g3349
  (
    n3369,
    n3366
  );


  buf
  g3350
  (
    n3372,
    n3365
  );


  buf
  g3351
  (
    n3367,
    n3366
  );


  or
  g3352
  (
    n3373,
    n3271,
    n3366
  );


  nand
  g3353
  (
    n3374,
    n3369,
    n3358,
    n3357,
    n3359
  );


  nand
  g3354
  (
    n3375,
    n3360,
    n3357,
    n3367
  );


  nor
  g3355
  (
    n3379,
    n3359,
    n3360,
    n3372
  );


  nand
  g3356
  (
    n3378,
    n3368,
    n3360,
    n3359
  );


  and
  g3357
  (
    n3376,
    n3358,
    n3358,
    n3357,
    n3371
  );


  nand
  g3358
  (
    n3377,
    n3358,
    n3356,
    n3370,
    n3305
  );


  or
  g3359
  (
    n3391,
    n3314,
    n3328,
    n3374,
    n3324
  );


  and
  g3360
  (
    n3390,
    n3313,
    n3322,
    n3315
  );


  xnor
  g3361
  (
    n3380,
    n3323,
    n3377,
    n3326
  );


  or
  g3362
  (
    n3397,
    n3328,
    n3319,
    n3320,
    n3327
  );


  xnor
  g3363
  (
    n3396,
    n3319,
    n3322,
    n3379,
    n3378
  );


  and
  g3364
  (
    n3389,
    n3318,
    n3329,
    n3323,
    n3316
  );


  xnor
  g3365
  (
    n3382,
    n3379,
    n3376,
    n3374,
    n3315
  );


  nand
  g3366
  (
    n3400,
    n3375,
    n3316,
    n3361,
    n3329
  );


  and
  g3367
  (
    n3401,
    n3328,
    n3362,
    n3325,
    n3319
  );


  nand
  g3368
  (
    n3398,
    n3379,
    n3323,
    n3326,
    n3322
  );


  nor
  g3369
  (
    n3395,
    n3379,
    n3325,
    n3018,
    n3378
  );


  nor
  g3370
  (
    n3392,
    n3329,
    n3318,
    n3314
  );


  xor
  g3371
  (
    n3388,
    n3315,
    n3327,
    n3317,
    n3324
  );


  or
  g3372
  (
    n3402,
    n3377,
    n3374,
    n3378,
    n3321
  );


  nand
  g3373
  (
    n3383,
    n3323,
    n3377,
    n3319
  );


  xnor
  g3374
  (
    n3386,
    n3376,
    n3318,
    n3329,
    n3320
  );


  xnor
  g3375
  (
    n3385,
    n3317,
    n3362,
    n3374,
    n3328
  );


  and
  g3376
  (
    n3381,
    n3321,
    n3325,
    n3314,
    n3317
  );


  xnor
  g3377
  (
    n3384,
    n3325,
    n3321,
    n3327,
    n3375
  );


  xor
  g3378
  (
    n3387,
    n3315,
    n3320,
    n3376,
    n3375
  );


  or
  g3379
  (
    n3403,
    n3317,
    n3375,
    n3321,
    n3320
  );


  xor
  g3380
  (
    n3399,
    n3324,
    n3378,
    n3326,
    n3316
  );


  nor
  g3381
  (
    n3394,
    n3018,
    n3314,
    n3316,
    n2167
  );


  or
  g3382
  (
    n3393,
    n3376,
    n3327,
    n3324,
    n2166
  );


  nand
  g3383
  (
    n3425,
    n3397,
    n2173,
    n3235,
    n3331
  );


  xnor
  g3384
  (
    n3423,
    n3393,
    n3403,
    n3235,
    n3234
  );


  nor
  g3385
  (
    n3414,
    n3384,
    n3403,
    n3386,
    n3387
  );


  xnor
  g3386
  (
    n3430,
    n3388,
    n3332,
    n2173,
    n3401
  );


  and
  g3387
  (
    n3428,
    n3332,
    n3397,
    n2683,
    n3236
  );


  and
  g3388
  (
    n3404,
    n3233,
    n3400,
    n3386,
    n3373
  );


  nor
  g3389
  (
    KeyWire_0_6,
    n2172,
    n3400,
    n2684,
    n2174
  );


  nand
  g3390
  (
    n3426,
    n2174,
    n3380,
    n3385,
    n3234
  );


  and
  g3391
  (
    n3424,
    n2170,
    n3237,
    n3391,
    n3396
  );


  or
  g3392
  (
    n3417,
    n3394,
    n3387,
    n3236,
    n3385
  );


  nor
  g3393
  (
    n3408,
    n3394,
    n3392,
    n2691,
    n3402
  );


  nor
  g3394
  (
    n3422,
    n3382,
    n3331,
    n3383,
    n3235
  );


  nor
  g3395
  (
    n3420,
    n3391,
    n3382,
    n3403,
    n3402
  );


  and
  g3396
  (
    n3411,
    n3392,
    n3393,
    n2172,
    n3390
  );


  nor
  g3397
  (
    n3412,
    n2693,
    n3395,
    n2685,
    n2168
  );


  xor
  g3398
  (
    n3406,
    n3398,
    n3232,
    n3399,
    n3333
  );


  xnor
  g3399
  (
    n3413,
    n2686,
    n3388,
    n3383,
    n3381
  );


  xor
  g3400
  (
    n3405,
    n3394,
    n3392,
    n3402,
    n2171
  );


  nand
  g3401
  (
    n3410,
    n3396,
    n2692,
    n3232,
    n3237
  );


  nor
  g3402
  (
    n3418,
    n3397,
    n3237,
    n2168,
    n3398
  );


  or
  g3403
  (
    n3415,
    n3398,
    n3399,
    n2171,
    n3331
  );


  or
  g3404
  (
    n3427,
    n2694,
    n2690,
    n3380,
    n3400
  );


  nand
  g3405
  (
    n3432,
    n2169,
    n3332,
    n3395,
    n3333
  );


  and
  g3406
  (
    n3409,
    n2688,
    n2687,
    n3391,
    n2170
  );


  and
  g3407
  (
    n3431,
    n2689,
    n3381,
    n3384,
    n3389
  );


  xnor
  g3408
  (
    n3421,
    n3236,
    n3332,
    n3401,
    n3231
  );


  nor
  g3409
  (
    n3416,
    n3396,
    n3393,
    n2167,
    n3401
  );


  nand
  g3410
  (
    n3429,
    n3233,
    n2169,
    n3389,
    n3399
  );


  nor
  g3411
  (
    n3407,
    n3390,
    n3395,
    n3333
  );


  not
  g3412
  (
    n3450,
    n3409
  );


  buf
  g3413
  (
    n3445,
    n3423
  );


  buf
  g3414
  (
    n3446,
    n3415
  );


  not
  g3415
  (
    n3439,
    n3419
  );


  not
  g3416
  (
    n3451,
    n3422
  );


  buf
  g3417
  (
    n3441,
    n3421
  );


  buf
  g3418
  (
    n3452,
    n3417
  );


  not
  g3419
  (
    n3443,
    n3405
  );


  not
  g3420
  (
    n3436,
    n3413
  );


  not
  g3421
  (
    n3448,
    n3416
  );


  buf
  g3422
  (
    n3437,
    n3420
  );


  not
  g3423
  (
    n3434,
    n3412
  );


  not
  g3424
  (
    n3447,
    n3404
  );


  not
  g3425
  (
    n3442,
    n3418
  );


  buf
  g3426
  (
    n3440,
    n3411
  );


  not
  g3427
  (
    n3444,
    n3407
  );


  not
  g3428
  (
    n3433,
    n3408
  );


  not
  g3429
  (
    n3449,
    n3410
  );


  buf
  g3430
  (
    n3438,
    n3414
  );


  not
  g3431
  (
    n3435,
    n3406
  );


  xnor
  g3432
  (
    n3460,
    n3435,
    n3424,
    n3426,
    n3436
  );


  nor
  g3433
  (
    n3455,
    n3442,
    n3425,
    n3427
  );


  xor
  g3434
  (
    n3456,
    n3428,
    n3436,
    n3437,
    n3427
  );


  nor
  g3435
  (
    n3458,
    n3442,
    n3443,
    n3437,
    n3425
  );


  xor
  g3436
  (
    n3454,
    n3428,
    n3438,
    n3426,
    n3440
  );


  or
  g3437
  (
    n3453,
    n3439,
    n3434,
    n3440,
    n3435
  );


  or
  g3438
  (
    n3457,
    n3427,
    n3424,
    n3441,
    n3426
  );


  xnor
  g3439
  (
    n3459,
    n3439,
    n3438,
    n3441,
    n3433
  );


  buf
  g3440
  (
    n3473,
    n3456
  );


  not
  g3441
  (
    n3468,
    n3453
  );


  not
  g3442
  (
    n3461,
    n3458
  );


  not
  g3443
  (
    n3470,
    n3453
  );


  not
  g3444
  (
    n3467,
    n3458
  );


  not
  g3445
  (
    n3472,
    n3454
  );


  buf
  g3446
  (
    n3466,
    n3457
  );


  buf
  g3447
  (
    n3465,
    n3455
  );


  buf
  g3448
  (
    n3463,
    n3455
  );


  not
  g3449
  (
    n3464,
    n3457
  );


  buf
  g3450
  (
    n3471,
    n3454
  );


  buf
  g3451
  (
    n3462,
    n3456
  );


  and
  g3452
  (
    n3469,
    n3458,
    n3459,
    n3457
  );


  nor
  g3453
  (
    n3483,
    n3468,
    n3466,
    n3465,
    n3472
  );


  xnor
  g3454
  (
    n3478,
    n3470,
    n3466,
    n3463
  );


  xnor
  g3455
  (
    n3476,
    n3469,
    n3469,
    n3468,
    n3464
  );


  nor
  g3456
  (
    n3482,
    n3472,
    n3464,
    n3467
  );


  nand
  g3457
  (
    n3475,
    n3473,
    n3472,
    n3467,
    n3470
  );


  or
  g3458
  (
    n3481,
    n3461,
    n3471,
    n3465
  );


  and
  g3459
  (
    n3477,
    n3467,
    n3466,
    n3464,
    n3468
  );


  nor
  g3460
  (
    n3474,
    n3467,
    n3462,
    n3469
  );


  xor
  g3461
  (
    n3485,
    n3471,
    n3466,
    n3472,
    n3469
  );


  xor
  g3462
  (
    n3484,
    n3465,
    n3461,
    n3470
  );


  xnor
  g3463
  (
    n3480,
    n3463,
    n3461,
    n3465,
    n3462
  );


  xnor
  g3464
  (
    n3479,
    n3471,
    n3473,
    n3468
  );


  nor
  g3465
  (
    n3486,
    n3474,
    n3459
  );


  nor
  g3466
  (
    n3487,
    n3429,
    n3430,
    n3428,
    n3486
  );


  xor
  g3467
  (
    n3488,
    n3486,
    n3430,
    n3429
  );


  not
  g3468
  (
    n3489,
    n3487
  );


  buf
  g3469
  (
    n3491,
    n3460
  );


  xnor
  g3470
  (
    n3490,
    n3460,
    n3489
  );


  and
  g3471
  (
    n3492,
    n3491,
    n2175
  );


  nor
  g3472
  (
    n3493,
    n3475,
    n3492,
    n3478
  );


  or
  g3473
  (
    n3494,
    n3477,
    n3479,
    n3480,
    n3476
  );


  or
  g3474
  (
    n3499,
    n3494,
    n3493,
    n3077,
    n3075
  );


  xnor
  g3475
  (
    n3498,
    n2698,
    n3494,
    n3078,
    n3076
  );


  xor
  g3476
  (
    n3495,
    n3075,
    n3494,
    n3493
  );


  xnor
  g3477
  (
    n3496,
    n3076,
    n2699,
    n2697,
    n3493
  );


  xor
  g3478
  (
    n3497,
    n3078,
    n2695,
    n3077,
    n2696
  );


  not
  g3479
  (
    n3509,
    n3499
  );


  buf
  g3480
  (
    n3517,
    n3495
  );


  buf
  g3481
  (
    n3501,
    n3498
  );


  buf
  g3482
  (
    n3510,
    n3497
  );


  not
  g3483
  (
    n3502,
    n3497
  );


  buf
  g3484
  (
    n3516,
    n3496
  );


  not
  g3485
  (
    n3508,
    n3498
  );


  not
  g3486
  (
    n3507,
    n3499
  );


  buf
  g3487
  (
    n3513,
    n3499
  );


  not
  g3488
  (
    n3506,
    n3499
  );


  not
  g3489
  (
    n3511,
    n3496
  );


  not
  g3490
  (
    n3515,
    n3495
  );


  buf
  g3491
  (
    n3514,
    n3496
  );


  not
  g3492
  (
    n3512,
    n3498
  );


  not
  g3493
  (
    n3503,
    n3497
  );


  not
  g3494
  (
    n3505,
    n3495
  );


  not
  g3495
  (
    n3504,
    n3497
  );


  not
  g3496
  (
    n3500,
    n3498
  );


  xor
  g3497
  (
    n3532,
    n2706,
    n3506,
    n2180,
    n2708
  );


  xnor
  g3498
  (
    n3522,
    n3446,
    n2178,
    n2176,
    n3505
  );


  xor
  g3499
  (
    n3523,
    n3444,
    n3509,
    n2180,
    n2705
  );


  nand
  g3500
  (
    n3531,
    n2179,
    n3503,
    n3512,
    n2707
  );


  or
  g3501
  (
    n3524,
    n2175,
    n2183,
    n3446,
    n3451
  );


  and
  g3502
  (
    n3526,
    n3444,
    n3447,
    n3511,
    n3448
  );


  and
  g3503
  (
    n3529,
    n2700,
    n3450,
    n2177
  );


  xor
  g3504
  (
    n3521,
    n3445,
    n3445,
    n3450,
    n3502
  );


  xor
  g3505
  (
    n3527,
    n3451,
    n2179,
    n2181,
    n2183
  );


  nand
  g3506
  (
    n3518,
    n2176,
    n3447,
    n3449,
    n3508
  );


  xnor
  g3507
  (
    n3519,
    n3452,
    n3513,
    n2701,
    n2704
  );


  or
  g3508
  (
    n3520,
    n2182,
    n3510,
    n2178,
    n3443
  );


  xnor
  g3509
  (
    n3525,
    n2702,
    n3452,
    n3504,
    n3507
  );


  and
  g3510
  (
    n3528,
    n3449,
    n3448,
    n2181,
    n3514
  );


  xor
  g3511
  (
    n3530,
    n3500,
    n2703,
    n2182,
    n3501
  );


  and
  g3512
  (
    n3533,
    n3525,
    n2184
  );


  and
  g3513
  (
    n3536,
    n2714,
    n2720,
    n3533,
    n2710
  );


  or
  g3514
  (
    n3534,
    n3533,
    n2717,
    n2715,
    n2712
  );


  xor
  g3515
  (
    n3537,
    n2719,
    n2709,
    n3533
  );


  and
  g3516
  (
    n3535,
    n2716,
    n2713,
    n2718,
    n2711
  );


  xor
  g3517
  (
    n3538,
    n3481,
    n3534,
    n3536
  );


  nand
  g3518
  (
    n3540,
    n3536,
    n3535,
    n3534
  );


  nor
  g3519
  (
    n3539,
    n3494,
    n3536,
    n3537
  );


  nand
  g3520
  (
    n3542,
    n3536,
    n3535
  );


  nor
  g3521
  (
    n3541,
    n3535,
    n3534,
    n3482
  );


  buf
  g3522
  (
    n3552,
    n3542
  );


  buf
  g3523
  (
    n3545,
    n3538
  );


  not
  g3524
  (
    n3554,
    n3538
  );


  not
  g3525
  (
    n3548,
    n3538
  );


  not
  g3526
  (
    n3547,
    n3540
  );


  buf
  g3527
  (
    n3544,
    n3538
  );


  not
  g3528
  (
    n3551,
    n3539
  );


  buf
  g3529
  (
    n3550,
    n3541
  );


  buf
  g3530
  (
    n3549,
    n3541
  );


  not
  g3531
  (
    n3546,
    n3539
  );


  xnor
  g3532
  (
    n3553,
    n3373,
    n3540,
    n3541
  );


  or
  g3533
  (
    n3543,
    n3540,
    n3541,
    n3539
  );


  buf
  g3534
  (
    n3555,
    n3543
  );


  nor
  g3535
  (
    n3556,
    n3528,
    n3530,
    n3526,
    n3555
  );


  nand
  g3536
  (
    n3557,
    n3483,
    n3527,
    n3555,
    n3529
  );


  not
  g3537
  (
    n3558,
    n3430
  );


  buf
  g3538
  (
    n3559,
    n3431
  );


  buf
  g3539
  (
    n3563,
    n3431
  );


  buf
  g3540
  (
    n3560,
    n3556
  );


  xor
  g3541
  (
    n3562,
    n3556,
    n3557
  );


  xor
  g3542
  (
    n3561,
    n3431,
    n3556,
    n3557
  );


  buf
  g3543
  (
    n3578,
    n2186
  );


  not
  g3544
  (
    n3585,
    n3558
  );


  not
  g3545
  (
    n3587,
    n3560
  );


  buf
  g3546
  (
    n3566,
    n3562
  );


  not
  g3547
  (
    n3579,
    n2188
  );


  buf
  g3548
  (
    n3564,
    n3558
  );


  buf
  g3549
  (
    n3581,
    n3559
  );


  buf
  g3550
  (
    n3580,
    n3558
  );


  buf
  g3551
  (
    n3569,
    n3563
  );


  buf
  g3552
  (
    n3584,
    n2187
  );


  buf
  g3553
  (
    n3567,
    n2186
  );


  buf
  g3554
  (
    n3572,
    n3558
  );


  not
  g3555
  (
    n3573,
    n3559
  );


  not
  g3556
  (
    n3575,
    n3561
  );


  buf
  g3557
  (
    n3568,
    n3561
  );


  not
  g3558
  (
    n3565,
    n3563
  );


  not
  g3559
  (
    n3583,
    n3563
  );


  buf
  g3560
  (
    n3574,
    n3561
  );


  xor
  g3561
  (
    n3582,
    n2188,
    n2187,
    n3560
  );


  nand
  g3562
  (
    n3570,
    n3559,
    n2184,
    n3562
  );


  nor
  g3563
  (
    n3577,
    n3563,
    n3560,
    n2185
  );


  xnor
  g3564
  (
    n3586,
    n3562,
    n2189,
    n2185
  );


  xnor
  g3565
  (
    n3576,
    n3561,
    n2190,
    n3562
  );


  and
  g3566
  (
    n3571,
    n3559,
    n2189,
    n3560
  );


  nor
  g3567
  (
    n3604,
    n2819,
    n2740,
    n3586,
    n2837
  );


  nand
  g3568
  (
    n3616,
    n2751,
    n2739,
    n2791,
    n2831
  );


  and
  g3569
  (
    n3618,
    n2746,
    n2796,
    n2725,
    n3579
  );


  nor
  g3570
  (
    n3607,
    n2764,
    n2836,
    n3571,
    n3585
  );


  nand
  g3571
  (
    n3617,
    n2741,
    n3584,
    n3570,
    n2732
  );


  nand
  g3572
  (
    n3602,
    n3581,
    n2813,
    n2808,
    n2765
  );


  or
  g3573
  (
    n3627,
    n3582,
    n2723,
    n3574,
    n3584
  );


  xnor
  g3574
  (
    n3588,
    n2767,
    n2822,
    n2770,
    n2777
  );


  nor
  g3575
  (
    n3595,
    n2797,
    n2781,
    n2763,
    n2736
  );


  xor
  g3576
  (
    n3593,
    n2840,
    n2820,
    n2832,
    n2795
  );


  nor
  g3577
  (
    n3596,
    n2726,
    n3564,
    n2766,
    n2757
  );


  and
  g3578
  (
    n3626,
    n2729,
    n2780,
    n2722,
    n2809
  );


  or
  g3579
  (
    n3589,
    n3568,
    n2825,
    n2754,
    n2727
  );


  and
  g3580
  (
    n3605,
    n3566,
    n2738,
    n2835,
    n2749
  );


  nand
  g3581
  (
    n3615,
    n2792,
    n2818,
    n2787,
    n3565
  );


  nand
  g3582
  (
    n3601,
    n2755,
    n2779,
    n2744,
    n2734
  );


  or
  g3583
  (
    n3612,
    n2805,
    n3587,
    n2758,
    n2826
  );


  nor
  g3584
  (
    n3592,
    n3567,
    n2752,
    n2829,
    n3573
  );


  nor
  g3585
  (
    n3606,
    n3576,
    n2802,
    n2743,
    n2784
  );


  or
  g3586
  (
    n3624,
    n2753,
    n2724,
    n2748,
    n3575
  );


  or
  g3587
  (
    n3619,
    n2775,
    n2810,
    n3575,
    n3572
  );


  nor
  g3588
  (
    n3620,
    n2745,
    n2814,
    n2839,
    n2761
  );


  or
  g3589
  (
    n3603,
    n2789,
    n2737,
    n3587,
    n3577
  );


  and
  g3590
  (
    n3597,
    n2772,
    n2811,
    n3586,
    n2823
  );


  xor
  g3591
  (
    n3594,
    n2742,
    n2833,
    n2799,
    n3574
  );


  xor
  g3592
  (
    n3625,
    n2774,
    n2834,
    n2801,
    n2800
  );


  xor
  g3593
  (
    n3599,
    n3583,
    n2815,
    n3576,
    n2762
  );


  xnor
  g3594
  (
    n3623,
    n2771,
    n2735,
    n2794,
    n2782
  );


  xor
  g3595
  (
    n3609,
    n3578,
    n2816,
    n2778,
    n2803
  );


  xor
  g3596
  (
    n3614,
    n2760,
    n2730,
    n2747,
    n3581
  );


  nand
  g3597
  (
    n3598,
    n2793,
    n2721,
    n2786,
    n3582
  );


  or
  g3598
  (
    n3611,
    n2731,
    n2788,
    n2812,
    n3577
  );


  and
  g3599
  (
    n3610,
    n3569,
    n2838,
    n2759,
    n2821
  );


  nand
  g3600
  (
    n3621,
    n2806,
    n3580,
    n2828,
    n2790
  );


  nand
  g3601
  (
    n3600,
    n2750,
    n3579,
    n3573,
    n2733
  );


  xnor
  g3602
  (
    n3608,
    n2728,
    n2785,
    n2830,
    n3578
  );


  nand
  g3603
  (
    n3591,
    n2776,
    n3583,
    n2807,
    n2773
  );


  nand
  g3604
  (
    n3622,
    n2827,
    n2824,
    n2783,
    n3580
  );


  nand
  g3605
  (
    n3590,
    n2798,
    n2804,
    n2768,
    n2769
  );


  xor
  g3606
  (
    n3613,
    n2817,
    n3572,
    n3585,
    n2756
  );


  buf
  g3607
  (
    n3628,
    n3608
  );


  buf
  g3608
  (
    n3637,
    n3612
  );


  not
  g3609
  (
    n3632,
    n3594
  );


  buf
  g3610
  (
    n3635,
    n3543
  );


  buf
  g3611
  (
    n3644,
    n3598
  );


  buf
  g3612
  (
    n3651,
    n3544
  );


  buf
  g3613
  (
    n3648,
    n3547
  );


  not
  g3614
  (
    n3650,
    n3596
  );


  buf
  g3615
  (
    n3638,
    n3613
  );


  not
  g3616
  (
    n3639,
    n3547
  );


  buf
  g3617
  (
    n3630,
    n3619
  );


  not
  g3618
  (
    n3631,
    n3617
  );


  not
  g3619
  (
    n3629,
    n3610
  );


  not
  g3620
  (
    n3640,
    n3588
  );


  buf
  g3621
  (
    n3652,
    n3545
  );


  buf
  g3622
  (
    n3647,
    n3546
  );


  not
  g3623
  (
    n3649,
    n3620
  );


  xor
  g3624
  (
    n3636,
    n3599,
    n3604,
    n3606
  );


  nor
  g3625
  (
    n3641,
    n3609,
    n3544,
    n3545,
    n3589
  );


  xor
  g3626
  (
    n3646,
    n3602,
    n3545,
    n3616,
    n3590
  );


  nand
  g3627
  (
    n3643,
    n3548,
    n3618,
    n3545,
    n3593
  );


  nand
  g3628
  (
    n3645,
    n3615,
    n3601,
    n3614,
    n3595
  );


  and
  g3629
  (
    n3633,
    n3544,
    n3546,
    n3473,
    n3592
  );


  and
  g3630
  (
    KeyWire_0_12,
    n3597,
    n3600,
    n3547,
    n3543
  );


  xnor
  g3631
  (
    n3653,
    n3605,
    n3547,
    n3611,
    n3591
  );


  or
  g3632
  (
    n3634,
    n3607,
    n3546,
    n3603
  );


  nand
  g3633
  (
    n3670,
    n3648,
    n3650,
    n2265,
    n2193
  );


  xor
  g3634
  (
    n3709,
    n3628,
    n2261,
    n3517,
    n2197
  );


  xnor
  g3635
  (
    n3664,
    n3516,
    n3643,
    n3636,
    n2239
  );


  or
  g3636
  (
    n3716,
    n3029,
    n3635,
    n3025,
    n2195
  );


  or
  g3637
  (
    n3702,
    n2234,
    n2254,
    n2265,
    n2228
  );


  nor
  g3638
  (
    n3673,
    n2251,
    n3651,
    n2198,
    n2203
  );


  and
  g3639
  (
    n3704,
    n3645,
    n2195,
    n3024,
    n2269
  );


  xor
  g3640
  (
    n3694,
    n3646,
    n2248,
    n2209,
    n3633
  );


  or
  g3641
  (
    n3660,
    n3639,
    n2214,
    n2194,
    n2285
  );


  or
  g3642
  (
    n3725,
    n3020,
    n2232,
    n2260,
    n2273
  );


  nand
  g3643
  (
    n3683,
    n2242,
    n2221,
    n2241,
    n2276
  );


  or
  g3644
  (
    n3731,
    n3645,
    n2201,
    n2202,
    n2280
  );


  xor
  g3645
  (
    n3690,
    n2267,
    n2208,
    n3644,
    n3027
  );


  or
  g3646
  (
    n3700,
    n2194,
    n3632,
    n3025,
    n2275
  );


  nor
  g3647
  (
    n3714,
    n2274,
    n3641,
    n2234,
    n3651
  );


  xor
  g3648
  (
    n3723,
    n3646,
    n2266,
    n2249,
    n2278
  );


  or
  g3649
  (
    n3662,
    n3641,
    n3018,
    n2212,
    n2281
  );


  nor
  g3650
  (
    n3661,
    n2280,
    n2216,
    n3632,
    n2266
  );


  nand
  g3651
  (
    n3686,
    n2284,
    n2210,
    n2245,
    n2228
  );


  xor
  g3652
  (
    n3678,
    n2255,
    n2220,
    n2268,
    n3640
  );


  nand
  g3653
  (
    n3718,
    n2282,
    n2218,
    n3028,
    n2235
  );


  and
  g3654
  (
    n3699,
    n2286,
    n3023,
    n3653,
    n3640
  );


  and
  g3655
  (
    n3677,
    n2209,
    n3029,
    n3025,
    n2264
  );


  nand
  g3656
  (
    n3698,
    n2247,
    n2193,
    n3648,
    n2241
  );


  nand
  g3657
  (
    n3703,
    n2238,
    n3637,
    n2213,
    n3631
  );


  xor
  g3658
  (
    n3720,
    n2242,
    n3020,
    n2284,
    n2196
  );


  xor
  g3659
  (
    n3696,
    n2197,
    n3648,
    n2244,
    n3653
  );


  and
  g3660
  (
    n3655,
    n2264,
    n3644,
    n2202,
    n3026
  );


  xnor
  g3661
  (
    n3707,
    n2259,
    n3637,
    n2196,
    n3026
  );


  nor
  g3662
  (
    n3671,
    n2252,
    n3022,
    n2285,
    n2247
  );


  or
  g3663
  (
    n3715,
    n2276,
    n2282,
    n2199,
    n3651
  );


  and
  g3664
  (
    n3654,
    n3632,
    n3636,
    n2210,
    n2288
  );


  nand
  g3665
  (
    n3669,
    n2190,
    n3019,
    n3642,
    n2235
  );


  and
  g3666
  (
    n3675,
    n3642,
    n3652,
    n2201,
    n2277
  );


  nor
  g3667
  (
    n3668,
    n2231,
    n3638,
    n2207,
    n3019
  );


  nor
  g3668
  (
    n3712,
    n2211,
    n2279,
    n3631,
    n2260
  );


  xor
  g3669
  (
    n3688,
    n2258,
    n3635,
    n2254,
    n3647
  );


  xnor
  g3670
  (
    n3730,
    n2275,
    n3646,
    n2243,
    n2257
  );


  and
  g3671
  (
    n3711,
    n2283,
    n2274,
    n3024,
    n2219
  );


  xor
  g3672
  (
    n3676,
    n3645,
    n2238,
    n3028,
    n2248
  );


  xor
  g3673
  (
    n3685,
    n3628,
    n3647,
    n2271,
    n3640
  );


  nor
  g3674
  (
    n3692,
    n2218,
    n3021,
    n2270,
    n3027
  );


  and
  g3675
  (
    n3689,
    n2225,
    n2231,
    n3649,
    n2219
  );


  nor
  g3676
  (
    n3656,
    n3643,
    n2226,
    n2191,
    n2278
  );


  or
  g3677
  (
    n3687,
    n3515,
    n2259,
    n2262,
    n2213
  );


  or
  g3678
  (
    n3722,
    n3634,
    n2257,
    n2222,
    n2233
  );


  nand
  g3679
  (
    n3726,
    n2223,
    n2288,
    n2289,
    n2239
  );


  xnor
  g3680
  (
    n3705,
    n2216,
    n2240,
    n2253,
    n2236
  );


  or
  g3681
  (
    n3719,
    n2249,
    n2222,
    n2229,
    n2272
  );


  nor
  g3682
  (
    KeyWire_0_7,
    n2232,
    n3629,
    n3650,
    n3028
  );


  xor
  g3683
  (
    n3710,
    n3633,
    n2236,
    n2224
  );


  xnor
  g3684
  (
    n3706,
    n2199,
    n3024,
    n3021,
    n2253
  );


  nand
  g3685
  (
    n3721,
    n3652,
    n2283,
    n2255,
    n3638
  );


  xnor
  g3686
  (
    n3658,
    n2277,
    n2198,
    n2227,
    n2225
  );


  nand
  g3687
  (
    n3695,
    n2237,
    n3635,
    n2203,
    n2246
  );


  and
  g3688
  (
    n3663,
    n3633,
    n3653,
    n2269,
    n2206
  );


  nor
  g3689
  (
    n3713,
    n2217,
    n3649,
    n2205,
    n2287
  );


  or
  g3690
  (
    n3680,
    n2230,
    n2272,
    n3023,
    n2200
  );


  xnor
  g3691
  (
    n3679,
    n2212,
    n3647,
    n2223,
    n2204
  );


  xnor
  g3692
  (
    n3728,
    n3650,
    n2229,
    n2227,
    n2273
  );


  or
  g3693
  (
    n3666,
    n2268,
    n2192,
    n2258,
    n2246
  );


  or
  g3694
  (
    n3684,
    n2261,
    n2281,
    n2243,
    n2206
  );


  nor
  g3695
  (
    n3727,
    n3021,
    n3629,
    n2267,
    n2207
  );


  xnor
  g3696
  (
    n3657,
    n3022,
    n2270,
    n2244,
    n2204
  );


  nor
  g3697
  (
    n3708,
    n3642,
    n2220,
    n2233,
    n3019
  );


  or
  g3698
  (
    n3717,
    n2250,
    n2262,
    n2252,
    n3638
  );


  or
  g3699
  (
    n3665,
    n2192,
    n2286,
    n3652,
    n3020
  );


  nor
  g3700
  (
    n3701,
    n2237,
    n3630,
    n2221,
    n3022
  );


  and
  g3701
  (
    n3659,
    n2256,
    n3641,
    n2208,
    n2251
  );


  or
  g3702
  (
    n3672,
    n3649,
    n3644,
    n3637,
    n2287
  );


  and
  g3703
  (
    n3681,
    n2245,
    n2214,
    n3634,
    n3639
  );


  xor
  g3704
  (
    n3682,
    n3639,
    n3026,
    n2215,
    n3636
  );


  xor
  g3705
  (
    n3667,
    n2271,
    n2230,
    n2205,
    n3628
  );


  nand
  g3706
  (
    n3674,
    n2191,
    n3631,
    n2250,
    n2256
  );


  xor
  g3707
  (
    n3691,
    n2211,
    n3023,
    n2200,
    n2217
  );


  xnor
  g3708
  (
    n3729,
    n3643,
    n3630,
    n2226,
    n2263
  );


  xor
  g3709
  (
    n3697,
    n3630,
    n2279,
    n2263,
    n3634
  );


  or
  g3710
  (
    n3693,
    n2240,
    n3027,
    n3629,
    n2215
  );


  nand
  g3711
  (
    n3747,
    n3685,
    n3713,
    n3662,
    n3704
  );


  xor
  g3712
  (
    n3769,
    n3690,
    n3659,
    n3699,
    n3664
  );


  xnor
  g3713
  (
    n3754,
    n3272,
    n3673,
    n3694,
    n3680
  );


  xnor
  g3714
  (
    n3778,
    n3699,
    n3665,
    n3666,
    n3724
  );


  and
  g3715
  (
    n3765,
    n3668,
    n3726,
    n3727,
    n3684
  );


  xnor
  g3716
  (
    n3773,
    n3726,
    n3692,
    n3711,
    n3716
  );


  nand
  g3717
  (
    n3762,
    n3708,
    n3714,
    n3719,
    n3725
  );


  xor
  g3718
  (
    n3772,
    n3711,
    n3683,
    n3707,
    n3671
  );


  or
  g3719
  (
    n3764,
    n3720,
    n3697,
    n3668,
    n3712
  );


  nand
  g3720
  (
    n3766,
    n3706,
    n3271,
    n3677,
    n3654
  );


  nand
  g3721
  (
    n3732,
    n3667,
    n3485,
    n3703,
    n3706
  );


  nor
  g3722
  (
    n3760,
    n3688,
    n3657,
    n3703,
    n3693
  );


  nor
  g3723
  (
    n3733,
    n3675,
    n3713,
    n3705,
    n3306
  );


  xnor
  g3724
  (
    n3750,
    n3683,
    n3666,
    n3660,
    n3657
  );


  nand
  g3725
  (
    n3748,
    n3678,
    n3663,
    n3701,
    n3707
  );


  nand
  g3726
  (
    n3735,
    n3671,
    n3711,
    n3726,
    n3665
  );


  or
  g3727
  (
    n3774,
    n3697,
    n3723,
    n3670,
    n3719
  );


  and
  g3728
  (
    n3761,
    n3669,
    n3694,
    n3484,
    n3307
  );


  or
  g3729
  (
    n3751,
    n3699,
    n3681,
    n3718,
    n3692
  );


  nand
  g3730
  (
    n3755,
    n3684,
    n3701,
    n3717,
    n3708
  );


  or
  g3731
  (
    n3744,
    n3719,
    n3667,
    n3678,
    n3704
  );


  xnor
  g3732
  (
    n3746,
    n3680,
    n3685,
    n3696,
    n3660
  );


  xor
  g3733
  (
    n3758,
    n3705,
    n3674,
    n3710,
    n3688
  );


  nand
  g3734
  (
    n3739,
    n3654,
    n3706,
    n3700,
    n3687
  );


  and
  g3735
  (
    n3768,
    n3712,
    n3723,
    n3691,
    n3682
  );


  nand
  g3736
  (
    n3771,
    n3691,
    n3689,
    n3696,
    n3305
  );


  nor
  g3737
  (
    n3742,
    n3693,
    n3661,
    n3725,
    n3702
  );


  xor
  g3738
  (
    n3776,
    n3722,
    n3662,
    n3713,
    n3709
  );


  nor
  g3739
  (
    n3763,
    n3700,
    n3718,
    n3698,
    n3306
  );


  xnor
  g3740
  (
    n3777,
    n3681,
    n3695,
    n3673,
    n3704
  );


  xnor
  g3741
  (
    n3757,
    n3705,
    n3672,
    n3717,
    n3701
  );


  nor
  g3742
  (
    n3779,
    n3722,
    n3715,
    n3687,
    n3682
  );


  nor
  g3743
  (
    n3738,
    n3695,
    n3716,
    n3672,
    n3720
  );


  nand
  g3744
  (
    n3743,
    n3664,
    n3720,
    n3724,
    n3679
  );


  nor
  g3745
  (
    n3734,
    n3709,
    n3702,
    n3724,
    n3655
  );


  xnor
  g3746
  (
    n3749,
    n3686,
    n3679,
    n3710,
    n3721
  );


  nor
  g3747
  (
    n3740,
    n3710,
    n3656,
    n3655,
    n3272
  );


  or
  g3748
  (
    n3753,
    n3714,
    n3661,
    n3717,
    n3656
  );


  xor
  g3749
  (
    n3745,
    n3709,
    n3663,
    n3658,
    n3712
  );


  nand
  g3750
  (
    n3770,
    n3677,
    n3307,
    n3670,
    n3689
  );


  or
  g3751
  (
    n3752,
    n3675,
    n3727,
    n3723,
    n3700
  );


  xor
  g3752
  (
    n3736,
    n3659,
    n3721,
    n3702,
    n3676
  );


  xnor
  g3753
  (
    n3759,
    n3271,
    n3715,
    n3669,
    n3718
  );


  nand
  g3754
  (
    n3767,
    n3716,
    n3722,
    n3707,
    n3714
  );


  nand
  g3755
  (
    n3737,
    n3721,
    n3698,
    n3697
  );


  and
  g3756
  (
    n3741,
    n3658,
    n3727,
    n3686,
    n3703
  );


  nor
  g3757
  (
    n3756,
    n3676,
    n3696,
    n3690,
    n3306
  );


  nor
  g3758
  (
    n3775,
    n3725,
    n3715,
    n3708,
    n3674
  );


  nor
  g3759
  (
    n3800,
    n3777,
    n3742,
    n3757,
    n3779
  );


  nor
  g3760
  (
    n3802,
    n3737,
    n2846,
    n3745
  );


  nor
  g3761
  (
    n3793,
    n3768,
    n3750,
    n2885,
    n3755
  );


  or
  g3762
  (
    n3842,
    n3749,
    n3747,
    n3748,
    n3757
  );


  nor
  g3763
  (
    n3792,
    n3741,
    n3753,
    n3487,
    n3769
  );


  or
  g3764
  (
    n3807,
    n3740,
    n3766,
    n3769
  );


  xnor
  g3765
  (
    n3844,
    n3747,
    n3767,
    n3766,
    n2883
  );


  nor
  g3766
  (
    n3789,
    n3755,
    n3748,
    n3749,
    n3746
  );


  nor
  g3767
  (
    n3796,
    n3752,
    n3756,
    n2886,
    n3746
  );


  xnor
  g3768
  (
    n3811,
    n3771,
    n2851,
    n2886,
    n3762
  );


  xnor
  g3769
  (
    n3825,
    n3746,
    n3762,
    n3730,
    n3778
  );


  or
  g3770
  (
    n3829,
    n3734,
    n3738,
    n3743,
    n3744
  );


  nor
  g3771
  (
    n3839,
    n2871,
    n3778,
    n3758
  );


  xnor
  g3772
  (
    n3804,
    n3774,
    n3734,
    n2861,
    n3750
  );


  nor
  g3773
  (
    n3785,
    n3775,
    n2875,
    n3773,
    n3771
  );


  xnor
  g3774
  (
    n3814,
    n3764,
    n2884,
    n3754,
    n3729
  );


  nor
  g3775
  (
    n3820,
    n3744,
    n2884,
    n2859,
    n3779
  );


  xnor
  g3776
  (
    n3803,
    n3776,
    n3771,
    n3770,
    n3736
  );


  xor
  g3777
  (
    n3809,
    n3752,
    n2865,
    n3768,
    n2856
  );


  xnor
  g3778
  (
    n3838,
    n3729,
    n3761,
    n3730,
    n3757
  );


  xnor
  g3779
  (
    n3805,
    n2847,
    n3745,
    n3755,
    n3769
  );


  xor
  g3780
  (
    n3837,
    n3777,
    n3770,
    n3733,
    n2885
  );


  and
  g3781
  (
    n3783,
    n2850,
    n3747,
    n3754,
    n2842
  );


  nand
  g3782
  (
    n3795,
    n2862,
    n3733,
    n2885,
    n2874
  );


  or
  g3783
  (
    n3791,
    n3739,
    n3728,
    n3748,
    n3734
  );


  xnor
  g3784
  (
    n3801,
    n3775,
    n3771,
    n3763,
    n2872
  );


  nor
  g3785
  (
    n3845,
    n3765,
    n2887,
    n3740,
    n3728
  );


  xor
  g3786
  (
    n3834,
    n3757,
    n2887,
    n3737,
    n3753
  );


  nand
  g3787
  (
    n3787,
    n3746,
    n2870,
    n2884,
    n3741
  );


  nand
  g3788
  (
    n3790,
    n3764,
    n3737,
    n2869,
    n3779
  );


  and
  g3789
  (
    n3810,
    n3779,
    n2864,
    n3755,
    n3743
  );


  xnor
  g3790
  (
    n3831,
    n3736,
    n3761,
    n3759,
    n3764
  );


  xor
  g3791
  (
    n3786,
    n3732,
    n2878,
    n3740,
    n3741
  );


  xnor
  g3792
  (
    n3830,
    n3488,
    n3749,
    n3770,
    n2854
  );


  nor
  g3793
  (
    n3822,
    n2852,
    n3776,
    n2867,
    n2863
  );


  nand
  g3794
  (
    n3781,
    n2873,
    n2857,
    n3772,
    n3738
  );


  nor
  g3795
  (
    n3841,
    n3759,
    n3750,
    n3735,
    n3770
  );


  nor
  g3796
  (
    KeyWire_0_5,
    n3730,
    n3763,
    n3775,
    n2844
  );


  and
  g3797
  (
    n3798,
    n3753,
    n2849,
    n2858,
    n3769
  );


  or
  g3798
  (
    n3846,
    n3731,
    n3756,
    n2845,
    n3754
  );


  nor
  g3799
  (
    n3833,
    n3741,
    n3742,
    n3739,
    n3765
  );


  xnor
  g3800
  (
    n3843,
    n3488,
    n3777,
    n3773,
    n3762
  );


  xor
  g3801
  (
    n3836,
    n3737,
    n2848,
    n2853,
    n3733
  );


  xnor
  g3802
  (
    n3797,
    n3773,
    n3735,
    n3751,
    n2881
  );


  xor
  g3803
  (
    n3823,
    n3743,
    n3738,
    n3753,
    n3765
  );


  xnor
  g3804
  (
    n3821,
    n3756,
    n2879,
    n2887,
    n2876
  );


  and
  g3805
  (
    n3827,
    n3743,
    n3739,
    n3756,
    n3776
  );


  or
  g3806
  (
    n3780,
    n3774,
    n3774,
    n3736,
    n3754
  );


  xnor
  g3807
  (
    n3794,
    n3760,
    n2880,
    n2855,
    n3762
  );


  or
  g3808
  (
    n3835,
    n3763,
    n3735,
    n2883,
    n3747
  );


  xor
  g3809
  (
    n3813,
    n3749,
    n2883,
    n3738,
    n3773
  );


  or
  g3810
  (
    n3819,
    n2843,
    n3766,
    n3772,
    n3778
  );


  or
  g3811
  (
    n3826,
    n3760,
    n3763,
    n2888
  );


  xor
  g3812
  (
    n3817,
    n2868,
    n2886,
    n3758,
    n3728
  );


  and
  g3813
  (
    n3824,
    n3732,
    n3768,
    n3750
  );


  xnor
  g3814
  (
    n3832,
    n3767,
    n3772,
    n3740,
    n3758
  );


  xor
  g3815
  (
    n3840,
    n3739,
    n3777,
    n3732,
    n3751
  );


  xnor
  g3816
  (
    n3784,
    n3764,
    n3775,
    n3729,
    n3734
  );


  xor
  g3817
  (
    n3788,
    n3760,
    n3488,
    n3752,
    n2888
  );


  xnor
  g3818
  (
    n3806,
    n3733,
    n3774,
    n3761,
    n3759
  );


  xor
  g3819
  (
    n3815,
    n3776,
    n3732,
    n2860,
    n3760
  );


  nand
  g3820
  (
    n3782,
    n3731,
    n2877,
    n3759,
    n3772
  );


  or
  g3821
  (
    n3816,
    n3752,
    n3745,
    n3742,
    n3735
  );


  xor
  g3822
  (
    n3808,
    n3731,
    n3765,
    n3748,
    n3767
  );


  and
  g3823
  (
    n3799,
    n3751,
    n3744,
    n3767,
    n2882
  );


  or
  g3824
  (
    n3828,
    n3761,
    n3742,
    n2841,
    n2866
  );


  or
  g3825
  (
    n3812,
    n3751,
    n3758,
    n3736,
    n3744
  );


  xor
  g3826
  (
    n3854,
    n3803,
    n3816,
    n3821,
    n3802
  );


  nor
  g3827
  (
    n3853,
    n3787,
    n3805,
    n3793,
    n3801
  );


  xor
  g3828
  (
    n3849,
    n3792,
    n3807,
    n3796,
    n3820
  );


  nand
  g3829
  (
    n3858,
    n3809,
    n3788,
    n3817,
    n3791
  );


  xor
  g3830
  (
    n3856,
    n3537,
    n3804,
    n3813,
    n3818
  );


  nand
  g3831
  (
    n3847,
    n3789,
    n3795,
    n3810,
    n3782
  );


  nand
  g3832
  (
    n3857,
    n19,
    n3785,
    n3819,
    n3537
  );


  xnor
  g3833
  (
    n3851,
    n3786,
    n3783,
    n3799,
    n3780
  );


  or
  g3834
  (
    n3855,
    n3797,
    n3814,
    n3781,
    n3798
  );


  and
  g3835
  (
    n3852,
    n3808,
    n3811,
    n3784,
    n3790
  );


  nand
  g3836
  (
    n3848,
    n3806,
    n20,
    n3537
  );


  nand
  g3837
  (
    n3850,
    n3800,
    n3794,
    n3812,
    n3815
  );


  buf
  g3838
  (
    n3865,
    n3856
  );


  not
  g3839
  (
    n3869,
    n20
  );


  not
  g3840
  (
    n3859,
    n3858
  );


  not
  g3841
  (
    n3861,
    n3626
  );


  not
  g3842
  (
    n3864,
    n3857
  );


  buf
  g3843
  (
    n3872,
    n3272
  );


  not
  g3844
  (
    n3862,
    n3542
  );


  not
  g3845
  (
    n3867,
    n3853
  );


  buf
  g3846
  (
    n3874,
    n3854
  );


  not
  g3847
  (
    n3866,
    n3855
  );


  xnor
  g3848
  (
    n3873,
    n3849,
    n3851,
    n3856
  );


  nand
  g3849
  (
    n3868,
    n3625,
    n3542,
    n3850
  );


  nand
  g3850
  (
    n3860,
    n3626,
    n3627,
    n3542,
    n3852
  );


  nand
  g3851
  (
    n3870,
    n3621,
    n3847,
    n3855,
    n3625
  );


  xnor
  g3852
  (
    n3871,
    n3623,
    n3858,
    n3622,
    n3624
  );


  xor
  g3853
  (
    n3863,
    n3857,
    n3627,
    n3848,
    n3822
  );


  xnor
  g3854
  (
    n3890,
    n20,
    n3866,
    n3551,
    n3308
  );


  xor
  g3855
  (
    n3877,
    n3872,
    n3865,
    n2291,
    n3552
  );


  nand
  g3856
  (
    n3894,
    n3549,
    n2292,
    n3871,
    n3550
  );


  xor
  g3857
  (
    n3893,
    n3871,
    n2290,
    n3551,
    n3872
  );


  nand
  g3858
  (
    n3887,
    n3873,
    n3554,
    n3307,
    n3868
  );


  xnor
  g3859
  (
    n3879,
    n3550,
    n2301,
    n3548,
    n3861
  );


  xnor
  g3860
  (
    n3880,
    n2298,
    n2301,
    n2293,
    n3870
  );


  nor
  g3861
  (
    n3882,
    n3309,
    n2299,
    n3554,
    n3551
  );


  or
  g3862
  (
    n3878,
    n3552,
    n2300,
    n3549,
    n2299
  );


  nand
  g3863
  (
    n3886,
    n2302,
    n2289,
    n3873,
    n3548
  );


  nand
  g3864
  (
    n3891,
    n2294,
    n3310,
    n3864,
    n2291
  );


  nand
  g3865
  (
    n3881,
    n3860,
    n2298,
    n2302,
    n3859
  );


  nor
  g3866
  (
    n3885,
    n3551,
    n2296,
    n3549,
    n3552
  );


  nor
  g3867
  (
    n3892,
    n3552,
    n3308,
    n2297,
    n3870
  );


  xor
  g3868
  (
    n3888,
    n3553,
    n3869,
    n3554,
    n3550
  );


  xnor
  g3869
  (
    n3876,
    n2294,
    n3874,
    n3310,
    n3554
  );


  xnor
  g3870
  (
    n3884,
    n3308,
    n3553,
    n3432,
    n3309
  );


  and
  g3871
  (
    n3883,
    n2293,
    n2300,
    n3432,
    n3553
  );


  xnor
  g3872
  (
    n3895,
    n2292,
    n3553,
    n3867,
    n3863
  );


  xor
  g3873
  (
    n3889,
    n3548,
    n2290,
    n3874,
    n3862
  );


  xnor
  g3874
  (
    n3875,
    n3309,
    n2295,
    n3549
  );


  nor
  g3875
  (
    n3896,
    n2296,
    n3869,
    n3550,
    n2297
  );


  buf
  g3876
  (
    n3897,
    n3875
  );


  xor
  g3877
  (
    n3898,
    n3897,
    n2889,
    n2890
  );


  nand
  g3878
  (
    n3899,
    n2889,
    n2890,
    n3897
  );


  xor
  g3879
  (
    n3904,
    n3826,
    n3830,
    n3898,
    n3840
  );


  xor
  g3880
  (
    n3903,
    n3841,
    n3824,
    n3899,
    n3829
  );


  nand
  g3881
  (
    n3906,
    n3837,
    n3898,
    n3899
  );


  xnor
  g3882
  (
    n3900,
    n3833,
    n3898,
    n3842,
    n3827
  );


  nand
  g3883
  (
    n3901,
    n3828,
    n3843,
    n3839,
    n3846
  );


  nor
  g3884
  (
    n3907,
    n3899,
    n3845,
    n3838,
    n3836
  );


  or
  g3885
  (
    n3905,
    n3831,
    n3899,
    n3834,
    n3832
  );


  nand
  g3886
  (
    n3902,
    n3825,
    n3844,
    n3823,
    n3835
  );


  xor
  g3887
  (
    n3918,
    n3902,
    n3889,
    n3906,
    n3904
  );


  xor
  g3888
  (
    n3909,
    n3888,
    n3906,
    n3905,
    n3030
  );


  xor
  g3889
  (
    n3913,
    n3903,
    n3878,
    n3432,
    n3907
  );


  xnor
  g3890
  (
    n3917,
    n3905,
    n3891,
    n3895,
    n3904
  );


  xnor
  g3891
  (
    n3911,
    n3894,
    n318,
    n3896,
    n3884
  );


  nand
  g3892
  (
    n3914,
    n3890,
    n318,
    n3877,
    n3896
  );


  nand
  g3893
  (
    n3912,
    n3882,
    n3907,
    n3887
  );


  nand
  g3894
  (
    n3908,
    n3892,
    n3893,
    n3885,
    n3880
  );


  xnor
  g3895
  (
    n3919,
    n3895,
    n3900,
    n108,
    n3906
  );


  nand
  g3896
  (
    n3920,
    n3886,
    n108,
    n3881,
    n3883
  );


  xnor
  g3897
  (
    n3910,
    n3532,
    n3030,
    n3901,
    n3894
  );


  and
  g3898
  (
    n3916,
    n3879,
    n3029,
    n318,
    n3876
  );


  nor
  g3899
  (
    n3915,
    n3030,
    n3904,
    n3531,
    n3905
  );


  xor
  g3900
  (
    n3924,
    n3913,
    n3909,
    n3920,
    n3912
  );


  and
  g3901
  (
    n3922,
    n3919,
    n3908,
    n3917,
    n108
  );


  or
  g3902
  (
    n3923,
    n108,
    n3914,
    n3915,
    n3918
  );


  nor
  g3903
  (
    n3921,
    n3310,
    n3916,
    n3911,
    n3910
  );


  xnor
  KeyGate_0_0
  (
    n1423,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n80,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n312,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1211,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1701,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n3818,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n3419,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n3724,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n2199,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n870,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n21,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n2790,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n3642,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1814,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n2058,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n57,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1672,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1160,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n679,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n327,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n387,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n786,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n2350,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n116,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n2474,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1221,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n285,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n3333,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n253,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n2257,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n2686,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n2958,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

