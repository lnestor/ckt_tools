

module Stat_1436_31_3
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n1241,
  n1303,
  n1310,
  n1313,
  n1305,
  n1306,
  n1309,
  n1311,
  n1301,
  n1367,
  n1357,
  n1355,
  n1363,
  n1353,
  n1358,
  n1366,
  n1370,
  n1368,
  n1359,
  n1462,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n1241;
  output n1303;
  output n1310;
  output n1313;
  output n1305;
  output n1306;
  output n1309;
  output n1311;
  output n1301;
  output n1367;
  output n1357;
  output n1355;
  output n1363;
  output n1353;
  output n1358;
  output n1366;
  output n1370;
  output n1368;
  output n1359;
  output n1462;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1302;
  wire n1304;
  wire n1307;
  wire n1308;
  wire n1312;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1354;
  wire n1356;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1364;
  wire n1365;
  wire n1369;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n96,
    n4
  );


  buf
  g1
  (
    n35,
    n26
  );


  not
  g2
  (
    n126,
    n2
  );


  not
  g3
  (
    n38,
    n10
  );


  not
  g4
  (
    n49,
    n5
  );


  buf
  g5
  (
    n108,
    n24
  );


  not
  g6
  (
    n82,
    n4
  );


  not
  g7
  (
    n98,
    n19
  );


  buf
  g8
  (
    n83,
    n26
  );


  not
  g9
  (
    n41,
    n23
  );


  not
  g10
  (
    n92,
    n11
  );


  buf
  g11
  (
    n52,
    n12
  );


  not
  g12
  (
    n53,
    n7
  );


  buf
  g13
  (
    KeyWire_0_52,
    n4
  );


  buf
  g14
  (
    n47,
    n15
  );


  buf
  g15
  (
    n91,
    n5
  );


  buf
  g16
  (
    n94,
    n18
  );


  buf
  g17
  (
    n33,
    n14
  );


  not
  g18
  (
    n62,
    n17
  );


  not
  g19
  (
    n70,
    n24
  );


  buf
  g20
  (
    n37,
    n24
  );


  not
  g21
  (
    n107,
    n2
  );


  buf
  g22
  (
    n34,
    n21
  );


  buf
  g23
  (
    n89,
    n16
  );


  buf
  g24
  (
    n60,
    n19
  );


  not
  g25
  (
    n28,
    n1
  );


  buf
  g26
  (
    n43,
    n25
  );


  buf
  g27
  (
    n90,
    n23
  );


  not
  g28
  (
    n128,
    n11
  );


  buf
  g29
  (
    n57,
    n9
  );


  not
  g30
  (
    n30,
    n24
  );


  not
  g31
  (
    n44,
    n18
  );


  not
  g32
  (
    n120,
    n7
  );


  buf
  g33
  (
    n95,
    n16
  );


  buf
  g34
  (
    n106,
    n9
  );


  not
  g35
  (
    n63,
    n19
  );


  buf
  g36
  (
    n127,
    n15
  );


  buf
  g37
  (
    n117,
    n10
  );


  buf
  g38
  (
    n122,
    n3
  );


  not
  g39
  (
    n125,
    n15
  );


  not
  g40
  (
    n99,
    n25
  );


  not
  g41
  (
    n58,
    n23
  );


  not
  g42
  (
    n66,
    n20
  );


  not
  g43
  (
    n65,
    n21
  );


  not
  g44
  (
    n112,
    n22
  );


  buf
  g45
  (
    n102,
    n21
  );


  buf
  g46
  (
    n29,
    n1
  );


  not
  g47
  (
    KeyWire_0_46,
    n14
  );


  buf
  g48
  (
    n85,
    n15
  );


  not
  g49
  (
    n76,
    n6
  );


  not
  g50
  (
    KeyWire_0_1,
    n12
  );


  buf
  g51
  (
    n74,
    n8
  );


  not
  g52
  (
    n32,
    n6
  );


  buf
  g53
  (
    n72,
    n20
  );


  buf
  g54
  (
    n64,
    n26
  );


  buf
  g55
  (
    n71,
    n8
  );


  not
  g56
  (
    n68,
    n22
  );


  not
  g57
  (
    n61,
    n11
  );


  not
  g58
  (
    n55,
    n3
  );


  not
  g59
  (
    n113,
    n5
  );


  buf
  g60
  (
    n111,
    n18
  );


  not
  g61
  (
    n97,
    n23
  );


  not
  g62
  (
    n88,
    n11
  );


  buf
  g63
  (
    n40,
    n3
  );


  not
  g64
  (
    n39,
    n10
  );


  buf
  g65
  (
    n86,
    n14
  );


  buf
  g66
  (
    n105,
    n14
  );


  buf
  g67
  (
    n118,
    n5
  );


  buf
  g68
  (
    n115,
    n6
  );


  not
  g69
  (
    n42,
    n1
  );


  buf
  g70
  (
    n50,
    n12
  );


  buf
  g71
  (
    n101,
    n19
  );


  not
  g72
  (
    n114,
    n22
  );


  buf
  g73
  (
    n79,
    n16
  );


  buf
  g74
  (
    n110,
    n17
  );


  buf
  g75
  (
    n103,
    n8
  );


  not
  g76
  (
    n109,
    n20
  );


  buf
  g77
  (
    n36,
    n8
  );


  not
  g78
  (
    n81,
    n10
  );


  not
  g79
  (
    n104,
    n9
  );


  buf
  g80
  (
    n93,
    n21
  );


  buf
  g81
  (
    n69,
    n25
  );


  buf
  g82
  (
    n124,
    n9
  );


  buf
  g83
  (
    n121,
    n13
  );


  not
  g84
  (
    n75,
    n17
  );


  not
  g85
  (
    n77,
    n1
  );


  buf
  g86
  (
    n59,
    n26
  );


  not
  g87
  (
    n80,
    n13
  );


  buf
  g88
  (
    n78,
    n18
  );


  not
  g89
  (
    n51,
    n25
  );


  buf
  g90
  (
    n116,
    n17
  );


  not
  g91
  (
    n129,
    n2
  );


  buf
  g92
  (
    KeyWire_0_7,
    n6
  );


  buf
  g93
  (
    n31,
    n3
  );


  not
  g94
  (
    n87,
    n7
  );


  not
  g95
  (
    n73,
    n13
  );


  buf
  g96
  (
    n54,
    n20
  );


  buf
  g97
  (
    n48,
    n12
  );


  not
  g98
  (
    n27,
    n2
  );


  buf
  g99
  (
    n119,
    n4
  );


  buf
  g100
  (
    n123,
    n13
  );


  buf
  g101
  (
    n56,
    n7
  );


  not
  g102
  (
    KeyWire_0_34,
    n22
  );


  buf
  g103
  (
    n130,
    n16
  );


  not
  g104
  (
    n394,
    n124
  );


  buf
  g105
  (
    n255,
    n70
  );


  buf
  g106
  (
    n515,
    n95
  );


  not
  g107
  (
    n299,
    n127
  );


  buf
  g108
  (
    n423,
    n69
  );


  not
  g109
  (
    n189,
    n65
  );


  buf
  g110
  (
    KeyWire_0_60,
    n39
  );


  buf
  g111
  (
    n187,
    n30
  );


  not
  g112
  (
    n356,
    n114
  );


  not
  g113
  (
    n155,
    n112
  );


  buf
  g114
  (
    n240,
    n73
  );


  buf
  g115
  (
    n320,
    n77
  );


  buf
  g116
  (
    n408,
    n129
  );


  buf
  g117
  (
    n263,
    n85
  );


  not
  g118
  (
    n289,
    n101
  );


  buf
  g119
  (
    n424,
    n85
  );


  buf
  g120
  (
    KeyWire_0_51,
    n48
  );


  not
  g121
  (
    n532,
    n50
  );


  buf
  g122
  (
    n524,
    n51
  );


  not
  g123
  (
    n301,
    n44
  );


  buf
  g124
  (
    n416,
    n43
  );


  not
  g125
  (
    n495,
    n119
  );


  buf
  g126
  (
    n164,
    n70
  );


  not
  g127
  (
    n251,
    n103
  );


  not
  g128
  (
    n428,
    n67
  );


  buf
  g129
  (
    n481,
    n127
  );


  not
  g130
  (
    n150,
    n87
  );


  not
  g131
  (
    KeyWire_0_25,
    n31
  );


  buf
  g132
  (
    n530,
    n62
  );


  buf
  g133
  (
    n201,
    n105
  );


  not
  g134
  (
    n279,
    n82
  );


  buf
  g135
  (
    n519,
    n97
  );


  buf
  g136
  (
    n329,
    n43
  );


  not
  g137
  (
    n304,
    n35
  );


  buf
  g138
  (
    n466,
    n29
  );


  buf
  g139
  (
    n435,
    n56
  );


  buf
  g140
  (
    n160,
    n44
  );


  buf
  g141
  (
    KeyWire_0_2,
    n51
  );


  buf
  g142
  (
    n199,
    n108
  );


  buf
  g143
  (
    n148,
    n33
  );


  buf
  g144
  (
    n206,
    n111
  );


  not
  g145
  (
    n382,
    n66
  );


  not
  g146
  (
    n285,
    n40
  );


  buf
  g147
  (
    KeyWire_0_30,
    n53
  );


  buf
  g148
  (
    n411,
    n65
  );


  not
  g149
  (
    n476,
    n101
  );


  not
  g150
  (
    n318,
    n98
  );


  buf
  g151
  (
    n173,
    n122
  );


  buf
  g152
  (
    n244,
    n113
  );


  buf
  g153
  (
    n236,
    n68
  );


  not
  g154
  (
    n305,
    n128
  );


  not
  g155
  (
    n259,
    n74
  );


  buf
  g156
  (
    n241,
    n30
  );


  not
  g157
  (
    n494,
    n110
  );


  not
  g158
  (
    n331,
    n40
  );


  not
  g159
  (
    n439,
    n82
  );


  buf
  g160
  (
    n312,
    n95
  );


  not
  g161
  (
    n385,
    n37
  );


  not
  g162
  (
    n488,
    n118
  );


  buf
  g163
  (
    KeyWire_0_54,
    n86
  );


  buf
  g164
  (
    n499,
    n130
  );


  not
  g165
  (
    n485,
    n91
  );


  buf
  g166
  (
    n195,
    n57
  );


  not
  g167
  (
    n307,
    n42
  );


  buf
  g168
  (
    n438,
    n87
  );


  not
  g169
  (
    n309,
    n105
  );


  not
  g170
  (
    n487,
    n50
  );


  buf
  g171
  (
    KeyWire_0_47,
    n28
  );


  not
  g172
  (
    n252,
    n80
  );


  not
  g173
  (
    n381,
    n59
  );


  buf
  g174
  (
    n321,
    n100
  );


  not
  g175
  (
    n174,
    n56
  );


  not
  g176
  (
    n194,
    n49
  );


  not
  g177
  (
    n256,
    n98
  );


  buf
  g178
  (
    n291,
    n74
  );


  not
  g179
  (
    n462,
    n64
  );


  not
  g180
  (
    n340,
    n79
  );


  buf
  g181
  (
    n429,
    n113
  );


  buf
  g182
  (
    n232,
    n100
  );


  not
  g183
  (
    n288,
    n55
  );


  not
  g184
  (
    n149,
    n122
  );


  not
  g185
  (
    n544,
    n61
  );


  buf
  g186
  (
    n358,
    n36
  );


  buf
  g187
  (
    n425,
    n47
  );


  not
  g188
  (
    n245,
    n89
  );


  buf
  g189
  (
    n175,
    n83
  );


  buf
  g190
  (
    n469,
    n94
  );


  buf
  g191
  (
    n342,
    n128
  );


  not
  g192
  (
    n351,
    n58
  );


  buf
  g193
  (
    n503,
    n72
  );


  buf
  g194
  (
    n498,
    n130
  );


  not
  g195
  (
    n354,
    n102
  );


  not
  g196
  (
    n242,
    n79
  );


  buf
  g197
  (
    n138,
    n67
  );


  buf
  g198
  (
    n541,
    n45
  );


  not
  g199
  (
    n396,
    n92
  );


  buf
  g200
  (
    n357,
    n64
  );


  not
  g201
  (
    n190,
    n49
  );


  buf
  g202
  (
    n296,
    n27
  );


  buf
  g203
  (
    n426,
    n62
  );


  buf
  g204
  (
    n414,
    n64
  );


  not
  g205
  (
    n472,
    n111
  );


  not
  g206
  (
    n520,
    n35
  );


  not
  g207
  (
    KeyWire_0_4,
    n109
  );


  buf
  g208
  (
    n336,
    n124
  );


  not
  g209
  (
    n440,
    n120
  );


  buf
  g210
  (
    n311,
    n61
  );


  not
  g211
  (
    n379,
    n54
  );


  buf
  g212
  (
    n167,
    n59
  );


  not
  g213
  (
    n225,
    n41
  );


  not
  g214
  (
    n389,
    n59
  );


  not
  g215
  (
    n172,
    n72
  );


  not
  g216
  (
    n535,
    n47
  );


  not
  g217
  (
    n516,
    n105
  );


  not
  g218
  (
    n538,
    n115
  );


  not
  g219
  (
    n184,
    n76
  );


  not
  g220
  (
    n243,
    n92
  );


  not
  g221
  (
    n412,
    n45
  );


  not
  g222
  (
    n274,
    n111
  );


  not
  g223
  (
    n267,
    n129
  );


  buf
  g224
  (
    n310,
    n129
  );


  buf
  g225
  (
    n334,
    n120
  );


  not
  g226
  (
    n161,
    n112
  );


  buf
  g227
  (
    n246,
    n116
  );


  not
  g228
  (
    n393,
    n117
  );


  not
  g229
  (
    n493,
    n75
  );


  not
  g230
  (
    n168,
    n115
  );


  buf
  g231
  (
    n355,
    n113
  );


  buf
  g232
  (
    n276,
    n28
  );


  buf
  g233
  (
    n534,
    n106
  );


  buf
  g234
  (
    n402,
    n125
  );


  not
  g235
  (
    n446,
    n121
  );


  not
  g236
  (
    KeyWire_0_17,
    n39
  );


  not
  g237
  (
    n217,
    n93
  );


  buf
  g238
  (
    n445,
    n70
  );


  buf
  g239
  (
    n509,
    n96
  );


  not
  g240
  (
    n459,
    n86
  );


  not
  g241
  (
    n457,
    n117
  );


  buf
  g242
  (
    n395,
    n93
  );


  not
  g243
  (
    n529,
    n34
  );


  buf
  g244
  (
    n480,
    n49
  );


  not
  g245
  (
    n448,
    n29
  );


  buf
  g246
  (
    n237,
    n121
  );


  not
  g247
  (
    n332,
    n100
  );


  not
  g248
  (
    n370,
    n93
  );


  not
  g249
  (
    n227,
    n40
  );


  buf
  g250
  (
    n341,
    n126
  );


  not
  g251
  (
    n271,
    n71
  );


  not
  g252
  (
    n364,
    n107
  );


  not
  g253
  (
    n328,
    n52
  );


  buf
  g254
  (
    n543,
    n102
  );


  not
  g255
  (
    n162,
    n60
  );


  buf
  g256
  (
    n359,
    n27
  );


  not
  g257
  (
    n501,
    n113
  );


  buf
  g258
  (
    n292,
    n57
  );


  not
  g259
  (
    n421,
    n37
  );


  buf
  g260
  (
    n514,
    n118
  );


  not
  g261
  (
    n221,
    n95
  );


  not
  g262
  (
    n506,
    n36
  );


  buf
  g263
  (
    n179,
    n119
  );


  buf
  g264
  (
    n399,
    n53
  );


  buf
  g265
  (
    n275,
    n66
  );


  buf
  g266
  (
    n250,
    n35
  );


  not
  g267
  (
    n171,
    n52
  );


  buf
  g268
  (
    n436,
    n73
  );


  buf
  g269
  (
    n343,
    n109
  );


  buf
  g270
  (
    n369,
    n41
  );


  buf
  g271
  (
    n204,
    n74
  );


  not
  g272
  (
    n239,
    n99
  );


  not
  g273
  (
    KeyWire_0_33,
    n46
  );


  not
  g274
  (
    n475,
    n85
  );


  not
  g275
  (
    n400,
    n109
  );


  not
  g276
  (
    n388,
    n29
  );


  buf
  g277
  (
    n461,
    n29
  );


  buf
  g278
  (
    n384,
    n50
  );


  buf
  g279
  (
    n234,
    n119
  );


  not
  g280
  (
    n387,
    n77
  );


  not
  g281
  (
    n193,
    n108
  );


  not
  g282
  (
    n365,
    n94
  );


  not
  g283
  (
    n492,
    n71
  );


  not
  g284
  (
    n235,
    n32
  );


  not
  g285
  (
    n473,
    n116
  );


  buf
  g286
  (
    n185,
    n119
  );


  buf
  g287
  (
    n135,
    n54
  );


  buf
  g288
  (
    n441,
    n27
  );


  not
  g289
  (
    n474,
    n91
  );


  buf
  g290
  (
    n390,
    n89
  );


  buf
  g291
  (
    n181,
    n111
  );


  buf
  g292
  (
    n373,
    n64
  );


  buf
  g293
  (
    n542,
    n103
  );


  buf
  g294
  (
    n319,
    n92
  );


  buf
  g295
  (
    n407,
    n74
  );


  not
  g296
  (
    n266,
    n48
  );


  not
  g297
  (
    n368,
    n99
  );


  buf
  g298
  (
    KeyWire_0_13,
    n75
  );


  buf
  g299
  (
    n419,
    n31
  );


  not
  g300
  (
    n417,
    n38
  );


  not
  g301
  (
    n497,
    n90
  );


  not
  g302
  (
    n323,
    n68
  );


  not
  g303
  (
    n418,
    n83
  );


  not
  g304
  (
    n208,
    n61
  );


  not
  g305
  (
    n460,
    n97
  );


  buf
  g306
  (
    n145,
    n46
  );


  not
  g307
  (
    n451,
    n89
  );


  buf
  g308
  (
    n360,
    n105
  );


  buf
  g309
  (
    n484,
    n81
  );


  buf
  g310
  (
    n152,
    n88
  );


  buf
  g311
  (
    n182,
    n95
  );


  buf
  g312
  (
    n437,
    n55
  );


  buf
  g313
  (
    n410,
    n122
  );


  not
  g314
  (
    n537,
    n110
  );


  not
  g315
  (
    n264,
    n36
  );


  buf
  g316
  (
    n531,
    n103
  );


  not
  g317
  (
    n447,
    n77
  );


  buf
  g318
  (
    n527,
    n125
  );


  not
  g319
  (
    n479,
    n45
  );


  not
  g320
  (
    n432,
    n94
  );


  buf
  g321
  (
    n482,
    n86
  );


  not
  g322
  (
    n330,
    n127
  );


  buf
  g323
  (
    n386,
    n75
  );


  buf
  g324
  (
    KeyWire_0_49,
    n115
  );


  not
  g325
  (
    n265,
    n54
  );


  not
  g326
  (
    n504,
    n63
  );


  buf
  g327
  (
    n324,
    n116
  );


  buf
  g328
  (
    n218,
    n114
  );


  not
  g329
  (
    n283,
    n97
  );


  not
  g330
  (
    n362,
    n78
  );


  not
  g331
  (
    n133,
    n32
  );


  buf
  g332
  (
    n261,
    n126
  );


  not
  g333
  (
    n219,
    n51
  );


  not
  g334
  (
    n147,
    n104
  );


  not
  g335
  (
    n545,
    n128
  );


  buf
  g336
  (
    n391,
    n84
  );


  buf
  g337
  (
    n293,
    n51
  );


  buf
  g338
  (
    n280,
    n104
  );


  buf
  g339
  (
    n202,
    n98
  );


  not
  g340
  (
    n380,
    n33
  );


  not
  g341
  (
    n361,
    n88
  );


  not
  g342
  (
    n348,
    n116
  );


  not
  g343
  (
    n282,
    n40
  );


  not
  g344
  (
    n143,
    n27
  );


  not
  g345
  (
    n372,
    n87
  );


  buf
  g346
  (
    n486,
    n96
  );


  buf
  g347
  (
    n277,
    n129
  );


  not
  g348
  (
    n403,
    n126
  );


  buf
  g349
  (
    n508,
    n54
  );


  not
  g350
  (
    n347,
    n48
  );


  buf
  g351
  (
    n231,
    n104
  );


  buf
  g352
  (
    n525,
    n81
  );


  not
  g353
  (
    n518,
    n124
  );


  not
  g354
  (
    n196,
    n78
  );


  not
  g355
  (
    n298,
    n32
  );


  not
  g356
  (
    KeyWire_0_10,
    n57
  );


  buf
  g357
  (
    n496,
    n127
  );


  buf
  g358
  (
    n316,
    n85
  );


  buf
  g359
  (
    n270,
    n102
  );


  not
  g360
  (
    n349,
    n91
  );


  buf
  g361
  (
    n197,
    n120
  );


  buf
  g362
  (
    n207,
    n88
  );


  not
  g363
  (
    n213,
    n106
  );


  buf
  g364
  (
    n546,
    n109
  );


  buf
  g365
  (
    n353,
    n28
  );


  buf
  g366
  (
    n502,
    n106
  );


  not
  g367
  (
    n450,
    n44
  );


  buf
  g368
  (
    n224,
    n82
  );


  not
  g369
  (
    n470,
    n38
  );


  buf
  g370
  (
    n272,
    n34
  );


  buf
  g371
  (
    KeyWire_0_19,
    n128
  );


  not
  g372
  (
    n281,
    n117
  );


  not
  g373
  (
    n183,
    n47
  );


  buf
  g374
  (
    n452,
    n86
  );


  not
  g375
  (
    n223,
    n94
  );


  buf
  g376
  (
    n464,
    n34
  );


  buf
  g377
  (
    n322,
    n50
  );


  buf
  g378
  (
    n521,
    n48
  );


  not
  g379
  (
    n453,
    n76
  );


  not
  g380
  (
    n352,
    n110
  );


  buf
  g381
  (
    n229,
    n58
  );


  not
  g382
  (
    n415,
    n123
  );


  not
  g383
  (
    n366,
    n39
  );


  not
  g384
  (
    KeyWire_0_35,
    n71
  );


  not
  g385
  (
    n404,
    n102
  );


  not
  g386
  (
    n378,
    n123
  );


  not
  g387
  (
    n420,
    n120
  );


  not
  g388
  (
    n203,
    n114
  );


  buf
  g389
  (
    n533,
    n121
  );


  buf
  g390
  (
    n490,
    n130
  );


  buf
  g391
  (
    n491,
    n90
  );


  not
  g392
  (
    n191,
    n38
  );


  buf
  g393
  (
    n159,
    n130
  );


  not
  g394
  (
    n401,
    n73
  );


  not
  g395
  (
    KeyWire_0_57,
    n83
  );


  not
  g396
  (
    n313,
    n80
  );


  buf
  g397
  (
    n434,
    n106
  );


  not
  g398
  (
    n295,
    n108
  );


  not
  g399
  (
    n297,
    n60
  );


  not
  g400
  (
    n338,
    n55
  );


  not
  g401
  (
    n214,
    n38
  );


  buf
  g402
  (
    n269,
    n87
  );


  buf
  g403
  (
    n489,
    n72
  );


  buf
  g404
  (
    n383,
    n36
  );


  not
  g405
  (
    n144,
    n117
  );


  buf
  g406
  (
    n463,
    n30
  );


  buf
  g407
  (
    n294,
    n96
  );


  not
  g408
  (
    n146,
    n52
  );


  not
  g409
  (
    n180,
    n69
  );


  buf
  g410
  (
    n216,
    n41
  );


  not
  g411
  (
    n539,
    n114
  );


  buf
  g412
  (
    n156,
    n107
  );


  buf
  g413
  (
    KeyWire_0_45,
    n99
  );


  buf
  g414
  (
    n376,
    n76
  );


  not
  g415
  (
    n248,
    n98
  );


  buf
  g416
  (
    n536,
    n62
  );


  buf
  g417
  (
    n517,
    n83
  );


  buf
  g418
  (
    n137,
    n80
  );


  buf
  g419
  (
    n230,
    n67
  );


  buf
  g420
  (
    KeyWire_0_0,
    n122
  );


  not
  g421
  (
    n317,
    n118
  );


  not
  g422
  (
    n131,
    n79
  );


  not
  g423
  (
    KeyWire_0_32,
    n66
  );


  not
  g424
  (
    n188,
    n53
  );


  not
  g425
  (
    KeyWire_0_28,
    n93
  );


  buf
  g426
  (
    n284,
    n84
  );


  buf
  g427
  (
    n468,
    n33
  );


  buf
  g428
  (
    n247,
    n97
  );


  buf
  g429
  (
    n507,
    n82
  );


  not
  g430
  (
    n513,
    n79
  );


  not
  g431
  (
    n153,
    n57
  );


  not
  g432
  (
    n132,
    n110
  );


  not
  g433
  (
    n178,
    n32
  );


  not
  g434
  (
    n170,
    n72
  );


  buf
  g435
  (
    n141,
    n60
  );


  buf
  g436
  (
    n290,
    n43
  );


  not
  g437
  (
    n413,
    n42
  );


  buf
  g438
  (
    n215,
    n42
  );


  buf
  g439
  (
    n158,
    n56
  );


  not
  g440
  (
    n306,
    n107
  );


  buf
  g441
  (
    n374,
    n69
  );


  not
  g442
  (
    n371,
    n78
  );


  not
  g443
  (
    n142,
    n77
  );


  buf
  g444
  (
    n210,
    n104
  );


  not
  g445
  (
    n262,
    n80
  );


  buf
  g446
  (
    n200,
    n60
  );


  buf
  g447
  (
    n136,
    n58
  );


  buf
  g448
  (
    KeyWire_0_26,
    n46
  );


  not
  g449
  (
    n166,
    n90
  );


  buf
  g450
  (
    n406,
    n53
  );


  not
  g451
  (
    n505,
    n30
  );


  not
  g452
  (
    n335,
    n35
  );


  not
  g453
  (
    n222,
    n33
  );


  buf
  g454
  (
    n163,
    n124
  );


  not
  g455
  (
    n367,
    n121
  );


  buf
  g456
  (
    n500,
    n107
  );


  not
  g457
  (
    n212,
    n81
  );


  buf
  g458
  (
    n327,
    n126
  );


  not
  g459
  (
    n444,
    n49
  );


  buf
  g460
  (
    n165,
    n84
  );


  not
  g461
  (
    n465,
    n112
  );


  buf
  g462
  (
    n430,
    n76
  );


  not
  g463
  (
    n422,
    n123
  );


  buf
  g464
  (
    n134,
    n63
  );


  buf
  g465
  (
    n169,
    n75
  );


  buf
  g466
  (
    n140,
    n103
  );


  not
  g467
  (
    n409,
    n66
  );


  buf
  g468
  (
    n375,
    n118
  );


  buf
  g469
  (
    n467,
    n91
  );


  not
  g470
  (
    n209,
    n34
  );


  not
  g471
  (
    n392,
    n55
  );


  not
  g472
  (
    n456,
    n52
  );


  buf
  g473
  (
    n257,
    n28
  );


  not
  g474
  (
    n337,
    n108
  );


  buf
  g475
  (
    n192,
    n58
  );


  buf
  g476
  (
    n302,
    n68
  );


  not
  g477
  (
    n471,
    n39
  );


  not
  g478
  (
    n238,
    n43
  );


  buf
  g479
  (
    n512,
    n63
  );


  not
  g480
  (
    KeyWire_0_58,
    n96
  );


  not
  g481
  (
    n249,
    n101
  );


  buf
  g482
  (
    n300,
    n73
  );


  buf
  g483
  (
    n540,
    n92
  );


  not
  g484
  (
    n431,
    n41
  );


  not
  g485
  (
    n398,
    n125
  );


  buf
  g486
  (
    n346,
    n88
  );


  buf
  g487
  (
    n177,
    n100
  );


  buf
  g488
  (
    n186,
    n44
  );


  not
  g489
  (
    n308,
    n84
  );


  buf
  g490
  (
    n278,
    n61
  );


  buf
  g491
  (
    n455,
    n37
  );


  not
  g492
  (
    n427,
    n125
  );


  buf
  g493
  (
    n314,
    n37
  );


  buf
  g494
  (
    n258,
    n47
  );


  not
  g495
  (
    n139,
    n31
  );


  not
  g496
  (
    n233,
    n101
  );


  not
  g497
  (
    n253,
    n46
  );


  not
  g498
  (
    n458,
    n42
  );


  buf
  g499
  (
    n325,
    n115
  );


  buf
  g500
  (
    n326,
    n59
  );


  buf
  g501
  (
    n198,
    n31
  );


  not
  g502
  (
    n510,
    n68
  );


  buf
  g503
  (
    n344,
    n112
  );


  buf
  g504
  (
    n405,
    n99
  );


  buf
  g505
  (
    n315,
    n70
  );


  not
  g506
  (
    n205,
    n62
  );


  not
  g507
  (
    n449,
    n45
  );


  buf
  g508
  (
    n220,
    n69
  );


  buf
  g509
  (
    n443,
    n78
  );


  buf
  g510
  (
    n303,
    n90
  );


  buf
  g511
  (
    n226,
    n71
  );


  buf
  g512
  (
    n154,
    n65
  );


  buf
  g513
  (
    n511,
    n65
  );


  not
  g514
  (
    n523,
    n67
  );


  not
  g515
  (
    n526,
    n81
  );


  not
  g516
  (
    n254,
    n89
  );


  buf
  g517
  (
    n397,
    n123
  );


  not
  g518
  (
    n442,
    n63
  );


  buf
  g519
  (
    n350,
    n56
  );


  not
  g520
  (
    n547,
    n134
  );


  buf
  g521
  (
    n550,
    n133
  );


  buf
  g522
  (
    n549,
    n131
  );


  buf
  g523
  (
    n548,
    n132
  );


  nor
  g524
  (
    n553,
    n140,
    n168,
    n181,
    n550
  );


  nand
  g525
  (
    n560,
    n142,
    n138,
    n548,
    n148
  );


  xor
  g526
  (
    KeyWire_0_50,
    n139,
    n151,
    n150,
    n165
  );


  nand
  g527
  (
    n565,
    n170,
    n163,
    n167,
    n147
  );


  xnor
  g528
  (
    n556,
    n550,
    n145,
    n164,
    n547
  );


  xor
  g529
  (
    n564,
    n160,
    n156,
    n161,
    n152
  );


  xor
  g530
  (
    n561,
    n166,
    n171,
    n143,
    n182
  );


  xnor
  g531
  (
    n551,
    n175,
    n550,
    n548,
    n179
  );


  xnor
  g532
  (
    KeyWire_0_40,
    n172,
    n153,
    n149,
    n169
  );


  nor
  g533
  (
    n558,
    n155,
    n549,
    n141
  );


  or
  g534
  (
    n563,
    n549,
    n548,
    n162,
    n146
  );


  xnor
  g535
  (
    n555,
    n144,
    n176,
    n549,
    n178
  );


  nor
  g536
  (
    n562,
    n135,
    n137,
    n180,
    n548
  );


  nand
  g537
  (
    n557,
    n173,
    n174,
    n158,
    n547
  );


  or
  g538
  (
    n566,
    n136,
    n547,
    n159
  );


  and
  g539
  (
    n552,
    n154,
    n550,
    n177,
    n157
  );


  buf
  g540
  (
    n587,
    n554
  );


  not
  g541
  (
    n578,
    n561
  );


  not
  g542
  (
    n576,
    n562
  );


  buf
  g543
  (
    n608,
    n551
  );


  not
  g544
  (
    n601,
    n557
  );


  not
  g545
  (
    KeyWire_0_6,
    n565
  );


  buf
  g546
  (
    n583,
    n558
  );


  buf
  g547
  (
    n597,
    n556
  );


  not
  g548
  (
    n616,
    n560
  );


  buf
  g549
  (
    n577,
    n556
  );


  not
  g550
  (
    KeyWire_0_11,
    n562
  );


  buf
  g551
  (
    n584,
    n559
  );


  not
  g552
  (
    n590,
    n563
  );


  buf
  g553
  (
    n607,
    n562
  );


  buf
  g554
  (
    n572,
    n565
  );


  not
  g555
  (
    n586,
    n558
  );


  not
  g556
  (
    n605,
    n555
  );


  buf
  g557
  (
    n606,
    n558
  );


  buf
  g558
  (
    n610,
    n555
  );


  not
  g559
  (
    n594,
    n565
  );


  buf
  g560
  (
    n588,
    n564
  );


  not
  g561
  (
    n580,
    n552
  );


  not
  g562
  (
    KeyWire_0_3,
    n553
  );


  not
  g563
  (
    n585,
    n557
  );


  buf
  g564
  (
    n600,
    n566
  );


  buf
  g565
  (
    n567,
    n183
  );


  buf
  g566
  (
    n579,
    n564
  );


  buf
  g567
  (
    n581,
    n557
  );


  not
  g568
  (
    n603,
    n565
  );


  buf
  g569
  (
    n582,
    n559
  );


  not
  g570
  (
    n593,
    n564
  );


  buf
  g571
  (
    n592,
    n563
  );


  not
  g572
  (
    n599,
    n566
  );


  buf
  g573
  (
    n571,
    n559
  );


  buf
  g574
  (
    n609,
    n557
  );


  buf
  g575
  (
    n602,
    n563
  );


  not
  g576
  (
    n604,
    n564
  );


  not
  g577
  (
    n598,
    n561
  );


  not
  g578
  (
    n615,
    n560
  );


  buf
  g579
  (
    n596,
    n563
  );


  buf
  g580
  (
    n575,
    n560
  );


  not
  g581
  (
    KeyWire_0_23,
    n561
  );


  not
  g582
  (
    n591,
    n561
  );


  not
  g583
  (
    n569,
    n556
  );


  not
  g584
  (
    n612,
    n562
  );


  buf
  g585
  (
    KeyWire_0_22,
    n559
  );


  not
  g586
  (
    n570,
    n566
  );


  buf
  g587
  (
    n568,
    n566
  );


  buf
  g588
  (
    n574,
    n558
  );


  xnor
  g589
  (
    n613,
    n556,
    n560
  );


  buf
  g590
  (
    n707,
    n611
  );


  not
  g591
  (
    n728,
    n276
  );


  buf
  g592
  (
    n665,
    n614
  );


  buf
  g593
  (
    n810,
    n584
  );


  buf
  g594
  (
    n736,
    n587
  );


  buf
  g595
  (
    n759,
    n206
  );


  buf
  g596
  (
    n708,
    n341
  );


  not
  g597
  (
    n706,
    n603
  );


  not
  g598
  (
    n625,
    n312
  );


  buf
  g599
  (
    n714,
    n187
  );


  buf
  g600
  (
    n619,
    n346
  );


  not
  g601
  (
    n727,
    n259
  );


  buf
  g602
  (
    n797,
    n610
  );


  not
  g603
  (
    n656,
    n227
  );


  not
  g604
  (
    n791,
    n243
  );


  buf
  g605
  (
    n778,
    n280
  );


  buf
  g606
  (
    n767,
    n256
  );


  not
  g607
  (
    KeyWire_0_39,
    n591
  );


  buf
  g608
  (
    n768,
    n592
  );


  buf
  g609
  (
    n765,
    n577
  );


  buf
  g610
  (
    n723,
    n580
  );


  not
  g611
  (
    n637,
    n609
  );


  not
  g612
  (
    n772,
    n596
  );


  buf
  g613
  (
    n648,
    n188
  );


  buf
  g614
  (
    n636,
    n198
  );


  not
  g615
  (
    n678,
    n260
  );


  not
  g616
  (
    n710,
    n201
  );


  not
  g617
  (
    n680,
    n594
  );


  not
  g618
  (
    n682,
    n572
  );


  not
  g619
  (
    n694,
    n569
  );


  not
  g620
  (
    n660,
    n607
  );


  not
  g621
  (
    n739,
    n615
  );


  buf
  g622
  (
    n807,
    n599
  );


  not
  g623
  (
    n734,
    n571
  );


  buf
  g624
  (
    n691,
    n586
  );


  not
  g625
  (
    n782,
    n599
  );


  not
  g626
  (
    n779,
    n612
  );


  buf
  g627
  (
    n679,
    n269
  );


  buf
  g628
  (
    n742,
    n330
  );


  buf
  g629
  (
    n649,
    n306
  );


  buf
  g630
  (
    n731,
    n602
  );


  not
  g631
  (
    n754,
    n342
  );


  not
  g632
  (
    n787,
    n610
  );


  not
  g633
  (
    n738,
    n345
  );


  buf
  g634
  (
    n816,
    n594
  );


  not
  g635
  (
    n662,
    n303
  );


  buf
  g636
  (
    n716,
    n257
  );


  buf
  g637
  (
    n666,
    n578
  );


  buf
  g638
  (
    n645,
    n574
  );


  buf
  g639
  (
    n766,
    n592
  );


  not
  g640
  (
    n774,
    n592
  );


  buf
  g641
  (
    n740,
    n604
  );


  not
  g642
  (
    n663,
    n570
  );


  buf
  g643
  (
    n659,
    n231
  );


  not
  g644
  (
    n721,
    n321
  );


  buf
  g645
  (
    n757,
    n229
  );


  buf
  g646
  (
    n802,
    n262
  );


  not
  g647
  (
    n642,
    n591
  );


  not
  g648
  (
    n681,
    n576
  );


  buf
  g649
  (
    n713,
    n598
  );


  not
  g650
  (
    n805,
    n203
  );


  buf
  g651
  (
    n755,
    n212
  );


  not
  g652
  (
    n704,
    n241
  );


  not
  g653
  (
    n777,
    n258
  );


  buf
  g654
  (
    n758,
    n576
  );


  buf
  g655
  (
    n812,
    n239
  );


  not
  g656
  (
    KeyWire_0_29,
    n595
  );


  not
  g657
  (
    n633,
    n591
  );


  buf
  g658
  (
    n654,
    n585
  );


  buf
  g659
  (
    n630,
    n611
  );


  not
  g660
  (
    n687,
    n593
  );


  not
  g661
  (
    n719,
    n613
  );


  buf
  g662
  (
    n617,
    n587
  );


  buf
  g663
  (
    n690,
    n582
  );


  not
  g664
  (
    n703,
    n214
  );


  buf
  g665
  (
    n650,
    n605
  );


  not
  g666
  (
    n792,
    n308
  );


  not
  g667
  (
    n638,
    n592
  );


  buf
  g668
  (
    n702,
    n249
  );


  buf
  g669
  (
    n788,
    n575
  );


  not
  g670
  (
    KeyWire_0_9,
    n602
  );


  not
  g671
  (
    n647,
    n573
  );


  not
  g672
  (
    n726,
    n568
  );


  not
  g673
  (
    n724,
    n254
  );


  buf
  g674
  (
    n790,
    n590
  );


  not
  g675
  (
    KeyWire_0_41,
    n583
  );


  not
  g676
  (
    n785,
    n575
  );


  not
  g677
  (
    n641,
    n284
  );


  buf
  g678
  (
    n770,
    n612
  );


  not
  g679
  (
    n798,
    n593
  );


  buf
  g680
  (
    n639,
    n317
  );


  not
  g681
  (
    n669,
    n261
  );


  not
  g682
  (
    n671,
    n577
  );


  buf
  g683
  (
    n741,
    n604
  );


  not
  g684
  (
    n756,
    n221
  );


  not
  g685
  (
    n764,
    n586
  );


  buf
  g686
  (
    n729,
    n574
  );


  not
  g687
  (
    n701,
    n602
  );


  not
  g688
  (
    n796,
    n235
  );


  not
  g689
  (
    KeyWire_0_20,
    n573
  );


  buf
  g690
  (
    n709,
    n304
  );


  not
  g691
  (
    n705,
    n607
  );


  buf
  g692
  (
    n771,
    n596
  );


  not
  g693
  (
    n711,
    n238
  );


  buf
  g694
  (
    n811,
    n608
  );


  not
  g695
  (
    n730,
    n323
  );


  not
  g696
  (
    KeyWire_0_5,
    n339
  );


  not
  g697
  (
    n717,
    n216
  );


  not
  g698
  (
    n676,
    n291
  );


  not
  g699
  (
    n698,
    n237
  );


  buf
  g700
  (
    n688,
    n287
  );


  buf
  g701
  (
    n808,
    n614
  );


  not
  g702
  (
    n794,
    n332
  );


  buf
  g703
  (
    n735,
    n598
  );


  not
  g704
  (
    n627,
    n596
  );


  not
  g705
  (
    n699,
    n575
  );


  buf
  g706
  (
    n786,
    n213
  );


  or
  g707
  (
    n628,
    n606,
    n570
  );


  nand
  g708
  (
    n799,
    n574,
    n603,
    n569
  );


  nor
  g709
  (
    n806,
    n185,
    n584,
    n211
  );


  xnor
  g710
  (
    n780,
    n275,
    n605,
    n616
  );


  nand
  g711
  (
    n763,
    n298,
    n589,
    n594
  );


  or
  g712
  (
    n652,
    n606,
    n569,
    n571
  );


  or
  g713
  (
    n775,
    n595,
    n322,
    n334
  );


  xnor
  g714
  (
    n675,
    n290,
    n593,
    n265
  );


  nor
  g715
  (
    n651,
    n193,
    n587,
    n604
  );


  or
  g716
  (
    n664,
    n293,
    n315,
    n569
  );


  nor
  g717
  (
    n658,
    n347,
    n590,
    n319
  );


  or
  g718
  (
    n684,
    n255,
    n210,
    n335
  );


  nand
  g719
  (
    n640,
    n578,
    n200,
    n307
  );


  nor
  g720
  (
    n635,
    n197,
    n208,
    n190
  );


  xnor
  g721
  (
    n769,
    n314,
    n266,
    n595
  );


  nand
  g722
  (
    n624,
    n340,
    n209,
    n590
  );


  or
  g723
  (
    n644,
    n612,
    n297,
    n609
  );


  xor
  g724
  (
    n720,
    n585,
    n184,
    n601
  );


  and
  g725
  (
    n693,
    n578,
    n600,
    n590
  );


  and
  g726
  (
    n745,
    n609,
    n616,
    n604
  );


  and
  g727
  (
    n631,
    n337,
    n348,
    n250
  );


  nor
  g728
  (
    n781,
    n300,
    n274,
    n302
  );


  nand
  g729
  (
    n661,
    n199,
    n588,
    n584
  );


  nand
  g730
  (
    n689,
    n600,
    n579,
    n202
  );


  and
  g731
  (
    n732,
    n615,
    n224,
    n582
  );


  nand
  g732
  (
    KeyWire_0_8,
    n603,
    n244,
    n586
  );


  nand
  g733
  (
    n773,
    n613,
    n585,
    n606
  );


  or
  g734
  (
    n683,
    n579,
    n233,
    n578
  );


  and
  g735
  (
    n750,
    n579,
    n272,
    n207
  );


  nand
  g736
  (
    n695,
    n246,
    n600,
    n324
  );


  nand
  g737
  (
    n718,
    n597,
    n325,
    n277
  );


  and
  g738
  (
    n621,
    n326,
    n616,
    n613
  );


  xor
  g739
  (
    n747,
    n205,
    n567
  );


  nor
  g740
  (
    n809,
    n316,
    n593,
    n226
  );


  xor
  g741
  (
    n804,
    n572,
    n584,
    n601
  );


  nand
  g742
  (
    n795,
    n311,
    n583,
    n573
  );


  nand
  g743
  (
    n783,
    n613,
    n299,
    n248
  );


  xor
  g744
  (
    n632,
    n601,
    n580,
    n264
  );


  or
  g745
  (
    n634,
    n580,
    n286,
    n581
  );


  xor
  g746
  (
    n801,
    n236,
    n570,
    n610
  );


  nor
  g747
  (
    n712,
    n338,
    n279,
    n327
  );


  xor
  g748
  (
    n629,
    n575,
    n587,
    n283
  );


  or
  g749
  (
    n618,
    n245,
    n615,
    n567
  );


  xnor
  g750
  (
    n749,
    n242,
    n574,
    n252
  );


  or
  g751
  (
    n653,
    n196,
    n582,
    n218
  );


  nor
  g752
  (
    n762,
    n596,
    n570,
    n610
  );


  xor
  g753
  (
    n753,
    n320,
    n605,
    n594
  );


  xor
  g754
  (
    n743,
    n285,
    n597,
    n189
  );


  or
  g755
  (
    n620,
    n599,
    n344,
    n568
  );


  xor
  g756
  (
    n670,
    n586,
    n568,
    n605
  );


  or
  g757
  (
    n751,
    n576,
    n278,
    n288
  );


  and
  g758
  (
    n668,
    n294,
    n606,
    n585
  );


  nand
  g759
  (
    KeyWire_0_24,
    n267,
    n607,
    n194
  );


  and
  g760
  (
    KeyWire_0_59,
    n295,
    n583,
    n331
  );


  or
  g761
  (
    n776,
    n270,
    n230,
    n580
  );


  nor
  g762
  (
    n815,
    n310,
    n318,
    n329
  );


  xnor
  g763
  (
    n643,
    n273,
    n577,
    n228
  );


  and
  g764
  (
    n626,
    n232,
    n268,
    n296
  );


  nor
  g765
  (
    n748,
    n333,
    n195,
    n271
  );


  xor
  g766
  (
    n692,
    n215,
    n282,
    n225
  );


  or
  g767
  (
    n646,
    n615,
    n598,
    n336
  );


  and
  g768
  (
    n686,
    n616,
    n600,
    n191
  );


  xnor
  g769
  (
    n746,
    n234,
    n220,
    n263
  );


  or
  g770
  (
    KeyWire_0_44,
    n597,
    n222,
    n611
  );


  xor
  g771
  (
    n744,
    n281,
    n614,
    n588
  );


  or
  g772
  (
    KeyWire_0_18,
    n253,
    n223,
    n599
  );


  nand
  g773
  (
    n700,
    n219,
    n589,
    n247
  );


  xnor
  g774
  (
    n674,
    n579,
    n589
  );


  nand
  g775
  (
    n737,
    n608,
    n595,
    n240
  );


  nor
  g776
  (
    n752,
    n591,
    n289,
    n582
  );


  xnor
  g777
  (
    n623,
    n581,
    n301,
    n292
  );


  or
  g778
  (
    n655,
    n609,
    n611,
    n572
  );


  and
  g779
  (
    n803,
    n577,
    n572,
    n217
  );


  and
  g780
  (
    n789,
    n305,
    n571,
    n614
  );


  and
  g781
  (
    n814,
    n607,
    n309,
    n204
  );


  xnor
  g782
  (
    n677,
    n583,
    n588,
    n573
  );


  and
  g783
  (
    n657,
    n608,
    n588,
    n612
  );


  xor
  g784
  (
    n761,
    n598,
    n597,
    n576
  );


  nand
  g785
  (
    n725,
    n192,
    n567,
    n571
  );


  xnor
  g786
  (
    n793,
    n602,
    n603,
    n251
  );


  nor
  g787
  (
    KeyWire_0_63,
    n581,
    n186,
    n328
  );


  nand
  g788
  (
    n722,
    n581,
    n343,
    n313
  );


  xor
  g789
  (
    n685,
    n568,
    n608,
    n601
  );


  not
  g790
  (
    KeyWire_0_27,
    n803
  );


  buf
  g791
  (
    n884,
    n675
  );


  buf
  g792
  (
    n998,
    n641
  );


  not
  g793
  (
    n1134,
    n639
  );


  buf
  g794
  (
    n1013,
    n791
  );


  not
  g795
  (
    n1109,
    n808
  );


  buf
  g796
  (
    n888,
    n759
  );


  buf
  g797
  (
    n1062,
    n701
  );


  not
  g798
  (
    n1161,
    n660
  );


  not
  g799
  (
    n864,
    n624
  );


  buf
  g800
  (
    n945,
    n807
  );


  buf
  g801
  (
    n1046,
    n711
  );


  buf
  g802
  (
    n1123,
    n623
  );


  not
  g803
  (
    n1101,
    n702
  );


  not
  g804
  (
    n970,
    n643
  );


  buf
  g805
  (
    n1120,
    n721
  );


  buf
  g806
  (
    n1107,
    n802
  );


  buf
  g807
  (
    n876,
    n751
  );


  not
  g808
  (
    n978,
    n763
  );


  not
  g809
  (
    n1130,
    n634
  );


  not
  g810
  (
    n880,
    n746
  );


  not
  g811
  (
    n841,
    n727
  );


  buf
  g812
  (
    n933,
    n638
  );


  buf
  g813
  (
    n829,
    n693
  );


  buf
  g814
  (
    n883,
    n729
  );


  buf
  g815
  (
    n1063,
    n689
  );


  buf
  g816
  (
    n999,
    n814
  );


  buf
  g817
  (
    n1100,
    n790
  );


  buf
  g818
  (
    n1069,
    n695
  );


  buf
  g819
  (
    n895,
    n807
  );


  not
  g820
  (
    n1086,
    n633
  );


  buf
  g821
  (
    n1111,
    n631
  );


  not
  g822
  (
    n832,
    n733
  );


  buf
  g823
  (
    n1164,
    n699
  );


  buf
  g824
  (
    n1000,
    n702
  );


  not
  g825
  (
    n937,
    n741
  );


  not
  g826
  (
    KeyWire_0_56,
    n650
  );


  not
  g827
  (
    n827,
    n645
  );


  not
  g828
  (
    n911,
    n782
  );


  not
  g829
  (
    n863,
    n658
  );


  buf
  g830
  (
    n1048,
    n664
  );


  buf
  g831
  (
    n965,
    n751
  );


  buf
  g832
  (
    n1117,
    n739
  );


  buf
  g833
  (
    n969,
    n640
  );


  buf
  g834
  (
    n1124,
    n730
  );


  buf
  g835
  (
    n861,
    n797
  );


  not
  g836
  (
    n1168,
    n796
  );


  buf
  g837
  (
    n878,
    n654
  );


  buf
  g838
  (
    KeyWire_0_36,
    n812
  );


  not
  g839
  (
    n1078,
    n678
  );


  buf
  g840
  (
    n957,
    n806
  );


  buf
  g841
  (
    n1053,
    n808
  );


  not
  g842
  (
    n1042,
    n730
  );


  buf
  g843
  (
    n1068,
    n775
  );


  not
  g844
  (
    n1080,
    n717
  );


  buf
  g845
  (
    n1035,
    n685
  );


  not
  g846
  (
    n1110,
    n683
  );


  buf
  g847
  (
    n1025,
    n793
  );


  not
  g848
  (
    n1137,
    n639
  );


  not
  g849
  (
    n1064,
    n803
  );


  not
  g850
  (
    n981,
    n788
  );


  not
  g851
  (
    n1088,
    n689
  );


  buf
  g852
  (
    n817,
    n735
  );


  not
  g853
  (
    n870,
    n799
  );


  not
  g854
  (
    n1039,
    n642
  );


  buf
  g855
  (
    n995,
    n809
  );


  not
  g856
  (
    KeyWire_0_15,
    n790
  );


  buf
  g857
  (
    n865,
    n723
  );


  buf
  g858
  (
    n1031,
    n793
  );


  not
  g859
  (
    n843,
    n685
  );


  not
  g860
  (
    n1082,
    n714
  );


  buf
  g861
  (
    n906,
    n770
  );


  not
  g862
  (
    n826,
    n729
  );


  buf
  g863
  (
    n979,
    n816
  );


  buf
  g864
  (
    n991,
    n794
  );


  not
  g865
  (
    n1043,
    n790
  );


  not
  g866
  (
    n1138,
    n686
  );


  not
  g867
  (
    n1136,
    n719
  );


  buf
  g868
  (
    n1028,
    n764
  );


  buf
  g869
  (
    n836,
    n747
  );


  buf
  g870
  (
    n925,
    n802
  );


  not
  g871
  (
    n1151,
    n810
  );


  buf
  g872
  (
    n1067,
    n724
  );


  buf
  g873
  (
    n1006,
    n750
  );


  buf
  g874
  (
    n856,
    n763
  );


  not
  g875
  (
    n894,
    n649
  );


  not
  g876
  (
    n1044,
    n745
  );


  buf
  g877
  (
    n875,
    n694
  );


  not
  g878
  (
    n907,
    n804
  );


  not
  g879
  (
    n931,
    n751
  );


  buf
  g880
  (
    n901,
    n681
  );


  not
  g881
  (
    n873,
    n752
  );


  buf
  g882
  (
    n1163,
    n719
  );


  not
  g883
  (
    n958,
    n646
  );


  not
  g884
  (
    n1089,
    n779
  );


  not
  g885
  (
    n1122,
    n713
  );


  not
  g886
  (
    n913,
    n770
  );


  not
  g887
  (
    n909,
    n653
  );


  buf
  g888
  (
    n1125,
    n656
  );


  not
  g889
  (
    n1114,
    n765
  );


  not
  g890
  (
    n908,
    n797
  );


  buf
  g891
  (
    n960,
    n697
  );


  not
  g892
  (
    n927,
    n666
  );


  not
  g893
  (
    n919,
    n764
  );


  buf
  g894
  (
    n1146,
    n815
  );


  not
  g895
  (
    n1020,
    n655
  );


  buf
  g896
  (
    n990,
    n666
  );


  buf
  g897
  (
    n834,
    n630
  );


  buf
  g898
  (
    n1143,
    n755
  );


  buf
  g899
  (
    n917,
    n705
  );


  buf
  g900
  (
    n892,
    n655
  );


  buf
  g901
  (
    n975,
    n628
  );


  not
  g902
  (
    n890,
    n681
  );


  not
  g903
  (
    n986,
    n779
  );


  buf
  g904
  (
    n1133,
    n718
  );


  not
  g905
  (
    n1083,
    n688
  );


  not
  g906
  (
    n1152,
    n804
  );


  buf
  g907
  (
    n882,
    n792
  );


  buf
  g908
  (
    n855,
    n816
  );


  not
  g909
  (
    n842,
    n733
  );


  not
  g910
  (
    n854,
    n637
  );


  not
  g911
  (
    n859,
    n351
  );


  buf
  g912
  (
    n889,
    n703
  );


  not
  g913
  (
    n1169,
    n661
  );


  not
  g914
  (
    n902,
    n736
  );


  buf
  g915
  (
    n887,
    n793
  );


  buf
  g916
  (
    n947,
    n671
  );


  not
  g917
  (
    n845,
    n674
  );


  not
  g918
  (
    n1144,
    n662
  );


  buf
  g919
  (
    n1149,
    n722
  );


  buf
  g920
  (
    n974,
    n692
  );


  buf
  g921
  (
    n1096,
    n756
  );


  buf
  g922
  (
    n1011,
    n691
  );


  buf
  g923
  (
    n1085,
    n750
  );


  not
  g924
  (
    n967,
    n731
  );


  buf
  g925
  (
    n1166,
    n716
  );


  not
  g926
  (
    n1059,
    n790
  );


  buf
  g927
  (
    n938,
    n664
  );


  not
  g928
  (
    n1016,
    n745
  );


  not
  g929
  (
    n953,
    n680
  );


  not
  g930
  (
    n1103,
    n715
  );


  buf
  g931
  (
    n1115,
    n795
  );


  buf
  g932
  (
    n932,
    n755
  );


  buf
  g933
  (
    n983,
    n786
  );


  buf
  g934
  (
    n1099,
    n767
  );


  buf
  g935
  (
    n1056,
    n803
  );


  not
  g936
  (
    n1104,
    n792
  );


  buf
  g937
  (
    n1036,
    n774
  );


  not
  g938
  (
    n837,
    n795
  );


  not
  g939
  (
    n982,
    n703
  );


  not
  g940
  (
    n1112,
    n754
  );


  not
  g941
  (
    n1172,
    n811
  );


  not
  g942
  (
    n1081,
    n630
  );


  buf
  g943
  (
    n1127,
    n768
  );


  not
  g944
  (
    n985,
    n733
  );


  not
  g945
  (
    n853,
    n649
  );


  buf
  g946
  (
    n1065,
    n648
  );


  buf
  g947
  (
    KeyWire_0_38,
    n684
  );


  not
  g948
  (
    n1105,
    n713
  );


  buf
  g949
  (
    n920,
    n798
  );


  buf
  g950
  (
    n858,
    n768
  );


  not
  g951
  (
    n1019,
    n668
  );


  buf
  g952
  (
    n1148,
    n743
  );


  not
  g953
  (
    n1090,
    n676
  );


  buf
  g954
  (
    n914,
    n691
  );


  not
  g955
  (
    n1029,
    n696
  );


  buf
  g956
  (
    n1070,
    n814
  );


  not
  g957
  (
    n1008,
    n737
  );


  buf
  g958
  (
    n954,
    n777
  );


  not
  g959
  (
    n1154,
    n763
  );


  buf
  g960
  (
    n848,
    n617
  );


  buf
  g961
  (
    n897,
    n671
  );


  not
  g962
  (
    n1034,
    n736
  );


  not
  g963
  (
    n891,
    n622
  );


  not
  g964
  (
    n1093,
    n707
  );


  buf
  g965
  (
    n893,
    n811
  );


  buf
  g966
  (
    KeyWire_0_42,
    n747
  );


  buf
  g967
  (
    n1098,
    n647
  );


  not
  g968
  (
    n1041,
    n744
  );


  buf
  g969
  (
    n852,
    n651
  );


  not
  g970
  (
    n903,
    n703
  );


  not
  g971
  (
    n846,
    n797
  );


  buf
  g972
  (
    n1061,
    n794
  );


  not
  g973
  (
    n851,
    n694
  );


  not
  g974
  (
    n963,
    n737
  );


  not
  g975
  (
    n1030,
    n794
  );


  buf
  g976
  (
    n879,
    n784
  );


  not
  g977
  (
    n1057,
    n733
  );


  buf
  g978
  (
    n819,
    n810
  );


  not
  g979
  (
    n899,
    n699
  );


  buf
  g980
  (
    n1076,
    n805
  );


  not
  g981
  (
    n1171,
    n695
  );


  not
  g982
  (
    KeyWire_0_53,
    n788
  );


  buf
  g983
  (
    n835,
    n644
  );


  not
  g984
  (
    n962,
    n669
  );


  not
  g985
  (
    n996,
    n657
  );


  not
  g986
  (
    KeyWire_0_16,
    n688
  );


  not
  g987
  (
    n988,
    n649
  );


  not
  g988
  (
    n1040,
    n748
  );


  buf
  g989
  (
    n1139,
    n686
  );


  not
  g990
  (
    n934,
    n754
  );


  not
  g991
  (
    n1058,
    n670
  );


  buf
  g992
  (
    n833,
    n783
  );


  not
  g993
  (
    n1026,
    n714
  );


  buf
  g994
  (
    n926,
    n663
  );


  not
  g995
  (
    n910,
    n761
  );


  not
  g996
  (
    n921,
    n656
  );


  buf
  g997
  (
    n993,
    n682
  );


  buf
  g998
  (
    n1170,
    n654
  );


  buf
  g999
  (
    n900,
    n628
  );


  not
  g1000
  (
    n940,
    n709
  );


  buf
  g1001
  (
    n1047,
    n757
  );


  nand
  g1002
  (
    n1119,
    n633,
    n654,
    n787,
    n680
  );


  xor
  g1003
  (
    n928,
    n696,
    n734,
    n760,
    n661
  );


  xnor
  g1004
  (
    n912,
    n801,
    n693,
    n762,
    n772
  );


  or
  g1005
  (
    n821,
    n750,
    n669,
    n639,
    n770
  );


  and
  g1006
  (
    n818,
    n781,
    n797,
    n774,
    n696
  );


  xor
  g1007
  (
    n942,
    n789,
    n796,
    n731,
    n721
  );


  nor
  g1008
  (
    n952,
    n692,
    n660,
    n364,
    n678
  );


  nor
  g1009
  (
    n944,
    n637,
    n767,
    n811,
    n659
  );


  nand
  g1010
  (
    n924,
    n666,
    n787,
    n639,
    n775
  );


  or
  g1011
  (
    n822,
    n670,
    n709,
    n722,
    n360
  );


  xnor
  g1012
  (
    n1045,
    n734,
    n656,
    n792,
    n354
  );


  xor
  g1013
  (
    n1017,
    n696,
    n730,
    n644,
    n811
  );


  and
  g1014
  (
    n1049,
    n647,
    n780,
    n721,
    n655
  );


  xnor
  g1015
  (
    n1001,
    n648,
    n798,
    n646,
    n704
  );


  xor
  g1016
  (
    n997,
    n669,
    n682,
    n782,
    n748
  );


  nor
  g1017
  (
    KeyWire_0_48,
    n349,
    n715,
    n648,
    n804
  );


  xor
  g1018
  (
    n966,
    n648,
    n668,
    n688,
    n722
  );


  or
  g1019
  (
    n930,
    n697,
    n725,
    n719,
    n708
  );


  nand
  g1020
  (
    n1052,
    n805,
    n693,
    n712,
    n357
  );


  and
  g1021
  (
    n1077,
    n717,
    n778,
    n692,
    n798
  );


  nor
  g1022
  (
    n918,
    n766,
    n747,
    n728,
    n716
  );


  and
  g1023
  (
    n1074,
    n728,
    n676,
    n699,
    n672
  );


  and
  g1024
  (
    n1003,
    n749,
    n709,
    n725,
    n798
  );


  nor
  g1025
  (
    n824,
    n706,
    n743,
    n739,
    n774
  );


  nor
  g1026
  (
    n1128,
    n684,
    n752,
    n748,
    n712
  );


  nor
  g1027
  (
    n1066,
    n629,
    n682,
    n670,
    n642
  );


  nand
  g1028
  (
    n1012,
    n796,
    n786,
    n631,
    n654
  );


  or
  g1029
  (
    n1097,
    n675,
    n638,
    n781,
    n767
  );


  nor
  g1030
  (
    n987,
    n695,
    n807,
    n638,
    n640
  );


  and
  g1031
  (
    n1005,
    n814,
    n743,
    n638,
    n716
  );


  or
  g1032
  (
    n968,
    n755,
    n641,
    n642,
    n715
  );


  nor
  g1033
  (
    n886,
    n634,
    n749,
    n361,
    n713
  );


  nand
  g1034
  (
    n1027,
    n665,
    n750,
    n663,
    n766
  );


  nand
  g1035
  (
    n959,
    n674,
    n632,
    n743,
    n718
  );


  and
  g1036
  (
    n830,
    n641,
    n757,
    n684,
    n628
  );


  xnor
  g1037
  (
    n964,
    n774,
    n753,
    n808,
    n684
  );


  nor
  g1038
  (
    n955,
    n792,
    n812,
    n742,
    n771
  );


  xnor
  g1039
  (
    n828,
    n629,
    n725,
    n791,
    n783
  );


  nand
  g1040
  (
    n820,
    n751,
    n765,
    n675,
    n737
  );


  xnor
  g1041
  (
    n869,
    n745,
    n712,
    n627,
    n731
  );


  and
  g1042
  (
    n850,
    n668,
    n796,
    n665,
    n746
  );


  and
  g1043
  (
    n973,
    n704,
    n761,
    n779,
    n672
  );


  or
  g1044
  (
    n1158,
    n703,
    n809,
    n739,
    n744
  );


  xnor
  g1045
  (
    n874,
    n715,
    n763,
    n662,
    n780
  );


  nand
  g1046
  (
    n1094,
    n643,
    n806,
    n780,
    n726
  );


  nand
  g1047
  (
    n972,
    n769,
    n711,
    n681,
    n666
  );


  xor
  g1048
  (
    n971,
    n730,
    n636,
    n689,
    n738
  );


  xor
  g1049
  (
    n1073,
    n707,
    n352,
    n717,
    n619
  );


  or
  g1050
  (
    n1167,
    n801,
    n732,
    n710,
    n740
  );


  nor
  g1051
  (
    n857,
    n700,
    n685,
    n778,
    n785
  );


  nor
  g1052
  (
    n1132,
    n672,
    n711,
    n800,
    n657
  );


  nand
  g1053
  (
    n976,
    n636,
    n627,
    n753,
    n754
  );


  or
  g1054
  (
    n1022,
    n679,
    n356,
    n769,
    n710
  );


  and
  g1055
  (
    n1118,
    n783,
    n772,
    n778,
    n660
  );


  nor
  g1056
  (
    n1162,
    n658,
    n816,
    n624,
    n664
  );


  nand
  g1057
  (
    n885,
    n765,
    n642,
    n769,
    n620
  );


  and
  g1058
  (
    n847,
    n630,
    n688,
    n772,
    n653
  );


  xor
  g1059
  (
    n1150,
    n626,
    n674,
    n732,
    n676
  );


  and
  g1060
  (
    n1014,
    n754,
    n784,
    n651,
    n671
  );


  nor
  g1061
  (
    n1092,
    n815,
    n744,
    n738,
    n745
  );


  and
  g1062
  (
    n989,
    n362,
    n744,
    n717,
    n801
  );


  and
  g1063
  (
    KeyWire_0_31,
    n789,
    n711,
    n746,
    n706
  );


  and
  g1064
  (
    n1004,
    n700,
    n705,
    n782,
    n718
  );


  and
  g1065
  (
    n1024,
    n752,
    n749,
    n651,
    n673
  );


  xnor
  g1066
  (
    n1009,
    n667,
    n775,
    n724,
    n762
  );


  xnor
  g1067
  (
    n877,
    n659,
    n640,
    n813,
    n637
  );


  or
  g1068
  (
    n1155,
    n813,
    n698,
    n707,
    n786
  );


  xor
  g1069
  (
    n868,
    n720,
    n624,
    n813,
    n697
  );


  or
  g1070
  (
    n936,
    n660,
    n777,
    n806,
    n625
  );


  or
  g1071
  (
    n994,
    n740,
    n629,
    n726,
    n793
  );


  nor
  g1072
  (
    n977,
    n677,
    n810,
    n766,
    n679
  );


  and
  g1073
  (
    n961,
    n726,
    n727,
    n771,
    n758
  );


  nand
  g1074
  (
    n980,
    n698,
    n634,
    n695,
    n770
  );


  nor
  g1075
  (
    n1054,
    n803,
    n678,
    n732,
    n767
  );


  xnor
  g1076
  (
    n838,
    n640,
    n800,
    n700
  );


  nor
  g1077
  (
    n949,
    n749,
    n759,
    n635
  );


  and
  g1078
  (
    n1165,
    n674,
    n724,
    n657,
    n644
  );


  xor
  g1079
  (
    n1126,
    n671,
    n759,
    n773,
    n736
  );


  nor
  g1080
  (
    n916,
    n776,
    n633,
    n742,
    n701
  );


  nor
  g1081
  (
    n1021,
    n773,
    n809,
    n687,
    n784
  );


  or
  g1082
  (
    n1091,
    n635,
    n768,
    n658,
    n800
  );


  xnor
  g1083
  (
    KeyWire_0_21,
    n704,
    n665,
    n788,
    n669
  );


  nor
  g1084
  (
    n1051,
    n761,
    n804,
    n662,
    n659
  );


  nor
  g1085
  (
    n1129,
    n718,
    n729,
    n690,
    n665
  );


  xnor
  g1086
  (
    n1050,
    n734,
    n704,
    n649,
    n791
  );


  nand
  g1087
  (
    n1159,
    n692,
    n701,
    n740,
    n813
  );


  nand
  g1088
  (
    n1157,
    n773,
    n721,
    n739,
    n787
  );


  xnor
  g1089
  (
    n839,
    n714,
    n728,
    n779,
    n756
  );


  xor
  g1090
  (
    n1087,
    n650,
    n653,
    n771,
    n673
  );


  nor
  g1091
  (
    n1147,
    n709,
    n723,
    n714,
    n753
  );


  and
  g1092
  (
    n956,
    n651,
    n794,
    n636,
    n652
  );


  or
  g1093
  (
    n1071,
    n689,
    n748,
    n355,
    n643
  );


  nor
  g1094
  (
    n823,
    n756,
    n708,
    n764,
    n702
  );


  xnor
  g1095
  (
    n1135,
    n683,
    n780,
    n645,
    n686
  );


  nor
  g1096
  (
    n860,
    n661,
    n816,
    n784,
    n752
  );


  or
  g1097
  (
    n896,
    n728,
    n720,
    n687,
    n760
  );


  or
  g1098
  (
    n1113,
    n809,
    n675,
    n656,
    n716
  );


  nor
  g1099
  (
    n1102,
    n634,
    n777,
    n667,
    n753
  );


  nand
  g1100
  (
    n1037,
    n741,
    n762,
    n623,
    n740
  );


  or
  g1101
  (
    n943,
    n782,
    n713,
    n802,
    n734
  );


  xor
  g1102
  (
    n946,
    n727,
    n636,
    n707,
    n677
  );


  nand
  g1103
  (
    n840,
    n359,
    n678,
    n781,
    n812
  );


  and
  g1104
  (
    n1131,
    n758,
    n668,
    n621,
    n736
  );


  and
  g1105
  (
    n950,
    n677,
    n647,
    n758,
    n637
  );


  nand
  g1106
  (
    n1075,
    n732,
    n663,
    n775,
    n785
  );


  nand
  g1107
  (
    n1145,
    n679,
    n787,
    n738,
    n801
  );


  or
  g1108
  (
    n1002,
    n737,
    n690,
    n757,
    n742
  );


  xnor
  g1109
  (
    n1095,
    n706,
    n653,
    n677,
    n663
  );


  and
  g1110
  (
    n1140,
    n720,
    n723,
    n694,
    n699
  );


  or
  g1111
  (
    n1023,
    n756,
    n785,
    n633,
    n710
  );


  and
  g1112
  (
    n1141,
    n776,
    n667,
    n682,
    n686
  );


  xnor
  g1113
  (
    n1079,
    n363,
    n710,
    n766,
    n789
  );


  xor
  g1114
  (
    n1018,
    n701,
    n776,
    n799,
    n781
  );


  xor
  g1115
  (
    n1033,
    n746,
    n685,
    n741,
    n795
  );


  and
  g1116
  (
    n1060,
    n708,
    n760,
    n627,
    n631
  );


  xnor
  g1117
  (
    n1116,
    n805,
    n643,
    n764,
    n652
  );


  nand
  g1118
  (
    n905,
    n723,
    n778,
    n658,
    n719
  );


  xor
  g1119
  (
    n941,
    n690,
    n741,
    n765,
    n657
  );


  or
  g1120
  (
    n1153,
    n762,
    n768,
    n673,
    n350
  );


  xnor
  g1121
  (
    n1121,
    n706,
    n805,
    n650,
    n799
  );


  nor
  g1122
  (
    n1142,
    n814,
    n738,
    n755,
    n687
  );


  xor
  g1123
  (
    n1015,
    n812,
    n769,
    n626,
    n786
  );


  xor
  g1124
  (
    n844,
    n724,
    n772,
    n691,
    n698
  );


  xor
  g1125
  (
    n825,
    n676,
    n680,
    n747,
    n806
  );


  xor
  g1126
  (
    n831,
    n712,
    n662,
    n641,
    n694
  );


  or
  g1127
  (
    n929,
    n726,
    n625,
    n785,
    n661
  );


  nand
  g1128
  (
    n871,
    n646,
    n720,
    n802,
    n679
  );


  and
  g1129
  (
    n904,
    n771,
    n650,
    n697,
    n729
  );


  nor
  g1130
  (
    n872,
    n683,
    n810,
    n632,
    n655
  );


  nor
  g1131
  (
    n1010,
    n700,
    n731,
    n791,
    n758
  );


  and
  g1132
  (
    n898,
    n789,
    n815,
    n795,
    n647
  );


  nand
  g1133
  (
    n992,
    n652,
    n708,
    n808,
    n644
  );


  xnor
  g1134
  (
    n915,
    n799,
    n646,
    n632,
    n777
  );


  nor
  g1135
  (
    n1038,
    n760,
    n645,
    n358,
    n776
  );


  nor
  g1136
  (
    n1160,
    n664,
    n698,
    n652,
    n687
  );


  and
  g1137
  (
    n1156,
    n673,
    n702,
    n735
  );


  nand
  g1138
  (
    n922,
    n690,
    n815,
    n618,
    n788
  );


  nor
  g1139
  (
    n1084,
    n807,
    n622,
    n705,
    n626
  );


  xnor
  g1140
  (
    n1055,
    n625,
    n645,
    n691,
    n759
  );


  xnor
  g1141
  (
    n1032,
    n672,
    n693,
    n722,
    n725
  );


  xor
  g1142
  (
    n1072,
    n680,
    n635,
    n705,
    n761
  );


  and
  g1143
  (
    n1108,
    n670,
    n683,
    n773,
    n742
  );


  nor
  g1144
  (
    n948,
    n667,
    n783,
    n757,
    n735
  );


  nand
  g1145
  (
    n951,
    n727,
    n681,
    n659,
    n353
  );


  not
  g1146
  (
    n1187,
    n817
  );


  buf
  g1147
  (
    n1179,
    n828
  );


  not
  g1148
  (
    n1176,
    n832
  );


  not
  g1149
  (
    n1183,
    n829
  );


  buf
  g1150
  (
    n1178,
    n826
  );


  buf
  g1151
  (
    n1182,
    n830
  );


  not
  g1152
  (
    n1177,
    n822
  );


  not
  g1153
  (
    n1173,
    n831
  );


  not
  g1154
  (
    n1185,
    n818
  );


  not
  g1155
  (
    n1174,
    n823
  );


  not
  g1156
  (
    n1186,
    n825
  );


  not
  g1157
  (
    n1181,
    n819
  );


  buf
  g1158
  (
    n1188,
    n820
  );


  buf
  g1159
  (
    n1180,
    n827
  );


  not
  g1160
  (
    n1184,
    n824
  );


  not
  g1161
  (
    n1175,
    n821
  );


  xnor
  g1162
  (
    n1189,
    n1178,
    n1177,
    n1174,
    n1179
  );


  xnor
  g1163
  (
    n1190,
    n833,
    n1176,
    n1173,
    n1175
  );


  buf
  g1164
  (
    n1191,
    n1190
  );


  not
  g1165
  (
    n1192,
    n1180
  );


  xor
  g1166
  (
    n1193,
    n1190,
    n1189
  );


  not
  g1167
  (
    n1200,
    n846
  );


  not
  g1168
  (
    n1195,
    n1191
  );


  nor
  g1169
  (
    n1202,
    n371,
    n1193
  );


  or
  g1170
  (
    n1201,
    n839,
    n367,
    n844,
    n847
  );


  xnor
  g1171
  (
    n1198,
    n838,
    n1192,
    n850
  );


  nor
  g1172
  (
    n1197,
    n1191,
    n372,
    n1193,
    n840
  );


  or
  g1173
  (
    n1199,
    n1181,
    n852,
    n843,
    n834
  );


  or
  g1174
  (
    n1203,
    n1191,
    n368,
    n849,
    n365
  );


  nor
  g1175
  (
    n1204,
    n845,
    n841,
    n837,
    n851
  );


  xor
  g1176
  (
    n1196,
    n1191,
    n848,
    n836,
    n366
  );


  xnor
  g1177
  (
    n1194,
    n1192,
    n370,
    n842,
    n1193
  );


  xnor
  g1178
  (
    n1205,
    n835,
    n1192,
    n369,
    n1193
  );


  nand
  g1179
  (
    n1238,
    n413,
    n452,
    n436,
    n458
  );


  or
  g1180
  (
    n1207,
    n394,
    n1199,
    n462,
    n473
  );


  xnor
  g1181
  (
    n1214,
    n423,
    n446,
    n1203,
    n380
  );


  xnor
  g1182
  (
    n1228,
    n442,
    n1205,
    n414,
    n392
  );


  xor
  g1183
  (
    n1225,
    n1204,
    n476,
    n454,
    n417
  );


  nand
  g1184
  (
    n1222,
    n374,
    n467,
    n1195,
    n404
  );


  xnor
  g1185
  (
    n1218,
    n441,
    n477,
    n464,
    n1198
  );


  and
  g1186
  (
    n1209,
    n449,
    n408,
    n470,
    n438
  );


  xor
  g1187
  (
    n1206,
    n450,
    n475,
    n424,
    n466
  );


  or
  g1188
  (
    n1239,
    n384,
    n402,
    n1202,
    n1204
  );


  nand
  g1189
  (
    n1236,
    n1201,
    n1200,
    n463,
    n397
  );


  and
  g1190
  (
    n1230,
    n1197,
    n431,
    n382,
    n399
  );


  xor
  g1191
  (
    n1220,
    n1199,
    n412,
    n383,
    n474
  );


  xor
  g1192
  (
    n1229,
    n439,
    n444,
    n409,
    n1204
  );


  and
  g1193
  (
    n1221,
    n451,
    n426,
    n447,
    n1203
  );


  xnor
  g1194
  (
    n1232,
    n387,
    n403,
    n1203,
    n448
  );


  and
  g1195
  (
    n1235,
    n386,
    n1202,
    n1200,
    n440
  );


  xor
  g1196
  (
    n1219,
    n1198,
    n427,
    n395,
    n1196
  );


  nand
  g1197
  (
    n1240,
    n381,
    n1197,
    n419,
    n1201
  );


  xnor
  g1198
  (
    n1210,
    n422,
    n469,
    n472,
    n391
  );


  and
  g1199
  (
    n1226,
    n1194,
    n420,
    n407,
    n456
  );


  or
  g1200
  (
    n1213,
    n421,
    n375,
    n400,
    n1205
  );


  nand
  g1201
  (
    n1223,
    n429,
    n418,
    n411,
    n459
  );


  xor
  g1202
  (
    n1208,
    n455,
    n457,
    n432,
    n388
  );


  nand
  g1203
  (
    n1212,
    n435,
    n1205,
    n1201,
    n377
  );


  and
  g1204
  (
    n1233,
    n1200,
    n1196,
    n471,
    n1204
  );


  nor
  g1205
  (
    n1211,
    n390,
    n430,
    n1205,
    n406
  );


  and
  g1206
  (
    n1231,
    n389,
    n1203,
    n443,
    n428
  );


  or
  g1207
  (
    n1215,
    n385,
    n468,
    n1195,
    n410
  );


  and
  g1208
  (
    n1224,
    n378,
    n437,
    n434,
    n396
  );


  and
  g1209
  (
    n1227,
    n379,
    n433,
    n398,
    n465
  );


  or
  g1210
  (
    n1216,
    n416,
    n1202,
    n376,
    n425
  );


  nand
  g1211
  (
    n1217,
    n393,
    n415,
    n1201,
    n461
  );


  nor
  g1212
  (
    n1234,
    n373,
    n453,
    n1202,
    n1200
  );


  xor
  g1213
  (
    n1237,
    n401,
    n460,
    n445,
    n405
  );


  xnor
  g1214
  (
    n1247,
    n1206,
    n1233,
    n1229,
    n1219
  );


  nor
  g1215
  (
    n1241,
    n1218,
    n1212,
    n1234,
    n1223
  );


  nand
  g1216
  (
    n1242,
    n1234,
    n1210,
    n1232,
    n1228
  );


  and
  g1217
  (
    n1245,
    n1214,
    n1230,
    n1225,
    n1227
  );


  xor
  g1218
  (
    n1250,
    n1229,
    n1231,
    n1208
  );


  nor
  g1219
  (
    n1246,
    n1220,
    n1232,
    n1221,
    n1217
  );


  xnor
  g1220
  (
    n1249,
    n1216,
    n1213,
    n1230,
    n1224
  );


  xor
  g1221
  (
    n1243,
    n1235,
    n1211,
    n1215,
    n1228
  );


  xor
  g1222
  (
    n1248,
    n1226,
    n1222,
    n1227,
    n1209
  );


  xnor
  g1223
  (
    n1244,
    n1226,
    n1233,
    n1235,
    n1207
  );


  buf
  g1224
  (
    n1254,
    n854
  );


  not
  g1225
  (
    n1253,
    n1244
  );


  buf
  g1226
  (
    n1257,
    n1250
  );


  buf
  g1227
  (
    n1255,
    n860
  );


  not
  g1228
  (
    n1259,
    n1246
  );


  buf
  g1229
  (
    n1256,
    n1243
  );


  or
  g1230
  (
    n1251,
    n856,
    n1242,
    n1249,
    n1245
  );


  or
  g1231
  (
    n1258,
    n853,
    n858,
    n859,
    n857
  );


  xnor
  g1232
  (
    n1252,
    n1248,
    n861,
    n855,
    n1247
  );


  buf
  g1233
  (
    n1260,
    n1251
  );


  buf
  g1234
  (
    n1261,
    n1251
  );


  buf
  g1235
  (
    n1263,
    n1252
  );


  buf
  g1236
  (
    n1262,
    n1251
  );


  nand
  g1237
  (
    n1270,
    n1252,
    n870,
    n1260,
    n865
  );


  and
  g1238
  (
    n1265,
    n1253,
    n1253,
    n863,
    n1261
  );


  xnor
  g1239
  (
    n1268,
    n864,
    n478,
    n1254,
    n873
  );


  xor
  g1240
  (
    n1266,
    n866,
    n868,
    n871,
    n1252
  );


  nor
  g1241
  (
    n1264,
    n867,
    n1261,
    n1263,
    n1262
  );


  nand
  g1242
  (
    n1269,
    n1253,
    n1253,
    n1252,
    n869
  );


  nor
  g1243
  (
    n1267,
    n1262,
    n872,
    n1263,
    n862
  );


  buf
  g1244
  (
    n1274,
    n1265
  );


  not
  g1245
  (
    n1273,
    n1264
  );


  buf
  g1246
  (
    n1272,
    n1265
  );


  buf
  g1247
  (
    n1271,
    n1264
  );


  buf
  g1248
  (
    n1277,
    n880
  );


  not
  g1249
  (
    n1276,
    n877
  );


  buf
  g1250
  (
    n1278,
    n1273
  );


  not
  g1251
  (
    n1282,
    n1272
  );


  buf
  g1252
  (
    n1280,
    n1274
  );


  or
  g1253
  (
    n1281,
    n879,
    n878,
    n1274
  );


  xnor
  g1254
  (
    n1275,
    n876,
    n874,
    n881,
    n1272
  );


  xor
  g1255
  (
    n1279,
    n1273,
    n1271,
    n875
  );


  nor
  g1256
  (
    n1296,
    n506,
    n487,
    n502,
    n481
  );


  nand
  g1257
  (
    n1283,
    n505,
    n1237,
    n508,
    n884
  );


  xnor
  g1258
  (
    n1289,
    n888,
    n1282,
    n482,
    n890
  );


  or
  g1259
  (
    n1288,
    n490,
    n483,
    n1182,
    n495
  );


  xnor
  g1260
  (
    n1295,
    n503,
    n491,
    n498,
    n497
  );


  nor
  g1261
  (
    n1300,
    n882,
    n1276,
    n1184,
    n1282
  );


  and
  g1262
  (
    n1287,
    n1282,
    n496,
    n1281
  );


  nand
  g1263
  (
    n1285,
    n1188,
    n504,
    n886,
    n480
  );


  xor
  g1264
  (
    n1292,
    n509,
    n510,
    n1278,
    n494
  );


  or
  g1265
  (
    KeyWire_0_37,
    n885,
    n484,
    n1277,
    n501
  );


  and
  g1266
  (
    n1293,
    n1279,
    n889,
    n1275,
    n1237
  );


  nand
  g1267
  (
    n1298,
    n887,
    n489,
    n1276,
    n492
  );


  nand
  g1268
  (
    n1284,
    n1183,
    n1275,
    n486,
    n500
  );


  xor
  g1269
  (
    n1297,
    n485,
    n883,
    n479,
    n1278
  );


  xor
  g1270
  (
    n1290,
    n1187,
    n1279,
    n507,
    n1277
  );


  and
  g1271
  (
    n1299,
    n488,
    n1281,
    n499,
    n1186
  );


  and
  g1272
  (
    n1286,
    n1280,
    n511,
    n493,
    n1236
  );


  or
  g1273
  (
    KeyWire_0_14,
    n1280,
    n1280,
    n1185,
    n1236
  );


  nand
  g1274
  (
    n1310,
    n894,
    n534,
    n517,
    n515
  );


  xor
  g1275
  (
    n1307,
    n1291,
    n1283,
    n1284,
    n891
  );


  or
  g1276
  (
    n1308,
    n535,
    n536,
    n520,
    n530
  );


  xnor
  g1277
  (
    n1311,
    n519,
    n533,
    n526,
    n1256
  );


  nand
  g1278
  (
    n1306,
    n537,
    n1255,
    n516,
    n1292
  );


  nand
  g1279
  (
    n1316,
    n1296,
    n1255,
    n529,
    n1300
  );


  and
  g1280
  (
    n1301,
    n538,
    n521,
    n892,
    n1299
  );


  or
  g1281
  (
    n1305,
    n895,
    n522,
    n527,
    n1294
  );


  and
  g1282
  (
    n1315,
    n1256,
    n1290,
    n1255,
    n1254
  );


  xnor
  g1283
  (
    n1304,
    n524,
    n525,
    n1254,
    n1298
  );


  or
  g1284
  (
    n1303,
    n1286,
    n1287,
    n539,
    n528
  );


  nand
  g1285
  (
    n1309,
    n1256,
    n1285,
    n1288,
    n513
  );


  nand
  g1286
  (
    n1313,
    n1295,
    n531,
    n532,
    n523
  );


  nor
  g1287
  (
    n1302,
    n1254,
    n897,
    n514,
    n1289
  );


  xnor
  g1288
  (
    n1314,
    n518,
    n896,
    n512,
    n898
  );


  xnor
  g1289
  (
    n1312,
    n1297,
    n893,
    n1293,
    n1255
  );


  buf
  g1290
  (
    n1317,
    n1313
  );


  not
  g1291
  (
    n1319,
    n900
  );


  buf
  g1292
  (
    n1323,
    n903
  );


  not
  g1293
  (
    n1320,
    n901
  );


  not
  g1294
  (
    KeyWire_0_12,
    n1309
  );


  xnor
  g1295
  (
    n1324,
    n1310,
    n906,
    n905
  );


  nand
  g1296
  (
    n1318,
    n1316,
    n904,
    n1314,
    n899
  );


  or
  g1297
  (
    n1321,
    n1311,
    n1312,
    n902,
    n1315
  );


  not
  g1298
  (
    n1326,
    n1319
  );


  buf
  g1299
  (
    n1327,
    n1318
  );


  buf
  g1300
  (
    n1333,
    n1318
  );


  buf
  g1301
  (
    n1329,
    n1320
  );


  buf
  g1302
  (
    n1330,
    n1319
  );


  buf
  g1303
  (
    n1335,
    n1317
  );


  buf
  g1304
  (
    n1331,
    n1320
  );


  not
  g1305
  (
    n1332,
    n1320
  );


  not
  g1306
  (
    n1325,
    n1317
  );


  xor
  g1307
  (
    n1328,
    n1320,
    n1318,
    n1319
  );


  nor
  g1308
  (
    n1334,
    n1318,
    n1317,
    n1319
  );


  xor
  g1309
  (
    n1344,
    n1332,
    n949,
    n944,
    n918
  );


  or
  g1310
  (
    n1342,
    n917,
    n914,
    n921,
    n1327
  );


  nor
  g1311
  (
    n1348,
    n1335,
    n1334,
    n951,
    n942
  );


  nor
  g1312
  (
    n1338,
    n919,
    n1326,
    n911,
    n945
  );


  xor
  g1313
  (
    n1351,
    n912,
    n952,
    n933,
    n943
  );


  nand
  g1314
  (
    n1350,
    n1331,
    n910,
    n927,
    n1334
  );


  xor
  g1315
  (
    n1336,
    n950,
    n940,
    n928,
    n931
  );


  xor
  g1316
  (
    n1340,
    n926,
    n1328,
    n908,
    n953
  );


  and
  g1317
  (
    n1343,
    n924,
    n920,
    n938,
    n909
  );


  nor
  g1318
  (
    n1349,
    n1325,
    n941,
    n1335,
    n937
  );


  nor
  g1319
  (
    n1337,
    n916,
    n1335,
    n925,
    n1330
  );


  xnor
  g1320
  (
    n1339,
    n932,
    n934,
    n1329,
    n929
  );


  xnor
  g1321
  (
    n1346,
    n913,
    n939,
    n923,
    n1333
  );


  or
  g1322
  (
    n1341,
    n947,
    n948,
    n954,
    n946
  );


  xnor
  g1323
  (
    n1347,
    n936,
    n915,
    n930,
    n1335
  );


  xor
  g1324
  (
    n1345,
    n907,
    n1334,
    n935,
    n922
  );


  or
  g1325
  (
    n1354,
    n970,
    n987,
    n964,
    n1348
  );


  xor
  g1326
  (
    n1364,
    n1347,
    n1344,
    n961,
    n963
  );


  nand
  g1327
  (
    n1369,
    n991,
    n1347,
    n997,
    n990
  );


  xnor
  g1328
  (
    n1355,
    n1343,
    n1336,
    n1346,
    n979
  );


  nor
  g1329
  (
    n1368,
    n992,
    n1345,
    n1337,
    n1341
  );


  or
  g1330
  (
    n1366,
    n966,
    n975,
    n1344,
    n962
  );


  xor
  g1331
  (
    n1353,
    n960,
    n984,
    n1346,
    n1343
  );


  or
  g1332
  (
    n1367,
    n973,
    n1346,
    n1343,
    n996
  );


  xnor
  g1333
  (
    n1359,
    n980,
    n968,
    n1338,
    n981
  );


  nand
  g1334
  (
    n1363,
    n985,
    n994,
    n974,
    n965
  );


  nand
  g1335
  (
    n1362,
    n1342,
    n959,
    n1340,
    n1345
  );


  xor
  g1336
  (
    n1361,
    n1344,
    n969,
    n978,
    n982
  );


  nor
  g1337
  (
    n1360,
    n1341,
    n956,
    n998,
    n1342
  );


  or
  g1338
  (
    n1358,
    n971,
    n989,
    n957,
    n1336
  );


  and
  g1339
  (
    n1352,
    n993,
    n1345,
    n976,
    n986
  );


  xor
  g1340
  (
    n1357,
    n972,
    n1348,
    n1337,
    n983
  );


  xor
  g1341
  (
    n1370,
    n955,
    n1339,
    n1338,
    n988
  );


  nand
  g1342
  (
    n1365,
    n958,
    n1340,
    n995,
    n1342
  );


  xor
  g1343
  (
    n1356,
    n1339,
    n967,
    n1347,
    n977
  );


  or
  g1344
  (
    n1371,
    n1004,
    n1002,
    n1020,
    n1018
  );


  xnor
  g1345
  (
    n1374,
    n1013,
    n1367,
    n1000,
    n1369
  );


  xor
  g1346
  (
    n1373,
    n1019,
    n1001,
    n1007,
    n1024
  );


  nor
  g1347
  (
    n1376,
    n1022,
    n1005,
    n1009,
    n1015
  );


  or
  g1348
  (
    n1375,
    n1014,
    n1366,
    n1370,
    n999
  );


  and
  g1349
  (
    n1378,
    n1025,
    n1016,
    n1012,
    n1368
  );


  nor
  g1350
  (
    KeyWire_0_55,
    n1362,
    n1023,
    n1011,
    n1003
  );


  nor
  g1351
  (
    n1379,
    n1008,
    n1006,
    n1017,
    n1010
  );


  and
  g1352
  (
    n1377,
    n1021,
    n1365,
    n1363,
    n1364
  );


  xor
  g1353
  (
    n1396,
    n1053,
    n1068,
    n1103,
    n545
  );


  or
  g1354
  (
    n1384,
    n1076,
    n1376,
    n1106,
    n1099
  );


  nand
  g1355
  (
    n1407,
    n1039,
    n1052,
    n1051,
    n1377
  );


  xnor
  g1356
  (
    n1403,
    n1082,
    n1038,
    n1373,
    n1379
  );


  xor
  g1357
  (
    n1398,
    n1375,
    n1372,
    n1058,
    n1121
  );


  xnor
  g1358
  (
    n1409,
    n1120,
    n1060,
    n1266,
    n1037
  );


  and
  g1359
  (
    n1386,
    n1054,
    n1044,
    n1375,
    n541
  );


  xnor
  g1360
  (
    n1395,
    n1100,
    n1371,
    n1108,
    n1116
  );


  or
  g1361
  (
    n1402,
    n1034,
    n543,
    n1036,
    n1029
  );


  nand
  g1362
  (
    n1388,
    n1073,
    n1374,
    n1069
  );


  nor
  g1363
  (
    n1408,
    n1096,
    n1372,
    n1041,
    n1378
  );


  nand
  g1364
  (
    n1412,
    n1375,
    n1055,
    n1118,
    n544
  );


  nor
  g1365
  (
    n1414,
    n1374,
    n1373,
    n1045,
    n1091
  );


  nand
  g1366
  (
    n1411,
    n1088,
    n1090,
    n1085,
    n1061
  );


  xnor
  g1367
  (
    n1400,
    n1372,
    n546,
    n1105,
    n1028
  );


  and
  g1368
  (
    n1410,
    n1084,
    n1075,
    n1070,
    n1378
  );


  or
  g1369
  (
    n1392,
    n542,
    n1114,
    n1374,
    n1040
  );


  nand
  g1370
  (
    n1380,
    n1077,
    n1094,
    n1074,
    n1062
  );


  xor
  g1371
  (
    n1391,
    n1050,
    n1373,
    n1372,
    n1072
  );


  xnor
  g1372
  (
    n1393,
    n1035,
    n1092,
    n1379,
    n1048
  );


  or
  g1373
  (
    n1413,
    n1046,
    n1102,
    n1087,
    n1376
  );


  or
  g1374
  (
    n1389,
    n1371,
    n540,
    n1111,
    n1375
  );


  xnor
  g1375
  (
    n1387,
    n1049,
    n1078,
    n1379,
    n1080
  );


  or
  g1376
  (
    n1405,
    n1026,
    n1110,
    n1115,
    n1030
  );


  nor
  g1377
  (
    n1397,
    n1378,
    n1047,
    n1064,
    n1377
  );


  or
  g1378
  (
    n1394,
    n1081,
    n1376,
    n1043,
    n1104
  );


  nor
  g1379
  (
    n1390,
    n1378,
    n1071,
    n1033,
    n1095
  );


  nor
  g1380
  (
    n1401,
    n1379,
    n1032,
    n1119,
    n1059
  );


  xor
  g1381
  (
    n1381,
    n1113,
    n1373,
    n1098,
    n1086
  );


  xnor
  g1382
  (
    n1406,
    n1027,
    n1097,
    n1067,
    n1109
  );


  nand
  g1383
  (
    n1399,
    n1063,
    n1089,
    n1056,
    n1065
  );


  nand
  g1384
  (
    n1383,
    n1101,
    n1107,
    n1079,
    n1117
  );


  xor
  g1385
  (
    n1385,
    n1112,
    n1266,
    n1376,
    n1031
  );


  nor
  g1386
  (
    n1382,
    n1093,
    n1377,
    n1042,
    n1066
  );


  or
  g1387
  (
    n1404,
    n1377,
    n1057,
    n1371,
    n1083
  );


  xor
  g1388
  (
    n1418,
    n1411,
    n1413,
    n1387,
    n1400
  );


  or
  g1389
  (
    n1419,
    n1383,
    n1409,
    n1391,
    n1408
  );


  nand
  g1390
  (
    n1426,
    n1406,
    n1397,
    n1268,
    n1414
  );


  and
  g1391
  (
    n1427,
    n1380,
    n1122,
    n1399,
    n1269
  );


  or
  g1392
  (
    n1424,
    n1410,
    n1395,
    n1381,
    n1398
  );


  and
  g1393
  (
    n1422,
    n1268,
    n1396,
    n1125,
    n1128
  );


  nand
  g1394
  (
    KeyWire_0_61,
    n1126,
    n1267,
    n1384
  );


  nor
  g1395
  (
    n1417,
    n1393,
    n1270,
    n1124,
    n1403
  );


  or
  g1396
  (
    n1420,
    n1412,
    n1269,
    n1385,
    n1386
  );


  nor
  g1397
  (
    n1415,
    n1129,
    n1392,
    n1390,
    n1402
  );


  nand
  g1398
  (
    KeyWire_0_43,
    n1401,
    n1270,
    n1394,
    n1127
  );


  nor
  g1399
  (
    n1416,
    n1270,
    n1407,
    n1388,
    n1382
  );


  xor
  g1400
  (
    n1425,
    n1389,
    n1404,
    n1405,
    n1123
  );


  nand
  g1401
  (
    n1434,
    n1150,
    n1424,
    n1132,
    n1418
  );


  nand
  g1402
  (
    n1440,
    n1142,
    n1133,
    n1151,
    n1427
  );


  nand
  g1403
  (
    n1439,
    n1168,
    n1165,
    n1426,
    n1140
  );


  nor
  g1404
  (
    n1436,
    n1167,
    n1131,
    n1154,
    n1415
  );


  and
  g1405
  (
    n1435,
    n1157,
    n1161,
    n1158,
    n1425
  );


  or
  g1406
  (
    n1441,
    n1416,
    n1171,
    n1419,
    n1135
  );


  and
  g1407
  (
    n1437,
    n1170,
    n1417,
    n1420,
    n1166
  );


  xor
  g1408
  (
    n1431,
    n1160,
    n1145,
    n1134,
    n1169
  );


  xor
  g1409
  (
    n1432,
    n1423,
    n1144,
    n1427,
    n1159
  );


  xnor
  g1410
  (
    n1428,
    n1422,
    n1152,
    n1141,
    n1421
  );


  xor
  g1411
  (
    n1433,
    n1137,
    n1162,
    n1163,
    n1139
  );


  or
  g1412
  (
    KeyWire_0_62,
    n1136,
    n1138,
    n1147,
    n1146
  );


  and
  g1413
  (
    n1430,
    n1156,
    n1155,
    n1164,
    n1148
  );


  and
  g1414
  (
    n1438,
    n1153,
    n1149,
    n1130,
    n1143
  );


  nand
  g1415
  (
    n1449,
    n1239,
    n1257,
    n1322
  );


  nand
  g1416
  (
    n1454,
    n1350,
    n1323,
    n1349,
    n1429
  );


  or
  g1417
  (
    n1446,
    n1438,
    n1322,
    n1351,
    n1324
  );


  xnor
  g1418
  (
    n1443,
    n1433,
    n1349,
    n1322,
    n1441
  );


  nor
  g1419
  (
    n1445,
    n1257,
    n1240,
    n1258,
    n1440
  );


  nor
  g1420
  (
    n1447,
    n1351,
    n1323,
    n1348,
    n1259
  );


  nand
  g1421
  (
    n1455,
    n1239,
    n1259,
    n1321,
    n1350
  );


  and
  g1422
  (
    n1451,
    n1321,
    n1258,
    n1257
  );


  xor
  g1423
  (
    n1456,
    n1350,
    n1435,
    n1259,
    n1172
  );


  nand
  g1424
  (
    n1448,
    n1436,
    n1434,
    n1321
  );


  or
  g1425
  (
    n1457,
    n1238,
    n1324,
    n1240
  );


  nand
  g1426
  (
    n1442,
    n1259,
    n1323,
    n1258,
    n1441
  );


  nand
  g1427
  (
    n1444,
    n1431,
    n1437,
    n1351,
    n1349
  );


  or
  g1428
  (
    n1452,
    n1256,
    n1432,
    n1240,
    n1323
  );


  or
  g1429
  (
    n1450,
    n1430,
    n1238,
    n1428,
    n1324
  );


  xnor
  g1430
  (
    n1453,
    n1440,
    n1240,
    n1258,
    n1439
  );


  nand
  g1431
  (
    n1458,
    n1455,
    n1447,
    n1454,
    n1456
  );


  and
  g1432
  (
    n1459,
    n1446,
    n1451,
    n1452,
    n1449
  );


  or
  g1433
  (
    n1460,
    n1453,
    n1450,
    n1445,
    n1443
  );


  xnor
  g1434
  (
    n1461,
    n1442,
    n1448,
    n1457,
    n1444
  );


  xor
  g1435
  (
    n1462,
    n1458,
    n1460,
    n1459,
    n1461
  );


  xnor
  KeyGate_0_0
  (
    n157,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n45,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n477,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n573,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n522,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n813,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n589,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n100,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n696,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n697,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n287,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n595,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1322,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n478,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1294,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1106,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n867,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n528,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n760,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n339,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n622,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n881,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n614,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n611,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n672,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n345,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n273,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n935,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n176,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n673,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n151,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1007,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n211,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n454,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n46,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n286,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n862,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n1291,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n939,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n667,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n554,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n733,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n984,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n1421,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n715,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n377,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n67,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n483,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n923,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n363,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n559,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n333,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n84,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n849,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n268,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n1372,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n866,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n433,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n260,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n800,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n228,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n1423,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n1429,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n784,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

