

module Stat_1577_23_10
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n389,
  n375,
  n382,
  n373,
  n1575,
  n1571,
  n1573,
  n1563,
  n1562,
  n1556,
  n1555,
  n1559,
  n1558,
  n1574,
  n1570,
  n1567,
  n1561,
  n1565,
  n1557,
  n1572,
  n1564,
  n1560,
  n1569,
  n1602,
  n1605,
  n1603,
  n1604,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n389;
  output n375;
  output n382;
  output n373;
  output n1575;
  output n1571;
  output n1573;
  output n1563;
  output n1562;
  output n1556;
  output n1555;
  output n1559;
  output n1558;
  output n1574;
  output n1570;
  output n1567;
  output n1561;
  output n1565;
  output n1557;
  output n1572;
  output n1564;
  output n1560;
  output n1569;
  output n1602;
  output n1605;
  output n1603;
  output n1604;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n374;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1566;
  wire n1568;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n48,
    n4
  );


  buf
  g1
  (
    n80,
    n20
  );


  buf
  g2
  (
    n74,
    n11
  );


  not
  g3
  (
    KeyWire_0_9,
    n7
  );


  not
  g4
  (
    n119,
    n12
  );


  buf
  g5
  (
    n112,
    n10
  );


  not
  g6
  (
    n63,
    n25
  );


  not
  g7
  (
    n134,
    n8
  );


  buf
  g8
  (
    n30,
    n19
  );


  not
  g9
  (
    n107,
    n1
  );


  not
  g10
  (
    n75,
    n22
  );


  not
  g11
  (
    n35,
    n2
  );


  not
  g12
  (
    n51,
    n18
  );


  buf
  g13
  (
    n117,
    n17
  );


  buf
  g14
  (
    n39,
    n6
  );


  not
  g15
  (
    n124,
    n19
  );


  buf
  g16
  (
    n136,
    n17
  );


  not
  g17
  (
    n87,
    n19
  );


  not
  g18
  (
    n77,
    n26
  );


  buf
  g19
  (
    n47,
    n12
  );


  buf
  g20
  (
    n123,
    n20
  );


  buf
  g21
  (
    n118,
    n3
  );


  buf
  g22
  (
    KeyWire_0_0,
    n10
  );


  buf
  g23
  (
    KeyWire_0_2,
    n17
  );


  buf
  g24
  (
    KeyWire_0_38,
    n26
  );


  not
  g25
  (
    n45,
    n6
  );


  buf
  g26
  (
    n120,
    n12
  );


  not
  g27
  (
    n129,
    n27
  );


  buf
  g28
  (
    n76,
    n9
  );


  not
  g29
  (
    KeyWire_0_21,
    n22
  );


  not
  g30
  (
    n56,
    n22
  );


  not
  g31
  (
    n37,
    n7
  );


  buf
  g32
  (
    n54,
    n23
  );


  buf
  g33
  (
    n82,
    n12
  );


  buf
  g34
  (
    n84,
    n11
  );


  buf
  g35
  (
    n73,
    n14
  );


  buf
  g36
  (
    n133,
    n20
  );


  buf
  g37
  (
    KeyWire_0_42,
    n27
  );


  not
  g38
  (
    n114,
    n20
  );


  buf
  g39
  (
    n59,
    n2
  );


  not
  g40
  (
    n99,
    n23
  );


  not
  g41
  (
    n83,
    n15
  );


  buf
  g42
  (
    n130,
    n16
  );


  buf
  g43
  (
    n52,
    n1
  );


  buf
  g44
  (
    n97,
    n9
  );


  not
  g45
  (
    n41,
    n16
  );


  not
  g46
  (
    n85,
    n15
  );


  buf
  g47
  (
    n89,
    n22
  );


  not
  g48
  (
    n126,
    n18
  );


  buf
  g49
  (
    n42,
    n13
  );


  not
  g50
  (
    n113,
    n14
  );


  buf
  g51
  (
    n110,
    n13
  );


  not
  g52
  (
    n67,
    n16
  );


  not
  g53
  (
    n111,
    n5
  );


  not
  g54
  (
    n33,
    n14
  );


  buf
  g55
  (
    n109,
    n21
  );


  not
  g56
  (
    n55,
    n27
  );


  buf
  g57
  (
    n34,
    n25
  );


  not
  g58
  (
    n101,
    n26
  );


  buf
  g59
  (
    n29,
    n2
  );


  buf
  g60
  (
    n72,
    n9
  );


  not
  g61
  (
    n132,
    n24
  );


  buf
  g62
  (
    n92,
    n1
  );


  not
  g63
  (
    n100,
    n19
  );


  buf
  g64
  (
    n93,
    n3
  );


  buf
  g65
  (
    n81,
    n14
  );


  buf
  g66
  (
    n127,
    n16
  );


  buf
  g67
  (
    n108,
    n7
  );


  not
  g68
  (
    n31,
    n15
  );


  buf
  g69
  (
    n95,
    n6
  );


  not
  g70
  (
    n86,
    n21
  );


  buf
  g71
  (
    n88,
    n8
  );


  buf
  g72
  (
    n104,
    n15
  );


  buf
  g73
  (
    n32,
    n25
  );


  buf
  g74
  (
    n122,
    n4
  );


  not
  g75
  (
    KeyWire_0_56,
    n1
  );


  not
  g76
  (
    n94,
    n9
  );


  not
  g77
  (
    n43,
    n25
  );


  not
  g78
  (
    n98,
    n10
  );


  buf
  g79
  (
    n91,
    n23
  );


  buf
  g80
  (
    n105,
    n6
  );


  not
  g81
  (
    n57,
    n18
  );


  buf
  g82
  (
    KeyWire_0_10,
    n8
  );


  buf
  g83
  (
    n79,
    n21
  );


  buf
  g84
  (
    n69,
    n18
  );


  not
  g85
  (
    n64,
    n4
  );


  buf
  g86
  (
    n40,
    n13
  );


  buf
  g87
  (
    n36,
    n2
  );


  not
  g88
  (
    n115,
    n5
  );


  buf
  g89
  (
    n70,
    n26
  );


  buf
  g90
  (
    n66,
    n5
  );


  not
  g91
  (
    n38,
    n8
  );


  not
  g92
  (
    n68,
    n11
  );


  not
  g93
  (
    n103,
    n27
  );


  buf
  g94
  (
    n121,
    n17
  );


  not
  g95
  (
    n106,
    n24
  );


  buf
  g96
  (
    n49,
    n11
  );


  not
  g97
  (
    n131,
    n3
  );


  not
  g98
  (
    n96,
    n4
  );


  buf
  g99
  (
    n50,
    n5
  );


  buf
  g100
  (
    n90,
    n23
  );


  buf
  g101
  (
    KeyWire_0_52,
    n24
  );


  not
  g102
  (
    n62,
    n24
  );


  not
  g103
  (
    n135,
    n21
  );


  buf
  g104
  (
    n58,
    n7
  );


  buf
  g105
  (
    n44,
    n13
  );


  buf
  g106
  (
    n46,
    n3
  );


  not
  g107
  (
    n102,
    n10
  );


  buf
  g108
  (
    n284,
    n92
  );


  not
  g109
  (
    n183,
    n42
  );


  not
  g110
  (
    n253,
    n49
  );


  not
  g111
  (
    n330,
    n100
  );


  not
  g112
  (
    n288,
    n67
  );


  buf
  g113
  (
    n353,
    n95
  );


  buf
  g114
  (
    n184,
    n34
  );


  not
  g115
  (
    n321,
    n35
  );


  buf
  g116
  (
    n153,
    n99
  );


  buf
  g117
  (
    n169,
    n90
  );


  buf
  g118
  (
    n144,
    n73
  );


  not
  g119
  (
    n150,
    n34
  );


  buf
  g120
  (
    n208,
    n66
  );


  buf
  g121
  (
    n293,
    n36
  );


  not
  g122
  (
    n248,
    n34
  );


  buf
  g123
  (
    n296,
    n94
  );


  not
  g124
  (
    n262,
    n31
  );


  not
  g125
  (
    n360,
    n99
  );


  buf
  g126
  (
    n333,
    n108
  );


  buf
  g127
  (
    n329,
    n60
  );


  buf
  g128
  (
    n200,
    n80
  );


  not
  g129
  (
    n260,
    n100
  );


  buf
  g130
  (
    n213,
    n119
  );


  buf
  g131
  (
    n261,
    n117
  );


  buf
  g132
  (
    n345,
    n81
  );


  not
  g133
  (
    n294,
    n35
  );


  not
  g134
  (
    n172,
    n85
  );


  not
  g135
  (
    n299,
    n88
  );


  not
  g136
  (
    n277,
    n81
  );


  buf
  g137
  (
    n164,
    n96
  );


  not
  g138
  (
    n203,
    n104
  );


  buf
  g139
  (
    n147,
    n94
  );


  not
  g140
  (
    n344,
    n49
  );


  buf
  g141
  (
    n290,
    n88
  );


  buf
  g142
  (
    n217,
    n66
  );


  buf
  g143
  (
    n197,
    n45
  );


  not
  g144
  (
    KeyWire_0_19,
    n110
  );


  not
  g145
  (
    n148,
    n117
  );


  buf
  g146
  (
    n282,
    n95
  );


  buf
  g147
  (
    n238,
    n35
  );


  buf
  g148
  (
    n181,
    n74
  );


  buf
  g149
  (
    n265,
    n58
  );


  not
  g150
  (
    n306,
    n110
  );


  buf
  g151
  (
    n241,
    n78
  );


  not
  g152
  (
    n231,
    n58
  );


  buf
  g153
  (
    n212,
    n109
  );


  not
  g154
  (
    n177,
    n53
  );


  buf
  g155
  (
    n185,
    n38
  );


  buf
  g156
  (
    n297,
    n103
  );


  not
  g157
  (
    n276,
    n48
  );


  not
  g158
  (
    n308,
    n42
  );


  buf
  g159
  (
    n180,
    n111
  );


  buf
  g160
  (
    n224,
    n105
  );


  buf
  g161
  (
    n140,
    n82
  );


  buf
  g162
  (
    n310,
    n105
  );


  not
  g163
  (
    n259,
    n57
  );


  not
  g164
  (
    n315,
    n90
  );


  not
  g165
  (
    n291,
    n29
  );


  buf
  g166
  (
    n195,
    n67
  );


  not
  g167
  (
    n194,
    n109
  );


  not
  g168
  (
    n222,
    n87
  );


  not
  g169
  (
    n305,
    n47
  );


  buf
  g170
  (
    n250,
    n34
  );


  not
  g171
  (
    n202,
    n74
  );


  buf
  g172
  (
    n314,
    n65
  );


  buf
  g173
  (
    n192,
    n65
  );


  not
  g174
  (
    n210,
    n100
  );


  not
  g175
  (
    n341,
    n90
  );


  buf
  g176
  (
    n255,
    n82
  );


  not
  g177
  (
    n313,
    n46
  );


  buf
  g178
  (
    n141,
    n32
  );


  buf
  g179
  (
    n201,
    n115
  );


  buf
  g180
  (
    n155,
    n46
  );


  buf
  g181
  (
    n274,
    n72
  );


  not
  g182
  (
    n190,
    n109
  );


  buf
  g183
  (
    n251,
    n116
  );


  buf
  g184
  (
    n176,
    n56
  );


  buf
  g185
  (
    n300,
    n43
  );


  not
  g186
  (
    n232,
    n46
  );


  not
  g187
  (
    n328,
    n111
  );


  buf
  g188
  (
    n216,
    n59
  );


  buf
  g189
  (
    n351,
    n116
  );


  not
  g190
  (
    n298,
    n36
  );


  not
  g191
  (
    n320,
    n108
  );


  not
  g192
  (
    n340,
    n60
  );


  not
  g193
  (
    n281,
    n68
  );


  buf
  g194
  (
    n168,
    n89
  );


  buf
  g195
  (
    n158,
    n89
  );


  buf
  g196
  (
    n356,
    n39
  );


  buf
  g197
  (
    n167,
    n106
  );


  buf
  g198
  (
    n145,
    n72
  );


  buf
  g199
  (
    n338,
    n30
  );


  not
  g200
  (
    n245,
    n47
  );


  buf
  g201
  (
    n348,
    n31
  );


  buf
  g202
  (
    n346,
    n43
  );


  not
  g203
  (
    n339,
    n117
  );


  not
  g204
  (
    KeyWire_0_44,
    n58
  );


  buf
  g205
  (
    n165,
    n118
  );


  buf
  g206
  (
    KeyWire_0_28,
    n72
  );


  buf
  g207
  (
    n178,
    n84
  );


  buf
  g208
  (
    KeyWire_0_35,
    n99
  );


  not
  g209
  (
    n207,
    n67
  );


  buf
  g210
  (
    n154,
    n94
  );


  not
  g211
  (
    n157,
    n56
  );


  buf
  g212
  (
    n322,
    n87
  );


  buf
  g213
  (
    n233,
    n42
  );


  not
  g214
  (
    n278,
    n29
  );


  buf
  g215
  (
    n191,
    n97
  );


  buf
  g216
  (
    n243,
    n78
  );


  not
  g217
  (
    n283,
    n74
  );


  not
  g218
  (
    n239,
    n108
  );


  buf
  g219
  (
    n163,
    n57
  );


  not
  g220
  (
    n237,
    n41
  );


  not
  g221
  (
    n179,
    n54
  );


  not
  g222
  (
    n295,
    n39
  );


  buf
  g223
  (
    n268,
    n102
  );


  buf
  g224
  (
    n254,
    n52
  );


  not
  g225
  (
    n264,
    n51
  );


  not
  g226
  (
    n137,
    n50
  );


  buf
  g227
  (
    KeyWire_0_45,
    n110
  );


  buf
  g228
  (
    n162,
    n52
  );


  not
  g229
  (
    n171,
    n84
  );


  not
  g230
  (
    n287,
    n99
  );


  not
  g231
  (
    n174,
    n107
  );


  buf
  g232
  (
    n143,
    n115
  );


  not
  g233
  (
    n311,
    n84
  );


  not
  g234
  (
    n186,
    n116
  );


  not
  g235
  (
    n156,
    n33
  );


  not
  g236
  (
    n204,
    n65
  );


  not
  g237
  (
    n247,
    n73
  );


  buf
  g238
  (
    n149,
    n56
  );


  buf
  g239
  (
    n175,
    n45
  );


  not
  g240
  (
    n323,
    n102
  );


  buf
  g241
  (
    n226,
    n92
  );


  not
  g242
  (
    n318,
    n83
  );


  not
  g243
  (
    n225,
    n36
  );


  not
  g244
  (
    n342,
    n115
  );


  buf
  g245
  (
    n316,
    n112
  );


  buf
  g246
  (
    n242,
    n77
  );


  buf
  g247
  (
    n280,
    n50
  );


  buf
  g248
  (
    n166,
    n91
  );


  buf
  g249
  (
    KeyWire_0_24,
    n54
  );


  not
  g250
  (
    n263,
    n106
  );


  buf
  g251
  (
    n347,
    n41
  );


  not
  g252
  (
    n160,
    n114
  );


  not
  g253
  (
    n337,
    n93
  );


  buf
  g254
  (
    n285,
    n51
  );


  not
  g255
  (
    n193,
    n66
  );


  buf
  g256
  (
    n359,
    n66
  );


  buf
  g257
  (
    n151,
    n80
  );


  not
  g258
  (
    n173,
    n47
  );


  not
  g259
  (
    n198,
    n69
  );


  buf
  g260
  (
    n286,
    n95
  );


  buf
  g261
  (
    n349,
    n69
  );


  buf
  g262
  (
    n357,
    n31
  );


  buf
  g263
  (
    n324,
    n104
  );


  not
  g264
  (
    n302,
    n48
  );


  buf
  g265
  (
    n301,
    n94
  );


  buf
  g266
  (
    n332,
    n96
  );


  buf
  g267
  (
    n257,
    n109
  );


  not
  g268
  (
    n138,
    n113
  );


  not
  g269
  (
    n289,
    n65
  );


  buf
  g270
  (
    n211,
    n110
  );


  not
  g271
  (
    n331,
    n68
  );


  not
  g272
  (
    n206,
    n98
  );


  buf
  g273
  (
    n317,
    n91
  );


  buf
  g274
  (
    n214,
    n62
  );


  not
  g275
  (
    n161,
    n31
  );


  buf
  g276
  (
    n307,
    n98
  );


  buf
  g277
  (
    n170,
    n30
  );


  not
  g278
  (
    n292,
    n76
  );


  buf
  g279
  (
    n258,
    n73
  );


  not
  g280
  (
    n235,
    n86
  );


  not
  g281
  (
    KeyWire_0_50,
    n37
  );


  buf
  g282
  (
    n219,
    n71
  );


  buf
  g283
  (
    n229,
    n29
  );


  buf
  g284
  (
    n236,
    n55
  );


  nand
  g285
  (
    n326,
    n88,
    n77
  );


  nor
  g286
  (
    n187,
    n114,
    n50
  );


  nor
  g287
  (
    n266,
    n44,
    n78,
    n79
  );


  nor
  g288
  (
    n209,
    n64,
    n102,
    n82,
    n90
  );


  and
  g289
  (
    n220,
    n53,
    n64,
    n41,
    n76
  );


  nor
  g290
  (
    KeyWire_0_5,
    n86,
    n95,
    n64,
    n40
  );


  nand
  g291
  (
    n188,
    n97,
    n30,
    n75,
    n62
  );


  xor
  g292
  (
    n309,
    n33,
    n32,
    n85,
    n89
  );


  nor
  g293
  (
    n199,
    n116,
    n61,
    n105,
    n86
  );


  xnor
  g294
  (
    n267,
    n88,
    n92,
    n75,
    n81
  );


  or
  g295
  (
    n230,
    n117,
    n51,
    n33,
    n39
  );


  xnor
  g296
  (
    n334,
    n107,
    n105,
    n60,
    n112
  );


  and
  g297
  (
    n350,
    n87,
    n40,
    n37,
    n104
  );


  xor
  g298
  (
    n159,
    n43,
    n75,
    n30,
    n93
  );


  xnor
  g299
  (
    n325,
    n62,
    n85,
    n45,
    n52
  );


  or
  g300
  (
    n249,
    n97,
    n118,
    n59,
    n111
  );


  or
  g301
  (
    n327,
    n71,
    n36,
    n44,
    n104
  );


  xnor
  g302
  (
    n215,
    n75,
    n38,
    n76,
    n55
  );


  xnor
  g303
  (
    n234,
    n52,
    n40,
    n63,
    n61
  );


  and
  g304
  (
    n146,
    n38,
    n51,
    n47,
    n79
  );


  nand
  g305
  (
    n304,
    n54,
    n71,
    n39,
    n46
  );


  nand
  g306
  (
    n271,
    n56,
    n118,
    n82,
    n64
  );


  and
  g307
  (
    KeyWire_0_12,
    n111,
    n101,
    n58,
    n96
  );


  or
  g308
  (
    n269,
    n69,
    n107,
    n70,
    n103
  );


  xnor
  g309
  (
    n228,
    n113,
    n38,
    n83,
    n69
  );


  nand
  g310
  (
    n221,
    n67,
    n112,
    n32
  );


  xnor
  g311
  (
    n189,
    n42,
    n93,
    n101
  );


  or
  g312
  (
    n336,
    n71,
    n93,
    n87,
    n68
  );


  nand
  g313
  (
    n355,
    n40,
    n98,
    n83,
    n44
  );


  or
  g314
  (
    n273,
    n77,
    n83,
    n89,
    n96
  );


  xor
  g315
  (
    n358,
    n62,
    n63,
    n57,
    n80
  );


  nor
  g316
  (
    n335,
    n113,
    n55,
    n44,
    n114
  );


  and
  g317
  (
    n152,
    n55,
    n63,
    n103,
    n29
  );


  or
  g318
  (
    n275,
    n98,
    n115,
    n48,
    n49
  );


  nor
  g319
  (
    n142,
    n60,
    n108,
    n72,
    n37
  );


  xnor
  g320
  (
    n272,
    n61,
    n50,
    n53,
    n76
  );


  nor
  g321
  (
    n343,
    n54,
    n114,
    n59,
    n68
  );


  nand
  g322
  (
    n244,
    n97,
    n32,
    n59,
    n91
  );


  xnor
  g323
  (
    n352,
    n118,
    n57,
    n35,
    n107
  );


  nor
  g324
  (
    n182,
    n106,
    n48,
    n41,
    n86
  );


  and
  g325
  (
    KeyWire_0_33,
    n79,
    n101,
    n45,
    n43
  );


  nor
  g326
  (
    n279,
    n73,
    n81,
    n100,
    n70
  );


  and
  g327
  (
    n240,
    n61,
    n70,
    n80
  );


  or
  g328
  (
    n256,
    n91,
    n79,
    n102,
    n84
  );


  or
  g329
  (
    n196,
    n53,
    n113,
    n63,
    n33
  );


  and
  g330
  (
    n270,
    n92,
    n74,
    n106,
    n85
  );


  or
  g331
  (
    n139,
    n77,
    n49,
    n37,
    n103
  );


  or
  g332
  (
    n362,
    n139,
    n144,
    n137,
    n138
  );


  xnor
  g333
  (
    n361,
    n141,
    n142,
    n140,
    n143
  );


  not
  g334
  (
    n364,
    n361
  );


  buf
  g335
  (
    n363,
    n362
  );


  xor
  g336
  (
    n365,
    n120,
    n124,
    n125,
    n363
  );


  xor
  g337
  (
    n369,
    n121,
    n364,
    n119,
    n123
  );


  nor
  g338
  (
    n370,
    n121,
    n122,
    n124
  );


  xnor
  g339
  (
    n367,
    n121,
    n364,
    n123,
    n124
  );


  or
  g340
  (
    n368,
    n364,
    n123,
    n363,
    n122
  );


  xor
  g341
  (
    n366,
    n120,
    n123,
    n121,
    n363
  );


  xnor
  g342
  (
    n372,
    n124,
    n119,
    n120,
    n364
  );


  xor
  g343
  (
    n371,
    n363,
    n119,
    n120,
    n122
  );


  or
  g344
  (
    n374,
    n370,
    n365,
    n366,
    n224
  );


  or
  g345
  (
    n402,
    n166,
    n169,
    n190,
    n229
  );


  xor
  g346
  (
    n382,
    n165,
    n368,
    n211,
    n171
  );


  xnor
  g347
  (
    n376,
    n156,
    n202,
    n367,
    n155
  );


  or
  g348
  (
    n373,
    n188,
    n195,
    n233,
    n182
  );


  or
  g349
  (
    n378,
    n231,
    n367,
    n196,
    n148
  );


  xnor
  g350
  (
    n388,
    n151,
    n369,
    n185,
    n367
  );


  xor
  g351
  (
    n398,
    n176,
    n232,
    n203,
    n170
  );


  nand
  g352
  (
    n387,
    n368,
    n157,
    n186,
    n199
  );


  nand
  g353
  (
    n395,
    n217,
    n177,
    n369,
    n367
  );


  xor
  g354
  (
    n377,
    n197,
    n236,
    n371,
    n370
  );


  or
  g355
  (
    n401,
    n369,
    n228,
    n180,
    n234
  );


  or
  g356
  (
    n396,
    n366,
    n154,
    n167,
    n173
  );


  xnor
  g357
  (
    n381,
    n189,
    n215,
    n365,
    n213
  );


  nor
  g358
  (
    n389,
    n146,
    n218,
    n145,
    n219
  );


  xnor
  g359
  (
    n394,
    n174,
    n160,
    n150,
    n153
  );


  and
  g360
  (
    n380,
    n210,
    n370,
    n368,
    n198
  );


  nor
  g361
  (
    n375,
    n164,
    n209,
    n212,
    n183
  );


  and
  g362
  (
    n384,
    n370,
    n207,
    n200,
    n159
  );


  nor
  g363
  (
    n390,
    n221,
    n369,
    n371,
    n201
  );


  and
  g364
  (
    n379,
    n192,
    n147,
    n162,
    n214
  );


  nand
  g365
  (
    n386,
    n158,
    n366,
    n371
  );


  or
  g366
  (
    n385,
    n149,
    n365,
    n372,
    n178
  );


  nand
  g367
  (
    n399,
    n237,
    n226,
    n194,
    n227
  );


  xnor
  g368
  (
    n400,
    n168,
    n225,
    n222,
    n223
  );


  or
  g369
  (
    n393,
    n368,
    n235,
    n371,
    n365
  );


  nor
  g370
  (
    n392,
    n187,
    n208,
    n372,
    n191
  );


  or
  g371
  (
    n397,
    n220,
    n175,
    n216,
    n206
  );


  and
  g372
  (
    n403,
    n193,
    n184,
    n172,
    n181
  );


  xor
  g373
  (
    n391,
    n204,
    n179,
    n163,
    n205
  );


  xnor
  g374
  (
    n383,
    n152,
    n161,
    n230,
    n372
  );


  buf
  g375
  (
    n429,
    n287
  );


  buf
  g376
  (
    n412,
    n385
  );


  not
  g377
  (
    n415,
    n396
  );


  not
  g378
  (
    n420,
    n397
  );


  not
  g379
  (
    n419,
    n251
  );


  buf
  g380
  (
    n405,
    n386
  );


  buf
  g381
  (
    n416,
    n249
  );


  not
  g382
  (
    n426,
    n377
  );


  xor
  g383
  (
    n410,
    n246,
    n390
  );


  nor
  g384
  (
    n406,
    n255,
    n284
  );


  and
  g385
  (
    n423,
    n392,
    n266,
    n286,
    n384
  );


  nand
  g386
  (
    KeyWire_0_18,
    n250,
    n391,
    n279,
    n381
  );


  xor
  g387
  (
    n418,
    n401,
    n389,
    n274,
    n399
  );


  and
  g388
  (
    n414,
    n273,
    n394,
    n282,
    n253
  );


  xnor
  g389
  (
    n428,
    n242,
    n402,
    n254,
    n278
  );


  nor
  g390
  (
    n422,
    n277,
    n280,
    n240,
    n262
  );


  xnor
  g391
  (
    n409,
    n283,
    n395,
    n247,
    n393
  );


  and
  g392
  (
    n425,
    n379,
    n271,
    n268,
    n270
  );


  nor
  g393
  (
    n408,
    n275,
    n252,
    n256,
    n387
  );


  xor
  g394
  (
    n417,
    n259,
    n239,
    n238,
    n241
  );


  nand
  g395
  (
    n427,
    n263,
    n260,
    n258,
    n398
  );


  or
  g396
  (
    n424,
    n276,
    n281,
    n400,
    n261
  );


  xor
  g397
  (
    n404,
    n380,
    n244,
    n382,
    n265
  );


  nor
  g398
  (
    n413,
    n272,
    n267,
    n388,
    n285
  );


  and
  g399
  (
    KeyWire_0_49,
    n243,
    n245,
    n248,
    n269
  );


  xnor
  g400
  (
    n421,
    n378,
    n257,
    n264,
    n383
  );


  not
  g401
  (
    KeyWire_0_43,
    n405
  );


  buf
  g402
  (
    n448,
    n410
  );


  buf
  g403
  (
    n449,
    n407
  );


  buf
  g404
  (
    n443,
    n406
  );


  buf
  g405
  (
    n435,
    n413
  );


  not
  g406
  (
    n436,
    n414
  );


  not
  g407
  (
    n432,
    n409
  );


  buf
  g408
  (
    n440,
    n408
  );


  buf
  g409
  (
    KeyWire_0_48,
    n418
  );


  buf
  g410
  (
    n431,
    n419
  );


  buf
  g411
  (
    n434,
    n412
  );


  not
  g412
  (
    n430,
    n411
  );


  buf
  g413
  (
    n439,
    n417
  );


  not
  g414
  (
    n446,
    n423
  );


  buf
  g415
  (
    n438,
    n416
  );


  buf
  g416
  (
    n445,
    n415
  );


  buf
  g417
  (
    n447,
    n421
  );


  buf
  g418
  (
    KeyWire_0_6,
    n422
  );


  buf
  g419
  (
    n444,
    n404
  );


  not
  g420
  (
    n437,
    n420
  );


  buf
  g421
  (
    n453,
    n449
  );


  buf
  g422
  (
    n486,
    n439
  );


  buf
  g423
  (
    n456,
    n437
  );


  not
  g424
  (
    n526,
    n436
  );


  buf
  g425
  (
    n468,
    n448
  );


  not
  g426
  (
    n452,
    n125
  );


  not
  g427
  (
    n458,
    n447
  );


  not
  g428
  (
    KeyWire_0_60,
    n403
  );


  buf
  g429
  (
    n487,
    n430
  );


  buf
  g430
  (
    n527,
    n442
  );


  not
  g431
  (
    n480,
    n440
  );


  buf
  g432
  (
    n469,
    n444
  );


  buf
  g433
  (
    n477,
    n443
  );


  not
  g434
  (
    n525,
    n436
  );


  buf
  g435
  (
    n522,
    n447
  );


  not
  g436
  (
    n495,
    n442
  );


  buf
  g437
  (
    n519,
    n446
  );


  not
  g438
  (
    n450,
    n434
  );


  buf
  g439
  (
    KeyWire_0_20,
    n446
  );


  buf
  g440
  (
    n490,
    n435
  );


  not
  g441
  (
    n497,
    n444
  );


  not
  g442
  (
    n454,
    n441
  );


  buf
  g443
  (
    n457,
    n430
  );


  buf
  g444
  (
    KeyWire_0_26,
    n445
  );


  buf
  g445
  (
    n518,
    n129
  );


  buf
  g446
  (
    n504,
    n447
  );


  buf
  g447
  (
    n500,
    n128
  );


  not
  g448
  (
    n514,
    n448
  );


  not
  g449
  (
    n494,
    n440
  );


  not
  g450
  (
    n515,
    n436
  );


  not
  g451
  (
    n508,
    n436
  );


  not
  g452
  (
    n520,
    n431
  );


  not
  g453
  (
    n463,
    n432
  );


  buf
  g454
  (
    n512,
    n444
  );


  buf
  g455
  (
    n524,
    n443
  );


  not
  g456
  (
    n464,
    n433
  );


  not
  g457
  (
    n466,
    n445
  );


  not
  g458
  (
    n451,
    n443
  );


  not
  g459
  (
    n521,
    n434
  );


  not
  g460
  (
    n481,
    n431
  );


  not
  g461
  (
    n498,
    n432
  );


  not
  g462
  (
    n462,
    n430
  );


  not
  g463
  (
    KeyWire_0_32,
    n442
  );


  not
  g464
  (
    n507,
    n126
  );


  not
  g465
  (
    n496,
    n128
  );


  not
  g466
  (
    n523,
    n430
  );


  buf
  g467
  (
    n476,
    n438
  );


  buf
  g468
  (
    n506,
    n437
  );


  buf
  g469
  (
    n475,
    n130
  );


  not
  g470
  (
    n505,
    n441
  );


  not
  g471
  (
    n509,
    n438
  );


  buf
  g472
  (
    n467,
    n435
  );


  not
  g473
  (
    n459,
    n432
  );


  buf
  g474
  (
    n479,
    n433
  );


  buf
  g475
  (
    n513,
    n441
  );


  buf
  g476
  (
    n516,
    n442
  );


  buf
  g477
  (
    n489,
    n437
  );


  not
  g478
  (
    n474,
    n432
  );


  not
  g479
  (
    n478,
    n439
  );


  buf
  g480
  (
    n502,
    n127
  );


  buf
  g481
  (
    n499,
    n431
  );


  not
  g482
  (
    n473,
    n449
  );


  buf
  g483
  (
    n517,
    n433
  );


  buf
  g484
  (
    n465,
    n448
  );


  not
  g485
  (
    n470,
    n125
  );


  buf
  g486
  (
    n460,
    n440
  );


  not
  g487
  (
    n488,
    n372
  );


  buf
  g488
  (
    n493,
    n127
  );


  buf
  g489
  (
    KeyWire_0_41,
    n431
  );


  not
  g490
  (
    n482,
    n435
  );


  xnor
  g491
  (
    n501,
    n446,
    n445
  );


  nand
  g492
  (
    n455,
    n438,
    n126,
    n439,
    n437
  );


  nor
  g493
  (
    n510,
    n440,
    n127,
    n434,
    n125
  );


  xnor
  g494
  (
    n491,
    n444,
    n443,
    n447,
    n128
  );


  xor
  g495
  (
    n461,
    n128,
    n126,
    n129,
    n446
  );


  xor
  g496
  (
    n471,
    n129,
    n445,
    n439,
    n127
  );


  xor
  g497
  (
    n483,
    n129,
    n126,
    n441,
    n434
  );


  xnor
  g498
  (
    n503,
    n435,
    n448,
    n438,
    n433
  );


  buf
  g499
  (
    n535,
    n484
  );


  not
  g500
  (
    n586,
    n511
  );


  not
  g501
  (
    n534,
    n501
  );


  buf
  g502
  (
    n680,
    n477
  );


  buf
  g503
  (
    n635,
    n476
  );


  not
  g504
  (
    n591,
    n485
  );


  buf
  g505
  (
    n711,
    n458
  );


  not
  g506
  (
    KeyWire_0_11,
    n479
  );


  buf
  g507
  (
    n599,
    n509
  );


  not
  g508
  (
    n679,
    n475
  );


  buf
  g509
  (
    n677,
    n504
  );


  buf
  g510
  (
    n549,
    n499
  );


  buf
  g511
  (
    n672,
    n498
  );


  not
  g512
  (
    n621,
    n494
  );


  buf
  g513
  (
    n612,
    n474
  );


  buf
  g514
  (
    n661,
    n463
  );


  buf
  g515
  (
    n648,
    n493
  );


  buf
  g516
  (
    n567,
    n456
  );


  buf
  g517
  (
    n710,
    n493
  );


  not
  g518
  (
    n542,
    n453
  );


  not
  g519
  (
    KeyWire_0_8,
    n512
  );


  not
  g520
  (
    n564,
    n503
  );


  not
  g521
  (
    n551,
    n508
  );


  buf
  g522
  (
    n556,
    n495
  );


  not
  g523
  (
    n618,
    n505
  );


  buf
  g524
  (
    n678,
    n501
  );


  buf
  g525
  (
    n708,
    n495
  );


  not
  g526
  (
    n596,
    n510
  );


  not
  g527
  (
    n714,
    n494
  );


  not
  g528
  (
    n583,
    n475
  );


  not
  g529
  (
    n566,
    n474
  );


  not
  g530
  (
    n683,
    n514
  );


  buf
  g531
  (
    n707,
    n497
  );


  not
  g532
  (
    n703,
    n496
  );


  buf
  g533
  (
    n706,
    n502
  );


  buf
  g534
  (
    n656,
    n512
  );


  buf
  g535
  (
    n585,
    n450
  );


  not
  g536
  (
    n624,
    n507
  );


  buf
  g537
  (
    n654,
    n479
  );


  buf
  g538
  (
    n643,
    n514
  );


  not
  g539
  (
    n589,
    n486
  );


  buf
  g540
  (
    n605,
    n468
  );


  buf
  g541
  (
    n616,
    n498
  );


  buf
  g542
  (
    n669,
    n477
  );


  not
  g543
  (
    n715,
    n491
  );


  not
  g544
  (
    n694,
    n512
  );


  buf
  g545
  (
    n613,
    n495
  );


  buf
  g546
  (
    n532,
    n484
  );


  buf
  g547
  (
    n653,
    n486
  );


  buf
  g548
  (
    n704,
    n498
  );


  not
  g549
  (
    n602,
    n491
  );


  not
  g550
  (
    n619,
    n481
  );


  not
  g551
  (
    n593,
    n482
  );


  buf
  g552
  (
    n636,
    n499
  );


  buf
  g553
  (
    n663,
    n494
  );


  buf
  g554
  (
    n692,
    n504
  );


  buf
  g555
  (
    n557,
    n484
  );


  not
  g556
  (
    n627,
    n471
  );


  not
  g557
  (
    KeyWire_0_39,
    n485
  );


  not
  g558
  (
    KeyWire_0_4,
    n508
  );


  buf
  g559
  (
    n530,
    n474
  );


  not
  g560
  (
    n670,
    n513
  );


  not
  g561
  (
    n685,
    n489
  );


  buf
  g562
  (
    n594,
    n513
  );


  buf
  g563
  (
    n699,
    n505
  );


  buf
  g564
  (
    n641,
    n491
  );


  not
  g565
  (
    n579,
    n484
  );


  buf
  g566
  (
    n600,
    n483
  );


  buf
  g567
  (
    n559,
    n497
  );


  not
  g568
  (
    n614,
    n510
  );


  not
  g569
  (
    n681,
    n498
  );


  not
  g570
  (
    n581,
    n504
  );


  buf
  g571
  (
    n665,
    n500
  );


  not
  g572
  (
    n701,
    n507
  );


  not
  g573
  (
    n697,
    n488
  );


  not
  g574
  (
    n646,
    n482
  );


  not
  g575
  (
    n705,
    n488
  );


  not
  g576
  (
    n541,
    n496
  );


  buf
  g577
  (
    n550,
    n483
  );


  not
  g578
  (
    KeyWire_0_61,
    n514
  );


  buf
  g579
  (
    n642,
    n490
  );


  not
  g580
  (
    n687,
    n461
  );


  buf
  g581
  (
    n623,
    n501
  );


  not
  g582
  (
    n552,
    n469
  );


  buf
  g583
  (
    n572,
    n485
  );


  buf
  g584
  (
    n634,
    n502
  );


  buf
  g585
  (
    n698,
    n478
  );


  buf
  g586
  (
    n644,
    n482
  );


  buf
  g587
  (
    n611,
    n509
  );


  not
  g588
  (
    n629,
    n452
  );


  buf
  g589
  (
    n676,
    n483
  );


  not
  g590
  (
    n649,
    n511
  );


  buf
  g591
  (
    n660,
    n490
  );


  not
  g592
  (
    n662,
    n497
  );


  not
  g593
  (
    n538,
    n507
  );


  buf
  g594
  (
    n647,
    n477
  );


  buf
  g595
  (
    n639,
    n476
  );


  buf
  g596
  (
    n632,
    n500
  );


  not
  g597
  (
    KeyWire_0_23,
    n493
  );


  not
  g598
  (
    n638,
    n472
  );


  buf
  g599
  (
    n582,
    n470
  );


  not
  g600
  (
    n592,
    n511
  );


  buf
  g601
  (
    n574,
    n478
  );


  buf
  g602
  (
    n597,
    n478
  );


  buf
  g603
  (
    n576,
    n483
  );


  buf
  g604
  (
    n543,
    n506
  );


  buf
  g605
  (
    n571,
    n466
  );


  buf
  g606
  (
    n555,
    n480
  );


  buf
  g607
  (
    n626,
    n486
  );


  buf
  g608
  (
    n658,
    n506
  );


  not
  g609
  (
    n617,
    n479
  );


  buf
  g610
  (
    n684,
    n492
  );


  not
  g611
  (
    n631,
    n473
  );


  buf
  g612
  (
    n713,
    n513
  );


  not
  g613
  (
    n558,
    n476
  );


  not
  g614
  (
    n547,
    n476
  );


  buf
  g615
  (
    n610,
    n504
  );


  buf
  g616
  (
    n544,
    n506
  );


  buf
  g617
  (
    n569,
    n485
  );


  buf
  g618
  (
    n563,
    n505
  );


  not
  g619
  (
    n625,
    n481
  );


  not
  g620
  (
    n709,
    n490
  );


  buf
  g621
  (
    n690,
    n459
  );


  buf
  g622
  (
    n688,
    n497
  );


  buf
  g623
  (
    n609,
    n462
  );


  not
  g624
  (
    n640,
    n509
  );


  not
  g625
  (
    n620,
    n474
  );


  not
  g626
  (
    n598,
    n506
  );


  buf
  g627
  (
    n560,
    n502
  );


  not
  g628
  (
    n673,
    n503
  );


  not
  g629
  (
    n531,
    n487
  );


  not
  g630
  (
    n584,
    n482
  );


  buf
  g631
  (
    n666,
    n514
  );


  not
  g632
  (
    n689,
    n490
  );


  buf
  g633
  (
    n533,
    n455
  );


  not
  g634
  (
    n545,
    n478
  );


  not
  g635
  (
    n659,
    n496
  );


  not
  g636
  (
    n607,
    n502
  );


  not
  g637
  (
    n712,
    n492
  );


  not
  g638
  (
    n615,
    n487
  );


  not
  g639
  (
    n575,
    n493
  );


  not
  g640
  (
    n570,
    n503
  );


  buf
  g641
  (
    n691,
    n500
  );


  not
  g642
  (
    n655,
    n489
  );


  buf
  g643
  (
    n603,
    n510
  );


  buf
  g644
  (
    n652,
    n480
  );


  not
  g645
  (
    n536,
    n475
  );


  buf
  g646
  (
    n601,
    n481
  );


  buf
  g647
  (
    n664,
    n480
  );


  buf
  g648
  (
    n637,
    n465
  );


  buf
  g649
  (
    n528,
    n492
  );


  buf
  g650
  (
    n695,
    n507
  );


  not
  g651
  (
    n693,
    n512
  );


  not
  g652
  (
    n628,
    n508
  );


  buf
  g653
  (
    n630,
    n496
  );


  buf
  g654
  (
    n671,
    n494
  );


  buf
  g655
  (
    n682,
    n492
  );


  buf
  g656
  (
    n675,
    n464
  );


  not
  g657
  (
    n587,
    n509
  );


  not
  g658
  (
    n546,
    n451
  );


  buf
  g659
  (
    n529,
    n499
  );


  not
  g660
  (
    n651,
    n508
  );


  buf
  g661
  (
    n700,
    n487
  );


  not
  g662
  (
    KeyWire_0_22,
    n487
  );


  buf
  g663
  (
    n578,
    n477
  );


  buf
  g664
  (
    n667,
    n454
  );


  not
  g665
  (
    n565,
    n503
  );


  not
  g666
  (
    KeyWire_0_3,
    n510
  );


  buf
  g667
  (
    n540,
    n460
  );


  not
  g668
  (
    n608,
    n489
  );


  buf
  g669
  (
    n561,
    n475
  );


  not
  g670
  (
    n645,
    n491
  );


  buf
  g671
  (
    n577,
    n479
  );


  not
  g672
  (
    n573,
    n488
  );


  buf
  g673
  (
    n622,
    n481
  );


  not
  g674
  (
    n606,
    n499
  );


  buf
  g675
  (
    n657,
    n489
  );


  buf
  g676
  (
    n562,
    n505
  );


  buf
  g677
  (
    n568,
    n480
  );


  buf
  g678
  (
    n650,
    n511
  );


  buf
  g679
  (
    n686,
    n488
  );


  not
  g680
  (
    n604,
    n513
  );


  buf
  g681
  (
    n702,
    n500
  );


  buf
  g682
  (
    n588,
    n486
  );


  buf
  g683
  (
    KeyWire_0_15,
    n457
  );


  buf
  g684
  (
    n595,
    n467
  );


  not
  g685
  (
    n590,
    n501
  );


  not
  g686
  (
    n580,
    n495
  );


  not
  g687
  (
    n1176,
    n624
  );


  buf
  g688
  (
    n1074,
    n560
  );


  not
  g689
  (
    n1120,
    n643
  );


  buf
  g690
  (
    n1147,
    n607
  );


  buf
  g691
  (
    n985,
    n607
  );


  buf
  g692
  (
    n1106,
    n556
  );


  buf
  g693
  (
    n771,
    n575
  );


  not
  g694
  (
    n1180,
    n593
  );


  buf
  g695
  (
    n1156,
    n612
  );


  buf
  g696
  (
    n728,
    n597
  );


  buf
  g697
  (
    n1056,
    n544
  );


  not
  g698
  (
    n1104,
    n558
  );


  not
  g699
  (
    n850,
    n649
  );


  buf
  g700
  (
    n769,
    n614
  );


  not
  g701
  (
    n1031,
    n632
  );


  not
  g702
  (
    n725,
    n590
  );


  not
  g703
  (
    KeyWire_0_59,
    n579
  );


  buf
  g704
  (
    n1177,
    n561
  );


  buf
  g705
  (
    n898,
    n619
  );


  not
  g706
  (
    n1050,
    n603
  );


  buf
  g707
  (
    n823,
    n621
  );


  buf
  g708
  (
    n984,
    n587
  );


  buf
  g709
  (
    n1146,
    n558
  );


  buf
  g710
  (
    n731,
    n609
  );


  not
  g711
  (
    n871,
    n605
  );


  not
  g712
  (
    n955,
    n568
  );


  not
  g713
  (
    n1200,
    n616
  );


  buf
  g714
  (
    n966,
    n650
  );


  not
  g715
  (
    n992,
    n594
  );


  buf
  g716
  (
    n958,
    n605
  );


  not
  g717
  (
    n1068,
    n639
  );


  not
  g718
  (
    n1126,
    n543
  );


  buf
  g719
  (
    n774,
    n553
  );


  not
  g720
  (
    n1015,
    n529
  );


  buf
  g721
  (
    n755,
    n627
  );


  not
  g722
  (
    n1211,
    n579
  );


  buf
  g723
  (
    n1095,
    n586
  );


  not
  g724
  (
    n1041,
    n565
  );


  buf
  g725
  (
    n859,
    n602
  );


  buf
  g726
  (
    n1210,
    n552
  );


  buf
  g727
  (
    n913,
    n530
  );


  buf
  g728
  (
    n949,
    n536
  );


  buf
  g729
  (
    n1030,
    n574
  );


  buf
  g730
  (
    n1206,
    n609
  );


  not
  g731
  (
    n720,
    n594
  );


  buf
  g732
  (
    n1174,
    n562
  );


  buf
  g733
  (
    n1117,
    n576
  );


  not
  g734
  (
    n874,
    n571
  );


  not
  g735
  (
    n877,
    n606
  );


  not
  g736
  (
    n905,
    n622
  );


  not
  g737
  (
    n937,
    n553
  );


  buf
  g738
  (
    n999,
    n637
  );


  buf
  g739
  (
    n788,
    n615
  );


  buf
  g740
  (
    n936,
    n595
  );


  not
  g741
  (
    n880,
    n529
  );


  buf
  g742
  (
    n977,
    n583
  );


  buf
  g743
  (
    n903,
    n621
  );


  not
  g744
  (
    n969,
    n571
  );


  not
  g745
  (
    n849,
    n622
  );


  not
  g746
  (
    n965,
    n541
  );


  buf
  g747
  (
    n734,
    n587
  );


  not
  g748
  (
    n1110,
    n639
  );


  not
  g749
  (
    n1158,
    n516
  );


  not
  g750
  (
    n1112,
    n578
  );


  not
  g751
  (
    n946,
    n519
  );


  buf
  g752
  (
    n972,
    n598
  );


  buf
  g753
  (
    n914,
    n585
  );


  not
  g754
  (
    n727,
    n570
  );


  not
  g755
  (
    n869,
    n578
  );


  buf
  g756
  (
    n1167,
    n564
  );


  not
  g757
  (
    n1090,
    n615
  );


  buf
  g758
  (
    n828,
    n591
  );


  not
  g759
  (
    n1119,
    n549
  );


  not
  g760
  (
    n978,
    n561
  );


  buf
  g761
  (
    n890,
    n532
  );


  not
  g762
  (
    n824,
    n567
  );


  not
  g763
  (
    n883,
    n599
  );


  buf
  g764
  (
    n820,
    n562
  );


  not
  g765
  (
    n1081,
    n594
  );


  buf
  g766
  (
    n741,
    n650
  );


  buf
  g767
  (
    n840,
    n606
  );


  not
  g768
  (
    n738,
    n576
  );


  not
  g769
  (
    n1209,
    n589
  );


  buf
  g770
  (
    n1017,
    n515
  );


  not
  g771
  (
    n736,
    n646
  );


  not
  g772
  (
    n835,
    n540
  );


  buf
  g773
  (
    n1212,
    n563
  );


  buf
  g774
  (
    n902,
    n557
  );


  not
  g775
  (
    n893,
    n645
  );


  buf
  g776
  (
    n799,
    n610
  );


  not
  g777
  (
    n1185,
    n538
  );


  not
  g778
  (
    n808,
    n559
  );


  not
  g779
  (
    n899,
    n577
  );


  not
  g780
  (
    n756,
    n556
  );


  not
  g781
  (
    n1152,
    n652
  );


  not
  g782
  (
    n794,
    n581
  );


  not
  g783
  (
    n717,
    n613
  );


  buf
  g784
  (
    n1183,
    n649
  );


  not
  g785
  (
    n1192,
    n609
  );


  buf
  g786
  (
    n956,
    n556
  );


  not
  g787
  (
    n852,
    n625
  );


  not
  g788
  (
    n1055,
    n573
  );


  buf
  g789
  (
    n730,
    n535
  );


  buf
  g790
  (
    n832,
    n580
  );


  not
  g791
  (
    KeyWire_0_36,
    n605
  );


  not
  g792
  (
    n1103,
    n593
  );


  buf
  g793
  (
    n1111,
    n598
  );


  not
  g794
  (
    n777,
    n623
  );


  not
  g795
  (
    n1082,
    n630
  );


  buf
  g796
  (
    n770,
    n600
  );


  not
  g797
  (
    n846,
    n648
  );


  buf
  g798
  (
    n900,
    n646
  );


  not
  g799
  (
    n1170,
    n624
  );


  buf
  g800
  (
    n960,
    n575
  );


  not
  g801
  (
    n930,
    n542
  );


  buf
  g802
  (
    n915,
    n550
  );


  not
  g803
  (
    n803,
    n603
  );


  buf
  g804
  (
    n753,
    n627
  );


  not
  g805
  (
    n876,
    n566
  );


  buf
  g806
  (
    n1198,
    n580
  );


  buf
  g807
  (
    n932,
    n579
  );


  buf
  g808
  (
    n754,
    n624
  );


  buf
  g809
  (
    n746,
    n643
  );


  not
  g810
  (
    n1182,
    n635
  );


  buf
  g811
  (
    n1065,
    n591
  );


  buf
  g812
  (
    n792,
    n605
  );


  not
  g813
  (
    n951,
    n538
  );


  buf
  g814
  (
    n924,
    n572
  );


  buf
  g815
  (
    n979,
    n515
  );


  buf
  g816
  (
    n864,
    n578
  );


  buf
  g817
  (
    n854,
    n622
  );


  buf
  g818
  (
    n740,
    n617
  );


  buf
  g819
  (
    n908,
    n585
  );


  not
  g820
  (
    n943,
    n568
  );


  not
  g821
  (
    n735,
    n588
  );


  buf
  g822
  (
    n1018,
    n584
  );


  buf
  g823
  (
    n749,
    n596
  );


  not
  g824
  (
    n775,
    n519
  );


  buf
  g825
  (
    n868,
    n646
  );


  not
  g826
  (
    n973,
    n608
  );


  buf
  g827
  (
    n1195,
    n611
  );


  buf
  g828
  (
    n1077,
    n612
  );


  not
  g829
  (
    n750,
    n534
  );


  buf
  g830
  (
    n830,
    n537
  );


  not
  g831
  (
    n1139,
    n424
  );


  buf
  g832
  (
    n1213,
    n537
  );


  buf
  g833
  (
    n804,
    n630
  );


  buf
  g834
  (
    n968,
    n614
  );


  not
  g835
  (
    n1022,
    n517
  );


  not
  g836
  (
    n940,
    n541
  );


  buf
  g837
  (
    n1070,
    n592
  );


  not
  g838
  (
    n1034,
    n595
  );


  not
  g839
  (
    n1133,
    n550
  );


  not
  g840
  (
    n950,
    n626
  );


  buf
  g841
  (
    n1127,
    n540
  );


  not
  g842
  (
    n1155,
    n596
  );


  not
  g843
  (
    n1088,
    n518
  );


  not
  g844
  (
    n1199,
    n570
  );


  not
  g845
  (
    n1140,
    n539
  );


  not
  g846
  (
    n981,
    n631
  );


  not
  g847
  (
    KeyWire_0_17,
    n555
  );


  not
  g848
  (
    n1004,
    n601
  );


  buf
  g849
  (
    n1010,
    n546
  );


  not
  g850
  (
    n765,
    n560
  );


  buf
  g851
  (
    n810,
    n569
  );


  not
  g852
  (
    n957,
    n585
  );


  not
  g853
  (
    n885,
    n625
  );


  not
  g854
  (
    n780,
    n557
  );


  not
  g855
  (
    KeyWire_0_57,
    n600
  );


  buf
  g856
  (
    n989,
    n637
  );


  not
  g857
  (
    n1016,
    n622
  );


  buf
  g858
  (
    n1179,
    n629
  );


  buf
  g859
  (
    n1025,
    n648
  );


  buf
  g860
  (
    n1105,
    n652
  );


  not
  g861
  (
    n1012,
    n645
  );


  buf
  g862
  (
    n1118,
    n588
  );


  buf
  g863
  (
    n1135,
    n611
  );


  buf
  g864
  (
    n1094,
    n629
  );


  not
  g865
  (
    n811,
    n650
  );


  buf
  g866
  (
    n1067,
    n516
  );


  not
  g867
  (
    n834,
    n538
  );


  buf
  g868
  (
    n1128,
    n630
  );


  buf
  g869
  (
    n1066,
    n641
  );


  not
  g870
  (
    n801,
    n608
  );


  buf
  g871
  (
    n716,
    n528
  );


  buf
  g872
  (
    n1148,
    n519
  );


  not
  g873
  (
    n1205,
    n539
  );


  not
  g874
  (
    n757,
    n529
  );


  not
  g875
  (
    n1172,
    n546
  );


  buf
  g876
  (
    n729,
    n562
  );


  not
  g877
  (
    n873,
    n635
  );


  buf
  g878
  (
    n1075,
    n591
  );


  buf
  g879
  (
    n1181,
    n603
  );


  buf
  g880
  (
    n813,
    n634
  );


  not
  g881
  (
    KeyWire_0_34,
    n621
  );


  not
  g882
  (
    n954,
    n533
  );


  not
  g883
  (
    n1026,
    n596
  );


  buf
  g884
  (
    KeyWire_0_1,
    n581
  );


  buf
  g885
  (
    n822,
    n638
  );


  not
  g886
  (
    n719,
    n623
  );


  buf
  g887
  (
    n1134,
    n588
  );


  buf
  g888
  (
    n1100,
    n542
  );


  not
  g889
  (
    n1084,
    n534
  );


  not
  g890
  (
    n1061,
    n632
  );


  not
  g891
  (
    n763,
    n580
  );


  not
  g892
  (
    KeyWire_0_31,
    n574
  );


  buf
  g893
  (
    n1149,
    n551
  );


  buf
  g894
  (
    n926,
    n554
  );


  not
  g895
  (
    n1024,
    n520
  );


  not
  g896
  (
    n844,
    n563
  );


  not
  g897
  (
    n1162,
    n593
  );


  not
  g898
  (
    n897,
    n540
  );


  not
  g899
  (
    n1000,
    n530
  );


  buf
  g900
  (
    n875,
    n584
  );


  buf
  g901
  (
    n1196,
    n555
  );


  buf
  g902
  (
    n962,
    n572
  );


  not
  g903
  (
    n1184,
    n599
  );


  buf
  g904
  (
    n904,
    n595
  );


  buf
  g905
  (
    n789,
    n578
  );


  buf
  g906
  (
    n845,
    n579
  );


  buf
  g907
  (
    n938,
    n563
  );


  not
  g908
  (
    n1151,
    n569
  );


  buf
  g909
  (
    n878,
    n638
  );


  not
  g910
  (
    n816,
    n607
  );


  not
  g911
  (
    n855,
    n632
  );


  buf
  g912
  (
    n1062,
    n565
  );


  buf
  g913
  (
    n1003,
    n582
  );


  buf
  g914
  (
    n1076,
    n573
  );


  buf
  g915
  (
    n783,
    n641
  );


  buf
  g916
  (
    n919,
    n572
  );


  not
  g917
  (
    n1020,
    n636
  );


  not
  g918
  (
    n861,
    n583
  );


  buf
  g919
  (
    n1164,
    n611
  );


  not
  g920
  (
    n1141,
    n584
  );


  buf
  g921
  (
    n994,
    n630
  );


  buf
  g922
  (
    n782,
    n602
  );


  buf
  g923
  (
    n764,
    n532
  );


  buf
  g924
  (
    n964,
    n623
  );


  buf
  g925
  (
    n825,
    n551
  );


  not
  g926
  (
    n991,
    n426
  );


  buf
  g927
  (
    n773,
    n574
  );


  not
  g928
  (
    n726,
    n633
  );


  not
  g929
  (
    n838,
    n638
  );


  not
  g930
  (
    n1087,
    n623
  );


  buf
  g931
  (
    KeyWire_0_51,
    n651
  );


  buf
  g932
  (
    n768,
    n590
  );


  not
  g933
  (
    n1040,
    n569
  );


  buf
  g934
  (
    n793,
    n533
  );


  not
  g935
  (
    n858,
    n553
  );


  not
  g936
  (
    n1005,
    n647
  );


  buf
  g937
  (
    n862,
    n629
  );


  buf
  g938
  (
    n896,
    n614
  );


  buf
  g939
  (
    n778,
    n535
  );


  not
  g940
  (
    n1114,
    n641
  );


  buf
  g941
  (
    n1042,
    n543
  );


  buf
  g942
  (
    n1098,
    n597
  );


  not
  g943
  (
    n922,
    n518
  );


  buf
  g944
  (
    n772,
    n518
  );


  buf
  g945
  (
    n851,
    n550
  );


  buf
  g946
  (
    n975,
    n566
  );


  buf
  g947
  (
    n1099,
    n562
  );


  not
  g948
  (
    n1130,
    n550
  );


  buf
  g949
  (
    n1059,
    n636
  );


  not
  g950
  (
    n721,
    n648
  );


  not
  g951
  (
    n1165,
    n640
  );


  buf
  g952
  (
    n781,
    n520
  );


  buf
  g953
  (
    n912,
    n639
  );


  not
  g954
  (
    n1060,
    n544
  );


  not
  g955
  (
    n1089,
    n571
  );


  not
  g956
  (
    n998,
    n589
  );


  buf
  g957
  (
    n1007,
    n620
  );


  not
  g958
  (
    n1116,
    n545
  );


  not
  g959
  (
    n929,
    n649
  );


  buf
  g960
  (
    n1129,
    n516
  );


  buf
  g961
  (
    n927,
    n618
  );


  not
  g962
  (
    n856,
    n531
  );


  not
  g963
  (
    n980,
    n626
  );


  not
  g964
  (
    n976,
    n598
  );


  not
  g965
  (
    n891,
    n577
  );


  buf
  g966
  (
    n784,
    n637
  );


  buf
  g967
  (
    n888,
    n645
  );


  buf
  g968
  (
    n923,
    n645
  );


  not
  g969
  (
    n907,
    n606
  );


  not
  g970
  (
    KeyWire_0_63,
    n616
  );


  buf
  g971
  (
    n1201,
    n621
  );


  not
  g972
  (
    n1071,
    n570
  );


  buf
  g973
  (
    n1092,
    n610
  );


  buf
  g974
  (
    n1123,
    n635
  );


  not
  g975
  (
    n921,
    n600
  );


  buf
  g976
  (
    n910,
    n546
  );


  not
  g977
  (
    n863,
    n631
  );


  buf
  g978
  (
    n831,
    n540
  );


  not
  g979
  (
    n931,
    n647
  );


  not
  g980
  (
    n800,
    n576
  );


  buf
  g981
  (
    n995,
    n547
  );


  not
  g982
  (
    n1036,
    n541
  );


  buf
  g983
  (
    n766,
    n647
  );


  not
  g984
  (
    n737,
    n604
  );


  not
  g985
  (
    n1091,
    n618
  );


  not
  g986
  (
    KeyWire_0_55,
    n575
  );


  buf
  g987
  (
    n1080,
    n607
  );


  buf
  g988
  (
    n879,
    n649
  );


  buf
  g989
  (
    n1014,
    n599
  );


  not
  g990
  (
    n1166,
    n589
  );


  not
  g991
  (
    n842,
    n528
  );


  buf
  g992
  (
    n829,
    n568
  );


  buf
  g993
  (
    n1150,
    n629
  );


  not
  g994
  (
    n724,
    n557
  );


  not
  g995
  (
    n894,
    n567
  );


  buf
  g996
  (
    n751,
    n428
  );


  buf
  g997
  (
    n1053,
    n571
  );


  not
  g998
  (
    n1101,
    n555
  );


  not
  g999
  (
    n733,
    n639
  );


  buf
  g1000
  (
    n1202,
    n576
  );


  buf
  g1001
  (
    n997,
    n642
  );


  buf
  g1002
  (
    n1145,
    n541
  );


  not
  g1003
  (
    n1011,
    n628
  );


  buf
  g1004
  (
    n1115,
    n535
  );


  not
  g1005
  (
    n959,
    n599
  );


  not
  g1006
  (
    n790,
    n548
  );


  buf
  g1007
  (
    n993,
    n564
  );


  buf
  g1008
  (
    n1168,
    n637
  );


  not
  g1009
  (
    n1009,
    n636
  );


  buf
  g1010
  (
    n971,
    n601
  );


  buf
  g1011
  (
    n1161,
    n549
  );


  not
  g1012
  (
    n747,
    n559
  );


  buf
  g1013
  (
    n1085,
    n566
  );


  buf
  g1014
  (
    n988,
    n613
  );


  buf
  g1015
  (
    n1194,
    n626
  );


  not
  g1016
  (
    n1163,
    n604
  );


  not
  g1017
  (
    n1121,
    n537
  );


  buf
  g1018
  (
    n867,
    n554
  );


  not
  g1019
  (
    n961,
    n589
  );


  not
  g1020
  (
    n881,
    n634
  );


  not
  g1021
  (
    KeyWire_0_54,
    n520
  );


  not
  g1022
  (
    n1047,
    n532
  );


  not
  g1023
  (
    n987,
    n530
  );


  not
  g1024
  (
    n815,
    n537
  );


  not
  g1025
  (
    n934,
    n547
  );


  not
  g1026
  (
    n1144,
    n561
  );


  buf
  g1027
  (
    n732,
    n552
  );


  buf
  g1028
  (
    n1019,
    n618
  );


  not
  g1029
  (
    n944,
    n595
  );


  not
  g1030
  (
    n1204,
    n650
  );


  not
  g1031
  (
    n1107,
    n636
  );


  not
  g1032
  (
    n759,
    n582
  );


  not
  g1033
  (
    n1008,
    n635
  );


  buf
  g1034
  (
    n1033,
    n545
  );


  buf
  g1035
  (
    n1208,
    n609
  );


  buf
  g1036
  (
    n935,
    n631
  );


  buf
  g1037
  (
    n911,
    n547
  );


  not
  g1038
  (
    n1054,
    n651
  );


  not
  g1039
  (
    n1197,
    n619
  );


  not
  g1040
  (
    n723,
    n548
  );


  buf
  g1041
  (
    n1002,
    n613
  );


  not
  g1042
  (
    n739,
    n648
  );


  not
  g1043
  (
    n1058,
    n628
  );


  buf
  g1044
  (
    n996,
    n533
  );


  buf
  g1045
  (
    n762,
    n515
  );


  not
  g1046
  (
    n906,
    n584
  );


  buf
  g1047
  (
    n1159,
    n517
  );


  not
  g1048
  (
    n1073,
    n615
  );


  not
  g1049
  (
    n1193,
    n606
  );


  not
  g1050
  (
    n1108,
    n618
  );


  buf
  g1051
  (
    n1039,
    n587
  );


  not
  g1052
  (
    n1029,
    n546
  );


  buf
  g1053
  (
    n1186,
    n642
  );


  buf
  g1054
  (
    n1189,
    n641
  );


  not
  g1055
  (
    n1057,
    n548
  );


  not
  g1056
  (
    n1086,
    n643
  );


  buf
  g1057
  (
    n1124,
    n567
  );


  not
  g1058
  (
    n866,
    n620
  );


  not
  g1059
  (
    n839,
    n612
  );


  not
  g1060
  (
    n1079,
    n633
  );


  not
  g1061
  (
    n952,
    n611
  );


  not
  g1062
  (
    n895,
    n551
  );


  buf
  g1063
  (
    n745,
    n646
  );


  not
  g1064
  (
    n916,
    n564
  );


  buf
  g1065
  (
    n752,
    n559
  );


  not
  g1066
  (
    n870,
    n529
  );


  not
  g1067
  (
    n798,
    n644
  );


  buf
  g1068
  (
    n901,
    n616
  );


  buf
  g1069
  (
    n872,
    n539
  );


  buf
  g1070
  (
    n1021,
    n592
  );


  not
  g1071
  (
    n761,
    n585
  );


  not
  g1072
  (
    n889,
    n569
  );


  not
  g1073
  (
    n1143,
    n594
  );


  buf
  g1074
  (
    n953,
    n517
  );


  not
  g1075
  (
    n843,
    n556
  );


  buf
  g1076
  (
    n1132,
    n528
  );


  not
  g1077
  (
    n795,
    n633
  );


  not
  g1078
  (
    n1097,
    n591
  );


  not
  g1079
  (
    n1045,
    n560
  );


  not
  g1080
  (
    n887,
    n640
  );


  not
  g1081
  (
    n882,
    n590
  );


  buf
  g1082
  (
    n760,
    n538
  );


  not
  g1083
  (
    n1113,
    n612
  );


  not
  g1084
  (
    n748,
    n608
  );


  buf
  g1085
  (
    n918,
    n542
  );


  buf
  g1086
  (
    n827,
    n632
  );


  buf
  g1087
  (
    n925,
    n551
  );


  not
  g1088
  (
    n920,
    n586
  );


  buf
  g1089
  (
    n1188,
    n628
  );


  not
  g1090
  (
    n1083,
    n530
  );


  buf
  g1091
  (
    n1006,
    n614
  );


  not
  g1092
  (
    n990,
    n553
  );


  buf
  g1093
  (
    n1131,
    n531
  );


  not
  g1094
  (
    n1173,
    n625
  );


  buf
  g1095
  (
    n1169,
    n593
  );


  buf
  g1096
  (
    n945,
    n565
  );


  buf
  g1097
  (
    n743,
    n616
  );


  buf
  g1098
  (
    n1154,
    n617
  );


  not
  g1099
  (
    n983,
    n619
  );


  buf
  g1100
  (
    n1122,
    n543
  );


  not
  g1101
  (
    n809,
    n536
  );


  buf
  g1102
  (
    n1137,
    n516
  );


  not
  g1103
  (
    n974,
    n520
  );


  not
  g1104
  (
    n1051,
    n573
  );


  not
  g1105
  (
    n718,
    n570
  );


  buf
  g1106
  (
    n819,
    n601
  );


  not
  g1107
  (
    n1064,
    n542
  );


  buf
  g1108
  (
    n1035,
    n613
  );


  not
  g1109
  (
    n1046,
    n586
  );


  not
  g1110
  (
    n742,
    n563
  );


  buf
  g1111
  (
    n767,
    n643
  );


  not
  g1112
  (
    n1125,
    n531
  );


  not
  g1113
  (
    n1028,
    n519
  );


  buf
  g1114
  (
    n837,
    n619
  );


  buf
  g1115
  (
    n836,
    n552
  );


  buf
  g1116
  (
    n1157,
    n624
  );


  not
  g1117
  (
    n982,
    n531
  );


  buf
  g1118
  (
    n758,
    n604
  );


  buf
  g1119
  (
    n1013,
    n651
  );


  not
  g1120
  (
    n1048,
    n582
  );


  buf
  g1121
  (
    n884,
    n566
  );


  not
  g1122
  (
    n970,
    n559
  );


  buf
  g1123
  (
    KeyWire_0_25,
    n604
  );


  not
  g1124
  (
    n1001,
    n573
  );


  not
  g1125
  (
    n814,
    n429
  );


  buf
  g1126
  (
    n826,
    n554
  );


  not
  g1127
  (
    n853,
    n583
  );


  buf
  g1128
  (
    n1203,
    n517
  );


  not
  g1129
  (
    n941,
    n554
  );


  not
  g1130
  (
    n776,
    n617
  );


  buf
  g1131
  (
    n909,
    n543
  );


  buf
  g1132
  (
    n1102,
    n600
  );


  not
  g1133
  (
    n860,
    n575
  );


  not
  g1134
  (
    n744,
    n555
  );


  not
  g1135
  (
    n807,
    n532
  );


  not
  g1136
  (
    n1191,
    n644
  );


  buf
  g1137
  (
    n802,
    n640
  );


  buf
  g1138
  (
    n917,
    n590
  );


  buf
  g1139
  (
    n1178,
    n582
  );


  buf
  g1140
  (
    n928,
    n627
  );


  buf
  g1141
  (
    n841,
    n567
  );


  buf
  g1142
  (
    n821,
    n620
  );


  buf
  g1143
  (
    KeyWire_0_53,
    n608
  );


  not
  g1144
  (
    n892,
    n617
  );


  buf
  g1145
  (
    n1052,
    n631
  );


  not
  g1146
  (
    n947,
    n633
  );


  buf
  g1147
  (
    n1043,
    n603
  );


  buf
  g1148
  (
    n785,
    n581
  );


  not
  g1149
  (
    n1207,
    n642
  );


  buf
  g1150
  (
    n942,
    n583
  );


  buf
  g1151
  (
    n1078,
    n597
  );


  buf
  g1152
  (
    n848,
    n547
  );


  buf
  g1153
  (
    n847,
    n539
  );


  buf
  g1154
  (
    n1136,
    n574
  );


  buf
  g1155
  (
    n786,
    n572
  );


  not
  g1156
  (
    n1187,
    n647
  );


  not
  g1157
  (
    n1175,
    n644
  );


  not
  g1158
  (
    n722,
    n602
  );


  not
  g1159
  (
    n1142,
    n544
  );


  not
  g1160
  (
    n1044,
    n528
  );


  buf
  g1161
  (
    KeyWire_0_29,
    n592
  );


  not
  g1162
  (
    n1160,
    n558
  );


  buf
  g1163
  (
    n1096,
    n592
  );


  not
  g1164
  (
    n779,
    n577
  );


  buf
  g1165
  (
    n1063,
    n577
  );


  not
  g1166
  (
    n805,
    n628
  );


  not
  g1167
  (
    n865,
    n515
  );


  buf
  g1168
  (
    n806,
    n534
  );


  buf
  g1169
  (
    n812,
    n561
  );


  buf
  g1170
  (
    n1069,
    n568
  );


  not
  g1171
  (
    n1049,
    n601
  );


  not
  g1172
  (
    n797,
    n627
  );


  buf
  g1173
  (
    n963,
    n536
  );


  not
  g1174
  (
    n939,
    n644
  );


  nand
  g1175
  (
    n933,
    n598,
    n651,
    n640,
    n610
  );


  xnor
  g1176
  (
    n787,
    n548,
    n518,
    n533,
    n545
  );


  xor
  g1177
  (
    n1093,
    n425,
    n625,
    n626,
    n580
  );


  nand
  g1178
  (
    n1023,
    n610,
    n564,
    n602,
    n597
  );


  and
  g1179
  (
    n986,
    n536,
    n596,
    n545,
    n544
  );


  or
  g1180
  (
    n1190,
    n549,
    n587,
    n565,
    n638
  );


  nor
  g1181
  (
    n1038,
    n560,
    n558,
    n586,
    n427
  );


  xnor
  g1182
  (
    n948,
    n634,
    n615,
    n534,
    n642
  );


  and
  g1183
  (
    n886,
    n588,
    n535,
    n549,
    n620
  );


  xor
  g1184
  (
    n1027,
    n552,
    n634,
    n581,
    n557
  );


  xnor
  g1185
  (
    n1220,
    n523,
    n524,
    n526,
    n135
  );


  xor
  g1186
  (
    n1218,
    n132,
    n130,
    n751,
    n524
  );


  or
  g1187
  (
    n1233,
    n762,
    n763,
    n290,
    n742
  );


  or
  g1188
  (
    n1216,
    n526,
    n733,
    n522
  );


  or
  g1189
  (
    n1219,
    n527,
    n757,
    n130,
    n737
  );


  or
  g1190
  (
    n1227,
    n134,
    n449,
    n524
  );


  xor
  g1191
  (
    n1221,
    n131,
    n740,
    n765,
    n133
  );


  nand
  g1192
  (
    n1229,
    n134,
    n133,
    n135,
    n130
  );


  and
  g1193
  (
    n1228,
    n525,
    n134,
    n723,
    n749
  );


  and
  g1194
  (
    n1226,
    n133,
    n761,
    n522,
    n759
  );


  and
  g1195
  (
    n1222,
    n132,
    n731,
    n722,
    n131
  );


  nor
  g1196
  (
    n1234,
    n131,
    n734,
    n526,
    n750
  );


  nand
  g1197
  (
    n1231,
    n739,
    n527,
    n131,
    n735
  );


  xnor
  g1198
  (
    n1239,
    n132,
    n716,
    n738,
    n525
  );


  or
  g1199
  (
    n1225,
    n288,
    n728,
    n521,
    n717
  );


  nor
  g1200
  (
    n1235,
    n764,
    n758,
    n523,
    n133
  );


  xnor
  g1201
  (
    n1230,
    n525,
    n727,
    n135,
    n755
  );


  or
  g1202
  (
    n1240,
    n525,
    n744,
    n136,
    n732
  );


  nor
  g1203
  (
    n1236,
    n719,
    n736,
    n521,
    n746
  );


  or
  g1204
  (
    n1215,
    n526,
    n134,
    n721,
    n725
  );


  xor
  g1205
  (
    n1214,
    n760,
    n747,
    n754,
    n523
  );


  xor
  g1206
  (
    n1237,
    n726,
    n741,
    n289,
    n521
  );


  xor
  g1207
  (
    n1224,
    n724,
    n523,
    n522,
    n524
  );


  xnor
  g1208
  (
    n1223,
    n753,
    n521,
    n729,
    n743
  );


  nor
  g1209
  (
    n1232,
    n718,
    n527,
    n748,
    n730
  );


  nor
  g1210
  (
    n1238,
    n745,
    n720,
    n132,
    n136
  );


  nor
  g1211
  (
    n1217,
    n752,
    n135,
    n756,
    n527
  );


  buf
  g1212
  (
    n1259,
    n1222
  );


  buf
  g1213
  (
    n1244,
    n1239
  );


  not
  g1214
  (
    n1250,
    n1234
  );


  buf
  g1215
  (
    n1266,
    n1235
  );


  not
  g1216
  (
    n1255,
    n1221
  );


  not
  g1217
  (
    n1242,
    n1228
  );


  not
  g1218
  (
    n1260,
    n1216
  );


  not
  g1219
  (
    n1247,
    n1238
  );


  not
  g1220
  (
    n1262,
    n1225
  );


  not
  g1221
  (
    n1249,
    n1231
  );


  buf
  g1222
  (
    n1248,
    n1226
  );


  buf
  g1223
  (
    n1256,
    n1223
  );


  not
  g1224
  (
    n1251,
    n1217
  );


  buf
  g1225
  (
    n1252,
    n1230
  );


  not
  g1226
  (
    n1245,
    n1215
  );


  buf
  g1227
  (
    n1264,
    n1224
  );


  not
  g1228
  (
    n1263,
    n1232
  );


  not
  g1229
  (
    n1253,
    n1220
  );


  not
  g1230
  (
    n1246,
    n1237
  );


  not
  g1231
  (
    n1243,
    n1219
  );


  buf
  g1232
  (
    n1261,
    n1229
  );


  not
  g1233
  (
    n1254,
    n1227
  );


  not
  g1234
  (
    n1265,
    n1236
  );


  buf
  g1235
  (
    n1258,
    n1233
  );


  not
  g1236
  (
    n1257,
    n1218
  );


  buf
  g1237
  (
    n1241,
    n1214
  );


  nand
  g1238
  (
    n1292,
    n679,
    n1261,
    n341,
    n684
  );


  xnor
  g1239
  (
    n1273,
    n342,
    n672,
    n701,
    n1263
  );


  and
  g1240
  (
    n1369,
    n713,
    n1240,
    n670,
    n1261
  );


  nor
  g1241
  (
    KeyWire_0_47,
    n1246,
    n679,
    n308,
    n674
  );


  nand
  g1242
  (
    n1353,
    n672,
    n712,
    n711,
    n675
  );


  xor
  g1243
  (
    n1346,
    n1245,
    n666,
    n677
  );


  or
  g1244
  (
    n1311,
    n699,
    n313,
    n694
  );


  or
  g1245
  (
    n1270,
    n673,
    n1257,
    n671,
    n325
  );


  xor
  g1246
  (
    n1367,
    n660,
    n673,
    n696,
    n655
  );


  or
  g1247
  (
    n1359,
    n1249,
    n660,
    n709,
    n1258
  );


  nor
  g1248
  (
    n1336,
    n1254,
    n712,
    n319,
    n690
  );


  xnor
  g1249
  (
    n1285,
    n301,
    n1264,
    n701,
    n320
  );


  nor
  g1250
  (
    n1325,
    n661,
    n682,
    n1255,
    n1257
  );


  and
  g1251
  (
    n1345,
    n335,
    n661,
    n1266
  );


  nor
  g1252
  (
    n1291,
    n654,
    n1241,
    n693,
    n1259
  );


  nand
  g1253
  (
    n1364,
    n685,
    n314,
    n1245,
    n703
  );


  nand
  g1254
  (
    n1269,
    n681,
    n298,
    n661,
    n696
  );


  xnor
  g1255
  (
    n1271,
    n324,
    n704,
    n1253,
    n659
  );


  nand
  g1256
  (
    n1334,
    n693,
    n653,
    n698,
    n687
  );


  xor
  g1257
  (
    n1338,
    n692,
    n681,
    n701,
    n714
  );


  or
  g1258
  (
    n1343,
    n692,
    n339,
    n676,
    n671
  );


  and
  g1259
  (
    n1355,
    n691,
    n292,
    n334,
    n681
  );


  nor
  g1260
  (
    n1289,
    n682,
    n677,
    n710,
    n687
  );


  xnor
  g1261
  (
    n1272,
    n658,
    n703,
    n1265,
    n340
  );


  or
  g1262
  (
    n1316,
    n1244,
    n713,
    n1264,
    n688
  );


  xor
  g1263
  (
    n1349,
    n665,
    n1258,
    n674,
    n28
  );


  nand
  g1264
  (
    n1288,
    n309,
    n708,
    n1253,
    n709
  );


  nand
  g1265
  (
    n1278,
    n704,
    n697,
    n690,
    n682
  );


  and
  g1266
  (
    n1276,
    n700,
    n665,
    n663,
    n697
  );


  xnor
  g1267
  (
    n1313,
    n1251,
    n669,
    n1253,
    n1241
  );


  xor
  g1268
  (
    n1333,
    n300,
    n663,
    n311,
    n695
  );


  xnor
  g1269
  (
    KeyWire_0_13,
    n303,
    n674,
    n667,
    n665
  );


  and
  g1270
  (
    n1279,
    n654,
    n696,
    n714,
    n706
  );


  nand
  g1271
  (
    n1361,
    n333,
    n1244,
    n295,
    n699
  );


  and
  g1272
  (
    n1296,
    n328,
    n666,
    n1250,
    n701
  );


  and
  g1273
  (
    n1282,
    n1248,
    n1258,
    n1257,
    n662
  );


  xor
  g1274
  (
    n1298,
    n700,
    n707,
    n1258,
    n318
  );


  or
  g1275
  (
    n1358,
    n1251,
    n711,
    n679,
    n659
  );


  nand
  g1276
  (
    n1331,
    n307,
    n1250,
    n705,
    n1249
  );


  or
  g1277
  (
    n1294,
    n655,
    n1247,
    n1249,
    n691
  );


  nor
  g1278
  (
    n1281,
    n293,
    n1259,
    n1263,
    n680
  );


  nand
  g1279
  (
    n1284,
    n677,
    n695,
    n1260,
    n697
  );


  xnor
  g1280
  (
    n1299,
    n1260,
    n710,
    n698,
    n655
  );


  nand
  g1281
  (
    n1312,
    n667,
    n703,
    n316,
    n655
  );


  nand
  g1282
  (
    n1307,
    n304,
    n692,
    n689,
    n1244
  );


  nor
  g1283
  (
    n1322,
    n1250,
    n658,
    n654,
    n662
  );


  or
  g1284
  (
    n1287,
    n666,
    n689,
    n706,
    n1242
  );


  xnor
  g1285
  (
    n1295,
    n691,
    n688,
    n656,
    n698
  );


  xor
  g1286
  (
    n1354,
    n1246,
    n686,
    n669,
    n678
  );


  xnor
  g1287
  (
    n1362,
    n667,
    n670,
    n1252,
    n685
  );


  xor
  g1288
  (
    n1357,
    n1260,
    n1256,
    n329,
    n705
  );


  nor
  g1289
  (
    n1317,
    n688,
    n657,
    n653,
    n683
  );


  nor
  g1290
  (
    n1340,
    n657,
    n708,
    n331,
    n1256
  );


  and
  g1291
  (
    n1348,
    n699,
    n687,
    n681,
    n682
  );


  nor
  g1292
  (
    n1297,
    n707,
    n664,
    n299,
    n653
  );


  or
  g1293
  (
    n1293,
    n706,
    n1265,
    n332,
    n661
  );


  and
  g1294
  (
    n1302,
    n291,
    n1262,
    n705,
    n715
  );


  nor
  g1295
  (
    n1344,
    n1262,
    n668,
    n712,
    n1259
  );


  nor
  g1296
  (
    n1286,
    n1245,
    n699,
    n703,
    n1257
  );


  or
  g1297
  (
    n1309,
    n664,
    n1255,
    n698,
    n695
  );


  or
  g1298
  (
    n1310,
    n326,
    n678,
    n317,
    n652
  );


  xnor
  g1299
  (
    n1306,
    n697,
    n695,
    n28,
    n336
  );


  and
  g1300
  (
    n1356,
    n312,
    n659,
    n338
  );


  nand
  g1301
  (
    KeyWire_0_30,
    n1262,
    n664,
    n1242,
    n297
  );


  nor
  g1302
  (
    n1341,
    n668,
    n1263,
    n708,
    n1255
  );


  xor
  g1303
  (
    n1352,
    n679,
    n710,
    n1248,
    n675
  );


  and
  g1304
  (
    n1308,
    n715,
    n305,
    n686,
    n678
  );


  xor
  g1305
  (
    n1335,
    n669,
    n1266,
    n323,
    n687
  );


  and
  g1306
  (
    n1280,
    n330,
    n1244,
    n675,
    n676
  );


  xor
  g1307
  (
    n1319,
    n662,
    n702,
    n1247,
    n1250
  );


  and
  g1308
  (
    n1360,
    n688,
    n1243,
    n710,
    n337
  );


  or
  g1309
  (
    KeyWire_0_14,
    n656,
    n702,
    n1249,
    n707
  );


  nand
  g1310
  (
    KeyWire_0_46,
    n1251,
    n660,
    n306,
    n322
  );


  and
  g1311
  (
    n1283,
    n674,
    n1254,
    n28,
    n671
  );


  nand
  g1312
  (
    n1368,
    n684,
    n684,
    n671,
    n310
  );


  and
  g1313
  (
    KeyWire_0_37,
    n1246,
    n693,
    n672,
    n680
  );


  and
  g1314
  (
    n1324,
    n1251,
    n700,
    n680,
    n1248
  );


  nor
  g1315
  (
    n1300,
    n668,
    n704,
    n702,
    n1243
  );


  and
  g1316
  (
    n1274,
    n657,
    n1264,
    n1246,
    n673
  );


  and
  g1317
  (
    n1366,
    n1247,
    n653,
    n1261,
    n676
  );


  nand
  g1318
  (
    n1275,
    n1262,
    n1248,
    n1265,
    n663
  );


  nand
  g1319
  (
    KeyWire_0_27,
    n700,
    n712,
    n1243,
    n702
  );


  xnor
  g1320
  (
    n1339,
    n680,
    n693,
    n656,
    n1243
  );


  xnor
  g1321
  (
    n1320,
    n665,
    n690,
    n705,
    n714
  );


  nor
  g1322
  (
    n1304,
    n1254,
    n321,
    n709,
    n683
  );


  xor
  g1323
  (
    n1350,
    n684,
    n711,
    n667,
    n1259
  );


  xnor
  g1324
  (
    n1318,
    n668,
    n709,
    n1254,
    n666
  );


  or
  g1325
  (
    n1330,
    n711,
    n686,
    n670,
    n302
  );


  or
  g1326
  (
    n1370,
    n690,
    n654,
    n1264,
    n1241
  );


  nand
  g1327
  (
    n1327,
    n715,
    n696,
    n675,
    n714
  );


  nand
  g1328
  (
    n1268,
    n706,
    n686,
    n672,
    n296
  );


  xnor
  g1329
  (
    n1326,
    n1263,
    n658,
    n1265,
    n685
  );


  nand
  g1330
  (
    n1351,
    n315,
    n691,
    n707,
    n663
  );


  xor
  g1331
  (
    n1315,
    n673,
    n343,
    n1241,
    n327
  );


  nand
  g1332
  (
    KeyWire_0_58,
    n1260,
    n656,
    n657,
    n658
  );


  or
  g1333
  (
    n1301,
    n689,
    n669,
    n683,
    n692
  );


  xor
  g1334
  (
    n1365,
    n662,
    n694,
    n1252,
    n704
  );


  and
  g1335
  (
    n1329,
    n294,
    n1256,
    n664,
    n713
  );


  xor
  g1336
  (
    n1347,
    n670,
    n678,
    n1266,
    n676
  );


  xnor
  g1337
  (
    n1305,
    n1242,
    n1261,
    n28,
    n685
  );


  and
  g1338
  (
    n1277,
    n1252,
    n708,
    n715,
    n1247
  );


  nor
  g1339
  (
    n1332,
    n652,
    n1245,
    n694,
    n683
  );


  nor
  g1340
  (
    n1363,
    n689,
    n1256,
    n713,
    n660
  );


  or
  g1341
  (
    n1321,
    n1242,
    n1255,
    n1252,
    n1253
  );


  or
  g1342
  (
    n1471,
    n1201,
    n799,
    n1204,
    n949
  );


  nor
  g1343
  (
    n1483,
    n844,
    n981,
    n1197,
    n936
  );


  nand
  g1344
  (
    n1500,
    n930,
    n1170,
    n1360,
    n1366
  );


  xnor
  g1345
  (
    n1433,
    n1156,
    n1345,
    n1179,
    n958
  );


  or
  g1346
  (
    n1443,
    n1134,
    n1370,
    n854,
    n1068
  );


  and
  g1347
  (
    n1518,
    n1369,
    n1166,
    n1308,
    n1009
  );


  xor
  g1348
  (
    n1474,
    n976,
    n778,
    n1290,
    n1034
  );


  xnor
  g1349
  (
    n1445,
    n1362,
    n870,
    n873,
    n983
  );


  nor
  g1350
  (
    n1409,
    n1368,
    n1295,
    n1074,
    n1181
  );


  nor
  g1351
  (
    n1455,
    n1312,
    n1362,
    n892,
    n886
  );


  or
  g1352
  (
    n1489,
    n1305,
    n1280,
    n1106,
    n1046
  );


  or
  g1353
  (
    n1478,
    n1357,
    n1111,
    n1339,
    n928
  );


  nor
  g1354
  (
    n1501,
    n1355,
    n1105,
    n797,
    n1103
  );


  nand
  g1355
  (
    n1431,
    n1118,
    n902,
    n1015,
    n826
  );


  or
  g1356
  (
    n1397,
    n990,
    n1272,
    n1365,
    n1340
  );


  xnor
  g1357
  (
    n1454,
    n1017,
    n1160,
    n1366,
    n1126
  );


  nand
  g1358
  (
    n1467,
    n1083,
    n1279,
    n1014,
    n1152
  );


  nor
  g1359
  (
    n1391,
    n1104,
    n1155,
    n1064,
    n859
  );


  xor
  g1360
  (
    n1402,
    n1069,
    n1012,
    n889,
    n787
  );


  xnor
  g1361
  (
    n1504,
    n954,
    n950,
    n1367,
    n777
  );


  nand
  g1362
  (
    n1435,
    n987,
    n1030,
    n1063,
    n841
  );


  xor
  g1363
  (
    n1516,
    n798,
    n1072,
    n966,
    n1333
  );


  or
  g1364
  (
    n1480,
    n1169,
    n1049,
    n875,
    n1370
  );


  nand
  g1365
  (
    n1487,
    n977,
    n1282,
    n776,
    n893
  );


  nor
  g1366
  (
    n1459,
    n1045,
    n957,
    n1291,
    n1041
  );


  xnor
  g1367
  (
    n1401,
    n1050,
    n1060,
    n1193,
    n1164
  );


  nand
  g1368
  (
    n1458,
    n807,
    n845,
    n1329,
    n1309
  );


  xnor
  g1369
  (
    n1515,
    n1327,
    n1143,
    n908,
    n786
  );


  and
  g1370
  (
    n1441,
    n1306,
    n1316,
    n964,
    n1191
  );


  and
  g1371
  (
    n1436,
    n931,
    n911,
    n1357,
    n866
  );


  nor
  g1372
  (
    n1372,
    n894,
    n1269,
    n1363,
    n785
  );


  nor
  g1373
  (
    n1451,
    n992,
    n1313,
    n774,
    n945
  );


  xnor
  g1374
  (
    n1395,
    n1149,
    n1205,
    n944,
    n1203
  );


  or
  g1375
  (
    n1492,
    n927,
    n802,
    n1213,
    n1364
  );


  xnor
  g1376
  (
    KeyWire_0_40,
    n960,
    n1370,
    n1325,
    n1328
  );


  or
  g1377
  (
    n1385,
    n874,
    n948,
    n923,
    n1364
  );


  or
  g1378
  (
    n1374,
    n968,
    n1359,
    n1366,
    n1056
  );


  or
  g1379
  (
    n1465,
    n813,
    n1349,
    n1032,
    n1367
  );


  nand
  g1380
  (
    n1371,
    n1212,
    n932,
    n1348,
    n1040
  );


  xor
  g1381
  (
    n1425,
    n924,
    n1292,
    n1358,
    n1035
  );


  and
  g1382
  (
    n1380,
    n1359,
    n1110,
    n1135,
    n910
  );


  nor
  g1383
  (
    n1427,
    n926,
    n1115,
    n898,
    n1132
  );


  or
  g1384
  (
    n1475,
    n1007,
    n836,
    n1289,
    n834
  );


  nor
  g1385
  (
    n1393,
    n955,
    n862,
    n1354,
    n1186
  );


  nor
  g1386
  (
    n1411,
    n851,
    n814,
    n1195,
    n793
  );


  nor
  g1387
  (
    n1508,
    n888,
    n909,
    n1303,
    n804
  );


  nor
  g1388
  (
    n1396,
    n1127,
    n962,
    n1028,
    n1341
  );


  or
  g1389
  (
    n1462,
    n1097,
    n1178,
    n877,
    n880
  );


  and
  g1390
  (
    n1509,
    n1315,
    n1057,
    n779,
    n1016
  );


  nand
  g1391
  (
    n1498,
    n1018,
    n991,
    n1274,
    n801
  );


  nand
  g1392
  (
    n1426,
    n1073,
    n1076,
    n789,
    n1116
  );


  nor
  g1393
  (
    n1511,
    n806,
    n878,
    n794,
    n946
  );


  nand
  g1394
  (
    n1408,
    n1002,
    n969,
    n1273,
    n1137
  );


  and
  g1395
  (
    n1449,
    n891,
    n1054,
    n833,
    n1140
  );


  or
  g1396
  (
    n1400,
    n795,
    n1368,
    n1285,
    n772
  );


  xnor
  g1397
  (
    n1382,
    n1102,
    n1095,
    n1369,
    n1337
  );


  and
  g1398
  (
    n1442,
    n1130,
    n846,
    n855,
    n1188
  );


  or
  g1399
  (
    n1488,
    n1363,
    n984,
    n1157,
    n837
  );


  xor
  g1400
  (
    n1437,
    n982,
    n842,
    n1322,
    n1120
  );


  xnor
  g1401
  (
    n1407,
    n905,
    n1100,
    n1023,
    n769
  );


  nor
  g1402
  (
    n1406,
    n1336,
    n1001,
    n848,
    n975
  );


  nand
  g1403
  (
    n1482,
    n1350,
    n1361,
    n811,
    n1067
  );


  xor
  g1404
  (
    n1383,
    n1062,
    n1202,
    n1196,
    n1091
  );


  or
  g1405
  (
    n1505,
    n825,
    n967,
    n1065,
    n1321
  );


  nor
  g1406
  (
    n1484,
    n1358,
    n1154,
    n879,
    n912
  );


  xnor
  g1407
  (
    n1430,
    n784,
    n899,
    n867,
    n1112
  );


  or
  g1408
  (
    n1416,
    n1286,
    n824,
    n767,
    n768
  );


  nor
  g1409
  (
    n1376,
    n791,
    n895,
    n890,
    n869
  );


  nand
  g1410
  (
    n1404,
    n1047,
    n843,
    n1363,
    n1085
  );


  xor
  g1411
  (
    n1399,
    n850,
    n1267,
    n827,
    n1167
  );


  nand
  g1412
  (
    n1453,
    n1208,
    n871,
    n831,
    n939
  );


  nor
  g1413
  (
    n1387,
    n800,
    n1061,
    n1353,
    n817
  );


  and
  g1414
  (
    n1429,
    n1361,
    n857,
    n1369,
    n805
  );


  nand
  g1415
  (
    n1485,
    n1128,
    n904,
    n1319,
    n809
  );


  xnor
  g1416
  (
    n1461,
    n906,
    n1165,
    n788,
    n995
  );


  or
  g1417
  (
    n1452,
    n1362,
    n1194,
    n1346,
    n876
  );


  and
  g1418
  (
    n1506,
    n1058,
    n1101,
    n861,
    n1171
  );


  xnor
  g1419
  (
    n1428,
    n1136,
    n885,
    n1020,
    n1187
  );


  or
  g1420
  (
    n1418,
    n1000,
    n1129,
    n1144,
    n1200
  );


  or
  g1421
  (
    n1403,
    n1361,
    n921,
    n1172,
    n1184
  );


  nor
  g1422
  (
    n1513,
    n1005,
    n951,
    n942,
    n941
  );


  xor
  g1423
  (
    KeyWire_0_62,
    n1052,
    n770,
    n980,
    n1334
  );


  xnor
  g1424
  (
    n1493,
    n1352,
    n952,
    n1275,
    n883
  );


  nor
  g1425
  (
    n1450,
    n1192,
    n1367,
    n933,
    n934
  );


  nor
  g1426
  (
    n1519,
    n796,
    n865,
    n989,
    n1153
  );


  xor
  g1427
  (
    n1481,
    n1123,
    n1119,
    n972,
    n1356
  );


  xor
  g1428
  (
    n1517,
    n1029,
    n965,
    n1121,
    n1093
  );


  nor
  g1429
  (
    n1438,
    n849,
    n1199,
    n1010,
    n943
  );


  nand
  g1430
  (
    n1477,
    n1173,
    n988,
    n887,
    n1175
  );


  nor
  g1431
  (
    n1398,
    n1177,
    n1320,
    n1026,
    n136
  );


  or
  g1432
  (
    n1388,
    n821,
    n1365,
    n1107,
    n1099
  );


  or
  g1433
  (
    n1464,
    n925,
    n1365,
    n1311,
    n1211
  );


  xor
  g1434
  (
    n1394,
    n970,
    n1098,
    n986,
    n1369
  );


  xnor
  g1435
  (
    n1444,
    n1025,
    n1351,
    n929,
    n1019
  );


  xnor
  g1436
  (
    n1410,
    n922,
    n828,
    n1182,
    n997
  );


  xnor
  g1437
  (
    n1392,
    n1124,
    n1370,
    n1044,
    n1358
  );


  xnor
  g1438
  (
    n1384,
    n1158,
    n1298,
    n1162,
    n1139
  );


  nand
  g1439
  (
    n1432,
    n1190,
    n1168,
    n884,
    n820
  );


  nand
  g1440
  (
    n1494,
    n1027,
    n985,
    n1031,
    n1363
  );


  nor
  g1441
  (
    n1434,
    n915,
    n1036,
    n1344,
    n1090
  );


  and
  g1442
  (
    n1463,
    n1150,
    n1125,
    n782,
    n1011
  );


  nor
  g1443
  (
    n1486,
    n816,
    n832,
    n830,
    n1151
  );


  and
  g1444
  (
    n1381,
    n829,
    n1368,
    n1276,
    n1359
  );


  nand
  g1445
  (
    n1470,
    n783,
    n900,
    n1053,
    n1096
  );


  xnor
  g1446
  (
    n1497,
    n1006,
    n1357,
    n1084,
    n1210
  );


  xnor
  g1447
  (
    n1378,
    n1283,
    n1042,
    n1330,
    n1087
  );


  or
  g1448
  (
    n1468,
    n1180,
    n1287,
    n1066,
    n822
  );


  nor
  g1449
  (
    n1389,
    n973,
    n1021,
    n1078,
    n993
  );


  and
  g1450
  (
    n1476,
    n1302,
    n1176,
    n940,
    n882
  );


  and
  g1451
  (
    n1412,
    n1364,
    n1332,
    n1297,
    n999
  );


  and
  g1452
  (
    n1473,
    n1318,
    n1331,
    n1284,
    n766
  );


  or
  g1453
  (
    n1413,
    n938,
    n914,
    n1089,
    n818
  );


  or
  g1454
  (
    n1447,
    n918,
    n1314,
    n978,
    n1183
  );


  or
  g1455
  (
    n1507,
    n919,
    n916,
    n840,
    n1024
  );


  or
  g1456
  (
    n1417,
    n1304,
    n1360,
    n1113,
    n1043
  );


  nor
  g1457
  (
    n1472,
    n907,
    n1147,
    n1075,
    n864
  );


  or
  g1458
  (
    n1424,
    n838,
    n994,
    n1361,
    n917
  );


  nand
  g1459
  (
    n1420,
    n1310,
    n863,
    n1335,
    n1270
  );


  xor
  g1460
  (
    n1510,
    n773,
    n856,
    n1059,
    n1080
  );


  nand
  g1461
  (
    n1422,
    n1299,
    n1355,
    n1206,
    n1003
  );


  nor
  g1462
  (
    n1512,
    n136,
    n881,
    n860,
    n1185
  );


  or
  g1463
  (
    n1419,
    n1296,
    n1114,
    n1109,
    n872
  );


  or
  g1464
  (
    n1496,
    n790,
    n1008,
    n819,
    n1338
  );


  or
  g1465
  (
    n1499,
    n897,
    n1022,
    n812,
    n1277
  );


  nor
  g1466
  (
    n1377,
    n935,
    n1038,
    n1356,
    n1081
  );


  nor
  g1467
  (
    n1520,
    n1138,
    n1288,
    n1324,
    n1174
  );


  and
  g1468
  (
    n1375,
    n971,
    n1071,
    n1356,
    n1360
  );


  xor
  g1469
  (
    n1514,
    n1161,
    n771,
    n961,
    n1300
  );


  xnor
  g1470
  (
    n1390,
    n1281,
    n901,
    n959,
    n1198
  );


  nor
  g1471
  (
    n1448,
    n853,
    n1077,
    n1189,
    n1117
  );


  and
  g1472
  (
    n1490,
    n896,
    n1145,
    n847,
    n963
  );


  and
  g1473
  (
    n1503,
    n1317,
    n1055,
    n1326,
    n1039
  );


  xor
  g1474
  (
    n1457,
    n781,
    n1108,
    n1133,
    n835
  );


  xor
  g1475
  (
    n1373,
    n1148,
    n1159,
    n1079,
    n1033
  );


  or
  g1476
  (
    n1405,
    n974,
    n858,
    n1207,
    n1301
  );


  xor
  g1477
  (
    n1479,
    n852,
    n1037,
    n1343,
    n979
  );


  and
  g1478
  (
    n1379,
    n1209,
    n1268,
    n1307,
    n1359
  );


  nor
  g1479
  (
    n1466,
    n920,
    n1356,
    n947,
    n953
  );


  nor
  g1480
  (
    KeyWire_0_16,
    n1362,
    n1271,
    n1364,
    n1358
  );


  or
  g1481
  (
    n1439,
    n1146,
    n1141,
    n913,
    n1323
  );


  nor
  g1482
  (
    n1446,
    n1278,
    n803,
    n780,
    n1070
  );


  and
  g1483
  (
    n1421,
    n1368,
    n775,
    n1013,
    n1131
  );


  xor
  g1484
  (
    n1456,
    n1092,
    n996,
    n956,
    n1347
  );


  xor
  g1485
  (
    n1386,
    n823,
    n1082,
    n1094,
    n810
  );


  nor
  g1486
  (
    n1469,
    n1367,
    n1293,
    n1360,
    n998
  );


  or
  g1487
  (
    n1440,
    n839,
    n1004,
    n1357,
    n868
  );


  nand
  g1488
  (
    n1502,
    n1122,
    n1366,
    n903,
    n1086
  );


  or
  g1489
  (
    n1460,
    n815,
    n1365,
    n1163,
    n1342
  );


  xor
  g1490
  (
    n1415,
    n1088,
    n792,
    n937,
    n1048
  );


  and
  g1491
  (
    n1414,
    n1294,
    n1051,
    n1142,
    n808
  );


  buf
  g1492
  (
    n1524,
    n1371
  );


  not
  g1493
  (
    n1522,
    n1374
  );


  buf
  g1494
  (
    n1523,
    n1373
  );


  not
  g1495
  (
    n1521,
    n1372
  );


  not
  g1496
  (
    n1530,
    n1522
  );


  buf
  g1497
  (
    n1527,
    n1522
  );


  not
  g1498
  (
    n1529,
    n1522
  );


  not
  g1499
  (
    n1525,
    n1521
  );


  buf
  g1500
  (
    n1526,
    n1521
  );


  not
  g1501
  (
    n1528,
    n1521
  );


  xor
  g1502
  (
    n1539,
    n1438,
    n1439,
    n1390,
    n1413
  );


  xor
  g1503
  (
    n1533,
    n1530,
    n1440,
    n1418,
    n1528
  );


  xnor
  g1504
  (
    n1540,
    n1525,
    n1397,
    n1434,
    n1383
  );


  or
  g1505
  (
    n1535,
    n1385,
    n1525,
    n1391,
    n1424
  );


  and
  g1506
  (
    n1548,
    n1384,
    n1406,
    n1404,
    n1529
  );


  xor
  g1507
  (
    n1547,
    n1526,
    n1530,
    n1528,
    n1415
  );


  xnor
  g1508
  (
    n1537,
    n1442,
    n1409,
    n1527,
    n1437
  );


  xor
  g1509
  (
    n1545,
    n1387,
    n1412,
    n1381,
    n1425
  );


  nand
  g1510
  (
    n1546,
    n1407,
    n1376,
    n1426,
    n1432
  );


  xor
  g1511
  (
    KeyWire_0_7,
    n1530,
    n1399,
    n1392,
    n1393
  );


  or
  g1512
  (
    n1534,
    n1420,
    n1445,
    n1389,
    n1388
  );


  xnor
  g1513
  (
    n1551,
    n1431,
    n1394,
    n1443,
    n1408
  );


  or
  g1514
  (
    n1550,
    n1396,
    n1419,
    n1429,
    n1395
  );


  and
  g1515
  (
    n1536,
    n1529,
    n1402,
    n1398,
    n1441
  );


  xor
  g1516
  (
    n1554,
    n1446,
    n1526,
    n1525,
    n1421
  );


  nor
  g1517
  (
    n1553,
    n1529,
    n1527,
    n1382,
    n1401
  );


  xnor
  g1518
  (
    n1543,
    n1403,
    n1411,
    n1428,
    n1527
  );


  nand
  g1519
  (
    n1549,
    n1530,
    n1379,
    n1414,
    n1444
  );


  or
  g1520
  (
    n1541,
    n1378,
    n1417,
    n1410,
    n1528
  );


  or
  g1521
  (
    n1544,
    n1529,
    n1433,
    n1400,
    n1423
  );


  nor
  g1522
  (
    n1531,
    n1386,
    n1435,
    n1436,
    n1526
  );


  or
  g1523
  (
    n1552,
    n1380,
    n1527,
    n1377,
    n1422
  );


  or
  g1524
  (
    n1542,
    n1375,
    n1526,
    n1416,
    n1405
  );


  and
  g1525
  (
    n1532,
    n1525,
    n1427,
    n1430,
    n1528
  );


  and
  g1526
  (
    n1569,
    n1489,
    n1507,
    n1466,
    n1499
  );


  and
  g1527
  (
    n1565,
    n1469,
    n1490,
    n1545,
    n1500
  );


  or
  g1528
  (
    n1572,
    n1462,
    n1482,
    n1468,
    n1543
  );


  and
  g1529
  (
    n1574,
    n1453,
    n1472,
    n1497,
    n1471
  );


  or
  g1530
  (
    n1573,
    n1544,
    n1448,
    n1496,
    n1538
  );


  xor
  g1531
  (
    n1559,
    n1452,
    n1447,
    n1461,
    n1537
  );


  and
  g1532
  (
    n1560,
    n1534,
    n1451,
    n1495,
    n1476
  );


  nor
  g1533
  (
    n1562,
    n1485,
    n1483,
    n1506,
    n1457
  );


  nand
  g1534
  (
    n1575,
    n1456,
    n1545,
    n1477,
    n1449
  );


  nand
  g1535
  (
    n1563,
    n1501,
    n1508,
    n1503,
    n1494
  );


  nor
  g1536
  (
    n1568,
    n1475,
    n1546,
    n1484,
    n1478
  );


  and
  g1537
  (
    n1558,
    n1467,
    n1465,
    n1491,
    n1464
  );


  xnor
  g1538
  (
    n1555,
    n1486,
    n1531,
    n1480,
    n1487
  );


  nand
  g1539
  (
    n1561,
    n1493,
    n1504,
    n1544,
    n1481
  );


  nand
  g1540
  (
    n1557,
    n1473,
    n1540,
    n1488,
    n1459
  );


  xnor
  g1541
  (
    n1570,
    n1535,
    n1454,
    n1502,
    n1545
  );


  nand
  g1542
  (
    n1564,
    n1533,
    n1544,
    n1492,
    n1458
  );


  xor
  g1543
  (
    n1571,
    n1541,
    n1463,
    n1474,
    n1460
  );


  xnor
  g1544
  (
    n1566,
    n1536,
    n1545,
    n1509,
    n1498
  );


  nand
  g1545
  (
    n1567,
    n1479,
    n1539,
    n1505,
    n1542
  );


  nor
  g1546
  (
    n1556,
    n1455,
    n1450,
    n1470,
    n1532
  );


  not
  g1547
  (
    n1576,
    n1575
  );


  not
  g1548
  (
    n1577,
    n1574
  );


  or
  g1549
  (
    n1580,
    n345,
    n346,
    n351,
    n349
  );


  nand
  g1550
  (
    n1578,
    n1524,
    n352,
    n1523,
    n1522
  );


  xor
  g1551
  (
    n1585,
    n1576,
    n1577,
    n1524
  );


  or
  g1552
  (
    n1584,
    n1523,
    n1524,
    n1510,
    n1576
  );


  nand
  g1553
  (
    n1581,
    n354,
    n1523,
    n1577,
    n344
  );


  xor
  g1554
  (
    n1583,
    n355,
    n1524,
    n347,
    n350
  );


  or
  g1555
  (
    n1579,
    n1576,
    n357,
    n1523,
    n348
  );


  or
  g1556
  (
    n1582,
    n1577,
    n1576,
    n356,
    n353
  );


  xnor
  g1557
  (
    n1592,
    n1547,
    n1548,
    n1519,
    n1553
  );


  nor
  g1558
  (
    n1588,
    n1520,
    n1548,
    n1584,
    n1580
  );


  and
  g1559
  (
    n1597,
    n1553,
    n1518,
    n358,
    n1582
  );


  nor
  g1560
  (
    n1600,
    n1550,
    n1513,
    n1584,
    n1581
  );


  nor
  g1561
  (
    n1591,
    n1554,
    n1550,
    n1583,
    n1548
  );


  xor
  g1562
  (
    n1589,
    n1552,
    n1579,
    n1549,
    n1553
  );


  or
  g1563
  (
    n1590,
    n1549,
    n1552,
    n1547,
    n1546
  );


  and
  g1564
  (
    n1594,
    n1551,
    n1553,
    n1583,
    n1548
  );


  xor
  g1565
  (
    n1601,
    n1515,
    n1517,
    n1549,
    n1514
  );


  nand
  g1566
  (
    n1587,
    n1552,
    n1584,
    n1546,
    n1554
  );


  nor
  g1567
  (
    n1599,
    n1554,
    n1546,
    n1585,
    n1551
  );


  nor
  g1568
  (
    n1595,
    n1578,
    n1585,
    n359,
    n1551
  );


  nor
  g1569
  (
    n1598,
    n1585,
    n1516,
    n1549,
    n1547
  );


  nor
  g1570
  (
    n1596,
    n1551,
    n360,
    n1511,
    n1550
  );


  and
  g1571
  (
    n1586,
    n1554,
    n1550,
    n1585,
    n1547
  );


  or
  g1572
  (
    n1593,
    n1584,
    n1512,
    n1552,
    n1583
  );


  nor
  g1573
  (
    n1605,
    n1596,
    n1590,
    n1595,
    n1599
  );


  xor
  g1574
  (
    n1604,
    n1586,
    n1598,
    n1587,
    n1588
  );


  or
  g1575
  (
    n1602,
    n1597,
    n1601,
    n1600,
    n1589
  );


  or
  g1576
  (
    n1603,
    n1592,
    n1591,
    n1593,
    n1594
  );


  xnor
  KeyGate_0_0
  (
    n71,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1153,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n60,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n668,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n633,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n252,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n433,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1538,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n696,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n125,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n53,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n553,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n246,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1303,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1328,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n537,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1423,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1109,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n411,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n205,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n472,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n128,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n539,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n548,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n319,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n818,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n484,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1342,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n354,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n796,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1337,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n967,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n485,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n312,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n1072,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n227,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1032,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n1290,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n116,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n674,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n1495,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n511,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n65,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n442,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n218,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n303,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n1323,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n1267,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n441,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n407,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n223,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n791,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n61,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1037,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n1171,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n833,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n78,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n857,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n1314,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n817,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n492,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n554,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n1491,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n1138,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

