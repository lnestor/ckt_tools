

module Stat_100_410
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n111,
  n106,
  n124,
  n110,
  n104,
  n132,
  n129,
  n125,
  n118,
  n119,
  n121,
  n108,
  n102,
  n109,
  n115,
  n112,
  n130,
  n123,
  n128,
  n101,
  n120,
  n131,
  n107,
  n103,
  n113,
  n117,
  n122,
  n126,
  n116,
  n105,
  n114,
  n127
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n111;output n106;output n124;output n110;output n104;output n132;output n129;output n125;output n118;output n119;output n121;output n108;output n102;output n109;output n115;output n112;output n130;output n123;output n128;output n101;output n120;output n131;output n107;output n103;output n113;output n117;output n122;output n126;output n116;output n105;output n114;output n127;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;

  buf
  g0
  (
    KeyWire_0_10,
    n1
  );


  buf
  g1
  (
    n34,
    n2
  );


  buf
  g2
  (
    n35,
    n2
  );


  buf
  g3
  (
    n33,
    n1
  );


  buf
  g4
  (
    n36,
    n1
  );


  buf
  g5
  (
    KeyWire_0_2,
    n34
  );


  not
  g6
  (
    KeyWire_0_6,
    n37
  );


  buf
  g7
  (
    n49,
    n34
  );


  buf
  g8
  (
    n50,
    n34
  );


  buf
  g9
  (
    n53,
    n35
  );


  not
  g10
  (
    n46,
    n33
  );


  not
  g11
  (
    n55,
    n36
  );


  buf
  g12
  (
    n44,
    n35
  );


  not
  g13
  (
    n52,
    n35
  );


  buf
  g14
  (
    n42,
    n33
  );


  buf
  g15
  (
    n48,
    n37
  );


  buf
  g16
  (
    n54,
    n36
  );


  buf
  g17
  (
    n45,
    n36
  );


  not
  g18
  (
    KeyWire_0_1,
    n36
  );


  buf
  g19
  (
    n39,
    n34
  );


  not
  g20
  (
    n51,
    n37
  );


  buf
  g21
  (
    n38,
    n35
  );


  buf
  g22
  (
    n43,
    n33
  );


  buf
  g23
  (
    n47,
    n37
  );


  buf
  g24
  (
    n96,
    n54
  );


  buf
  g25
  (
    n94,
    n40
  );


  not
  g26
  (
    n93,
    n54
  );


  not
  g27
  (
    KeyWire_0_15,
    n45
  );


  buf
  g28
  (
    KeyWire_0_9,
    n9
  );


  buf
  g29
  (
    n60,
    n26
  );


  xnor
  g30
  (
    n61,
    n31,
    n47,
    n48
  );


  nor
  g31
  (
    KeyWire_0_13,
    n28,
    n31,
    n18,
    n4
  );


  xor
  g32
  (
    n88,
    n28,
    n38,
    n16,
    n48
  );


  xnor
  g33
  (
    n98,
    n53,
    n29,
    n14,
    n25
  );


  xor
  g34
  (
    KeyWire_0_11,
    n16,
    n5,
    n28,
    n43
  );


  or
  g35
  (
    KeyWire_0_4,
    n22,
    n19,
    n6,
    n21
  );


  xnor
  g36
  (
    n57,
    n52,
    n10,
    n7,
    n18
  );


  xor
  g37
  (
    n71,
    n22,
    n9,
    n42,
    n26
  );


  xnor
  g38
  (
    n63,
    n44,
    n6,
    n32,
    n55
  );


  nor
  g39
  (
    n64,
    n38,
    n25,
    n4,
    n41
  );


  xnor
  g40
  (
    KeyWire_0_7,
    n39,
    n46,
    n49,
    n13
  );


  nor
  g41
  (
    n95,
    n27,
    n27,
    n21,
    n46
  );


  and
  g42
  (
    n99,
    n25,
    n47,
    n23,
    n3
  );


  nor
  g43
  (
    KeyWire_0_3,
    n46,
    n23,
    n49,
    n19
  );


  and
  g44
  (
    n58,
    n43,
    n13,
    n53,
    n2
  );


  or
  g45
  (
    n87,
    n5,
    n12,
    n25,
    n56
  );


  and
  g46
  (
    n69,
    n50,
    n55,
    n40,
    n29
  );


  nand
  g47
  (
    n89,
    n7,
    n13,
    n39,
    n52
  );


  nand
  g48
  (
    n80,
    n17,
    n32,
    n30
  );


  nor
  g49
  (
    n81,
    n18,
    n51,
    n45,
    n12
  );


  nand
  g50
  (
    n67,
    n6,
    n24,
    n30,
    n28
  );


  nand
  g51
  (
    n86,
    n24,
    n49,
    n27,
    n56
  );


  nand
  g52
  (
    n76,
    n14,
    n11,
    n3,
    n26
  );


  and
  g53
  (
    n83,
    n17,
    n27,
    n9,
    n41
  );


  nand
  g54
  (
    n59,
    n12,
    n41,
    n3,
    n8
  );


  and
  g55
  (
    KeyWire_0_12,
    n53,
    n47,
    n51,
    n44
  );


  and
  g56
  (
    n100,
    n8,
    n44,
    n56,
    n24
  );


  nor
  g57
  (
    n77,
    n19,
    n17,
    n15,
    n31
  );


  and
  g58
  (
    n68,
    n14,
    n15,
    n30,
    n20
  );


  xor
  g59
  (
    n90,
    n23,
    n32,
    n8,
    n20
  );


  or
  g60
  (
    n91,
    n31,
    n43,
    n42,
    n10
  );


  and
  g61
  (
    n74,
    n38,
    n51,
    n55,
    n11
  );


  xnor
  g62
  (
    n62,
    n29,
    n54,
    n50,
    n52
  );


  nor
  g63
  (
    KeyWire_0_14,
    n26,
    n16,
    n5,
    n15
  );


  or
  g64
  (
    n65,
    n40,
    n39,
    n7,
    n10
  );


  xnor
  g65
  (
    n75,
    n32,
    n24,
    n22,
    n48
  );


  xnor
  g66
  (
    n66,
    n50,
    n21,
    n29,
    n4
  );


  nand
  g67
  (
    n97,
    n20,
    n42,
    n11,
    n45
  );


  xnor
  g68
  (
    n104,
    n72,
    n78,
    n92,
    n59
  );


  nor
  g69
  (
    n117,
    n81,
    n93,
    n80,
    n85
  );


  or
  g70
  (
    n115,
    n59,
    n74,
    n65,
    n93
  );


  xor
  g71
  (
    n106,
    n80,
    n95,
    n67,
    n97
  );


  xor
  g72
  (
    n118,
    n100,
    n84,
    n76,
    n71
  );


  nor
  g73
  (
    n124,
    n86,
    n62,
    n90,
    n59
  );


  and
  g74
  (
    n131,
    n77,
    n72,
    n70,
    n63
  );


  nor
  g75
  (
    n116,
    n97,
    n83,
    n95
  );


  or
  g76
  (
    n105,
    n76,
    n64,
    n80,
    n96
  );


  xnor
  g77
  (
    n103,
    n91,
    n66,
    n58,
    n98
  );


  or
  g78
  (
    n129,
    n70,
    n69,
    n62,
    n81
  );


  xnor
  g79
  (
    n101,
    n98,
    n60,
    n100,
    n78
  );


  xnor
  g80
  (
    n109,
    n99,
    n70,
    n85,
    n87
  );


  xnor
  g81
  (
    n121,
    n88,
    n61,
    n65,
    n77
  );


  and
  g82
  (
    n102,
    n73,
    n67,
    n89,
    n63
  );


  and
  g83
  (
    n111,
    n90,
    n73,
    n78,
    n72
  );


  and
  g84
  (
    n127,
    n87,
    n92,
    n68,
    n79
  );


  xor
  g85
  (
    n119,
    n94,
    n75,
    n74,
    n91
  );


  xor
  g86
  (
    n113,
    n87,
    n96,
    n92,
    n71
  );


  xnor
  g87
  (
    n110,
    n67,
    n75,
    n94,
    n73
  );


  nor
  g88
  (
    n114,
    n64,
    n71,
    n89,
    n79
  );


  or
  g89
  (
    n107,
    n63,
    n83,
    n85,
    n65
  );


  xnor
  g90
  (
    n112,
    n77,
    n74,
    n88,
    n68
  );


  nor
  g91
  (
    n120,
    n99,
    n60,
    n86,
    n75
  );


  nand
  g92
  (
    n128,
    n99,
    n86,
    n95,
    n66
  );


  nand
  g93
  (
    KeyWire_0_0,
    n96,
    n81,
    n57,
    n62
  );


  nor
  g94
  (
    n132,
    n82,
    n84,
    n88,
    n91
  );


  xnor
  g95
  (
    KeyWire_0_5,
    n61,
    n98,
    n90,
    n69
  );


  and
  g96
  (
    n125,
    n64,
    n61,
    n66,
    n84
  );


  xnor
  g97
  (
    KeyWire_0_8,
    n60,
    n69,
    n76,
    n68
  );


  xnor
  g98
  (
    n126,
    n93,
    n79,
    n97,
    n82
  );


  xor
  g99
  (
    n108,
    n89,
    n100,
    n82,
    n94
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n123,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n41,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n40,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n78,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n82,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n122,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n56,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n70,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n130,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n85,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n37,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n92,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n84,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n79,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n73,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n72,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


