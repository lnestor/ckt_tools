

module Stat_100_63
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n43,
  n115,
  n88,
  n103,
  n96,
  n97,
  n80,
  n100,
  n66,
  n77,
  n102,
  n75,
  n65,
  n111,
  n78,
  n95,
  n82,
  n106,
  n129,
  n123,
  n121,
  n119,
  n124,
  n125,
  n120,
  n122,
  n127,
  n126,
  n128,
  n132,
  n131,
  n130
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n43;output n115;output n88;output n103;output n96;output n97;output n80;output n100;output n66;output n77;output n102;output n75;output n65;output n111;output n78;output n95;output n82;output n106;output n129;output n123;output n121;output n119;output n124;output n125;output n120;output n122;output n127;output n126;output n128;output n132;output n131;output n130;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n76;wire n79;wire n81;wire n83;wire n84;wire n85;wire n86;wire n87;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n98;wire n99;wire n101;wire n104;wire n105;wire n107;wire n108;wire n109;wire n110;wire n112;wire n113;wire n114;wire n116;wire n117;wire n118;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n35,
    n1
  );


  buf
  g1
  (
    n36,
    n2
  );


  buf
  g2
  (
    n33,
    n1
  );


  not
  g3
  (
    n37,
    n1
  );


  buf
  g4
  (
    n38,
    n1
  );


  not
  g5
  (
    KeyWire_0_20,
    n2
  );


  not
  g6
  (
    KeyWire_0_22,
    n37
  );


  not
  g7
  (
    n41,
    n37
  );


  buf
  g8
  (
    n42,
    n2
  );


  buf
  g9
  (
    n43,
    n3
  );


  nand
  g10
  (
    n39,
    n2,
    n36
  );


  not
  g11
  (
    n44,
    n43
  );


  buf
  g12
  (
    KeyWire_0_29,
    n40
  );


  buf
  g13
  (
    n47,
    n41
  );


  not
  g14
  (
    KeyWire_0_0,
    n42
  );


  buf
  g15
  (
    n61,
    n44
  );


  buf
  g16
  (
    n58,
    n44
  );


  buf
  g17
  (
    KeyWire_0_11,
    n4
  );


  not
  g18
  (
    KeyWire_0_5,
    n5
  );


  buf
  g19
  (
    n56,
    n47
  );


  buf
  g20
  (
    KeyWire_0_18,
    n45
  );


  buf
  g21
  (
    KeyWire_0_21,
    n4
  );


  buf
  g22
  (
    KeyWire_0_7,
    n46
  );


  buf
  g23
  (
    n55,
    n6
  );


  buf
  g24
  (
    n62,
    n3
  );


  buf
  g25
  (
    n52,
    n46
  );


  buf
  g26
  (
    n53,
    n46
  );


  nor
  g27
  (
    n60,
    n45,
    n4,
    n5,
    n46
  );


  nor
  g28
  (
    n57,
    n45,
    n47,
    n44
  );


  xnor
  g29
  (
    KeyWire_0_24,
    n44,
    n5,
    n3,
    n4
  );


  or
  g30
  (
    n51,
    n47,
    n45,
    n5,
    n3
  );


  not
  g31
  (
    n110,
    n9
  );


  buf
  g32
  (
    n100,
    n7
  );


  buf
  g33
  (
    n80,
    n59
  );


  buf
  g34
  (
    KeyWire_0_26,
    n52
  );


  not
  g35
  (
    n117,
    n26
  );


  not
  g36
  (
    n73,
    n23
  );


  buf
  g37
  (
    n94,
    n19
  );


  not
  g38
  (
    n86,
    n50
  );


  buf
  g39
  (
    KeyWire_0_25,
    n38
  );


  not
  g40
  (
    KeyWire_0_31,
    n20
  );


  not
  g41
  (
    n107,
    n60
  );


  not
  g42
  (
    n72,
    n6
  );


  not
  g43
  (
    KeyWire_0_9,
    n9
  );


  buf
  g44
  (
    KeyWire_0_14,
    n8
  );


  not
  g45
  (
    KeyWire_0_15,
    n28
  );


  xor
  g46
  (
    n66,
    n20,
    n61,
    n10
  );


  xnor
  g47
  (
    n105,
    n8,
    n14,
    n18,
    n28
  );


  nor
  g48
  (
    n88,
    n57,
    n56,
    n58,
    n31
  );


  xnor
  g49
  (
    n67,
    n51,
    n56,
    n11,
    n13
  );


  xnor
  g50
  (
    n84,
    n18,
    n61,
    n27,
    n60
  );


  nand
  g51
  (
    n103,
    n53,
    n18,
    n62
  );


  and
  g52
  (
    KeyWire_0_2,
    n14,
    n48,
    n31,
    n7
  );


  xor
  g53
  (
    KeyWire_0_4,
    n28,
    n57,
    n60,
    n49
  );


  nor
  g54
  (
    n95,
    n16,
    n32,
    n15,
    n57
  );


  nor
  g55
  (
    n118,
    n26,
    n12,
    n31,
    n27
  );


  xnor
  g56
  (
    n109,
    n21,
    n12,
    n49,
    n32
  );


  nor
  g57
  (
    n102,
    n28,
    n30,
    n14,
    n16
  );


  xnor
  g58
  (
    n78,
    n32,
    n11,
    n15,
    n54
  );


  or
  g59
  (
    n71,
    n16,
    n63,
    n18,
    n25
  );


  nor
  g60
  (
    KeyWire_0_28,
    n53,
    n14,
    n51,
    n57
  );


  nand
  g61
  (
    n93,
    n22,
    n30,
    n63,
    n58
  );


  xor
  g62
  (
    n74,
    n23,
    n10,
    n37,
    n27
  );


  xor
  g63
  (
    n85,
    n60,
    n29,
    n6,
    n27
  );


  xor
  g64
  (
    KeyWire_0_13,
    n55,
    n53,
    n12,
    n13
  );


  xnor
  g65
  (
    KeyWire_0_16,
    n52,
    n52,
    n21,
    n16
  );


  and
  g66
  (
    n106,
    n25,
    n19,
    n23,
    n55
  );


  or
  g67
  (
    KeyWire_0_27,
    n26,
    n55,
    n63,
    n29
  );


  xnor
  g68
  (
    n87,
    n59,
    n52,
    n50,
    n13
  );


  or
  g69
  (
    KeyWire_0_23,
    n53,
    n15,
    n19,
    n24
  );


  or
  g70
  (
    n116,
    n58,
    n29,
    n56,
    n62
  );


  and
  g71
  (
    n104,
    n21,
    n38,
    n22,
    n17
  );


  nand
  g72
  (
    n82,
    n23,
    n10,
    n48,
    n51
  );


  xnor
  g73
  (
    n65,
    n20,
    n48,
    n9,
    n13
  );


  and
  g74
  (
    n76,
    n6,
    n63,
    n49,
    n10
  );


  and
  g75
  (
    KeyWire_0_3,
    n24,
    n50,
    n7,
    n59
  );


  nor
  g76
  (
    KeyWire_0_30,
    n21,
    n24,
    n30
  );


  nand
  g77
  (
    KeyWire_0_6,
    n51,
    n54,
    n8,
    n56
  );


  xnor
  g78
  (
    n98,
    n8,
    n22,
    n9,
    n26
  );


  nand
  g79
  (
    n101,
    n20,
    n59,
    n54,
    n17
  );


  nand
  g80
  (
    n77,
    n49,
    n25,
    n29,
    n61
  );


  nor
  g81
  (
    KeyWire_0_12,
    n15,
    n31,
    n19,
    n12
  );


  and
  g82
  (
    n90,
    n38,
    n58,
    n22,
    n11
  );


  and
  g83
  (
    KeyWire_0_8,
    n55,
    n32,
    n62,
    n48
  );


  nand
  g84
  (
    KeyWire_0_1,
    n7,
    n50,
    n25,
    n54
  );


  or
  g85
  (
    n70,
    n11,
    n30,
    n17
  );


  xnor
  g86
  (
    KeyWire_0_10,
    n118,
    n101,
    n107,
    n115
  );


  xnor
  g87
  (
    n122,
    n95,
    n110,
    n113,
    n103
  );


  xor
  g88
  (
    KeyWire_0_19,
    n115,
    n111,
    n116,
    n118
  );


  xnor
  g89
  (
    n119,
    n86,
    n106,
    n100,
    n84
  );


  nor
  g90
  (
    n132,
    n112,
    n99,
    n94,
    n82
  );


  xnor
  g91
  (
    n120,
    n80,
    n77,
    n117,
    n93
  );


  and
  g92
  (
    n124,
    n117,
    n97,
    n116,
    n115
  );


  or
  g93
  (
    KeyWire_0_17,
    n117,
    n89,
    n104,
    n98
  );


  and
  g94
  (
    n126,
    n114,
    n116,
    n88,
    n87
  );


  nand
  g95
  (
    n125,
    n105,
    n113,
    n96,
    n92
  );


  nor
  g96
  (
    n127,
    n85,
    n109,
    n102,
    n78
  );


  nand
  g97
  (
    n129,
    n112,
    n114,
    n90,
    n113
  );


  and
  g98
  (
    n123,
    n79,
    n108,
    n114,
    n112
  );


  and
  g99
  (
    n121,
    n83,
    n118,
    n81,
    n91
  );


  xnor
  KeyGate_0_0
  (
    n45,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n114,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n79,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n113,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n89,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n50,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n112,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n63,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n92,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n68,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n130,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n59,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n111,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n69,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n115,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n81,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n99,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n128,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n54,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n131,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n34,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n49,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n40,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n91,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n48,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n75,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n108,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n64,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n96,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n46,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n83,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n97,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


