// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_59 written by SynthGen on 2021/04/05 11:22:31
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_59 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n90, n113, n105, n89, n92, n114, n94, n118,
 n82, n88, n111, n102, n95, n119, n110, n93,
 n101, n87, n91, n97, n86, n98, n107, n106,
 n112, n117, n123, n130, n132, n128, n131, n129);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n90, n113, n105, n89, n92, n114, n94, n118,
 n82, n88, n111, n102, n95, n119, n110, n93,
 n101, n87, n91, n97, n86, n98, n107, n106,
 n112, n117, n123, n130, n132, n128, n131, n129;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n83, n84, n85, n96, n99, n100, n103,
 n104, n108, n109, n115, n116, n120, n121, n122,
 n124, n125, n126, n127;

not  g0 (n68, n17);
buf  g1 (n58, n30);
buf  g2 (n55, n30);
buf  g3 (n34, n6);
not  g4 (n53, n31);
not  g5 (n64, n14);
buf  g6 (n63, n11);
not  g7 (n35, n26);
buf  g8 (n42, n31);
buf  g9 (n37, n5);
not  g10 (n36, n24);
buf  g11 (n61, n23);
buf  g12 (n51, n32);
not  g13 (n54, n9);
not  g14 (n38, n18);
buf  g15 (n71, n8);
buf  g16 (n44, n21);
buf  g17 (n65, n7);
buf  g18 (n40, n20);
not  g19 (n56, n31);
not  g20 (n66, n15);
not  g21 (n49, n32);
buf  g22 (n50, n28);
buf  g23 (n62, n10);
not  g24 (n33, n13);
buf  g25 (n52, n12);
not  g26 (n43, n4);
not  g27 (n70, n22);
buf  g28 (n67, n2);
buf  g29 (n59, n19);
not  g30 (n41, n29);
buf  g31 (n47, n25);
not  g32 (n46, n30);
not  g33 (n60, n3);
not  g34 (n39, n1);
buf  g35 (n57, n27);
buf  g36 (n45, n31);
buf  g37 (n48, n32);
buf  g38 (n69, n16);
not  g39 (n73, n35);
not  g40 (n76, n37);
not  g41 (n75, n37);
not  g42 (n80, n34);
not  g43 (n78, n36);
not  g44 (n77, n37);
not  g45 (n81, n33);
not  g46 (n74, n36);
buf  g47 (n72, n38);
not  g48 (n79, n36);
or   g49 (n91, n76, n60, n72, n59);
xor  g50 (n92, n60, n75, n80, n48);
or   g51 (n106, n57, n56, n42, n74);
and  g52 (n84, n57, n74, n65, n44);
nand g53 (n88, n43, n47, n41, n46);
or   g54 (n103, n57, n79, n80, n58);
xor  g55 (n82, n66, n73, n46, n40);
nand g56 (n86, n39, n58, n55, n78);
xnor g57 (n115, n63, n54, n56, n46);
xor  g58 (n105, n66, n42, n62, n77);
nand g59 (n120, n50, n47, n40, n79);
xnor g60 (n87, n44, n47, n56, n49);
nor  g61 (n114, n78, n81, n48, n40);
or   g62 (n95, n51, n43, n48, n64);
or   g63 (n108, n43, n66, n77, n42);
xor  g64 (n117, n55, n57, n74, n47);
nand g65 (n97, n58, n63, n53, n51);
nand g66 (n113, n56, n52, n45, n75);
nor  g67 (n112, n61, n53, n39, n54);
or   g68 (n90, n50, n78, n41, n73);
nor  g69 (n83, n46, n80, n58, n49);
nor  g70 (n119, n67, n78, n81, n49);
xor  g71 (n104, n48, n53, n67);
xor  g72 (n110, n77, n60, n76, n44);
xor  g73 (n99, n63, n50, n64, n39);
and  g74 (n94, n79, n79, n40, n72);
xor  g75 (n121, n44, n39, n67, n66);
or   g76 (n107, n49, n73, n54, n77);
or   g77 (n98, n61, n81, n72);
nand g78 (n116, n74, n42, n45, n38);
xor  g79 (n93, n55, n52, n68, n75);
or   g80 (n100, n67, n50, n55, n72);
and  g81 (n111, n65, n52, n45, n38);
xnor g82 (n89, n80, n59, n64, n75);
or   g83 (n109, n76, n61, n63, n38);
and  g84 (n96, n76, n65, n59, n41);
nor  g85 (n102, n65, n61, n62, n59);
xor  g86 (n118, n51, n43, n64, n54);
nor  g87 (n101, n62, n62, n73, n51);
nand g88 (n85, n60, n41, n45, n52);
not  g89 (n122, n116);
not  g90 (n123, n120);
not  g91 (n126, n118);
nand g92 (n124, n117, n32, n119, n110);
and  g93 (n125, n113, n109, n121, n115);
nor  g94 (n127, n112, n114, n111, n108);
nand g95 (n130, n69, n71, n126, n125);
or   g96 (n131, n71, n69);
or   g97 (n128, n68, n70, n123, n69);
xor  g98 (n132, n71, n68, n70);
and  g99 (n129, n124, n70, n68, n127);
endmodule
