// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_403_1822 written by SynthGen on 2021/05/24 19:47:35
module Stat_403_1822( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19,
 n193, n210, n211, n204, n189, n202, n212, n364,
 n368, n367, n371, n372, n377, n375, n418, n421,
 n417, n419, n422, n420);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19;

output n193, n210, n211, n204, n189, n202, n212, n364,
 n368, n367, n371, n372, n377, n375, n418, n421,
 n417, n419, n422, n420;

wire n20, n21, n22, n23, n24, n25, n26, n27,
 n28, n29, n30, n31, n32, n33, n34, n35,
 n36, n37, n38, n39, n40, n41, n42, n43,
 n44, n45, n46, n47, n48, n49, n50, n51,
 n52, n53, n54, n55, n56, n57, n58, n59,
 n60, n61, n62, n63, n64, n65, n66, n67,
 n68, n69, n70, n71, n72, n73, n74, n75,
 n76, n77, n78, n79, n80, n81, n82, n83,
 n84, n85, n86, n87, n88, n89, n90, n91,
 n92, n93, n94, n95, n96, n97, n98, n99,
 n100, n101, n102, n103, n104, n105, n106, n107,
 n108, n109, n110, n111, n112, n113, n114, n115,
 n116, n117, n118, n119, n120, n121, n122, n123,
 n124, n125, n126, n127, n128, n129, n130, n131,
 n132, n133, n134, n135, n136, n137, n138, n139,
 n140, n141, n142, n143, n144, n145, n146, n147,
 n148, n149, n150, n151, n152, n153, n154, n155,
 n156, n157, n158, n159, n160, n161, n162, n163,
 n164, n165, n166, n167, n168, n169, n170, n171,
 n172, n173, n174, n175, n176, n177, n178, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n190, n191, n192, n194, n195, n196, n197,
 n198, n199, n200, n201, n203, n205, n206, n207,
 n208, n209, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n365, n366, n369, n370, n373, n374, n376,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416;

buf  g0 (n39, n12);
not  g1 (n94, n1);
buf  g2 (n32, n17);
buf  g3 (n73, n8);
buf  g4 (n78, n3);
buf  g5 (n22, n19);
not  g6 (n59, n1);
buf  g7 (n27, n11);
not  g8 (n89, n18);
not  g9 (n40, n14);
buf  g10 (n20, n18);
buf  g11 (n74, n9);
buf  g12 (n82, n5);
not  g13 (n63, n8);
buf  g14 (n42, n9);
not  g15 (n43, n17);
buf  g16 (n80, n10);
not  g17 (n35, n2);
buf  g18 (n67, n10);
not  g19 (n56, n8);
buf  g20 (n50, n3);
not  g21 (n70, n5);
buf  g22 (n44, n16);
buf  g23 (n68, n6);
not  g24 (n81, n4);
not  g25 (n41, n9);
not  g26 (n26, n2);
buf  g27 (n53, n13);
buf  g28 (n29, n5);
buf  g29 (n88, n16);
not  g30 (n38, n18);
buf  g31 (n51, n3);
not  g32 (n46, n18);
not  g33 (n90, n13);
buf  g34 (n49, n1);
not  g35 (n25, n8);
not  g36 (n31, n9);
not  g37 (n34, n5);
not  g38 (n58, n3);
buf  g39 (n71, n13);
not  g40 (n37, n7);
not  g41 (n47, n13);
buf  g42 (n93, n19);
buf  g43 (n86, n2);
not  g44 (n91, n6);
buf  g45 (n45, n12);
buf  g46 (n55, n17);
buf  g47 (n61, n11);
buf  g48 (n33, n14);
buf  g49 (n83, n17);
not  g50 (n79, n1);
not  g51 (n24, n10);
buf  g52 (n87, n11);
not  g53 (n62, n16);
buf  g54 (n77, n12);
not  g55 (n69, n7);
not  g56 (n92, n15);
buf  g57 (n60, n7);
buf  g58 (n28, n10);
buf  g59 (n76, n15);
buf  g60 (n65, n16);
buf  g61 (n84, n2);
buf  g62 (n95, n19);
buf  g63 (n21, n6);
not  g64 (n30, n14);
not  g65 (n64, n4);
not  g66 (n23, n11);
not  g67 (n72, n4);
not  g68 (n36, n15);
buf  g69 (n54, n12);
not  g70 (n48, n14);
not  g71 (n85, n4);
not  g72 (n52, n15);
not  g73 (n75, n19);
buf  g74 (n57, n6);
buf  g75 (n66, n7);
not  g76 (n115, n36);
buf  g77 (n124, n47);
not  g78 (n156, n37);
buf  g79 (n123, n37);
buf  g80 (n152, n57);
buf  g81 (n168, n57);
buf  g82 (n153, n54);
not  g83 (n137, n33);
buf  g84 (n159, n30);
not  g85 (n132, n34);
not  g86 (n136, n53);
not  g87 (n148, n33);
buf  g88 (n135, n29);
buf  g89 (n130, n23);
not  g90 (n160, n39);
buf  g91 (n141, n26);
buf  g92 (n133, n53);
buf  g93 (n112, n34);
buf  g94 (n181, n47);
buf  g95 (n107, n21);
not  g96 (n151, n41);
not  g97 (n171, n40);
buf  g98 (n158, n45);
buf  g99 (n169, n52);
buf  g100 (n176, n50);
buf  g101 (n125, n30);
not  g102 (n108, n59);
buf  g103 (n175, n44);
buf  g104 (n119, n43);
not  g105 (n116, n46);
not  g106 (n161, n26);
buf  g107 (n157, n51);
not  g108 (n105, n42);
buf  g109 (n163, n48);
not  g110 (n99, n22);
buf  g111 (n179, n60);
buf  g112 (n117, n49);
buf  g113 (n178, n50);
not  g114 (n102, n49);
buf  g115 (n131, n51);
buf  g116 (n182, n36);
buf  g117 (n165, n27);
not  g118 (n166, n30);
buf  g119 (n167, n24);
buf  g120 (n113, n55);
buf  g121 (n188, n50);
buf  g122 (n172, n61);
buf  g123 (n177, n42);
buf  g124 (n147, n58);
not  g125 (n185, n48);
not  g126 (n98, n27);
buf  g127 (n111, n41);
not  g128 (n122, n60);
buf  g129 (n164, n60);
not  g130 (n120, n29);
not  g131 (n101, n60);
buf  g132 (n104, n31);
not  g133 (n145, n57);
not  g134 (n110, n61);
buf  g135 (n106, n59);
buf  g136 (n126, n43);
buf  g137 (n128, n53);
not  g138 (n121, n35);
buf  g139 (n154, n35);
buf  g140 (n114, n20);
not  g141 (n187, n52);
buf  g142 (n96, n44);
buf  g143 (n186, n38);
not  g144 (n146, n56);
not  g145 (n180, n51);
not  g146 (n155, n28);
not  g147 (n144, n55);
nor  g148 (n134, n42, n61);
nor  g149 (n162, n25, n46, n40, n50);
xnor g150 (n97, n48, n58, n40, n56);
xor  g151 (n183, n28, n28, n38, n55);
nor  g152 (n143, n36, n49, n35, n37);
nand g153 (n139, n56, n54, n27, n55);
xor  g154 (n184, n52, n53, n32, n58);
nor  g155 (n140, n47, n34, n32, n46);
xnor g156 (n109, n52, n56, n22, n45);
nor  g157 (n127, n33, n54, n42, n59);
nand g158 (n150, n41, n21, n59, n40);
xnor g159 (n142, n28, n47, n48, n41);
xnor g160 (n149, n38, n32, n25, n61);
xor  g161 (n173, n44, n43, n58, n31);
xnor g162 (n138, n31, n39, n45, n57);
xnor g163 (n118, n45, n32, n30, n37);
nor  g164 (n103, n23, n24, n20, n44);
nor  g165 (n129, n31, n38, n34, n46);
xor  g166 (n100, n49, n35, n33, n51);
nand g167 (n174, n29, n29, n39, n36);
or   g168 (n170, n43, n54, n27, n39);
xor  g169 (n191, n75, n100, n64, n70);
xnor g170 (n204, n63, n125, n71, n97);
nand g171 (n199, n104, n72, n98, n74);
xnor g172 (n196, n101, n111, n115, n76);
and  g173 (n189, n65, n124, n106, n129);
and  g174 (n203, n65, n77, n74);
xor  g175 (n208, n96, n126, n120, n122);
xor  g176 (n192, n68, n119, n65, n113);
xor  g177 (n190, n70, n99, n67);
nand g178 (n197, n76, n71, n77, n107);
nor  g179 (n205, n127, n62, n68, n66);
nor  g180 (n201, n65, n62, n73, n117);
or   g181 (n206, n76, n69, n123, n71);
and  g182 (n207, n67, n75, n118, n108);
nand g183 (n210, n69, n72, n64, n78);
nor  g184 (n194, n73, n73, n63, n75);
or   g185 (n211, n128, n63, n72, n110);
and  g186 (n200, n72, n74, n64, n69);
nand g187 (n195, n105, n66, n77, n62);
and  g188 (n213, n70, n74, n68, n62);
and  g189 (n202, n102, n112, n121, n66);
and  g190 (n193, n116, n109, n63, n66);
or   g191 (n209, n114, n68, n78, n73);
nor  g192 (n198, n64, n70, n69, n76);
xnor g193 (n212, n67, n71, n103, n75);
buf  g194 (n223, n205);
buf  g195 (n225, n197);
not  g196 (n219, n145);
buf  g197 (n221, n137);
not  g198 (n217, n138);
buf  g199 (n214, n135);
xor  g200 (n220, n131, n196);
xnor g201 (n215, n207, n136, n201, n130);
and  g202 (n222, n202, n140, n198, n203);
and  g203 (n224, n142, n139, n133, n200);
xor  g204 (n216, n144, n143, n199, n206);
nand g205 (n218, n204, n141, n132, n134);
buf  g206 (n246, n220);
not  g207 (n232, n214);
buf  g208 (n242, n217);
buf  g209 (n241, n225);
not  g210 (n227, n210);
not  g211 (n226, n225);
buf  g212 (n240, n221);
buf  g213 (n236, n218);
not  g214 (n235, n223);
buf  g215 (n231, n215);
buf  g216 (n234, n224);
buf  g217 (n239, n222);
buf  g218 (n228, n224);
not  g219 (n243, n222);
buf  g220 (n233, n221);
buf  g221 (n247, n208);
not  g222 (n245, n216);
not  g223 (n244, n219);
buf  g224 (n237, n220);
buf  g225 (n238, n216);
buf  g226 (n230, n223);
xor  g227 (n229, n217, n218, n209, n219);
not  g228 (n250, n230);
not  g229 (n255, n232);
buf  g230 (n254, n227);
buf  g231 (n253, n226);
not  g232 (n265, n229);
buf  g233 (n258, n229);
buf  g234 (n249, n232);
buf  g235 (n260, n233);
buf  g236 (n259, n230);
buf  g237 (n263, n232);
not  g238 (n256, n231);
buf  g239 (n264, n232);
not  g240 (n266, n228);
not  g241 (n251, n231);
buf  g242 (n252, n231);
buf  g243 (n261, n226);
not  g244 (n262, n228);
buf  g245 (n248, n231);
not  g246 (n257, n227);
and  g247 (n291, n149, n147, n234, n253);
nor  g248 (n274, n166, n235, n236, n168);
nor  g249 (n279, n255, n252, n153, n233);
nand g250 (n270, n241, n243, n239, n257);
nor  g251 (n277, n160, n241, n249);
xnor g252 (n286, n256, n254, n179, n173);
nand g253 (n290, n250, n248, n253, n239);
xor  g254 (n268, n243, n237, n250, n236);
nand g255 (n281, n167, n238, n161, n239);
nand g256 (n282, n242, n242, n234, n238);
xor  g257 (n267, n235, n233, n163, n236);
or   g258 (n271, n169, n237, n248, n254);
xnor g259 (n292, n146, n256, n251, n158);
nand g260 (n273, n157, n174, n243, n162);
xnor g261 (n284, n171, n176, n155, n256);
xor  g262 (n278, n257, n152, n175, n178);
xnor g263 (n272, n254, n256, n177, n255);
nor  g264 (n283, n255, n252, n240, n235);
and  g265 (n269, n239, n151, n236, n165);
or   g266 (n276, n159, n251, n164, n255);
or   g267 (n280, n243, n238, n249, n241);
xnor g268 (n275, n235, n242, n233, n150);
nor  g269 (n288, n240, n170, n172, n238);
nor  g270 (n285, n234, n242, n240, n254);
xnor g271 (n289, n237, n154, n257, n240);
nand g272 (n287, n156, n237, n148, n234);
or   g273 (n295, n257, n269, n270, n259);
nor  g274 (n296, n268, n260, n258);
or   g275 (n293, n259, n274, n272, n271);
or   g276 (n297, n267, n258, n273);
nor  g277 (n294, n260, n259);
buf  g278 (n304, n294);
not  g279 (n308, n297);
buf  g280 (n309, n297);
not  g281 (n311, n275);
not  g282 (n301, n295);
not  g283 (n310, n295);
not  g284 (n307, n296);
not  g285 (n305, n294);
not  g286 (n300, n295);
not  g287 (n303, n293);
buf  g288 (n298, n278);
buf  g289 (n306, n296);
buf  g290 (n313, n297);
buf  g291 (n312, n296);
and  g292 (n299, n276, n277);
or   g293 (n302, n293, n295, n296, n297);
not  g294 (n315, n78);
xnor g295 (n321, n284, n245);
xor  g296 (n330, n300, n313, n80, n247);
nor  g297 (n331, n244, n310, n213, n312);
xor  g298 (n326, n244, n78, n79, n311);
and  g299 (n328, n301, n290, n313, n79);
or   g300 (n316, n279, n286, n312, n280);
xnor g301 (n332, n245, n212, n303, n310);
and  g302 (n325, n246, n82, n81, n307);
nor  g303 (n323, n285, n82, n81, n80);
nand g304 (n314, n247, n298, n306, n309);
or   g305 (n329, n79, n302, n247, n82);
xor  g306 (n322, n311, n246, n289, n79);
xor  g307 (n317, n245, n83, n246, n288);
or   g308 (n320, n304, n281, n287, n80);
nor  g309 (n324, n244, n308, n246, n291);
nand g310 (n318, n80, n211, n83, n282);
and  g311 (n327, n299, n81, n247, n244);
nor  g312 (n319, n305, n82, n81, n283);
not  g313 (n347, n315);
buf  g314 (n339, n318);
not  g315 (n344, n318);
not  g316 (n337, n317);
not  g317 (n350, n322);
buf  g318 (n340, n314);
buf  g319 (n351, n316);
buf  g320 (n349, n319);
buf  g321 (n341, n321);
buf  g322 (n345, n322);
not  g323 (n346, n322);
buf  g324 (n333, n315);
buf  g325 (n342, n319);
buf  g326 (n352, n314);
not  g327 (n335, n316);
not  g328 (n338, n320);
buf  g329 (n348, n322);
not  g330 (n336, n320);
not  g331 (n334, n321);
not  g332 (n343, n317);
and  g333 (n355, n335, n333, n326, n327);
and  g334 (n353, n327, n328, n324, n323);
xnor g335 (n359, n335, n328, n334, n329);
or   g336 (n354, n328, n323, n327, n326);
and  g337 (n361, n336, n324, n325);
xor  g338 (n357, n326, n333, n334, n328);
or   g339 (n356, n329, n323, n324, n335);
and  g340 (n360, n324, n327, n325, n336);
xor  g341 (n358, n325, n335, n323, n326);
or   g342 (n368, n342, n341, n356, n338);
nor  g343 (n365, n353, n360, n342, n341);
nand g344 (n370, n337, n337, n343, n342);
xor  g345 (n366, n343, n340);
nand g346 (n369, n337, n339, n338);
and  g347 (n371, n336, n339, n337);
and  g348 (n364, n359, n343, n358, n342);
xor  g349 (n367, n355, n338, n361);
xor  g350 (n363, n338, n340, n354, n357);
nor  g351 (n362, n336, n341, n343);
nor  g352 (n375, n85, n85, n369, n368);
nand g353 (n372, n83, n85, n87);
xor  g354 (n376, n86, n84);
nor  g355 (n377, n87, n86, n371, n370);
and  g356 (n373, n84, n366, n367, n83);
xnor g357 (n374, n292, n85, n86);
nand g358 (n380, n188, n185, n182, n183);
xor  g359 (n378, n186, n184, n375, n180);
nand g360 (n379, n376, n187, n181, n377);
or   g361 (n381, n352, n379, n347, n345);
xnor g362 (n383, n352, n345, n348, n349);
and  g363 (n390, n349, n345, n380, n379);
or   g364 (n391, n379, n347, n380, n378);
and  g365 (n389, n346, n352, n351, n344);
xnor g366 (n392, n379, n346, n378);
xnor g367 (n387, n378, n380, n346, n350);
xor  g368 (n386, n344, n349, n351, n348);
or   g369 (n382, n345, n378, n344, n349);
and  g370 (n388, n380, n350, n351);
nand g371 (n384, n348, n344, n347, n351);
xnor g372 (n385, n348, n350, n352, n347);
xnor g373 (n399, n263, n332, n89, n95);
nand g374 (n414, n91, n332, n264, n94);
nor  g375 (n406, n266, n262, n261, n391);
xnor g376 (n410, n91, n386, n388, n93);
xor  g377 (n396, n264, n330, n261, n93);
or   g378 (n405, n389, n382, n262, n386);
nor  g379 (n401, n93, n88, n94, n95);
nor  g380 (n395, n383, n92, n331, n94);
nor  g381 (n400, n260, n266, n88, n92);
and  g382 (n394, n382, n90, n264, n332);
and  g383 (n415, n389, n265, n261, n387);
xor  g384 (n407, n330, n88, n263);
xnor g385 (n403, n266, n90, n390, n392);
nor  g386 (n398, n329, n89, n90, n261);
nor  g387 (n393, n332, n387, n263, n91);
or   g388 (n397, n265, n330, n331, n390);
and  g389 (n408, n95, n392, n92, n89);
xor  g390 (n402, n263, n331, n262, n384);
xor  g391 (n413, n381, n329, n331, n262);
xor  g392 (n409, n385, n95, n90, n89);
xnor g393 (n411, n265, n381, n385, n94);
nand g394 (n416, n383, n391, n92, n265);
and  g395 (n412, n330, n87, n266, n91);
xor  g396 (n404, n93, n264, n388, n384);
and  g397 (n420, n412, n400, n398, n413);
nand g398 (n421, n405, n415, n397, n409);
nor  g399 (n419, n403, n393, n408, n411);
xnor g400 (n418, n396, n406, n401, n416);
and  g401 (n422, n414, n394, n399, n402);
and  g402 (n417, n407, n410, n404, n395);
endmodule
