// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1639_37_8 written by SynthGen on 2021/05/24 19:45:40
module Stat_1639_37_8( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17,
 n1393, n1395, n1402, n1392, n1376, n1379, n1387, n1381,
 n1390, n1380, n1399, n1388, n1386, n1374, n1445, n1449,
 n1467, n1656);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17;

output n1393, n1395, n1402, n1392, n1376, n1379, n1387, n1381,
 n1390, n1380, n1399, n1388, n1386, n1374, n1445, n1449,
 n1467, n1656;

wire n18, n19, n20, n21, n22, n23, n24, n25,
 n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
 n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
 n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
 n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
 n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
 n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
 n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
 n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
 n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
 n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
 n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
 n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
 n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
 n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
 n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
 n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
 n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
 n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
 n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
 n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
 n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
 n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
 n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
 n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
 n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
 n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
 n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
 n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
 n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
 n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
 n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
 n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
 n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
 n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
 n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
 n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
 n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
 n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
 n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
 n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
 n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
 n1370, n1371, n1372, n1373, n1375, n1377, n1378, n1382,
 n1383, n1384, n1385, n1389, n1391, n1394, n1396, n1397,
 n1398, n1400, n1401, n1403, n1404, n1405, n1406, n1407,
 n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
 n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
 n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
 n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
 n1440, n1441, n1442, n1443, n1444, n1446, n1447, n1448,
 n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
 n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
 n1466, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655;

not  g0 (n83, n11);
not  g1 (n43, n12);
buf  g2 (n67, n13);
not  g3 (n68, n16);
buf  g4 (n49, n16);
buf  g5 (n51, n4);
not  g6 (n42, n15);
not  g7 (n58, n9);
buf  g8 (n31, n9);
not  g9 (n45, n11);
not  g10 (n69, n6);
not  g11 (n82, n11);
buf  g12 (n30, n7);
buf  g13 (n46, n5);
buf  g14 (n41, n4);
not  g15 (n22, n5);
not  g16 (n60, n11);
not  g17 (n35, n7);
not  g18 (n72, n13);
not  g19 (n47, n3);
buf  g20 (n57, n6);
buf  g21 (n38, n10);
buf  g22 (n37, n1);
buf  g23 (n62, n15);
buf  g24 (n40, n4);
not  g25 (n36, n1);
buf  g26 (n54, n14);
not  g27 (n23, n14);
not  g28 (n32, n6);
buf  g29 (n63, n8);
not  g30 (n76, n16);
not  g31 (n71, n14);
buf  g32 (n53, n16);
not  g33 (n70, n3);
not  g34 (n65, n17);
buf  g35 (n50, n13);
buf  g36 (n19, n1);
buf  g37 (n27, n15);
buf  g38 (n85, n6);
buf  g39 (n61, n12);
not  g40 (n29, n14);
buf  g41 (n48, n9);
not  g42 (n66, n13);
buf  g43 (n28, n12);
buf  g44 (n56, n10);
not  g45 (n33, n12);
not  g46 (n79, n15);
not  g47 (n25, n10);
buf  g48 (n26, n10);
buf  g49 (n20, n17);
buf  g50 (n39, n2);
not  g51 (n55, n4);
not  g52 (n64, n7);
not  g53 (n81, n2);
not  g54 (n59, n3);
not  g55 (n84, n3);
buf  g56 (n18, n17);
not  g57 (n80, n1);
buf  g58 (n73, n8);
buf  g59 (n44, n8);
buf  g60 (n21, n5);
buf  g61 (n34, n8);
not  g62 (n77, n9);
buf  g63 (n78, n5);
buf  g64 (n75, n17);
not  g65 (n24, n2);
not  g66 (n52, n7);
not  g67 (n74, n2);
buf  g68 (n250, n35);
not  g69 (n170, n38);
buf  g70 (n131, n27);
not  g71 (n295, n47);
not  g72 (n189, n49);
buf  g73 (n160, n50);
buf  g74 (n280, n45);
not  g75 (n242, n26);
not  g76 (n212, n55);
buf  g77 (n210, n34);
buf  g78 (n149, n60);
not  g79 (n183, n68);
buf  g80 (n220, n38);
buf  g81 (n256, n39);
buf  g82 (n224, n23);
buf  g83 (n180, n46);
buf  g84 (n285, n31);
buf  g85 (n252, n33);
buf  g86 (n209, n57);
not  g87 (n119, n29);
buf  g88 (n182, n22);
not  g89 (n264, n60);
not  g90 (n243, n52);
buf  g91 (n88, n67);
not  g92 (n269, n69);
buf  g93 (n96, n44);
buf  g94 (n187, n44);
not  g95 (n266, n52);
not  g96 (n117, n59);
not  g97 (n239, n45);
buf  g98 (n112, n23);
not  g99 (n270, n37);
buf  g100 (n142, n65);
not  g101 (n110, n30);
not  g102 (n143, n69);
not  g103 (n144, n36);
buf  g104 (n120, n36);
not  g105 (n116, n68);
not  g106 (n244, n59);
not  g107 (n139, n30);
not  g108 (n291, n48);
buf  g109 (n275, n39);
buf  g110 (n192, n42);
buf  g111 (n289, n57);
not  g112 (n129, n65);
not  g113 (n225, n35);
buf  g114 (n154, n61);
not  g115 (n146, n41);
buf  g116 (n113, n29);
not  g117 (n229, n53);
not  g118 (n161, n48);
not  g119 (n249, n41);
not  g120 (n196, n31);
buf  g121 (n228, n56);
not  g122 (n136, n34);
not  g123 (n157, n46);
buf  g124 (n206, n43);
buf  g125 (n99, n30);
not  g126 (n86, n49);
buf  g127 (n150, n26);
buf  g128 (n151, n48);
not  g129 (n167, n70);
not  g130 (n272, n46);
not  g131 (n191, n29);
buf  g132 (n185, n40);
buf  g133 (n287, n19);
buf  g134 (n273, n69);
not  g135 (n231, n27);
not  g136 (n194, n58);
buf  g137 (n169, n62);
buf  g138 (n234, n19);
not  g139 (n171, n49);
buf  g140 (n259, n37);
not  g141 (n162, n19);
not  g142 (n248, n32);
not  g143 (n195, n32);
buf  g144 (n122, n64);
buf  g145 (n89, n28);
not  g146 (n271, n65);
buf  g147 (n147, n62);
not  g148 (n125, n25);
buf  g149 (n178, n26);
not  g150 (n104, n38);
buf  g151 (n199, n63);
not  g152 (n121, n50);
not  g153 (n101, n55);
buf  g154 (n155, n43);
buf  g155 (n230, n66);
buf  g156 (n100, n27);
not  g157 (n245, n25);
buf  g158 (n90, n54);
buf  g159 (n216, n39);
buf  g160 (n254, n33);
buf  g161 (n204, n31);
not  g162 (n260, n18);
not  g163 (n102, n68);
not  g164 (n276, n18);
not  g165 (n237, n51);
not  g166 (n98, n51);
not  g167 (n241, n29);
buf  g168 (n141, n67);
buf  g169 (n223, n58);
buf  g170 (n168, n63);
not  g171 (n94, n42);
buf  g172 (n135, n43);
not  g173 (n261, n28);
buf  g174 (n284, n63);
not  g175 (n173, n43);
not  g176 (n222, n22);
not  g177 (n140, n64);
buf  g178 (n277, n63);
buf  g179 (n97, n37);
not  g180 (n200, n36);
buf  g181 (n207, n69);
not  g182 (n197, n47);
buf  g183 (n106, n61);
not  g184 (n214, n62);
not  g185 (n91, n23);
buf  g186 (n172, n57);
not  g187 (n267, n21);
not  g188 (n188, n20);
not  g189 (n174, n48);
not  g190 (n114, n41);
buf  g191 (n293, n61);
buf  g192 (n283, n33);
buf  g193 (n247, n20);
not  g194 (n246, n40);
buf  g195 (n124, n24);
buf  g196 (n263, n34);
not  g197 (n240, n60);
not  g198 (n215, n66);
buf  g199 (n115, n33);
not  g200 (n133, n49);
buf  g201 (n132, n52);
buf  g202 (n92, n45);
buf  g203 (n213, n21);
not  g204 (n255, n44);
not  g205 (n176, n24);
buf  g206 (n111, n70);
not  g207 (n288, n57);
buf  g208 (n175, n39);
not  g209 (n202, n50);
buf  g210 (n274, n53);
not  g211 (n265, n21);
not  g212 (n292, n21);
buf  g213 (n190, n24);
buf  g214 (n153, n53);
buf  g215 (n152, n22);
buf  g216 (n227, n67);
not  g217 (n268, n24);
not  g218 (n184, n54);
not  g219 (n208, n58);
not  g220 (n105, n36);
buf  g221 (n257, n42);
not  g222 (n232, n27);
not  g223 (n217, n30);
not  g224 (n109, n22);
not  g225 (n87, n40);
buf  g226 (n164, n64);
buf  g227 (n258, n64);
buf  g228 (n108, n25);
buf  g229 (n262, n50);
buf  g230 (n201, n66);
not  g231 (n156, n51);
buf  g232 (n221, n25);
buf  g233 (n107, n55);
not  g234 (n126, n56);
buf  g235 (n95, n23);
buf  g236 (n159, n34);
buf  g237 (n251, n59);
buf  g238 (n137, n28);
not  g239 (n186, n67);
not  g240 (n103, n56);
not  g241 (n279, n54);
not  g242 (n179, n55);
not  g243 (n236, n58);
buf  g244 (n123, n47);
not  g245 (n203, n41);
buf  g246 (n294, n52);
buf  g247 (n130, n31);
buf  g248 (n278, n26);
buf  g249 (n138, n54);
not  g250 (n226, n44);
buf  g251 (n290, n38);
not  g252 (n218, n45);
not  g253 (n118, n68);
buf  g254 (n158, n65);
buf  g255 (n286, n51);
buf  g256 (n177, n19);
buf  g257 (n219, n62);
not  g258 (n163, n35);
not  g259 (n134, n18);
not  g260 (n145, n32);
buf  g261 (n181, n53);
buf  g262 (n128, n61);
not  g263 (n281, n60);
buf  g264 (n235, n32);
buf  g265 (n166, n47);
buf  g266 (n165, n37);
buf  g267 (n198, n35);
buf  g268 (n233, n20);
not  g269 (n193, n59);
buf  g270 (n93, n40);
not  g271 (n282, n46);
not  g272 (n127, n18);
not  g273 (n211, n28);
not  g274 (n253, n42);
buf  g275 (n148, n20);
not  g276 (n238, n56);
buf  g277 (n205, n66);
not  g278 (n1000, n197);
buf  g279 (n351, n291);
not  g280 (n670, n282);
buf  g281 (n621, n133);
not  g282 (n360, n266);
buf  g283 (n455, n156);
not  g284 (n1037, n131);
buf  g285 (n936, n278);
buf  g286 (n620, n86);
not  g287 (n655, n188);
buf  g288 (n638, n122);
buf  g289 (n744, n222);
not  g290 (n952, n196);
buf  g291 (n1009, n143);
buf  g292 (n1011, n262);
buf  g293 (n297, n135);
not  g294 (n1042, n120);
not  g295 (n357, n205);
not  g296 (n468, n152);
not  g297 (n431, n115);
not  g298 (n964, n182);
not  g299 (n754, n90);
buf  g300 (n732, n189);
not  g301 (n579, n260);
buf  g302 (n520, n101);
not  g303 (n984, n107);
buf  g304 (n944, n138);
buf  g305 (n731, n177);
not  g306 (n920, n209);
not  g307 (n750, n276);
not  g308 (n826, n141);
buf  g309 (n828, n286);
not  g310 (n302, n193);
not  g311 (n786, n150);
buf  g312 (n667, n179);
buf  g313 (n449, n241);
not  g314 (n582, n147);
not  g315 (n562, n200);
not  g316 (n861, n288);
not  g317 (n906, n259);
not  g318 (n590, n281);
buf  g319 (n969, n191);
buf  g320 (n1048, n234);
buf  g321 (n1047, n103);
not  g322 (n589, n214);
buf  g323 (n927, n254);
not  g324 (n1054, n201);
not  g325 (n488, n246);
not  g326 (n618, n143);
buf  g327 (n1058, n179);
not  g328 (n834, n88);
buf  g329 (n997, n248);
buf  g330 (n1010, n216);
not  g331 (n342, n210);
not  g332 (n914, n143);
not  g333 (n540, n171);
buf  g334 (n462, n150);
buf  g335 (n672, n182);
buf  g336 (n661, n183);
not  g337 (n660, n244);
buf  g338 (n332, n264);
not  g339 (n546, n226);
not  g340 (n950, n291);
not  g341 (n532, n87);
not  g342 (n598, n265);
buf  g343 (n447, n170);
not  g344 (n921, n291);
buf  g345 (n989, n141);
not  g346 (n939, n166);
buf  g347 (n885, n175);
not  g348 (n1035, n236);
not  g349 (n690, n161);
not  g350 (n572, n289);
not  g351 (n413, n292);
buf  g352 (n869, n273);
buf  g353 (n668, n264);
not  g354 (n391, n233);
buf  g355 (n912, n110);
not  g356 (n634, n223);
not  g357 (n985, n188);
not  g358 (n894, n167);
buf  g359 (n507, n228);
buf  g360 (n979, n270);
not  g361 (n784, n252);
buf  g362 (n677, n278);
not  g363 (n626, n254);
not  g364 (n785, n286);
buf  g365 (n816, n286);
buf  g366 (n791, n191);
not  g367 (n533, n234);
not  g368 (n593, n117);
not  g369 (n900, n166);
buf  g370 (n755, n222);
not  g371 (n477, n230);
not  g372 (n712, n203);
not  g373 (n902, n231);
not  g374 (n1021, n290);
buf  g375 (n1041, n246);
buf  g376 (n519, n124);
buf  g377 (n474, n206);
buf  g378 (n949, n182);
buf  g379 (n487, n237);
buf  g380 (n646, n176);
buf  g381 (n630, n279);
not  g382 (n359, n162);
not  g383 (n873, n125);
not  g384 (n1014, n204);
not  g385 (n597, n124);
buf  g386 (n794, n262);
not  g387 (n945, n220);
buf  g388 (n525, n230);
not  g389 (n693, n258);
not  g390 (n876, n203);
buf  g391 (n535, n91);
buf  g392 (n851, n186);
not  g393 (n448, n125);
buf  g394 (n790, n247);
buf  g395 (n314, n259);
not  g396 (n820, n199);
not  g397 (n671, n110);
buf  g398 (n575, n266);
not  g399 (n502, n197);
buf  g400 (n508, n214);
buf  g401 (n493, n184);
buf  g402 (n767, n268);
buf  g403 (n1017, n167);
not  g404 (n1016, n213);
not  g405 (n406, n179);
buf  g406 (n963, n250);
not  g407 (n547, n201);
buf  g408 (n913, n238);
not  g409 (n639, n163);
not  g410 (n722, n248);
not  g411 (n980, n120);
not  g412 (n1051, n148);
not  g413 (n930, n229);
buf  g414 (n938, n237);
buf  g415 (n743, n172);
not  g416 (n1044, n263);
buf  g417 (n560, n259);
not  g418 (n889, n129);
buf  g419 (n537, n227);
buf  g420 (n830, n147);
buf  g421 (n498, n150);
not  g422 (n724, n237);
buf  g423 (n496, n285);
buf  g424 (n922, n284);
not  g425 (n865, n147);
not  g426 (n511, n180);
buf  g427 (n401, n123);
not  g428 (n1059, n122);
not  g429 (n955, n263);
buf  g430 (n435, n232);
not  g431 (n764, n98);
not  g432 (n821, n124);
not  g433 (n962, n281);
buf  g434 (n749, n284);
buf  g435 (n399, n228);
buf  g436 (n599, n266);
buf  g437 (n381, n98);
buf  g438 (n499, n173);
not  g439 (n362, n265);
not  g440 (n315, n167);
not  g441 (n832, n102);
not  g442 (n684, n279);
buf  g443 (n741, n254);
buf  g444 (n891, n212);
buf  g445 (n1004, n249);
buf  g446 (n375, n162);
buf  g447 (n747, n199);
buf  g448 (n926, n172);
not  g449 (n862, n149);
buf  g450 (n321, n237);
buf  g451 (n787, n228);
buf  g452 (n728, n118);
not  g453 (n908, n116);
not  g454 (n471, n206);
not  g455 (n494, n164);
not  g456 (n421, n120);
buf  g457 (n772, n130);
buf  g458 (n654, n261);
not  g459 (n866, n219);
buf  g460 (n319, n136);
not  g461 (n890, n265);
not  g462 (n662, n289);
buf  g463 (n941, n199);
not  g464 (n602, n178);
not  g465 (n358, n124);
not  g466 (n354, n274);
not  g467 (n640, n227);
buf  g468 (n402, n161);
not  g469 (n1036, n184);
not  g470 (n703, n236);
buf  g471 (n298, n152);
not  g472 (n965, n103);
not  g473 (n692, n281);
buf  g474 (n418, n189);
not  g475 (n622, n230);
buf  g476 (n1034, n136);
buf  g477 (n363, n280);
not  g478 (n367, n277);
not  g479 (n714, n125);
buf  g480 (n542, n177);
not  g481 (n858, n233);
buf  g482 (n443, n176);
buf  g483 (n611, n164);
buf  g484 (n932, n231);
buf  g485 (n849, n120);
not  g486 (n991, n130);
not  g487 (n460, n215);
buf  g488 (n669, n140);
not  g489 (n387, n244);
buf  g490 (n616, n215);
buf  g491 (n549, n246);
not  g492 (n553, n86);
buf  g493 (n458, n186);
buf  g494 (n1024, n191);
buf  g495 (n839, n255);
buf  g496 (n1056, n157);
not  g497 (n1022, n115);
not  g498 (n355, n209);
not  g499 (n423, n182);
buf  g500 (n735, n106);
not  g501 (n683, n128);
not  g502 (n696, n213);
buf  g503 (n781, n262);
buf  g504 (n937, n109);
not  g505 (n442, n282);
buf  g506 (n842, n280);
not  g507 (n751, n135);
not  g508 (n925, n108);
buf  g509 (n419, n245);
buf  g510 (n469, n257);
buf  g511 (n464, n279);
not  g512 (n570, n158);
buf  g513 (n329, n134);
not  g514 (n472, n203);
buf  g515 (n960, n272);
not  g516 (n623, n91);
not  g517 (n859, n89);
buf  g518 (n372, n229);
not  g519 (n994, n227);
not  g520 (n734, n276);
not  g521 (n860, n189);
not  g522 (n420, n151);
not  g523 (n365, n219);
buf  g524 (n1057, n123);
buf  g525 (n393, n212);
not  g526 (n489, n140);
not  g527 (n574, n162);
buf  g528 (n336, n146);
buf  g529 (n877, n173);
not  g530 (n948, n156);
not  g531 (n765, n218);
not  g532 (n933, n206);
buf  g533 (n361, n89);
buf  g534 (n1033, n255);
buf  g535 (n721, n240);
not  g536 (n601, n119);
not  g537 (n919, n271);
buf  g538 (n648, n111);
not  g539 (n716, n217);
buf  g540 (n335, n231);
buf  g541 (n588, n248);
buf  g542 (n910, n250);
buf  g543 (n817, n283);
buf  g544 (n380, n99);
buf  g545 (n343, n239);
buf  g546 (n776, n185);
buf  g547 (n710, n251);
buf  g548 (n774, n166);
buf  g549 (n430, n154);
buf  g550 (n641, n269);
buf  g551 (n345, n261);
not  g552 (n461, n102);
buf  g553 (n495, n139);
not  g554 (n675, n173);
buf  g555 (n658, n190);
buf  g556 (n608, n292);
not  g557 (n567, n253);
buf  g558 (n674, n241);
buf  g559 (n799, n175);
not  g560 (n739, n165);
buf  g561 (n306, n158);
buf  g562 (n768, n196);
not  g563 (n895, n293);
not  g564 (n304, n111);
not  g565 (n452, n274);
buf  g566 (n673, n274);
buf  g567 (n580, n260);
buf  g568 (n628, n236);
not  g569 (n417, n170);
buf  g570 (n709, n252);
not  g571 (n565, n276);
not  g572 (n901, n195);
buf  g573 (n564, n293);
buf  g574 (n935, n211);
buf  g575 (n454, n139);
buf  g576 (n1031, n247);
not  g577 (n529, n241);
buf  g578 (n797, n155);
buf  g579 (n441, n267);
buf  g580 (n967, n232);
buf  g581 (n436, n290);
not  g582 (n522, n199);
not  g583 (n353, n225);
buf  g584 (n917, n289);
not  g585 (n649, n242);
not  g586 (n946, n277);
not  g587 (n451, n251);
not  g588 (n301, n194);
not  g589 (n923, n201);
not  g590 (n867, n223);
not  g591 (n528, n279);
not  g592 (n470, n271);
buf  g593 (n656, n208);
buf  g594 (n727, n151);
buf  g595 (n465, n207);
not  g596 (n808, n96);
not  g597 (n536, n266);
not  g598 (n689, n162);
buf  g599 (n303, n207);
buf  g600 (n534, n204);
buf  g601 (n491, n153);
not  g602 (n550, n161);
not  g603 (n390, n153);
buf  g604 (n338, n195);
not  g605 (n814, n202);
not  g606 (n717, n251);
not  g607 (n940, n92);
buf  g608 (n513, n144);
not  g609 (n317, n242);
not  g610 (n956, n243);
buf  g611 (n569, n168);
not  g612 (n676, n210);
buf  g613 (n551, n287);
buf  g614 (n1029, n208);
buf  g615 (n957, n211);
buf  g616 (n591, n168);
not  g617 (n323, n127);
buf  g618 (n538, n263);
buf  g619 (n825, n221);
not  g620 (n878, n220);
buf  g621 (n778, n88);
not  g622 (n340, n177);
not  g623 (n915, n275);
not  g624 (n339, n119);
buf  g625 (n539, n223);
buf  g626 (n833, n181);
not  g627 (n934, n246);
buf  g628 (n823, n188);
not  g629 (n379, n269);
not  g630 (n752, n174);
not  g631 (n356, n219);
buf  g632 (n679, n138);
not  g633 (n327, n243);
not  g634 (n871, n216);
not  g635 (n476, n202);
not  g636 (n446, n215);
buf  g637 (n863, n163);
not  g638 (n897, n292);
not  g639 (n713, n198);
not  g640 (n485, n244);
buf  g641 (n974, n264);
buf  g642 (n831, n181);
buf  g643 (n617, n150);
not  g644 (n411, n143);
not  g645 (n612, n154);
buf  g646 (n1053, n264);
buf  g647 (n389, n123);
buf  g648 (n993, n158);
buf  g649 (n978, n96);
not  g650 (n384, n113);
buf  g651 (n886, n208);
buf  g652 (n615, n170);
buf  g653 (n746, n249);
not  g654 (n879, n105);
buf  g655 (n310, n97);
not  g656 (n619, n145);
buf  g657 (n635, n280);
not  g658 (n771, n196);
not  g659 (n483, n267);
buf  g660 (n970, n192);
not  g661 (n490, n104);
buf  g662 (n584, n243);
not  g663 (n299, n107);
buf  g664 (n1055, n292);
not  g665 (n976, n220);
buf  g666 (n947, n113);
buf  g667 (n1015, n136);
not  g668 (n457, n226);
buf  g669 (n691, n263);
not  g670 (n531, n178);
buf  g671 (n653, n209);
not  g672 (n973, n269);
buf  g673 (n334, n244);
buf  g674 (n903, n235);
not  g675 (n857, n169);
buf  g676 (n603, n253);
not  g677 (n586, n252);
buf  g678 (n811, n130);
not  g679 (n311, n207);
buf  g680 (n800, n206);
not  g681 (n840, n239);
not  g682 (n835, n216);
buf  g683 (n426, n256);
not  g684 (n806, n135);
not  g685 (n606, n272);
not  g686 (n337, n119);
not  g687 (n514, n152);
not  g688 (n308, n232);
not  g689 (n497, n253);
buf  g690 (n783, n204);
buf  g691 (n422, n198);
not  g692 (n990, n138);
not  g693 (n1007, n238);
not  g694 (n898, n202);
not  g695 (n500, n200);
not  g696 (n804, n172);
buf  g697 (n459, n164);
buf  g698 (n300, n142);
not  g699 (n809, n207);
not  g700 (n1045, n174);
not  g701 (n510, n278);
buf  g702 (n347, n190);
buf  g703 (n466, n145);
not  g704 (n374, n87);
not  g705 (n523, n258);
buf  g706 (n405, n114);
buf  g707 (n296, n221);
not  g708 (n796, n163);
not  g709 (n792, n226);
not  g710 (n313, n183);
buf  g711 (n366, n153);
buf  g712 (n893, n149);
not  g713 (n704, n255);
not  g714 (n845, n285);
buf  g715 (n1050, n274);
not  g716 (n1005, n267);
buf  g717 (n410, n291);
not  g718 (n988, n192);
not  g719 (n408, n121);
not  g720 (n371, n222);
buf  g721 (n445, n186);
not  g722 (n942, n225);
not  g723 (n1028, n201);
not  g724 (n370, n176);
buf  g725 (n382, n151);
not  g726 (n836, n140);
buf  g727 (n999, n171);
buf  g728 (n557, n216);
buf  g729 (n899, n197);
not  g730 (n951, n165);
not  g731 (n720, n134);
not  g732 (n650, n194);
buf  g733 (n518, n145);
buf  g734 (n700, n195);
buf  g735 (n394, n95);
not  g736 (n665, n137);
buf  g737 (n972, n160);
buf  g738 (n473, n144);
not  g739 (n1008, n257);
buf  g740 (n305, n187);
not  g741 (n813, n137);
buf  g742 (n943, n209);
not  g743 (n916, n128);
buf  g744 (n484, n208);
buf  g745 (n812, n260);
buf  g746 (n456, n187);
not  g747 (n853, n99);
not  g748 (n911, n234);
buf  g749 (n856, n93);
not  g750 (n516, n259);
not  g751 (n707, n154);
not  g752 (n909, n212);
not  g753 (n847, n164);
not  g754 (n779, n190);
not  g755 (n624, n268);
not  g756 (n663, n136);
not  g757 (n782, n225);
not  g758 (n827, n159);
buf  g759 (n986, n181);
buf  g760 (n872, n168);
not  g761 (n726, n277);
buf  g762 (n733, n138);
buf  g763 (n388, n282);
not  g764 (n438, n157);
not  g765 (n924, n200);
buf  g766 (n810, n241);
not  g767 (n307, n146);
buf  g768 (n770, n255);
buf  g769 (n555, n240);
buf  g770 (n1002, n245);
not  g771 (n864, n116);
buf  g772 (n368, n129);
buf  g773 (n718, n93);
not  g774 (n742, n127);
buf  g775 (n659, n183);
not  g776 (n706, n290);
not  g777 (n753, n160);
not  g778 (n711, n174);
not  g779 (n666, n127);
buf  g780 (n541, n215);
buf  g781 (n705, n239);
buf  g782 (n854, n261);
not  g783 (n1012, n273);
buf  g784 (n759, n172);
not  g785 (n631, n118);
buf  g786 (n467, n104);
buf  g787 (n1023, n187);
buf  g788 (n837, n117);
not  g789 (n330, n196);
not  g790 (n364, n130);
not  g791 (n571, n152);
buf  g792 (n838, n160);
buf  g793 (n479, n236);
buf  g794 (n407, n149);
not  g795 (n352, n275);
buf  g796 (n633, n287);
not  g797 (n585, n142);
buf  g798 (n708, n262);
buf  g799 (n376, n224);
not  g800 (n982, n146);
buf  g801 (n758, n287);
buf  g802 (n773, n210);
not  g803 (n587, n249);
buf  g804 (n1027, n283);
not  g805 (n576, n224);
buf  g806 (n801, n225);
buf  g807 (n882, n284);
not  g808 (n995, n140);
buf  g809 (n1043, n132);
not  g810 (n512, n126);
buf  g811 (n918, n232);
buf  g812 (n775, n218);
not  g813 (n645, n214);
buf  g814 (n841, n258);
not  g815 (n651, n217);
not  g816 (n719, n186);
not  g817 (n780, n121);
buf  g818 (n501, n178);
not  g819 (n1038, n185);
buf  g820 (n740, n213);
not  g821 (n492, n289);
not  g822 (n760, n191);
buf  g823 (n762, n247);
buf  g824 (n843, n251);
not  g825 (n552, n155);
buf  g826 (n425, n121);
not  g827 (n530, n221);
not  g828 (n953, n156);
not  g829 (n998, n132);
not  g830 (n429, n258);
buf  g831 (n604, n286);
not  g832 (n344, n131);
buf  g833 (n412, n284);
not  g834 (n798, n229);
not  g835 (n524, n288);
buf  g836 (n395, n185);
buf  g837 (n341, n133);
buf  g838 (n1039, n193);
buf  g839 (n766, n195);
buf  g840 (n453, n151);
not  g841 (n561, n256);
buf  g842 (n803, n148);
not  g843 (n819, n183);
not  g844 (n807, n105);
buf  g845 (n600, n272);
not  g846 (n888, n272);
not  g847 (n605, n248);
not  g848 (n688, n135);
buf  g849 (n657, n125);
not  g850 (n416, n212);
not  g851 (n829, n166);
buf  g852 (n398, n227);
not  g853 (n1013, n271);
buf  g854 (n404, n167);
not  g855 (n996, n218);
not  g856 (n573, n275);
not  g857 (n795, n245);
buf  g858 (n958, n188);
buf  g859 (n777, n106);
buf  g860 (n369, n256);
buf  g861 (n992, n134);
buf  g862 (n527, n122);
buf  g863 (n1001, n127);
not  g864 (n971, n265);
not  g865 (n1025, n169);
not  g866 (n350, n217);
buf  g867 (n378, n141);
buf  g868 (n577, n92);
buf  g869 (n647, n250);
buf  g870 (n789, n175);
not  g871 (n439, n290);
not  g872 (n409, n133);
buf  g873 (n333, n210);
buf  g874 (n987, n276);
buf  g875 (n581, n147);
not  g876 (n961, n287);
not  g877 (n558, n165);
buf  g878 (n1046, n181);
not  g879 (n848, n94);
buf  g880 (n349, n145);
buf  g881 (n1019, n288);
buf  g882 (n424, n171);
buf  g883 (n385, n211);
not  g884 (n870, n283);
not  g885 (n463, n108);
not  g886 (n968, n192);
not  g887 (n324, n194);
not  g888 (n444, n119);
buf  g889 (n875, n187);
not  g890 (n373, n250);
not  g891 (n644, n202);
buf  g892 (n977, n249);
not  g893 (n757, n220);
not  g894 (n482, n197);
not  g895 (n642, n132);
buf  g896 (n824, n268);
not  g897 (n694, n205);
buf  g898 (n904, n205);
not  g899 (n983, n122);
buf  g900 (n543, n198);
not  g901 (n852, n175);
buf  g902 (n844, n180);
not  g903 (n607, n189);
not  g904 (n594, n128);
not  g905 (n1020, n177);
buf  g906 (n769, n142);
buf  g907 (n954, n185);
not  g908 (n521, n242);
buf  g909 (n846, n100);
buf  g910 (n805, n224);
not  g911 (n905, n156);
buf  g912 (n818, n268);
buf  g913 (n383, n240);
buf  g914 (n907, n142);
not  g915 (n1026, n90);
not  g916 (n392, n235);
buf  g917 (n309, n184);
not  g918 (n931, n126);
not  g919 (n312, n261);
not  g920 (n815, n238);
buf  g921 (n745, n282);
not  g922 (n883, n137);
not  g923 (n678, n94);
buf  g924 (n929, n247);
buf  g925 (n437, n193);
buf  g926 (n583, n154);
buf  g927 (n1049, n270);
buf  g928 (n884, n132);
buf  g929 (n475, n285);
buf  g930 (n715, n277);
not  g931 (n346, n252);
not  g932 (n737, n243);
not  g933 (n440, n101);
buf  g934 (n788, n180);
not  g935 (n386, n273);
buf  g936 (n548, n173);
buf  g937 (n966, n238);
buf  g938 (n316, n288);
not  g939 (n855, n153);
buf  g940 (n554, n178);
buf  g941 (n563, n217);
not  g942 (n556, n157);
buf  g943 (n729, n139);
buf  g944 (n544, n148);
buf  g945 (n503, n285);
buf  g946 (n478, n174);
not  g947 (n328, n155);
buf  g948 (n761, n213);
buf  g949 (n517, n193);
buf  g950 (n725, n270);
not  g951 (n730, n170);
not  g952 (n959, n205);
not  g953 (n480, n129);
not  g954 (n566, n233);
buf  g955 (n643, n155);
not  g956 (n509, n222);
buf  g957 (n1018, n144);
buf  g958 (n578, n223);
not  g959 (n515, n235);
buf  g960 (n559, n214);
not  g961 (n625, n240);
not  g962 (n686, n160);
buf  g963 (n636, n231);
buf  g964 (n325, n194);
buf  g965 (n793, n126);
buf  g966 (n428, n168);
not  g967 (n1003, n131);
not  g968 (n331, n275);
buf  g969 (n736, n278);
not  g970 (n756, n234);
not  g971 (n433, n242);
buf  g972 (n723, n131);
not  g973 (n738, n157);
buf  g974 (n637, n176);
buf  g975 (n629, n179);
buf  g976 (n981, n180);
buf  g977 (n1052, n141);
not  g978 (n652, n123);
buf  g979 (n613, n200);
buf  g980 (n415, n283);
not  g981 (n822, n148);
not  g982 (n627, n269);
buf  g983 (n896, n184);
buf  g984 (n763, n128);
not  g985 (n892, n235);
buf  g986 (n504, n219);
not  g987 (n434, n280);
not  g988 (n568, n270);
buf  g989 (n596, n273);
buf  g990 (n1030, n129);
buf  g991 (n377, n190);
buf  g992 (n400, n204);
not  g993 (n396, n139);
buf  g994 (n506, n134);
buf  g995 (n664, n158);
buf  g996 (n1032, n198);
not  g997 (n348, n112);
not  g998 (n687, n95);
not  g999 (n595, n260);
not  g1000 (n326, n254);
buf  g1001 (n748, n137);
buf  g1002 (n320, n203);
buf  g1003 (n632, n257);
buf  g1004 (n695, n192);
buf  g1005 (n682, n267);
buf  g1006 (n702, n228);
not  g1007 (n486, n256);
not  g1008 (n701, n171);
not  g1009 (n322, n126);
not  g1010 (n881, n144);
not  g1011 (n880, n159);
not  g1012 (n427, n163);
not  g1013 (n685, n239);
buf  g1014 (n802, n149);
buf  g1015 (n610, n100);
not  g1016 (n850, n224);
buf  g1017 (n614, n161);
buf  g1018 (n887, n253);
buf  g1019 (n481, n159);
buf  g1020 (n698, n281);
buf  g1021 (n397, n159);
buf  g1022 (n928, n257);
not  g1023 (n403, n133);
buf  g1024 (n592, n230);
not  g1025 (n874, n169);
buf  g1026 (n545, n165);
not  g1027 (n868, n112);
not  g1028 (n699, n169);
buf  g1029 (n681, n211);
buf  g1030 (n1040, n233);
buf  g1031 (n680, n218);
not  g1032 (n450, n271);
buf  g1033 (n609, n226);
buf  g1034 (n1006, n114);
buf  g1035 (n505, n229);
buf  g1036 (n526, n245);
not  g1037 (n697, n146);
buf  g1038 (n975, n97);
buf  g1039 (n432, n109);
not  g1040 (n414, n121);
not  g1041 (n318, n221);
xnor g1042 (n1254, n907, n647, n878, n963);
nand g1043 (n1133, n525, n355, n1005, n910);
xor  g1044 (n1145, n1021, n922, n946, n642);
xnor g1045 (n1294, n780, n778, n822, n875);
and  g1046 (n1299, n842, n947, n982, n863);
nor  g1047 (n1227, n755, n466, n849, n400);
or   g1048 (n1184, n894, n998, n403, n937);
xnor g1049 (n1114, n943, n992, n407, n897);
or   g1050 (n1136, n486, n663, n981, n1042);
nand g1051 (n1200, n601, n541, n590, n747);
nand g1052 (n1181, n477, n438, n851, n420);
and  g1053 (n1206, n979, n587, n876, n1018);
or   g1054 (n1230, n373, n955, n894, n928);
and  g1055 (n1126, n808, n1022, n361, n905);
xnor g1056 (n1279, n391, n449, n775, n451);
xnor g1057 (n1228, n873, n1029, n726, n654);
or   g1058 (n1298, n966, n481, n501, n1040);
nand g1059 (n1288, n995, n961, n344, n882);
xor  g1060 (n1118, n425, n903, n574, n896);
xor  g1061 (n1141, n368, n820, n898, n746);
xor  g1062 (n1068, n356, n860, n799, n510);
xnor g1063 (n1215, n872, n1036, n932, n821);
nand g1064 (n1165, n624, n976, n431, n867);
xnor g1065 (n1073, n741, n460, n395, n433);
nand g1066 (n1255, n508, n914, n1037, n524);
and  g1067 (n1175, n596, n514, n729, n763);
nand g1068 (n1143, n1009, n488, n826, n606);
xnor g1069 (n1237, n877, n823, n986, n1027);
nand g1070 (n1224, n677, n968, n318, n956);
nor  g1071 (n1067, n838, n1011, n644, n689);
xnor g1072 (n1235, n929, n1010, n963, n618);
xor  g1073 (n1193, n354, n699, n887, n444);
xor  g1074 (n1214, n389, n1019, n367, n896);
or   g1075 (n1261, n927, n529, n1000, n837);
nand g1076 (n1185, n558, n804, n803, n650);
nand g1077 (n1265, n921, n952, n936, n907);
nand g1078 (n1125, n1038, n846, n475, n450);
xnor g1079 (n1166, n539, n523, n1013, n620);
xnor g1080 (n1198, n997, n424, n551, n685);
nand g1081 (n1240, n600, n374, n405, n994);
nor  g1082 (n1088, n652, n597, n393, n352);
nor  g1083 (n1163, n678, n435, n1021, n879);
xor  g1084 (n1069, n987, n917, n519, n521);
or   g1085 (n1177, n462, n379, n483, n629);
nor  g1086 (n1062, n404, n1038, n446, n940);
nand g1087 (n1195, n975, n711, n691, n714);
or   g1088 (n1078, n968, n897, n831, n977);
nand g1089 (n1225, n871, n864, n572, n437);
nand g1090 (n1098, n912, n550, n298, n909);
xor  g1091 (n1092, n308, n328, n735, n672);
and  g1092 (n1223, n948, n1002, n967, n633);
or   g1093 (n1296, n398, n553, n957, n910);
and  g1094 (n1282, n320, n683, n1037, n964);
and  g1095 (n1239, n545, n901, n439, n826);
and  g1096 (n1274, n1006, n409, n332, n536);
xor  g1097 (n1113, n845, n939, n737, n970);
xor  g1098 (n1196, n839, n951, n700, n632);
nand g1099 (n1293, n487, n987, n1025, n829);
or   g1100 (n1263, n309, n936, n376, n930);
or   g1101 (n1083, n675, n923, n717, n532);
xor  g1102 (n1251, n421, n863, n776, n810);
nor  g1103 (n1060, n1008, n338, n1026, n748);
xnor g1104 (n1104, n578, n478, n615, n313);
or   g1105 (n1176, n1033, n331, n866, n534);
nor  g1106 (n1247, n311, n838, n415, n771);
xor  g1107 (n1065, n891, n622, n814, n779);
or   g1108 (n1142, n892, n651, n324, n441);
xnor g1109 (n1300, n859, n933, n966, n670);
xnor g1110 (n1151, n883, n975, n855, n599);
and  g1111 (n1269, n453, n761, n640, n941);
xor  g1112 (n1156, n698, n458, n323, n718);
or   g1113 (n1134, n588, n312, n1012, n934);
or   g1114 (n1087, n386, n1003, n759, n476);
xor  g1115 (n1302, n544, n563, n962, n862);
and  g1116 (n1174, n649, n315, n831, n317);
or   g1117 (n1187, n631, n984, n972, n1035);
and  g1118 (n1250, n540, n1005, n730, n1010);
xnor g1119 (n1116, n768, n870, n1018, n859);
xor  g1120 (n1095, n823, n489, n865, n888);
xor  g1121 (n1154, n837, n621, n962, n866);
nand g1122 (n1268, n656, n394, n739, n555);
nor  g1123 (n1271, n911, n904, n1034, n1001);
and  g1124 (n1130, n949, n673, n794, n360);
xnor g1125 (n1106, n750, n410, n971, n990);
xnor g1126 (n1218, n925, n983, n695, n522);
and  g1127 (n1289, n720, n1041, n719, n375);
xnor g1128 (n1257, n999, n505, n549, n772);
xnor g1129 (n1284, n942, n918, n392, n842);
and  g1130 (n1276, n874, n853, n297, n947);
xor  g1131 (n1186, n1008, n858, n445, n382);
and  g1132 (n1097, n970, n713, n828, n503);
or   g1133 (n1122, n800, n855, n591, n1025);
nor  g1134 (n1081, n628, n661, n762, n1032);
or   g1135 (n1148, n335, n547, n731, n482);
xnor g1136 (n1260, n740, n704, n494, n961);
xnor g1137 (n1192, n881, n872, n686, n834);
or   g1138 (n1270, n875, n949, n571, n364);
and  g1139 (n1281, n326, n978, n1016, n913);
nand g1140 (n1219, n758, n844, n358, n781);
xor  g1141 (n1086, n997, n369, n377, n690);
and  g1142 (n1094, n414, n793, n898, n818);
nor  g1143 (n1074, n371, n565, n416, n824);
nand g1144 (n1120, n1026, n751, n914, n638);
or   g1145 (n1117, n822, n959, n579, n960);
nand g1146 (n1064, n850, n434, n589, n383);
and  g1147 (n1217, n902, n347, n999, n378);
nor  g1148 (n1267, n497, n911, n492, n1030);
nor  g1149 (n1084, n319, n608, n680, n901);
or   g1150 (n1241, n868, n862, n417, n797);
nor  g1151 (n1101, n1002, n1031, n890, n852);
nor  g1152 (n1061, n915, n1020, n934, n296);
xor  g1153 (n1258, n969, n783, n1004, n345);
nand g1154 (n1209, n385, n725, n840, n708);
and  g1155 (n1194, n958, n457, n527, n945);
xor  g1156 (n1286, n307, n986, n769, n805);
xnor g1157 (n1155, n535, n890, n1035, n646);
xor  g1158 (n1210, n428, n641, n491, n515);
xnor g1159 (n1158, n899, n372, n869, n390);
nor  g1160 (n1202, n305, n625, n411, n350);
xor  g1161 (n1278, n639, n658, n557, n893);
or   g1162 (n1207, n959, n339, n496, n770);
nor  g1163 (n1205, n611, n880, n448, n607);
xor  g1164 (n1275, n811, n506, n353, n856);
xnor g1165 (n1301, n542, n471, n917, n452);
nand g1166 (n1180, n301, n357, n852, n697);
xnor g1167 (n1246, n990, n655, n942, n812);
xnor g1168 (n1220, n594, n692, n736, n732);
and  g1169 (n1182, n888, n696, n988, n329);
or   g1170 (n1204, n766, n325, n693, n929);
or   g1171 (n1183, n556, n1016, n773, n412);
xnor g1172 (n1256, n554, n705, n790, n971);
xor  g1173 (n1164, n703, n743, n977, n348);
xnor g1174 (n1201, n575, n485, n994, n470);
and  g1175 (n1221, n548, n653, n1032, n912);
or   g1176 (n1243, n760, n919, n848, n945);
or   g1177 (n1124, n604, n978, n876, n722);
xnor g1178 (n1160, n951, n517, n880, n370);
and  g1179 (n1208, n351, n728, n499, n363);
nand g1180 (n1197, n791, n564, n334, n1014);
nand g1181 (n1103, n566, n878, n995, n459);
and  g1182 (n1168, n464, n1028, n1029, n668);
xor  g1183 (n1262, n844, n526, n935, n342);
or   g1184 (n1093, n909, n809, n903, n388);
or   g1185 (n1090, n682, n955, n733, n724);
xor  g1186 (n1127, n512, n932, n938, n973);
and  g1187 (n1236, n889, n1007, n832, n974);
nor  g1188 (n1099, n516, n442, n681, n537);
or   g1189 (n1077, n504, n1012, n518, n833);
nor  g1190 (n1085, n687, n851, n996, n463);
nand g1191 (n1102, n669, n427, n861, n1007);
nor  g1192 (n1129, n454, n576, n965, n617);
and  g1193 (n1238, n782, n406, n847, n795);
xor  g1194 (n1100, n1020, n796, n980, n1042);
xnor g1195 (n1242, n349, n340, n1027, n937);
or   g1196 (n1280, n956, n840, n712, n627);
or   g1197 (n1253, n1019, n1028, n752, n1014);
xor  g1198 (n1229, n304, n957, n546, n785);
nand g1199 (n1082, n1039, n303, n694, n841);
and  g1200 (n1121, n365, n306, n857, n923);
or   g1201 (n1119, n813, n396, n983, n456);
nor  g1202 (n1292, n461, n1024, n568, n613);
nand g1203 (n1283, n992, n530, n467, n853);
nor  g1204 (n1203, n806, n902, n958, n916);
xor  g1205 (n1199, n850, n927, n980, n1017);
nand g1206 (n1089, n1015, n583, n996, n343);
nor  g1207 (n1273, n715, n721, n895, n336);
xnor g1208 (n1231, n1024, n819, n559, n327);
nor  g1209 (n1259, n520, n1033, n920, n1031);
nand g1210 (n1290, n674, n419, n528, n614);
xnor g1211 (n1110, n418, n786, n314, n832);
and  g1212 (n1138, n948, n884, n882, n507);
xnor g1213 (n1277, n399, n834, n801, n824);
xor  g1214 (n1107, n836, n1000, n1015, n648);
xnor g1215 (n1149, n798, n619, n605, n870);
or   g1216 (n1232, n662, n322, n401, n828);
nand g1217 (n1291, n710, n734, n592, n1003);
xor  g1218 (n1096, n905, n988, n843, n408);
xnor g1219 (n1070, n952, n561, n688, n754);
and  g1220 (n1297, n965, n889, n792, n854);
and  g1221 (n1146, n381, n538, n765, n946);
nor  g1222 (n1108, n447, n940, n436, n969);
nor  g1223 (n1135, n468, n744, n981, n742);
xor  g1224 (n1128, n933, n610, n764, n474);
nand g1225 (n1188, n849, n426, n827, n586);
xor  g1226 (n1153, n854, n702, n817, n835);
xnor g1227 (n1264, n429, n500, n684, n989);
nor  g1228 (n1171, n667, n816, n1013, n915);
nand g1229 (n1137, n954, n919, n362, n879);
nand g1230 (n1169, n387, n774, n953, n581);
nor  g1231 (n1245, n569, n665, n943, n967);
nand g1232 (n1066, n833, n964, n1036, n479);
nand g1233 (n1272, n300, n921, n580, n777);
and  g1234 (n1109, n893, n455, n830, n938);
and  g1235 (n1152, n676, n533, n380, n868);
xor  g1236 (n1249, n637, n659, n1001, n993);
xnor g1237 (n1080, n384, n636, n706, n493);
nand g1238 (n1075, n891, n593, n920, n502);
xor  g1239 (n1266, n480, n626, n321, n858);
nor  g1240 (n1091, n861, n885, n603, n820);
nand g1241 (n1287, n979, n830, n825, n660);
and  g1242 (n1190, n609, n973, n570, n998);
and  g1243 (n1123, n821, n886, n954, n860);
nand g1244 (n1159, n916, n789, n630, n757);
xor  g1245 (n1170, n974, n657, n939, n1009);
and  g1246 (n1140, n857, n869, n925, n616);
nand g1247 (n1172, n598, n359, n931, n666);
and  g1248 (n1248, n908, n341, n944, n922);
and  g1249 (n1072, n848, n982, n825, n885);
or   g1250 (n1112, n788, n723, n490, n1040);
xor  g1251 (n1105, n337, n900, n935, n422);
nand g1252 (n1173, n865, n498, n423, n873);
nor  g1253 (n1115, n924, n612, n784, n930);
or   g1254 (n1132, n991, n513, n1004, n472);
xor  g1255 (n1216, n843, n960, n991, n443);
or   g1256 (n1295, n874, n1043, n484, n432);
xor  g1257 (n1189, n552, n543, n884, n819);
xor  g1258 (n1063, n871, n926, n511);
xor  g1259 (n1226, n531, n430, n1039, n767);
nand g1260 (n1167, n867, n972, n815, n440);
xnor g1261 (n1252, n886, n756, n573, n716);
and  g1262 (n1213, n560, n299, n709, n595);
xor  g1263 (n1191, n1022, n701, n366, n856);
or   g1264 (n1244, n906, n953, n671, n918);
xnor g1265 (n1157, n738, n931, n1041, n877);
or   g1266 (n1178, n1034, n465, n835, n302);
nand g1267 (n1150, n509, n906, n864, n941);
xor  g1268 (n1234, n908, n913, n1023, n495);
or   g1269 (n1147, n807, n582, n928, n469);
nor  g1270 (n1211, n664, n802, n847, n836);
nor  g1271 (n1139, n745, n944, n333, n787);
nor  g1272 (n1161, n839, n899, n1006, n984);
nor  g1273 (n1076, n892, n1023, n634, n904);
xor  g1274 (n1131, n643, n1030, n985, n635);
and  g1275 (n1212, n827, n316, n346, n895);
and  g1276 (n1285, n330, n753, n985, n402);
nand g1277 (n1079, n883, n585, n881, n397);
nor  g1278 (n1111, n707, n413, n749, n950);
and  g1279 (n1233, n829, n584, n976, n841);
nand g1280 (n1071, n562, n577, n1017, n602);
nor  g1281 (n1179, n887, n567, n950, n924);
and  g1282 (n1222, n993, n623, n1011, n846);
and  g1283 (n1162, n989, n473, n845, n310);
and  g1284 (n1144, n900, n679, n645, n727);
xnor g1285 (n1307, n1148, n1162, n1177, n1146);
and  g1286 (n1333, n1149, n1078, n1181, n1132);
nor  g1287 (n1314, n1188, n1153, n1186, n1066);
xor  g1288 (n1326, n1139, n1080, n1169, n1196);
nor  g1289 (n1308, n1077, n1131, n1060, n1156);
xor  g1290 (n1330, n1081, n1145, n1084, n1191);
xor  g1291 (n1318, n1127, n1100, n1160, n1172);
nand g1292 (n1316, n1094, n1122, n1069, n1194);
nand g1293 (n1310, n1125, n1110, n1075, n1114);
xor  g1294 (n1306, n1165, n1157, n1120, n1092);
xnor g1295 (n1305, n1087, n1199, n1068, n1182);
xnor g1296 (n1311, n1159, n1121, n1175, n1103);
xor  g1297 (n1329, n1083, n1130, n1150, n1093);
and  g1298 (n1331, n1198, n1115, n1174, n1171);
nand g1299 (n1328, n1117, n1101, n1197, n1187);
or   g1300 (n1337, n1063, n1190, n1065, n1062);
nor  g1301 (n1321, n1189, n1129, n1070, n1089);
and  g1302 (n1332, n1135, n1099, n1123, n1167);
nand g1303 (n1334, n1163, n1128, n1090, n1088);
nor  g1304 (n1304, n1195, n1107, n1124, n1111);
nand g1305 (n1323, n1147, n1192, n1091, n1161);
or   g1306 (n1335, n1073, n1061, n1098, n1142);
nor  g1307 (n1303, n1097, n1180, n1116, n1102);
xor  g1308 (n1324, n1144, n1179, n1118, n1152);
xor  g1309 (n1312, n1106, n1178, n1071, n1096);
nor  g1310 (n1336, n1133, n1136, n1140, n1170);
xnor g1311 (n1327, n1104, n1126, n1113, n1166);
xor  g1312 (n1315, n1137, n1074, n1155, n1067);
xor  g1313 (n1320, n1119, n1072, n1158, n1085);
nand g1314 (n1325, n1076, n1183, n1105, n1064);
and  g1315 (n1313, n1082, n1168, n1108, n1184);
and  g1316 (n1322, n1109, n1095, n1164, n1185);
nor  g1317 (n1309, n1138, n1086, n1141, n1143);
nor  g1318 (n1319, n1151, n1079, n1193, n1173);
and  g1319 (n1317, n1134, n1176, n1154, n1112);
not  g1320 (n1344, n1209);
buf  g1321 (n1340, n1309);
xor  g1322 (n1343, n1204, n1307, n1208, n1211);
nor  g1323 (n1339, n1210, n1207, n1202, n1304);
nand g1324 (n1338, n1201, n1205, n1305, n1213);
and  g1325 (n1342, n1206, n1306, n1308, n1200);
xor  g1326 (n1341, n1203, n1303, n1214, n1212);
not  g1327 (n1361, n1341);
buf  g1328 (n1349, n1344);
not  g1329 (n1355, n1342);
buf  g1330 (n1367, n1342);
not  g1331 (n1353, n1341);
buf  g1332 (n1358, n1339);
buf  g1333 (n1362, n1341);
not  g1334 (n1359, n1339);
buf  g1335 (n1366, n1344);
buf  g1336 (n1350, n1338);
buf  g1337 (n1371, n1338);
buf  g1338 (n1347, n1344);
buf  g1339 (n1360, n1340);
not  g1340 (n1364, n1343);
buf  g1341 (n1370, n1341);
buf  g1342 (n1365, n1338);
buf  g1343 (n1368, n1344);
not  g1344 (n1345, n1340);
buf  g1345 (n1369, n1343);
not  g1346 (n1346, n1342);
buf  g1347 (n1357, n1342);
buf  g1348 (n1372, n1215);
buf  g1349 (n1356, n1340);
buf  g1350 (n1352, n1339);
buf  g1351 (n1354, n1340);
buf  g1352 (n1351, n1338);
buf  g1353 (n1363, n1216);
nor  g1354 (n1348, n1339, n1343);
xor  g1355 (n1389, n1354, n1351, n1363, n1230);
or   g1356 (n1387, n1351, n1367, n1361, n1368);
nor  g1357 (n1381, n1226, n1371, n1352, n1365);
and  g1358 (n1376, n1359, n1348, n1043, n1356);
nor  g1359 (n1396, n1370, n1360, n1362, n1367);
nand g1360 (n1393, n1217, n293, n1369, n1347);
or   g1361 (n1374, n1369, n1372, n1366, n1364);
nand g1362 (n1384, n1353, n1370, n1045, n1046);
and  g1363 (n1398, n1356, n1362, n1367, n1220);
or   g1364 (n1375, n1358, n1355, n1371, n1360);
and  g1365 (n1379, n1361, n1045, n1357, n1368);
nor  g1366 (n1380, n1371, n1369, n1355, n1358);
or   g1367 (n1395, n1364, n1368, n1218, n1357);
xnor g1368 (n1399, n1368, n1352, n1370, n1354);
nor  g1369 (n1386, n1348, n1358, n1347, n1359);
nand g1370 (n1391, n1221, n1365, n1219, n1222);
or   g1371 (n1402, n1359, n1371, n1346, n1364);
xnor g1372 (n1397, n1345, n1367, n1355, n1357);
xor  g1373 (n1401, n1361, n1351, n1360, n1224);
or   g1374 (n1383, n1362, n1360, n1359, n1231);
xnor g1375 (n1392, n1372, n1366, n1363, n1346);
nand g1376 (n1394, n1350, n1372, n1228, n1358);
nand g1377 (n1382, n1354, n1356, n1365);
xor  g1378 (n1378, n1363, n1372, n1370, n1350);
and  g1379 (n1390, n1366, n1356, n1364, n1353);
xnor g1380 (n1400, n1362, n1044, n1363, n1349);
or   g1381 (n1385, n1366, n1369, n1352, n1345);
nand g1382 (n1377, n1225, n1354, n1227, n1353);
nand g1383 (n1373, n1357, n1223, n1355, n1229);
nand g1384 (n1388, n1361, n1044, n1349, n1353);
buf  g1385 (n1403, n1387);
and  g1386 (n1404, n1391, n1392, n1239, n1237);
xor  g1387 (n1407, n1240, n1235, n1238, n1388);
xnor g1388 (n1406, n1236, n1393, n1234, n1241);
nand g1389 (n1405, n1389, n1233, n1232, n1390);
xnor g1390 (n1410, n1243, n1246, n1403, n1244);
or   g1391 (n1409, n1404, n1245, n1250, n1248);
or   g1392 (n1408, n1247, n1242, n1403, n1249);
nand g1393 (n1411, n1252, n1409, n1049, n1053);
nor  g1394 (n1418, n1048, n1255, n1408, n1052);
or   g1395 (n1415, n1410, n1257, n1046, n1055);
and  g1396 (n1419, n1056, n1410, n1251, n1408);
xor  g1397 (n1412, n1408, n1054, n1256, n1409);
xor  g1398 (n1420, n1052, n1253, n1254, n1409);
xnor g1399 (n1414, n1409, n1050, n1047, n1053);
nor  g1400 (n1416, n1050, n1054, n1051, n1408);
nor  g1401 (n1413, n1258, n1051, n1259, n1049);
nand g1402 (n1417, n1056, n1047, n1055, n1048);
not  g1403 (n1425, n1260);
buf  g1404 (n1423, n1411);
not  g1405 (n1424, n1413);
not  g1406 (n1422, n1412);
buf  g1407 (n1426, n1414);
buf  g1408 (n1427, n1413);
not  g1409 (n1428, n1413);
xnor g1410 (n1421, n1411, n1261, n1412);
nand g1411 (n1430, n1266, n1421, n1265, n1262);
xor  g1412 (n1429, n1264, n1421, n1263, n1267);
buf  g1413 (n1434, n1429);
not  g1414 (n1432, n1430);
buf  g1415 (n1433, n1430);
not  g1416 (n1431, n1429);
and  g1417 (n1435, n1273, n1271, n1269, n1431);
nand g1418 (n1436, n1268, n1270, n1272, n1431);
or   g1419 (n1437, n1435, n1276, n1275, n1274);
not  g1420 (n1439, n1277);
or   g1421 (n1438, n1278, n1437);
buf  g1422 (n1440, n1438);
buf  g1423 (n1441, n1279);
buf  g1424 (n1442, n1438);
not  g1425 (n1443, n1440);
and  g1426 (n1446, n1423, n1443, n1422);
and  g1427 (n1445, n1443, n1423, n1422);
or   g1428 (n1444, n1422, n1421);
not  g1429 (n1447, n1445);
not  g1430 (n1448, n1446);
or   g1431 (n1452, n1282, n1432, n1286);
xnor g1432 (n1454, n1433, n1280, n1431);
xnor g1433 (n1456, n1281, n1433, n1431);
xor  g1434 (n1455, n1447, n1410, n1434, n1283);
xor  g1435 (n1449, n1448, n1448, n1433, n1284);
xor  g1436 (n1450, n1285, n1448, n1447);
or   g1437 (n1451, n1434, n1432);
nand g1438 (n1453, n1410, n1447, n1434);
and  g1439 (n1462, n1423, n1396, n1436, n1424);
or   g1440 (n1461, n1397, n1425, n1453, n1455);
nand g1441 (n1458, n1454, n1450, n1402, n1425);
or   g1442 (n1459, n1452, n1424, n1436);
and  g1443 (n1457, n1394, n1398, n1400, n1451);
xor  g1444 (n1460, n1399, n1424, n1401, n1395);
and  g1445 (n1463, n1427, n1426, n1459);
or   g1446 (n1465, n1426, n1425, n1458);
xor  g1447 (n1464, n1426, n1427, n1457);
nor  g1448 (n1467, n1465, n1465, n1289, n1428);
nor  g1449 (n1468, n1428, n1463, n1464, n1427);
nand g1450 (n1466, n1288, n1293, n1290, n1291);
or   g1451 (n1469, n1428, n1428, n1287, n1292);
xor  g1452 (n1470, n1467, n1058, n1057);
nand g1453 (n1473, n1294, n1300, n1296, n1301);
nand g1454 (n1471, n1295, n1298, n1297, n1302);
and  g1455 (n1472, n1299, n1470);
buf  g1456 (n1477, n1472);
not  g1457 (n1476, n1473);
not  g1458 (n1475, n1471);
not  g1459 (n1474, n1473);
nor  g1460 (n1481, n1477, n1442, n1440, n1434);
and  g1461 (n1479, n1476, n294, n295);
nor  g1462 (n1478, n1474, n294, n1477);
and  g1463 (n1482, n1441, n1441, n295, n1442);
xnor g1464 (n1480, n295, n294, n293, n1475);
not  g1465 (n1485, n1482);
not  g1466 (n1483, n1480);
buf  g1467 (n1484, n1059);
not  g1468 (n1488, n1059);
nand g1469 (n1487, n1482, n1481);
xnor g1470 (n1486, n1478, n1479, n1058);
not  g1471 (n1490, n1487);
not  g1472 (n1497, n1486);
not  g1473 (n1489, n1488);
buf  g1474 (n1493, n1483);
buf  g1475 (n1492, n1486);
not  g1476 (n1496, n1484);
not  g1477 (n1495, n1488);
not  g1478 (n1494, n1485);
not  g1479 (n1491, n1487);
buf  g1480 (n1506, n1493);
not  g1481 (n1526, n1496);
not  g1482 (n1531, n1329);
buf  g1483 (n1514, n1439);
not  g1484 (n1524, n1493);
not  g1485 (n1517, n1490);
not  g1486 (n1520, n1327);
buf  g1487 (n1511, n1404);
not  g1488 (n1525, n1310);
buf  g1489 (n1519, n1311);
not  g1490 (n1529, n1334);
not  g1491 (n1515, n1496);
not  g1492 (n1518, n1493);
buf  g1493 (n1513, n1492);
buf  g1494 (n1530, n1333);
buf  g1495 (n1505, n1497);
not  g1496 (n1527, n1495);
buf  g1497 (n1507, n1336);
not  g1498 (n1503, n1405);
not  g1499 (n1523, n1495);
and  g1500 (n1512, n1407, n1337, n1494, n1497);
and  g1501 (n1516, n1494, n1496, n1312, n1495);
xnor g1502 (n1508, n1322, n1489, n1318, n1491);
and  g1503 (n1501, n1405, n1406, n1497, n1313);
and  g1504 (n1522, n1323, n1497, n1491, n1494);
nor  g1505 (n1521, n1439, n1491, n1325, n1494);
nand g1506 (n1528, n1317, n1489, n1493, n1326);
nor  g1507 (n1509, n1335, n1491, n1438, n1332);
nand g1508 (n1504, n1490, n1324, n1314, n1489);
nor  g1509 (n1498, n1489, n1492, n1316);
xnor g1510 (n1510, n1490, n1330, n1439, n1492);
xor  g1511 (n1500, n1321, n1495, n1490, n1331);
xnor g1512 (n1499, n1320, n1319, n1496, n1406);
xnor g1513 (n1502, n1439, n1407, n1315, n1328);
not  g1514 (n1563, n1521);
buf  g1515 (n1533, n1500);
not  g1516 (n1548, n1501);
buf  g1517 (n1535, n1504);
not  g1518 (n1569, n1525);
buf  g1519 (n1537, n1527);
buf  g1520 (n1568, n1531);
buf  g1521 (n1549, n1510);
buf  g1522 (n1540, n1519);
not  g1523 (n1543, n1503);
buf  g1524 (n1566, n1523);
buf  g1525 (n1558, n1530);
buf  g1526 (n1560, n1522);
not  g1527 (n1559, n1513);
not  g1528 (n1564, n1531);
not  g1529 (n1534, n1517);
not  g1530 (n1555, n1499);
not  g1531 (n1547, n1509);
buf  g1532 (n1565, n1530);
buf  g1533 (n1557, n1528);
not  g1534 (n1546, n1529);
buf  g1535 (n1551, n1512);
not  g1536 (n1545, n1498);
not  g1537 (n1570, n1527);
buf  g1538 (n1541, n1502);
buf  g1539 (n1562, n1506);
not  g1540 (n1538, n1518);
not  g1541 (n1544, n1508);
buf  g1542 (n1536, n1507);
not  g1543 (n1553, n1529);
buf  g1544 (n1554, n1526);
buf  g1545 (n1556, n1511);
not  g1546 (n1561, n1515);
buf  g1547 (n1550, n1514);
buf  g1548 (n1532, n1516);
not  g1549 (n1539, n1520);
not  g1550 (n1552, n1505);
not  g1551 (n1571, n1528);
buf  g1552 (n1542, n1524);
buf  g1553 (n1567, n1526);
nor  g1554 (n1629, n1419, n1559, n1418);
or   g1555 (n1610, n1539, n1418, n1417, n1468);
xnor g1556 (n1590, n1549, n73, n1416, n1418);
and  g1557 (n1574, n1534, n71, n73, n1535);
xor  g1558 (n1612, n1565, n1561, n81, n1539);
nand g1559 (n1606, n1539, n1558, n1542, n80);
xor  g1560 (n1622, n1547, n1543, n1566);
nor  g1561 (n1585, n75, n81, n1566, n1419);
xor  g1562 (n1587, n1547, n77, n1420);
xnor g1563 (n1626, n1565, n1551, n1547, n1554);
xor  g1564 (n1578, n81, n1416, n1563, n1540);
xnor g1565 (n1600, n1541, n1534, n1545, n1546);
and  g1566 (n1630, n1570, n1545, n1456, n1420);
or   g1567 (n1580, n84, n79, n1414, n83);
nand g1568 (n1602, n1540, n1558, n1538, n74);
nand g1569 (n1591, n1414, n1443, n1566, n1541);
xor  g1570 (n1593, n1553, n1562, n1560, n1416);
nand g1571 (n1618, n72, n70, n1533, n1542);
xnor g1572 (n1615, n1543, n1556, n1532, n1553);
nand g1573 (n1596, n1557, n1558, n72, n1556);
or   g1574 (n1598, n74, n84, n1567, n70);
or   g1575 (n1589, n1557, n78, n1569, n81);
nand g1576 (n1597, n85, n1544, n1549, n83);
and  g1577 (n1631, n1570, n82, n1569, n1461);
xnor g1578 (n1614, n1550, n75, n1414, n1543);
and  g1579 (n1620, n76, n1550, n1418, n1563);
xnor g1580 (n1628, n1557, n76, n1550, n1555);
nor  g1581 (n1625, n1555, n1543, n1536, n1542);
xor  g1582 (n1583, n1554, n85, n1415, n1536);
or   g1583 (n1584, n1535, n73, n1544, n1538);
nand g1584 (n1603, n1551, n1541, n1571, n1532);
and  g1585 (n1621, n1571, n1563, n1567, n1534);
nand g1586 (n1604, n1567, n1552, n78, n1554);
or   g1587 (n1623, n76, n79, n1541, n1564);
xor  g1588 (n1611, n1545, n1549, n1552);
xor  g1589 (n1616, n1567, n1569, n1533, n85);
xor  g1590 (n1607, n85, n1558, n1537);
xnor g1591 (n1579, n80, n83, n1420, n1547);
xor  g1592 (n1605, n1417, n75, n1550, n1534);
nand g1593 (n1575, n1568, n1571, n73, n1564);
xor  g1594 (n1635, n1419, n1571, n79, n1569);
and  g1595 (n1627, n1546, n80, n1415, n1539);
xnor g1596 (n1581, n1565, n1540, n1538, n1553);
nor  g1597 (n1592, n1532, n1570, n84, n1556);
nor  g1598 (n1633, n1561, n1536, n1548, n74);
xor  g1599 (n1608, n1557, n1554, n1537, n1551);
and  g1600 (n1572, n1536, n1565, n1552, n1556);
xnor g1601 (n1609, n1417, n1537, n1564, n1548);
xnor g1602 (n1595, n1553, n1555, n1562, n1546);
xor  g1603 (n1577, n82, n1560, n1420, n1532);
xor  g1604 (n1601, n1415, n1544, n1561, n71);
nor  g1605 (n1617, n82, n1568, n1548, n1562);
and  g1606 (n1573, n1545, n1416, n1564, n1562);
and  g1607 (n1619, n1560, n1417, n72, n77);
xor  g1608 (n1594, n1535, n79, n78, n1548);
xor  g1609 (n1632, n1535, n1533, n1546, n83);
and  g1610 (n1588, n1469, n1563, n76, n1568);
xor  g1611 (n1582, n1559, n78, n71, n82);
nand g1612 (n1634, n1540, n77, n1561, n1460);
nand g1613 (n1613, n72, n1538, n1555, n75);
or   g1614 (n1624, n1568, n74, n1570, n1419);
nand g1615 (n1586, n1533, n1462, n1415, n80);
nor  g1616 (n1576, n1551, n71, n84, n1559);
nand g1617 (n1599, n1542, n1544, n1549, n1560);
and  g1618 (n1650, n1596, n1587, n1629, n1594);
nand g1619 (n1636, n1612, n1618, n1579, n1600);
nor  g1620 (n1648, n1603, n1619, n1607, n1624);
and  g1621 (n1645, n1614, n1604, n1609, n1626);
and  g1622 (n1651, n1633, n1631, n1635, n1632);
xnor g1623 (n1649, n1634, n1584, n1576, n1601);
and  g1624 (n1642, n1581, n1617, n1595, n1583);
nor  g1625 (n1643, n1591, n1610, n1582, n1625);
nor  g1626 (n1637, n1589, n1593, n1586, n1606);
and  g1627 (n1646, n1580, n1588, n1574, n1616);
and  g1628 (n1638, n1605, n1597, n1627, n1575);
nor  g1629 (n1647, n1620, n1598, n1615, n1628);
nor  g1630 (n1641, n1592, n1622, n1572, n1599);
xor  g1631 (n1640, n1613, n1608, n1602, n1630);
and  g1632 (n1639, n1611, n1621, n1573, n1578);
xnor g1633 (n1644, n1590, n1623, n1585, n1577);
nor  g1634 (n1655, n1651, n1642, n1640, n1637);
nand g1635 (n1653, n1650, n1636, n1644, n1643);
or   g1636 (n1654, n1646, n1639, n1641, n1638);
xor  g1637 (n1652, n1649, n1648, n1645, n1647);
xor  g1638 (n1656, n1655, n1653, n1652, n1654);
endmodule
