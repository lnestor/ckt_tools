

module Stat_100_59
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n90,
  n113,
  n105,
  n89,
  n92,
  n114,
  n94,
  n118,
  n82,
  n88,
  n111,
  n102,
  n95,
  n119,
  n110,
  n93,
  n101,
  n87,
  n91,
  n97,
  n86,
  n98,
  n107,
  n106,
  n112,
  n117,
  n123,
  n130,
  n132,
  n128,
  n131,
  n129,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n90;
  output n113;
  output n105;
  output n89;
  output n92;
  output n114;
  output n94;
  output n118;
  output n82;
  output n88;
  output n111;
  output n102;
  output n95;
  output n119;
  output n110;
  output n93;
  output n101;
  output n87;
  output n91;
  output n97;
  output n86;
  output n98;
  output n107;
  output n106;
  output n112;
  output n117;
  output n123;
  output n130;
  output n132;
  output n128;
  output n131;
  output n129;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n83;
  wire n84;
  wire n85;
  wire n96;
  wire n99;
  wire n100;
  wire n103;
  wire n104;
  wire n108;
  wire n109;
  wire n115;
  wire n116;
  wire n120;
  wire n121;
  wire n122;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n68,
    n17
  );


  buf
  g1
  (
    n58,
    n30
  );


  buf
  g2
  (
    n55,
    n30
  );


  buf
  g3
  (
    n34,
    n6
  );


  not
  g4
  (
    n53,
    n31
  );


  not
  g5
  (
    n64,
    n14
  );


  buf
  g6
  (
    n63,
    n11
  );


  not
  g7
  (
    n35,
    n26
  );


  buf
  g8
  (
    KeyWire_0_13,
    n31
  );


  buf
  g9
  (
    n37,
    n5
  );


  not
  g10
  (
    n36,
    n24
  );


  buf
  g11
  (
    n61,
    n23
  );


  buf
  g12
  (
    n51,
    n32
  );


  not
  g13
  (
    n54,
    n9
  );


  not
  g14
  (
    n38,
    n18
  );


  buf
  g15
  (
    KeyWire_0_0,
    n8
  );


  buf
  g16
  (
    n44,
    n21
  );


  buf
  g17
  (
    n65,
    n7
  );


  buf
  g18
  (
    n40,
    n20
  );


  not
  g19
  (
    n56,
    n31
  );


  not
  g20
  (
    n66,
    n15
  );


  not
  g21
  (
    n49,
    n32
  );


  buf
  g22
  (
    KeyWire_0_1,
    n28
  );


  buf
  g23
  (
    n62,
    n10
  );


  not
  g24
  (
    n33,
    n13
  );


  buf
  g25
  (
    n52,
    n12
  );


  not
  g26
  (
    n43,
    n4
  );


  not
  g27
  (
    n70,
    n22
  );


  buf
  g28
  (
    n67,
    n2
  );


  buf
  g29
  (
    n59,
    n19
  );


  not
  g30
  (
    n41,
    n29
  );


  buf
  g31
  (
    n47,
    n25
  );


  not
  g32
  (
    n46,
    n30
  );


  not
  g33
  (
    n60,
    n3
  );


  not
  g34
  (
    KeyWire_0_6,
    n1
  );


  buf
  g35
  (
    n57,
    n27
  );


  buf
  g36
  (
    n45,
    n31
  );


  buf
  g37
  (
    n48,
    n32
  );


  buf
  g38
  (
    n69,
    n16
  );


  not
  g39
  (
    n73,
    n35
  );


  not
  g40
  (
    n76,
    n37
  );


  not
  g41
  (
    n75,
    n37
  );


  not
  g42
  (
    KeyWire_0_11,
    n34
  );


  not
  g43
  (
    KeyWire_0_12,
    n36
  );


  not
  g44
  (
    n77,
    n37
  );


  not
  g45
  (
    n81,
    n33
  );


  not
  g46
  (
    KeyWire_0_9,
    n36
  );


  buf
  g47
  (
    KeyWire_0_5,
    n38
  );


  not
  g48
  (
    n79,
    n36
  );


  or
  g49
  (
    n91,
    n76,
    n60,
    n72,
    n59
  );


  xor
  g50
  (
    n92,
    n60,
    n75,
    n80,
    n48
  );


  or
  g51
  (
    n106,
    n57,
    n56,
    n42,
    n74
  );


  and
  g52
  (
    KeyWire_0_8,
    n57,
    n74,
    n65,
    n44
  );


  nand
  g53
  (
    n88,
    n43,
    n47,
    n41,
    n46
  );


  or
  g54
  (
    n103,
    n57,
    n79,
    n80,
    n58
  );


  xor
  g55
  (
    n82,
    n66,
    n73,
    n46,
    n40
  );


  nand
  g56
  (
    KeyWire_0_3,
    n39,
    n58,
    n55,
    n78
  );


  xnor
  g57
  (
    n115,
    n63,
    n54,
    n56,
    n46
  );


  xor
  g58
  (
    n105,
    n66,
    n42,
    n62,
    n77
  );


  nand
  g59
  (
    n120,
    n50,
    n47,
    n40,
    n79
  );


  xnor
  g60
  (
    n87,
    n44,
    n47,
    n56,
    n49
  );


  nor
  g61
  (
    n114,
    n78,
    n81,
    n48,
    n40
  );


  or
  g62
  (
    n95,
    n51,
    n43,
    n48,
    n64
  );


  or
  g63
  (
    n108,
    n43,
    n66,
    n77,
    n42
  );


  xor
  g64
  (
    KeyWire_0_10,
    n55,
    n57,
    n74,
    n47
  );


  nand
  g65
  (
    KeyWire_0_7,
    n58,
    n63,
    n53,
    n51
  );


  nand
  g66
  (
    n113,
    n56,
    n52,
    n45,
    n75
  );


  nor
  g67
  (
    n112,
    n61,
    n53,
    n39,
    n54
  );


  or
  g68
  (
    n90,
    n50,
    n78,
    n41,
    n73
  );


  nor
  g69
  (
    KeyWire_0_15,
    n46,
    n80,
    n58,
    n49
  );


  nor
  g70
  (
    n119,
    n67,
    n78,
    n81,
    n49
  );


  xor
  g71
  (
    KeyWire_0_14,
    n48,
    n53,
    n67
  );


  xor
  g72
  (
    n110,
    n77,
    n60,
    n76,
    n44
  );


  xor
  g73
  (
    n99,
    n63,
    n50,
    n64,
    n39
  );


  and
  g74
  (
    n94,
    n79,
    n79,
    n40,
    n72
  );


  xor
  g75
  (
    n121,
    n44,
    n39,
    n67,
    n66
  );


  or
  g76
  (
    n107,
    n49,
    n73,
    n54,
    n77
  );


  or
  g77
  (
    n98,
    n61,
    n81,
    n72
  );


  nand
  g78
  (
    KeyWire_0_4,
    n74,
    n42,
    n45,
    n38
  );


  xor
  g79
  (
    n93,
    n55,
    n52,
    n68,
    n75
  );


  or
  g80
  (
    n100,
    n67,
    n50,
    n55,
    n72
  );


  and
  g81
  (
    n111,
    n65,
    n52,
    n45,
    n38
  );


  xnor
  g82
  (
    n89,
    n80,
    n59,
    n64,
    n75
  );


  or
  g83
  (
    n109,
    n76,
    n61,
    n63,
    n38
  );


  and
  g84
  (
    n96,
    n76,
    n65,
    n59,
    n41
  );


  nor
  g85
  (
    n102,
    n65,
    n61,
    n62,
    n59
  );


  xor
  g86
  (
    n118,
    n51,
    n43,
    n64,
    n54
  );


  nor
  g87
  (
    n101,
    n62,
    n62,
    n73,
    n51
  );


  nand
  g88
  (
    n85,
    n60,
    n41,
    n45,
    n52
  );


  not
  g89
  (
    n122,
    n116
  );


  not
  g90
  (
    n123,
    n120
  );


  not
  g91
  (
    KeyWire_0_2,
    n118
  );


  nand
  g92
  (
    n124,
    n117,
    n32,
    n119,
    n110
  );


  and
  g93
  (
    n125,
    n113,
    n109,
    n121,
    n115
  );


  nor
  g94
  (
    n127,
    n112,
    n114,
    n111,
    n108
  );


  nand
  g95
  (
    n130,
    n69,
    n71,
    n126,
    n125
  );


  or
  g96
  (
    n131,
    n71,
    n69
  );


  or
  g97
  (
    n128,
    n68,
    n70,
    n123,
    n69
  );


  xor
  g98
  (
    n132,
    n71,
    n68,
    n70
  );


  and
  g99
  (
    n129,
    n124,
    n70,
    n68,
    n127
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n71,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n50,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n126,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n86,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n116,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n72,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n39,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n97,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n84,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n74,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n117,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n80,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n78,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n42,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n104,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n83,
    KeyNOTWire_0_15
  );


endmodule

