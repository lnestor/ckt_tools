

module Stat_175_832
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n99,
  n113,
  n104,
  n108,
  n121,
  n116,
  n115,
  n109,
  n111,
  n107,
  n103,
  n120,
  n118,
  n185,
  n178,
  n188,
  n189,
  n192,
  n196,
  n186,
  n194,
  n193,
  n195,
  n187,
  n182,
  n179,
  n183,
  n181,
  n180,
  n190,
  n191,
  n184
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n99;output n113;output n104;output n108;output n121;output n116;output n115;output n109;output n111;output n107;output n103;output n120;output n118;output n185;output n178;output n188;output n189;output n192;output n196;output n186;output n194;output n193;output n195;output n187;output n182;output n179;output n183;output n181;output n180;output n190;output n191;output n184;
  wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n100;wire n101;wire n102;wire n105;wire n106;wire n110;wire n112;wire n114;wire n117;wire n119;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n47,
    n1
  );


  buf
  g1
  (
    n34,
    n2
  );


  not
  g2
  (
    n40,
    n2
  );


  buf
  g3
  (
    KeyWire_0_25,
    n3
  );


  buf
  g4
  (
    n43,
    n3
  );


  buf
  g5
  (
    KeyWire_0_11,
    n1
  );


  not
  g6
  (
    KeyWire_0_7,
    n7
  );


  buf
  g7
  (
    n35,
    n7
  );


  not
  g8
  (
    n28,
    n5
  );


  not
  g9
  (
    n42,
    n7
  );


  buf
  g10
  (
    KeyWire_0_24,
    n1
  );


  buf
  g11
  (
    n45,
    n8
  );


  buf
  g12
  (
    KeyWire_0_5,
    n1
  );


  buf
  g13
  (
    n23,
    n4
  );


  buf
  g14
  (
    n30,
    n4
  );


  buf
  g15
  (
    n38,
    n6
  );


  buf
  g16
  (
    KeyWire_0_15,
    n3
  );


  buf
  g17
  (
    n27,
    n6
  );


  buf
  g18
  (
    n36,
    n3
  );


  buf
  g19
  (
    n41,
    n2
  );


  not
  g20
  (
    n48,
    n4
  );


  not
  g21
  (
    n37,
    n2
  );


  not
  g22
  (
    n33,
    n5
  );


  buf
  g23
  (
    KeyWire_0_2,
    n5
  );


  not
  g24
  (
    n51,
    n5
  );


  buf
  g25
  (
    KeyWire_0_31,
    n6
  );


  not
  g26
  (
    n22,
    n4
  );


  buf
  g27
  (
    n39,
    n7
  );


  not
  g28
  (
    n29,
    n8
  );


  not
  g29
  (
    n24,
    n6
  );


  buf
  g30
  (
    n71,
    n24
  );


  not
  g31
  (
    n57,
    n22
  );


  nor
  g32
  (
    n55,
    n44,
    n42,
    n24,
    n45
  );


  xnor
  g33
  (
    n74,
    n34,
    n38,
    n37,
    n43
  );


  and
  g34
  (
    n65,
    n46,
    n23,
    n39,
    n45
  );


  and
  g35
  (
    n53,
    n24,
    n26,
    n22,
    n25
  );


  nand
  g36
  (
    n63,
    n30,
    n36,
    n46,
    n35
  );


  nor
  g37
  (
    n76,
    n23,
    n41,
    n43,
    n25
  );


  nand
  g38
  (
    n75,
    n31,
    n23,
    n38,
    n29
  );


  nand
  g39
  (
    n68,
    n47,
    n25,
    n22,
    n27
  );


  xnor
  g40
  (
    n56,
    n32,
    n33,
    n44,
    n36
  );


  or
  g41
  (
    n77,
    n26,
    n43,
    n35
  );


  and
  g42
  (
    n72,
    n48,
    n28,
    n24,
    n39
  );


  nor
  g43
  (
    n58,
    n39,
    n40,
    n47,
    n42
  );


  nand
  g44
  (
    n79,
    n30,
    n37,
    n42,
    n41
  );


  and
  g45
  (
    n78,
    n45,
    n33,
    n38,
    n29
  );


  xor
  g46
  (
    n52,
    n30,
    n26,
    n40,
    n36
  );


  xnor
  g47
  (
    n64,
    n48,
    n31,
    n36,
    n30
  );


  or
  g48
  (
    n59,
    n38,
    n43,
    n41,
    n46
  );


  xor
  g49
  (
    n54,
    n39,
    n31,
    n28,
    n22
  );


  nand
  g50
  (
    n61,
    n34,
    n27,
    n47,
    n23
  );


  xnor
  g51
  (
    n67,
    n47,
    n32,
    n33,
    n41
  );


  nand
  g52
  (
    KeyWire_0_23,
    n44,
    n46,
    n28,
    n45
  );


  xor
  g53
  (
    n70,
    n34,
    n44,
    n29,
    n37
  );


  xor
  g54
  (
    n69,
    n31,
    n33,
    n27
  );


  and
  g55
  (
    n60,
    n29,
    n34,
    n40,
    n32
  );


  and
  g56
  (
    n66,
    n32,
    n28,
    n25,
    n37
  );


  or
  g57
  (
    n62,
    n40,
    n26,
    n42,
    n35
  );


  not
  g58
  (
    n84,
    n69
  );


  buf
  g59
  (
    n99,
    n65
  );


  not
  g60
  (
    n80,
    n52
  );


  buf
  g61
  (
    n101,
    n67
  );


  not
  g62
  (
    KeyWire_0_26,
    n66
  );


  not
  g63
  (
    n91,
    n64
  );


  buf
  g64
  (
    n92,
    n59
  );


  buf
  g65
  (
    n83,
    n68
  );


  buf
  g66
  (
    KeyWire_0_21,
    n60
  );


  not
  g67
  (
    n85,
    n63
  );


  not
  g68
  (
    n81,
    n69
  );


  not
  g69
  (
    n86,
    n55
  );


  not
  g70
  (
    n87,
    n67
  );


  buf
  g71
  (
    n89,
    n56
  );


  buf
  g72
  (
    KeyWire_0_22,
    n62
  );


  not
  g73
  (
    n95,
    n61
  );


  buf
  g74
  (
    n97,
    n57
  );


  buf
  g75
  (
    n98,
    n70
  );


  buf
  g76
  (
    n100,
    n54
  );


  not
  g77
  (
    KeyWire_0_8,
    n53
  );


  not
  g78
  (
    KeyWire_0_17,
    n68
  );


  buf
  g79
  (
    n94,
    n58
  );


  not
  g80
  (
    n109,
    n49
  );


  buf
  g81
  (
    n104,
    n49
  );


  not
  g82
  (
    n121,
    n90
  );


  not
  g83
  (
    n102,
    n96
  );


  buf
  g84
  (
    n105,
    n89
  );


  buf
  g85
  (
    n111,
    n101
  );


  buf
  g86
  (
    KeyWire_0_18,
    n100
  );


  buf
  g87
  (
    KeyWire_0_20,
    n48
  );


  buf
  g88
  (
    n113,
    n92
  );


  buf
  g89
  (
    n114,
    n99
  );


  not
  g90
  (
    n115,
    n95
  );


  not
  g91
  (
    n106,
    n50
  );


  not
  g92
  (
    n110,
    n48
  );


  buf
  g93
  (
    n119,
    n82
  );


  not
  g94
  (
    n118,
    n85
  );


  not
  g95
  (
    n120,
    n81
  );


  not
  g96
  (
    n108,
    n98
  );


  not
  g97
  (
    n122,
    n97
  );


  xor
  g98
  (
    n103,
    n84,
    n49
  );


  xor
  g99
  (
    n107,
    n83,
    n91,
    n93,
    n87
  );


  and
  g100
  (
    n117,
    n94,
    n49,
    n86,
    n88
  );


  not
  g101
  (
    n138,
    n70
  );


  buf
  g102
  (
    n140,
    n8
  );


  buf
  g103
  (
    n139,
    n102
  );


  not
  g104
  (
    n135,
    n79
  );


  buf
  g105
  (
    n123,
    n78
  );


  not
  g106
  (
    n132,
    n106
  );


  buf
  g107
  (
    KeyWire_0_29,
    n118
  );


  buf
  g108
  (
    n131,
    n76
  );


  nor
  g109
  (
    n126,
    n78,
    n109,
    n77,
    n72
  );


  or
  g110
  (
    KeyWire_0_1,
    n10,
    n71,
    n107
  );


  or
  g111
  (
    n127,
    n104,
    n112,
    n8,
    n10
  );


  nor
  g112
  (
    n142,
    n120,
    n9
  );


  nand
  g113
  (
    n134,
    n73,
    n117,
    n75,
    n10
  );


  xor
  g114
  (
    KeyWire_0_27,
    n113,
    n78,
    n116,
    n77
  );


  and
  g115
  (
    n133,
    n9,
    n76,
    n103,
    n115
  );


  and
  g116
  (
    n141,
    n76,
    n76,
    n79,
    n111
  );


  or
  g117
  (
    n129,
    n114,
    n79,
    n74,
    n121
  );


  nor
  g118
  (
    n136,
    n77,
    n108,
    n78,
    n79
  );


  and
  g119
  (
    n137,
    n73,
    n74,
    n72,
    n105
  );


  and
  g120
  (
    n124,
    n75,
    n119,
    n77,
    n110
  );


  buf
  g121
  (
    n144,
    n51
  );


  nand
  g122
  (
    n151,
    n50,
    n51,
    n140
  );


  nor
  g123
  (
    n149,
    n136,
    n132,
    n135,
    n131
  );


  and
  g124
  (
    n157,
    n140,
    n137,
    n130,
    n136
  );


  xnor
  g125
  (
    KeyWire_0_19,
    n133,
    n51,
    n134,
    n138
  );


  or
  g126
  (
    n153,
    n131,
    n132,
    n137,
    n130
  );


  xnor
  g127
  (
    KeyWire_0_14,
    n131,
    n129,
    n51
  );


  xnor
  g128
  (
    n156,
    n50,
    n134,
    n139,
    n135
  );


  xor
  g129
  (
    KeyWire_0_10,
    n141,
    n137,
    n139,
    n127
  );


  xor
  g130
  (
    n159,
    n134,
    n130,
    n138,
    n125
  );


  or
  g131
  (
    KeyWire_0_4,
    n137,
    n129,
    n139,
    n132
  );


  xor
  g132
  (
    KeyWire_0_28,
    n134,
    n133,
    n131
  );


  nor
  g133
  (
    KeyWire_0_12,
    n130,
    n123,
    n136,
    n141
  );


  or
  g134
  (
    n155,
    n132,
    n124,
    n138,
    n141
  );


  nand
  g135
  (
    n147,
    n128,
    n135,
    n126
  );


  or
  g136
  (
    n150,
    n136,
    n50,
    n141,
    n129
  );


  xnor
  g137
  (
    n158,
    n133,
    n140,
    n139,
    n138
  );


  buf
  g138
  (
    n161,
    n157
  );


  nor
  g139
  (
    n164,
    n151,
    n159,
    n21
  );


  xnor
  g140
  (
    n176,
    n18,
    n15,
    n17
  );


  nand
  g141
  (
    KeyWire_0_13,
    n11,
    n150,
    n20
  );


  xor
  g142
  (
    n177,
    n149,
    n143,
    n158,
    n148
  );


  nor
  g143
  (
    n166,
    n155,
    n156,
    n157,
    n19
  );


  nor
  g144
  (
    KeyWire_0_30,
    n13,
    n11,
    n19,
    n155
  );


  xor
  g145
  (
    n167,
    n14,
    n13,
    n21,
    n147
  );


  xor
  g146
  (
    n170,
    n11,
    n12,
    n145
  );


  or
  g147
  (
    n171,
    n14,
    n13,
    n20,
    n15
  );


  xnor
  g148
  (
    KeyWire_0_0,
    n153,
    n19,
    n15,
    n16
  );


  xnor
  g149
  (
    n160,
    n159,
    n14,
    n18,
    n156
  );


  nor
  g150
  (
    n169,
    n12,
    n16,
    n152,
    n21
  );


  or
  g151
  (
    n172,
    n15,
    n158,
    n16,
    n12
  );


  nand
  g152
  (
    n175,
    n11,
    n19,
    n17,
    n13
  );


  nand
  g153
  (
    n163,
    n146,
    n16,
    n17,
    n21
  );


  xor
  g154
  (
    n162,
    n10,
    n18,
    n122
  );


  xnor
  g155
  (
    n168,
    n144,
    n14,
    n20,
    n154
  );


  nor
  g156
  (
    n180,
    n162,
    n167,
    n165,
    n170
  );


  xor
  g157
  (
    n187,
    n177,
    n166,
    n163,
    n169
  );


  or
  g158
  (
    n193,
    n169,
    n173,
    n174,
    n176
  );


  and
  g159
  (
    n183,
    n162,
    n172,
    n164,
    n142
  );


  xnor
  g160
  (
    n186,
    n164,
    n167,
    n171,
    n174
  );


  nor
  g161
  (
    n191,
    n162,
    n166,
    n175
  );


  xor
  g162
  (
    n181,
    n176,
    n165,
    n177,
    n171
  );


  nand
  g163
  (
    n192,
    n163,
    n160,
    n167
  );


  xor
  g164
  (
    n189,
    n175,
    n176,
    n171,
    n160
  );


  nor
  g165
  (
    n195,
    n170,
    n165,
    n172,
    n142
  );


  nor
  g166
  (
    KeyWire_0_6,
    n174,
    n142,
    n170,
    n172
  );


  nand
  g167
  (
    n188,
    n171,
    n165,
    n168,
    n161
  );


  xnor
  g168
  (
    KeyWire_0_9,
    n173,
    n160,
    n172,
    n175
  );


  xnor
  g169
  (
    n185,
    n168,
    n170,
    n169,
    n174
  );


  or
  g170
  (
    n179,
    n173,
    n164,
    n168
  );


  nand
  g171
  (
    n182,
    n175,
    n177,
    n161,
    n167
  );


  nand
  g172
  (
    KeyWire_0_3,
    n168,
    n162,
    n163,
    n173
  );


  xor
  g173
  (
    KeyWire_0_16,
    n161,
    n161,
    n166,
    n169
  );


  nand
  g174
  (
    n190,
    n177,
    n163,
    n176,
    n142
  );


  xor
  KeyGate_0_0
  (
    n174,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n125,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n49,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n194,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n143,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n25,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n178,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n32,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n82,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n196,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n145,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n46,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n146,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n173,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n154,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n44,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n184,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n88,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n112,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n148,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n116,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n93,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n96,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n73,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n50,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n26,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n90,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n130,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n152,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n128,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n165,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n31,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


