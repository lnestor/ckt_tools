

module Stat_1647_33_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n1129,
  n1121,
  n1189,
  n1199,
  n1204,
  n1213,
  n1202,
  n1211,
  n1206,
  n1205,
  n1208,
  n1210,
  n1200,
  n1209,
  n1252,
  n1250,
  n1251,
  n1665,
  n1664,
  n1662,
  n1663,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n1129;
  output n1121;
  output n1189;
  output n1199;
  output n1204;
  output n1213;
  output n1202;
  output n1211;
  output n1206;
  output n1205;
  output n1208;
  output n1210;
  output n1200;
  output n1209;
  output n1252;
  output n1250;
  output n1251;
  output n1665;
  output n1664;
  output n1662;
  output n1663;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1201;
  wire n1203;
  wire n1207;
  wire n1212;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    n32,
    n2
  );


  not
  g1
  (
    n28,
    n4
  );


  not
  g2
  (
    n77,
    n17
  );


  not
  g3
  (
    n90,
    n15
  );


  buf
  g4
  (
    n27,
    n16
  );


  buf
  g5
  (
    n26,
    n5
  );


  buf
  g6
  (
    n56,
    n9
  );


  not
  g7
  (
    n23,
    n10
  );


  buf
  g8
  (
    n69,
    n1
  );


  buf
  g9
  (
    n30,
    n6
  );


  not
  g10
  (
    n43,
    n18
  );


  not
  g11
  (
    n39,
    n10
  );


  buf
  g12
  (
    n70,
    n14
  );


  buf
  g13
  (
    n41,
    n14
  );


  buf
  g14
  (
    n80,
    n15
  );


  not
  g15
  (
    n40,
    n3
  );


  buf
  g16
  (
    n87,
    n7
  );


  not
  g17
  (
    n86,
    n4
  );


  buf
  g18
  (
    n37,
    n12
  );


  buf
  g19
  (
    n34,
    n5
  );


  buf
  g20
  (
    n79,
    n18
  );


  buf
  g21
  (
    n57,
    n13
  );


  buf
  g22
  (
    n76,
    n13
  );


  buf
  g23
  (
    n82,
    n10
  );


  buf
  g24
  (
    n60,
    n12
  );


  not
  g25
  (
    n49,
    n16
  );


  not
  g26
  (
    n19,
    n18
  );


  buf
  g27
  (
    n21,
    n17
  );


  not
  g28
  (
    n81,
    n11
  );


  buf
  g29
  (
    n45,
    n8
  );


  buf
  g30
  (
    n42,
    n16
  );


  buf
  g31
  (
    n51,
    n2
  );


  not
  g32
  (
    n84,
    n7
  );


  not
  g33
  (
    n55,
    n7
  );


  not
  g34
  (
    n33,
    n12
  );


  not
  g35
  (
    n20,
    n11
  );


  buf
  g36
  (
    n50,
    n6
  );


  not
  g37
  (
    n73,
    n8
  );


  not
  g38
  (
    n66,
    n15
  );


  buf
  g39
  (
    n36,
    n5
  );


  not
  g40
  (
    n67,
    n5
  );


  not
  g41
  (
    n85,
    n3
  );


  buf
  g42
  (
    n31,
    n17
  );


  buf
  g43
  (
    n62,
    n6
  );


  buf
  g44
  (
    n47,
    n9
  );


  buf
  g45
  (
    n25,
    n11
  );


  not
  g46
  (
    n38,
    n10
  );


  buf
  g47
  (
    n65,
    n6
  );


  not
  g48
  (
    n35,
    n12
  );


  buf
  g49
  (
    n68,
    n14
  );


  buf
  g50
  (
    n22,
    n16
  );


  buf
  g51
  (
    KeyWire_0_12,
    n15
  );


  buf
  g52
  (
    n52,
    n1
  );


  buf
  g53
  (
    n89,
    n3
  );


  not
  g54
  (
    n46,
    n4
  );


  not
  g55
  (
    n72,
    n1
  );


  buf
  g56
  (
    n53,
    n8
  );


  buf
  g57
  (
    KeyWire_0_45,
    n17
  );


  buf
  g58
  (
    n74,
    n13
  );


  not
  g59
  (
    n61,
    n4
  );


  not
  g60
  (
    n48,
    n18
  );


  buf
  g61
  (
    n44,
    n9
  );


  not
  g62
  (
    n64,
    n11
  );


  buf
  g63
  (
    n75,
    n2
  );


  buf
  g64
  (
    n58,
    n2
  );


  not
  g65
  (
    n71,
    n3
  );


  not
  g66
  (
    n54,
    n13
  );


  buf
  g67
  (
    n88,
    n14
  );


  buf
  g68
  (
    n24,
    n7
  );


  not
  g69
  (
    n63,
    n8
  );


  not
  g70
  (
    n78,
    n9
  );


  not
  g71
  (
    n83,
    n1
  );


  buf
  g72
  (
    n337,
    n55
  );


  not
  g73
  (
    n230,
    n23
  );


  buf
  g74
  (
    n276,
    n43
  );


  buf
  g75
  (
    n115,
    n82
  );


  not
  g76
  (
    n199,
    n64
  );


  not
  g77
  (
    n211,
    n85
  );


  not
  g78
  (
    n328,
    n76
  );


  buf
  g79
  (
    n253,
    n56
  );


  buf
  g80
  (
    n270,
    n59
  );


  not
  g81
  (
    n356,
    n47
  );


  buf
  g82
  (
    n171,
    n89
  );


  buf
  g83
  (
    n235,
    n42
  );


  not
  g84
  (
    n279,
    n77
  );


  not
  g85
  (
    n301,
    n55
  );


  buf
  g86
  (
    n358,
    n42
  );


  buf
  g87
  (
    n272,
    n89
  );


  not
  g88
  (
    KeyWire_0_25,
    n48
  );


  buf
  g89
  (
    n158,
    n66
  );


  not
  g90
  (
    n225,
    n27
  );


  not
  g91
  (
    n333,
    n60
  );


  buf
  g92
  (
    KeyWire_0_19,
    n34
  );


  buf
  g93
  (
    n334,
    n87
  );


  not
  g94
  (
    n317,
    n37
  );


  buf
  g95
  (
    n169,
    n66
  );


  buf
  g96
  (
    n273,
    n20
  );


  not
  g97
  (
    n193,
    n32
  );


  not
  g98
  (
    n331,
    n75
  );


  buf
  g99
  (
    n179,
    n67
  );


  buf
  g100
  (
    n101,
    n77
  );


  buf
  g101
  (
    n350,
    n63
  );


  not
  g102
  (
    n281,
    n82
  );


  not
  g103
  (
    n265,
    n58
  );


  buf
  g104
  (
    n91,
    n58
  );


  not
  g105
  (
    n367,
    n26
  );


  buf
  g106
  (
    n113,
    n73
  );


  not
  g107
  (
    n355,
    n77
  );


  not
  g108
  (
    n156,
    n27
  );


  buf
  g109
  (
    n251,
    n66
  );


  buf
  g110
  (
    n345,
    n40
  );


  buf
  g111
  (
    n292,
    n41
  );


  buf
  g112
  (
    n255,
    n67
  );


  not
  g113
  (
    n238,
    n78
  );


  not
  g114
  (
    n149,
    n61
  );


  not
  g115
  (
    n141,
    n69
  );


  buf
  g116
  (
    n336,
    n46
  );


  not
  g117
  (
    n216,
    n87
  );


  not
  g118
  (
    n252,
    n19
  );


  buf
  g119
  (
    n243,
    n44
  );


  buf
  g120
  (
    n326,
    n61
  );


  not
  g121
  (
    n342,
    n80
  );


  not
  g122
  (
    n201,
    n51
  );


  not
  g123
  (
    n363,
    n50
  );


  buf
  g124
  (
    n283,
    n47
  );


  buf
  g125
  (
    n286,
    n43
  );


  not
  g126
  (
    n239,
    n38
  );


  not
  g127
  (
    n190,
    n19
  );


  not
  g128
  (
    n200,
    n62
  );


  not
  g129
  (
    KeyWire_0_15,
    n86
  );


  not
  g130
  (
    n232,
    n50
  );


  not
  g131
  (
    n366,
    n71
  );


  not
  g132
  (
    n347,
    n81
  );


  buf
  g133
  (
    n204,
    n45
  );


  buf
  g134
  (
    n118,
    n47
  );


  not
  g135
  (
    n185,
    n83
  );


  not
  g136
  (
    n268,
    n37
  );


  not
  g137
  (
    n192,
    n42
  );


  buf
  g138
  (
    n96,
    n89
  );


  buf
  g139
  (
    n145,
    n32
  );


  not
  g140
  (
    n140,
    n36
  );


  buf
  g141
  (
    n175,
    n34
  );


  buf
  g142
  (
    n344,
    n37
  );


  buf
  g143
  (
    KeyWire_0_41,
    n87
  );


  not
  g144
  (
    n189,
    n40
  );


  not
  g145
  (
    n330,
    n47
  );


  not
  g146
  (
    n92,
    n49
  );


  buf
  g147
  (
    n123,
    n39
  );


  not
  g148
  (
    n137,
    n28
  );


  not
  g149
  (
    n332,
    n79
  );


  buf
  g150
  (
    n129,
    n68
  );


  buf
  g151
  (
    n150,
    n84
  );


  not
  g152
  (
    n100,
    n24
  );


  buf
  g153
  (
    n320,
    n21
  );


  not
  g154
  (
    n260,
    n46
  );


  buf
  g155
  (
    KeyWire_0_46,
    n75
  );


  not
  g156
  (
    n146,
    n30
  );


  not
  g157
  (
    n148,
    n60
  );


  buf
  g158
  (
    n289,
    n71
  );


  not
  g159
  (
    n98,
    n49
  );


  buf
  g160
  (
    n215,
    n72
  );


  not
  g161
  (
    n119,
    n48
  );


  buf
  g162
  (
    n109,
    n64
  );


  buf
  g163
  (
    n174,
    n90
  );


  buf
  g164
  (
    n304,
    n52
  );


  buf
  g165
  (
    n284,
    n59
  );


  not
  g166
  (
    n288,
    n62
  );


  not
  g167
  (
    KeyWire_0_63,
    n34
  );


  buf
  g168
  (
    n209,
    n40
  );


  not
  g169
  (
    n138,
    n60
  );


  not
  g170
  (
    n143,
    n45
  );


  not
  g171
  (
    n324,
    n72
  );


  not
  g172
  (
    n142,
    n50
  );


  buf
  g173
  (
    n133,
    n38
  );


  not
  g174
  (
    n349,
    n84
  );


  buf
  g175
  (
    n340,
    n76
  );


  buf
  g176
  (
    n160,
    n33
  );


  buf
  g177
  (
    n130,
    n45
  );


  not
  g178
  (
    n110,
    n30
  );


  not
  g179
  (
    n343,
    n80
  );


  not
  g180
  (
    n97,
    n74
  );


  not
  g181
  (
    n170,
    n56
  );


  not
  g182
  (
    n357,
    n70
  );


  not
  g183
  (
    n106,
    n69
  );


  buf
  g184
  (
    n335,
    n20
  );


  buf
  g185
  (
    n147,
    n79
  );


  buf
  g186
  (
    n229,
    n35
  );


  buf
  g187
  (
    n151,
    n49
  );


  buf
  g188
  (
    n233,
    n58
  );


  buf
  g189
  (
    n315,
    n86
  );


  buf
  g190
  (
    n261,
    n88
  );


  not
  g191
  (
    n371,
    n79
  );


  buf
  g192
  (
    n295,
    n37
  );


  not
  g193
  (
    n221,
    n43
  );


  not
  g194
  (
    n132,
    n32
  );


  buf
  g195
  (
    n307,
    n84
  );


  not
  g196
  (
    n325,
    n23
  );


  not
  g197
  (
    n236,
    n85
  );


  buf
  g198
  (
    n165,
    n63
  );


  buf
  g199
  (
    n202,
    n73
  );


  not
  g200
  (
    n114,
    n85
  );


  not
  g201
  (
    n181,
    n40
  );


  not
  g202
  (
    n302,
    n72
  );


  buf
  g203
  (
    n353,
    n69
  );


  buf
  g204
  (
    n122,
    n62
  );


  not
  g205
  (
    n254,
    n76
  );


  not
  g206
  (
    n184,
    n33
  );


  buf
  g207
  (
    n212,
    n65
  );


  buf
  g208
  (
    n362,
    n22
  );


  not
  g209
  (
    n319,
    n76
  );


  buf
  g210
  (
    n213,
    n84
  );


  not
  g211
  (
    n197,
    n75
  );


  not
  g212
  (
    n188,
    n51
  );


  not
  g213
  (
    n274,
    n50
  );


  buf
  g214
  (
    n364,
    n65
  );


  not
  g215
  (
    n378,
    n27
  );


  buf
  g216
  (
    n126,
    n24
  );


  buf
  g217
  (
    n178,
    n38
  );


  buf
  g218
  (
    n368,
    n75
  );


  not
  g219
  (
    n285,
    n70
  );


  not
  g220
  (
    n127,
    n20
  );


  buf
  g221
  (
    n280,
    n28
  );


  not
  g222
  (
    n191,
    n19
  );


  buf
  g223
  (
    n168,
    n61
  );


  buf
  g224
  (
    n316,
    n83
  );


  buf
  g225
  (
    n256,
    n57
  );


  not
  g226
  (
    n308,
    n74
  );


  not
  g227
  (
    n154,
    n54
  );


  buf
  g228
  (
    n300,
    n39
  );


  buf
  g229
  (
    n263,
    n33
  );


  buf
  g230
  (
    n278,
    n36
  );


  buf
  g231
  (
    n206,
    n65
  );


  not
  g232
  (
    n266,
    n32
  );


  buf
  g233
  (
    n242,
    n83
  );


  buf
  g234
  (
    n205,
    n26
  );


  not
  g235
  (
    n176,
    n30
  );


  not
  g236
  (
    n282,
    n67
  );


  not
  g237
  (
    n348,
    n81
  );


  not
  g238
  (
    n103,
    n31
  );


  buf
  g239
  (
    n359,
    n51
  );


  not
  g240
  (
    n291,
    n62
  );


  buf
  g241
  (
    n155,
    n26
  );


  buf
  g242
  (
    n226,
    n88
  );


  buf
  g243
  (
    n218,
    n53
  );


  not
  g244
  (
    KeyWire_0_51,
    n89
  );


  not
  g245
  (
    n246,
    n73
  );


  not
  g246
  (
    n93,
    n44
  );


  not
  g247
  (
    n370,
    n68
  );


  buf
  g248
  (
    n102,
    n80
  );


  buf
  g249
  (
    n214,
    n23
  );


  not
  g250
  (
    n167,
    n52
  );


  not
  g251
  (
    n157,
    n78
  );


  buf
  g252
  (
    n352,
    n21
  );


  not
  g253
  (
    n94,
    n44
  );


  buf
  g254
  (
    n241,
    n56
  );


  buf
  g255
  (
    n135,
    n54
  );


  buf
  g256
  (
    n108,
    n73
  );


  buf
  g257
  (
    n271,
    n63
  );


  not
  g258
  (
    n309,
    n69
  );


  not
  g259
  (
    n318,
    n29
  );


  buf
  g260
  (
    n163,
    n55
  );


  not
  g261
  (
    n338,
    n44
  );


  not
  g262
  (
    n240,
    n46
  );


  buf
  g263
  (
    n104,
    n82
  );


  buf
  g264
  (
    n322,
    n25
  );


  not
  g265
  (
    n267,
    n64
  );


  buf
  g266
  (
    n287,
    n60
  );


  buf
  g267
  (
    n296,
    n45
  );


  not
  g268
  (
    n245,
    n30
  );


  buf
  g269
  (
    n258,
    n35
  );


  buf
  g270
  (
    n365,
    n57
  );


  buf
  g271
  (
    n196,
    n21
  );


  buf
  g272
  (
    n327,
    n23
  );


  not
  g273
  (
    n161,
    n71
  );


  buf
  g274
  (
    n231,
    n59
  );


  not
  g275
  (
    n220,
    n28
  );


  not
  g276
  (
    n227,
    n88
  );


  buf
  g277
  (
    n341,
    n27
  );


  not
  g278
  (
    n298,
    n81
  );


  not
  g279
  (
    n257,
    n74
  );


  not
  g280
  (
    n360,
    n66
  );


  buf
  g281
  (
    n290,
    n80
  );


  not
  g282
  (
    n259,
    n39
  );


  not
  g283
  (
    n248,
    n74
  );


  buf
  g284
  (
    n262,
    n36
  );


  buf
  g285
  (
    n210,
    n72
  );


  not
  g286
  (
    n346,
    n38
  );


  buf
  g287
  (
    n306,
    n68
  );


  buf
  g288
  (
    n173,
    n77
  );


  buf
  g289
  (
    n303,
    n31
  );


  buf
  g290
  (
    n269,
    n19
  );


  not
  g291
  (
    n310,
    n34
  );


  not
  g292
  (
    n124,
    n53
  );


  buf
  g293
  (
    n152,
    n90
  );


  buf
  g294
  (
    n139,
    n82
  );


  buf
  g295
  (
    n217,
    n88
  );


  buf
  g296
  (
    n117,
    n68
  );


  not
  g297
  (
    n120,
    n54
  );


  buf
  g298
  (
    n186,
    n35
  );


  not
  g299
  (
    n264,
    n25
  );


  buf
  g300
  (
    n195,
    n24
  );


  buf
  g301
  (
    n329,
    n90
  );


  buf
  g302
  (
    n321,
    n25
  );


  buf
  g303
  (
    n159,
    n57
  );


  not
  g304
  (
    n111,
    n24
  );


  not
  g305
  (
    n228,
    n28
  );


  not
  g306
  (
    n237,
    n85
  );


  not
  g307
  (
    n361,
    n29
  );


  not
  g308
  (
    n105,
    n41
  );


  not
  g309
  (
    KeyWire_0_28,
    n43
  );


  not
  g310
  (
    n224,
    n53
  );


  buf
  g311
  (
    n112,
    n26
  );


  not
  g312
  (
    n277,
    n39
  );


  not
  g313
  (
    n323,
    n56
  );


  buf
  g314
  (
    n275,
    n41
  );


  not
  g315
  (
    n183,
    n48
  );


  buf
  g316
  (
    n297,
    n53
  );


  buf
  g317
  (
    n95,
    n35
  );


  buf
  g318
  (
    KeyWire_0_1,
    n33
  );


  not
  g319
  (
    n131,
    n86
  );


  buf
  g320
  (
    n377,
    n65
  );


  buf
  g321
  (
    n299,
    n63
  );


  not
  g322
  (
    KeyWire_0_21,
    n48
  );


  buf
  g323
  (
    n250,
    n21
  );


  not
  g324
  (
    n194,
    n29
  );


  not
  g325
  (
    n164,
    n57
  );


  buf
  g326
  (
    n373,
    n29
  );


  buf
  g327
  (
    n312,
    n42
  );


  not
  g328
  (
    n134,
    n22
  );


  not
  g329
  (
    n153,
    n31
  );


  not
  g330
  (
    n187,
    n59
  );


  buf
  g331
  (
    KeyWire_0_35,
    n25
  );


  not
  g332
  (
    n172,
    n22
  );


  buf
  g333
  (
    n351,
    n41
  );


  not
  g334
  (
    n116,
    n71
  );


  not
  g335
  (
    n293,
    n58
  );


  not
  g336
  (
    n203,
    n83
  );


  not
  g337
  (
    n219,
    n61
  );


  not
  g338
  (
    n374,
    n90
  );


  not
  g339
  (
    n162,
    n67
  );


  not
  g340
  (
    n311,
    n46
  );


  buf
  g341
  (
    n166,
    n51
  );


  buf
  g342
  (
    n294,
    n86
  );


  not
  g343
  (
    n180,
    n64
  );


  not
  g344
  (
    n244,
    n20
  );


  buf
  g345
  (
    n208,
    n81
  );


  not
  g346
  (
    n198,
    n22
  );


  buf
  g347
  (
    n372,
    n78
  );


  buf
  g348
  (
    n247,
    n52
  );


  not
  g349
  (
    n182,
    n78
  );


  buf
  g350
  (
    n177,
    n70
  );


  buf
  g351
  (
    n305,
    n79
  );


  buf
  g352
  (
    n314,
    n70
  );


  not
  g353
  (
    n375,
    n54
  );


  buf
  g354
  (
    n128,
    n31
  );


  not
  g355
  (
    n144,
    n49
  );


  buf
  g356
  (
    n121,
    n55
  );


  not
  g357
  (
    n376,
    n87
  );


  buf
  g358
  (
    n222,
    n52
  );


  buf
  g359
  (
    n99,
    n36
  );


  nand
  g360
  (
    n599,
    n232,
    n112,
    n241,
    n289
  );


  xnor
  g361
  (
    n382,
    n289,
    n256,
    n237,
    n206
  );


  nand
  g362
  (
    n495,
    n204,
    n309,
    n176,
    n290
  );


  nand
  g363
  (
    KeyWire_0_16,
    n140,
    n145,
    n245,
    n364
  );


  nand
  g364
  (
    n551,
    n366,
    n252,
    n351,
    n247
  );


  nor
  g365
  (
    n535,
    n197,
    n217,
    n315,
    n151
  );


  nand
  g366
  (
    n416,
    n166,
    n169,
    n250,
    n91
  );


  nand
  g367
  (
    n480,
    n235,
    n143,
    n199,
    n179
  );


  or
  g368
  (
    n554,
    n319,
    n192,
    n295,
    n115
  );


  nand
  g369
  (
    n544,
    n124,
    n320,
    n255,
    n160
  );


  nor
  g370
  (
    n543,
    n199,
    n93,
    n277,
    n286
  );


  nand
  g371
  (
    n542,
    n339,
    n207,
    n103,
    n248
  );


  and
  g372
  (
    n386,
    n295,
    n226,
    n232,
    n254
  );


  xor
  g373
  (
    n379,
    n308,
    n113,
    n259,
    n327
  );


  and
  g374
  (
    n408,
    n355,
    n341,
    n208,
    n360
  );


  and
  g375
  (
    n517,
    n257,
    n125,
    n322,
    n263
  );


  xor
  g376
  (
    n385,
    n363,
    n290,
    n244,
    n96
  );


  xor
  g377
  (
    n510,
    n264,
    n345,
    n359,
    n193
  );


  or
  g378
  (
    n552,
    n120,
    n304,
    n336,
    n279
  );


  nand
  g379
  (
    n420,
    n210,
    n296,
    n219,
    n285
  );


  nand
  g380
  (
    n598,
    n139,
    n258,
    n206,
    n211
  );


  and
  g381
  (
    n575,
    n311,
    n187,
    n274,
    n278
  );


  nand
  g382
  (
    n567,
    n216,
    n355,
    n327,
    n361
  );


  nor
  g383
  (
    n566,
    n353,
    n271,
    n98,
    n122
  );


  nand
  g384
  (
    n569,
    n288,
    n348,
    n350,
    n234
  );


  xnor
  g385
  (
    n450,
    n267,
    n361,
    n111,
    n100
  );


  or
  g386
  (
    n458,
    n333,
    n230,
    n95,
    n215
  );


  xnor
  g387
  (
    n426,
    n231,
    n216,
    n335,
    n341
  );


  or
  g388
  (
    n391,
    n354,
    n271,
    n230,
    n109
  );


  nand
  g389
  (
    n445,
    n175,
    n199,
    n287,
    n260
  );


  nand
  g390
  (
    n577,
    n257,
    n332,
    n340,
    n178
  );


  nor
  g391
  (
    n568,
    n167,
    n228,
    n196,
    n349
  );


  or
  g392
  (
    n380,
    n203,
    n242,
    n236,
    n271
  );


  and
  g393
  (
    n425,
    n326,
    n286,
    n212,
    n201
  );


  xor
  g394
  (
    n438,
    n225,
    n138,
    n243,
    n272
  );


  xor
  g395
  (
    n466,
    n168,
    n264,
    n311,
    n196
  );


  xnor
  g396
  (
    n455,
    n297,
    n346,
    n218,
    n349
  );


  xor
  g397
  (
    n459,
    n260,
    n232,
    n316,
    n194
  );


  and
  g398
  (
    n484,
    n198,
    n343,
    n312,
    n239
  );


  and
  g399
  (
    n605,
    n102,
    n161,
    n213,
    n324
  );


  nor
  g400
  (
    n468,
    n273,
    n249,
    n278,
    n229
  );


  or
  g401
  (
    n550,
    n135,
    n349,
    n119,
    n316
  );


  xnor
  g402
  (
    n487,
    n349,
    n330,
    n367,
    n240
  );


  xor
  g403
  (
    n584,
    n317,
    n165,
    n229,
    n219
  );


  xnor
  g404
  (
    n483,
    n229,
    n325,
    n285,
    n338
  );


  and
  g405
  (
    n574,
    n297,
    n133,
    n278,
    n197
  );


  nand
  g406
  (
    n443,
    n262,
    n156,
    n323,
    n300
  );


  nand
  g407
  (
    n448,
    n227,
    n346,
    n182,
    n264
  );


  xnor
  g408
  (
    n580,
    n191,
    n200,
    n294,
    n338
  );


  xnor
  g409
  (
    n496,
    n142,
    n301,
    n344,
    n139
  );


  xnor
  g410
  (
    n406,
    n358,
    n231,
    n266,
    n162
  );


  and
  g411
  (
    n430,
    n280,
    n264,
    n331,
    n279
  );


  or
  g412
  (
    n428,
    n312,
    n155,
    n116,
    n173
  );


  nor
  g413
  (
    n515,
    n347,
    n355,
    n131,
    n315
  );


  or
  g414
  (
    n431,
    n100,
    n247,
    n108,
    n334
  );


  xor
  g415
  (
    n593,
    n313,
    n222,
    n273,
    n279
  );


  xor
  g416
  (
    n446,
    n328,
    n280,
    n167,
    n230
  );


  nor
  g417
  (
    n507,
    n135,
    n99,
    n359,
    n257
  );


  xor
  g418
  (
    n525,
    n361,
    n270,
    n251,
    n303
  );


  xnor
  g419
  (
    n427,
    n203,
    n95,
    n313,
    n284
  );


  xor
  g420
  (
    n573,
    n294,
    n308,
    n200,
    n272
  );


  nor
  g421
  (
    n475,
    n154,
    n364,
    n262,
    n328
  );


  xor
  g422
  (
    n479,
    n289,
    n266,
    n187,
    n104
  );


  nor
  g423
  (
    n418,
    n283,
    n333,
    n336,
    n302
  );


  nand
  g424
  (
    n444,
    n282,
    n272,
    n292,
    n353
  );


  xor
  g425
  (
    n583,
    n204,
    n203,
    n312,
    n294
  );


  nand
  g426
  (
    n541,
    n283,
    n346,
    n157,
    n344
  );


  nand
  g427
  (
    n465,
    n309,
    n185,
    n276,
    n366
  );


  nor
  g428
  (
    n493,
    n297,
    n363,
    n321,
    n288
  );


  xnor
  g429
  (
    n460,
    n255,
    n350,
    n235,
    n180
  );


  and
  g430
  (
    n595,
    n205,
    n207,
    n194,
    n145
  );


  xnor
  g431
  (
    n486,
    n171,
    n244,
    n172,
    n207
  );


  nand
  g432
  (
    n502,
    n132,
    n365,
    n243,
    n191
  );


  xor
  g433
  (
    n530,
    n342,
    n144,
    n152,
    n107
  );


  nor
  g434
  (
    n451,
    n152,
    n189,
    n195,
    n257
  );


  xor
  g435
  (
    n539,
    n227,
    n354,
    n113,
    n105
  );


  or
  g436
  (
    n453,
    n325,
    n178,
    n316,
    n210
  );


  xnor
  g437
  (
    n531,
    n116,
    n334,
    n207,
    n298
  );


  nor
  g438
  (
    n399,
    n210,
    n218,
    n293,
    n198
  );


  nor
  g439
  (
    n547,
    n327,
    n296,
    n293,
    n231
  );


  or
  g440
  (
    n602,
    n193,
    n341,
    n360,
    n265
  );


  or
  g441
  (
    n508,
    n110,
    n220,
    n228,
    n241
  );


  nor
  g442
  (
    n601,
    n240,
    n233,
    n177,
    n222
  );


  and
  g443
  (
    n402,
    n281,
    n193,
    n190,
    n208
  );


  nand
  g444
  (
    n506,
    n194,
    n293,
    n131,
    n249
  );


  and
  g445
  (
    n536,
    n158,
    n269,
    n295,
    n136
  );


  or
  g446
  (
    n590,
    n310,
    n147,
    n261,
    n196
  );


  nand
  g447
  (
    n589,
    n284,
    n118,
    n242,
    n164
  );


  or
  g448
  (
    n548,
    n314,
    n322,
    n117,
    n142
  );


  nor
  g449
  (
    n457,
    n158,
    n215,
    n317,
    n305
  );


  xnor
  g450
  (
    n404,
    n268,
    n216,
    n305,
    n103
  );


  xnor
  g451
  (
    n560,
    n224,
    n220,
    n261,
    n251
  );


  nand
  g452
  (
    n557,
    n271,
    n272,
    n275,
    n159
  );


  or
  g453
  (
    n519,
    n237,
    n343,
    n323,
    n290
  );


  or
  g454
  (
    n534,
    n297,
    n315,
    n223,
    n119
  );


  xor
  g455
  (
    n389,
    n326,
    n362,
    n233,
    n241
  );


  xor
  g456
  (
    n415,
    n284,
    n277,
    n228,
    n120
  );


  nor
  g457
  (
    n556,
    n296,
    n110,
    n308,
    n214
  );


  xor
  g458
  (
    n527,
    n236,
    n97,
    n192,
    n324
  );


  nand
  g459
  (
    n481,
    n303,
    n331,
    n246,
    n202
  );


  xor
  g460
  (
    n395,
    n192,
    n356,
    n220,
    n300
  );


  and
  g461
  (
    n565,
    n327,
    n286,
    n197,
    n209
  );


  xnor
  g462
  (
    n434,
    n305,
    n200,
    n265,
    n101
  );


  xor
  g463
  (
    n478,
    n317,
    n300,
    n241,
    n206
  );


  or
  g464
  (
    n520,
    n310,
    n183,
    n141,
    n247
  );


  xnor
  g465
  (
    n581,
    n115,
    n277,
    n240,
    n237
  );


  xnor
  g466
  (
    n410,
    n195,
    n185,
    n225,
    n334
  );


  and
  g467
  (
    n473,
    n226,
    n251,
    n302,
    n270
  );


  or
  g468
  (
    n436,
    n348,
    n329,
    n188,
    n209
  );


  nand
  g469
  (
    n559,
    n219,
    n326,
    n200,
    n176
  );


  or
  g470
  (
    n488,
    n318,
    n329,
    n285,
    n210
  );


  nor
  g471
  (
    n526,
    n223,
    n248,
    n243,
    n268
  );


  nand
  g472
  (
    n503,
    n284,
    n275,
    n184,
    n269
  );


  nand
  g473
  (
    n498,
    n125,
    n320,
    n340,
    n238
  );


  xor
  g474
  (
    KeyWire_0_18,
    n347,
    n235,
    n276,
    n304
  );


  nor
  g475
  (
    n537,
    n223,
    n212,
    n340,
    n129
  );


  or
  g476
  (
    n513,
    n330,
    n151,
    n281,
    n305
  );


  and
  g477
  (
    n523,
    n337,
    n215,
    n333,
    n208
  );


  xnor
  g478
  (
    KeyWire_0_6,
    n196,
    n365,
    n287,
    n231
  );


  xnor
  g479
  (
    n586,
    n230,
    n267,
    n337,
    n299
  );


  or
  g480
  (
    n529,
    n109,
    n214,
    n306,
    n208
  );


  nor
  g481
  (
    n509,
    n367,
    n189,
    n306,
    n209
  );


  nand
  g482
  (
    n400,
    n287,
    n328,
    n335
  );


  xor
  g483
  (
    n491,
    n218,
    n291,
    n107,
    n122
  );


  and
  g484
  (
    n411,
    n348,
    n302,
    n338,
    n227
  );


  or
  g485
  (
    n570,
    n276,
    n313,
    n259,
    n221
  );


  xor
  g486
  (
    n471,
    n314,
    n203,
    n353,
    n320
  );


  xor
  g487
  (
    n424,
    n236,
    n263,
    n276,
    n222
  );


  xnor
  g488
  (
    KeyWire_0_57,
    n312,
    n314,
    n307,
    n256
  );


  xor
  g489
  (
    n572,
    n274,
    n226,
    n329,
    n102
  );


  and
  g490
  (
    n521,
    n221,
    n147,
    n325,
    n287
  );


  nand
  g491
  (
    n417,
    n123,
    n163,
    n274,
    n345
  );


  nor
  g492
  (
    n464,
    n337,
    n342,
    n356,
    n205
  );


  nand
  g493
  (
    n499,
    n235,
    n191,
    n211,
    n364
  );


  or
  g494
  (
    n596,
    n253,
    n322,
    n181,
    n273
  );


  and
  g495
  (
    n579,
    n317,
    n364,
    n252,
    n319
  );


  or
  g496
  (
    n388,
    n351,
    n357,
    n205,
    n211
  );


  xnor
  g497
  (
    n545,
    n261,
    n308,
    n240,
    n106
  );


  nor
  g498
  (
    n562,
    n190,
    n238,
    n336,
    n123
  );


  xor
  g499
  (
    n381,
    n128,
    n250,
    n265,
    n299
  );


  or
  g500
  (
    n413,
    n344,
    n265,
    n335,
    n291
  );


  nand
  g501
  (
    n518,
    n132,
    n361,
    n275
  );


  and
  g502
  (
    n432,
    n266,
    n354,
    n228,
    n213
  );


  and
  g503
  (
    n403,
    n254,
    n161,
    n315,
    n239
  );


  nor
  g504
  (
    n578,
    n299,
    n362,
    n310,
    n281
  );


  nand
  g505
  (
    n504,
    n274,
    n316,
    n182,
    n137
  );


  nand
  g506
  (
    n447,
    n260,
    n217,
    n201,
    n124
  );


  nor
  g507
  (
    n588,
    n313,
    n331,
    n295,
    n281
  );


  nor
  g508
  (
    n384,
    n202,
    n146,
    n236,
    n249
  );


  and
  g509
  (
    KeyWire_0_2,
    n165,
    n215,
    n249,
    n216
  );


  or
  g510
  (
    n490,
    n358,
    n353,
    n134,
    n160
  );


  or
  g511
  (
    n512,
    n309,
    n96,
    n358,
    n360
  );


  nand
  g512
  (
    n383,
    n175,
    n166,
    n321,
    n350
  );


  nand
  g513
  (
    n600,
    n324,
    n213,
    n234,
    n266
  );


  xor
  g514
  (
    n405,
    n141,
    n259,
    n99,
    n345
  );


  xor
  g515
  (
    n433,
    n290,
    n352,
    n248,
    n328
  );


  nand
  g516
  (
    n561,
    n277,
    n259,
    n174,
    n322
  );


  or
  g517
  (
    n524,
    n157,
    n351,
    n357,
    n198
  );


  xor
  g518
  (
    n394,
    n323,
    n144,
    n250,
    n106
  );


  xnor
  g519
  (
    n522,
    n242,
    n298,
    n303,
    n366
  );


  xnor
  g520
  (
    n494,
    n319,
    n341,
    n148,
    n163
  );


  or
  g521
  (
    n463,
    n94,
    n214,
    n252,
    n280
  );


  nand
  g522
  (
    n456,
    n268,
    n321,
    n117,
    n283
  );


  or
  g523
  (
    n440,
    n245,
    n260,
    n234,
    n195
  );


  or
  g524
  (
    n485,
    n98,
    n214,
    n227,
    n173
  );


  xnor
  g525
  (
    n482,
    n246,
    n244,
    n352,
    n337
  );


  and
  g526
  (
    n449,
    n224,
    n105,
    n256,
    n307
  );


  nand
  g527
  (
    n563,
    n254,
    n253,
    n238,
    n224
  );


  nor
  g528
  (
    n558,
    n201,
    n183,
    n253,
    n127
  );


  nand
  g529
  (
    n454,
    n301,
    n282,
    n292,
    n111
  );


  and
  g530
  (
    n489,
    n321,
    n363,
    n150,
    n149
  );


  xnor
  g531
  (
    n393,
    n226,
    n92,
    n248,
    n159
  );


  and
  g532
  (
    n603,
    n330,
    n285,
    n209,
    n347
  );


  xnor
  g533
  (
    n452,
    n202,
    n242,
    n153,
    n347
  );


  nand
  g534
  (
    n501,
    n177,
    n301,
    n263,
    n330
  );


  nor
  g535
  (
    n421,
    n292,
    n191,
    n140,
    n197
  );


  and
  g536
  (
    KeyWire_0_32,
    n234,
    n303,
    n363,
    n280
  );


  xor
  g537
  (
    n461,
    n356,
    n134,
    n199,
    n298
  );


  or
  g538
  (
    n472,
    n293,
    n223,
    n291,
    n155
  );


  nand
  g539
  (
    n564,
    n169,
    n255,
    n93,
    n172
  );


  nor
  g540
  (
    n514,
    n193,
    n288,
    n222,
    n314
  );


  nor
  g541
  (
    n409,
    n318,
    n298,
    n311,
    n224
  );


  xnor
  g542
  (
    n387,
    n186,
    n262,
    n258,
    n294
  );


  or
  g543
  (
    n422,
    n352,
    n342,
    n245,
    n256
  );


  xnor
  g544
  (
    n553,
    n254,
    n114,
    n332,
    n237
  );


  and
  g545
  (
    n412,
    n126,
    n288,
    n339,
    n343
  );


  nand
  g546
  (
    n435,
    n244,
    n267,
    n194,
    n350
  );


  nor
  g547
  (
    n555,
    n268,
    n114,
    n232,
    n137
  );


  nor
  g548
  (
    n582,
    n188,
    n278,
    n334,
    n146
  );


  xnor
  g549
  (
    n414,
    n359,
    n282,
    n233,
    n291
  );


  nor
  g550
  (
    n437,
    n263,
    n304,
    n346,
    n239
  );


  nand
  g551
  (
    n546,
    n340,
    n247,
    n362,
    n245
  );


  nand
  g552
  (
    n528,
    n97,
    n324,
    n220,
    n304
  );


  and
  g553
  (
    n397,
    n118,
    n246,
    n358,
    n121
  );


  and
  g554
  (
    n540,
    n150,
    n153,
    n333,
    n130
  );


  xnor
  g555
  (
    n442,
    n306,
    n219,
    n336,
    n352
  );


  nor
  g556
  (
    n469,
    n92,
    n148,
    n365,
    n218
  );


  or
  g557
  (
    n470,
    n136,
    n206,
    n296,
    n101
  );


  nand
  g558
  (
    n591,
    n345,
    n356,
    n323,
    n128
  );


  nand
  g559
  (
    n597,
    n270,
    n299,
    n269,
    n331
  );


  or
  g560
  (
    n439,
    n127,
    n213,
    n332,
    n192
  );


  nand
  g561
  (
    n441,
    n362,
    n181,
    n252,
    n184
  );


  xor
  g562
  (
    n474,
    n149,
    n343,
    n121,
    n112
  );


  nor
  g563
  (
    n511,
    n270,
    n365,
    n170,
    n301
  );


  or
  g564
  (
    n392,
    n279,
    n211,
    n357,
    n243
  );


  nand
  g565
  (
    n423,
    n171,
    n238,
    n180,
    n212
  );


  and
  g566
  (
    KeyWire_0_54,
    n357,
    n359,
    n126,
    n186
  );


  nor
  g567
  (
    n585,
    n204,
    n307,
    n195
  );


  nor
  g568
  (
    n592,
    n320,
    n258,
    n292,
    n311
  );


  and
  g569
  (
    n497,
    n202,
    n205,
    n217,
    n360
  );


  and
  g570
  (
    n538,
    n204,
    n344,
    n229,
    n217
  );


  xor
  g571
  (
    n576,
    n319,
    n309,
    n338,
    n300
  );


  or
  g572
  (
    n429,
    n138,
    n246,
    n156,
    n94
  );


  xnor
  g573
  (
    n462,
    n129,
    n190,
    n221,
    n255
  );


  or
  g574
  (
    n604,
    n233,
    n289,
    n174,
    n212
  );


  xnor
  g575
  (
    n492,
    n318,
    n366,
    n339,
    n283
  );


  xor
  g576
  (
    n505,
    n179,
    n318,
    n339,
    n198
  );


  nor
  g577
  (
    n398,
    n221,
    n250,
    n286,
    n164
  );


  xor
  g578
  (
    KeyWire_0_49,
    n332,
    n325,
    n367,
    n306
  );


  nor
  g579
  (
    n390,
    n326,
    n143,
    n351,
    n329
  );


  nor
  g580
  (
    n532,
    n108,
    n267,
    n251,
    n162
  );


  nor
  g581
  (
    n549,
    n154,
    n168,
    n133,
    n104
  );


  or
  g582
  (
    n396,
    n225,
    n190,
    n310,
    n342
  );


  or
  g583
  (
    n571,
    n239,
    n273,
    n355,
    n258
  );


  and
  g584
  (
    n500,
    n201,
    n130,
    n225,
    n253
  );


  or
  g585
  (
    n533,
    n354,
    n302,
    n348,
    n269
  );


  or
  g586
  (
    n476,
    n261,
    n282,
    n170,
    n262
  );


  buf
  g587
  (
    n633,
    n516
  );


  buf
  g588
  (
    n776,
    n496
  );


  not
  g589
  (
    n678,
    n434
  );


  not
  g590
  (
    n606,
    n572
  );


  buf
  g591
  (
    n613,
    n407
  );


  not
  g592
  (
    n789,
    n550
  );


  not
  g593
  (
    n798,
    n542
  );


  not
  g594
  (
    n627,
    n382
  );


  not
  g595
  (
    n729,
    n379
  );


  buf
  g596
  (
    n692,
    n563
  );


  buf
  g597
  (
    n716,
    n439
  );


  not
  g598
  (
    n750,
    n462
  );


  not
  g599
  (
    n720,
    n530
  );


  buf
  g600
  (
    n764,
    n497
  );


  not
  g601
  (
    n809,
    n416
  );


  not
  g602
  (
    n609,
    n513
  );


  not
  g603
  (
    n682,
    n454
  );


  buf
  g604
  (
    n792,
    n500
  );


  not
  g605
  (
    n691,
    n482
  );


  not
  g606
  (
    n812,
    n387
  );


  not
  g607
  (
    n641,
    n491
  );


  not
  g608
  (
    n672,
    n435
  );


  buf
  g609
  (
    n730,
    n527
  );


  not
  g610
  (
    n710,
    n570
  );


  buf
  g611
  (
    KeyWire_0_59,
    n488
  );


  not
  g612
  (
    n654,
    n477
  );


  not
  g613
  (
    n656,
    n507
  );


  buf
  g614
  (
    n788,
    n538
  );


  buf
  g615
  (
    n695,
    n539
  );


  not
  g616
  (
    n608,
    n395
  );


  not
  g617
  (
    n801,
    n418
  );


  buf
  g618
  (
    n615,
    n546
  );


  not
  g619
  (
    n762,
    n438
  );


  not
  g620
  (
    n763,
    n514
  );


  not
  g621
  (
    n616,
    n429
  );


  not
  g622
  (
    n647,
    n489
  );


  buf
  g623
  (
    n810,
    n493
  );


  not
  g624
  (
    n701,
    n545
  );


  buf
  g625
  (
    n621,
    n520
  );


  not
  g626
  (
    n617,
    n455
  );


  not
  g627
  (
    n804,
    n490
  );


  not
  g628
  (
    n696,
    n498
  );


  not
  g629
  (
    n742,
    n544
  );


  not
  g630
  (
    n658,
    n381
  );


  buf
  g631
  (
    n785,
    n463
  );


  buf
  g632
  (
    n775,
    n577
  );


  not
  g633
  (
    n739,
    n412
  );


  not
  g634
  (
    n738,
    n494
  );


  not
  g635
  (
    n699,
    n447
  );


  buf
  g636
  (
    n644,
    n502
  );


  not
  g637
  (
    n632,
    n471
  );


  buf
  g638
  (
    n705,
    n401
  );


  buf
  g639
  (
    n784,
    n464
  );


  not
  g640
  (
    n813,
    n451
  );


  not
  g641
  (
    n796,
    n510
  );


  buf
  g642
  (
    n618,
    n430
  );


  not
  g643
  (
    n657,
    n433
  );


  not
  g644
  (
    KeyWire_0_56,
    n571
  );


  not
  g645
  (
    n625,
    n585
  );


  buf
  g646
  (
    n740,
    n388
  );


  not
  g647
  (
    KeyWire_0_3,
    n472
  );


  buf
  g648
  (
    n637,
    n541
  );


  not
  g649
  (
    n797,
    n526
  );


  not
  g650
  (
    n639,
    n413
  );


  not
  g651
  (
    n686,
    n554
  );


  buf
  g652
  (
    n714,
    n560
  );


  not
  g653
  (
    n806,
    n522
  );


  buf
  g654
  (
    n752,
    n564
  );


  not
  g655
  (
    n757,
    n406
  );


  not
  g656
  (
    n794,
    n420
  );


  not
  g657
  (
    n663,
    n385
  );


  buf
  g658
  (
    n807,
    n529
  );


  not
  g659
  (
    n693,
    n431
  );


  buf
  g660
  (
    n646,
    n409
  );


  buf
  g661
  (
    n765,
    n393
  );


  buf
  g662
  (
    n704,
    n414
  );


  buf
  g663
  (
    n760,
    n553
  );


  not
  g664
  (
    n808,
    n415
  );


  buf
  g665
  (
    n707,
    n573
  );


  buf
  g666
  (
    n718,
    n524
  );


  not
  g667
  (
    n689,
    n453
  );


  buf
  g668
  (
    n643,
    n558
  );


  not
  g669
  (
    KeyWire_0_0,
    n436
  );


  buf
  g670
  (
    n790,
    n466
  );


  not
  g671
  (
    n624,
    n534
  );


  buf
  g672
  (
    n690,
    n532
  );


  not
  g673
  (
    n635,
    n384
  );


  buf
  g674
  (
    n661,
    n556
  );


  not
  g675
  (
    n681,
    n400
  );


  not
  g676
  (
    n640,
    n584
  );


  not
  g677
  (
    n759,
    n394
  );


  not
  g678
  (
    n630,
    n391
  );


  buf
  g679
  (
    n766,
    n479
  );


  buf
  g680
  (
    n726,
    n410
  );


  not
  g681
  (
    n767,
    n480
  );


  not
  g682
  (
    n782,
    n487
  );


  buf
  g683
  (
    n793,
    n555
  );


  not
  g684
  (
    n652,
    n459
  );


  not
  g685
  (
    n715,
    n422
  );


  buf
  g686
  (
    n778,
    n442
  );


  buf
  g687
  (
    n741,
    n411
  );


  buf
  g688
  (
    KeyWire_0_44,
    n586
  );


  not
  g689
  (
    n727,
    n469
  );


  buf
  g690
  (
    n683,
    n389
  );


  buf
  g691
  (
    n722,
    n565
  );


  buf
  g692
  (
    n773,
    n423
  );


  buf
  g693
  (
    n736,
    n399
  );


  buf
  g694
  (
    n747,
    n427
  );


  not
  g695
  (
    n702,
    n458
  );


  not
  g696
  (
    n719,
    n537
  );


  buf
  g697
  (
    n669,
    n547
  );


  not
  g698
  (
    n733,
    n484
  );


  not
  g699
  (
    n675,
    n552
  );


  buf
  g700
  (
    n803,
    n398
  );


  buf
  g701
  (
    n706,
    n499
  );


  not
  g702
  (
    KeyWire_0_9,
    n408
  );


  not
  g703
  (
    n774,
    n540
  );


  buf
  g704
  (
    n645,
    n517
  );


  buf
  g705
  (
    n667,
    n583
  );


  buf
  g706
  (
    n732,
    n465
  );


  not
  g707
  (
    n680,
    n505
  );


  not
  g708
  (
    n651,
    n452
  );


  not
  g709
  (
    n700,
    n444
  );


  not
  g710
  (
    n671,
    n533
  );


  buf
  g711
  (
    n628,
    n404
  );


  buf
  g712
  (
    n623,
    n523
  );


  not
  g713
  (
    KeyWire_0_7,
    n543
  );


  buf
  g714
  (
    n779,
    n467
  );


  buf
  g715
  (
    n665,
    n475
  );


  not
  g716
  (
    n650,
    n474
  );


  not
  g717
  (
    n612,
    n512
  );


  buf
  g718
  (
    n694,
    n449
  );


  not
  g719
  (
    n799,
    n448
  );


  not
  g720
  (
    n697,
    n383
  );


  not
  g721
  (
    n748,
    n461
  );


  not
  g722
  (
    n674,
    n580
  );


  buf
  g723
  (
    n744,
    n443
  );


  not
  g724
  (
    n655,
    n428
  );


  buf
  g725
  (
    n745,
    n437
  );


  buf
  g726
  (
    n677,
    n386
  );


  not
  g727
  (
    n769,
    n432
  );


  buf
  g728
  (
    n768,
    n468
  );


  buf
  g729
  (
    n755,
    n566
  );


  buf
  g730
  (
    n662,
    n568
  );


  not
  g731
  (
    n619,
    n486
  );


  buf
  g732
  (
    n724,
    n569
  );


  buf
  g733
  (
    n811,
    n518
  );


  not
  g734
  (
    n642,
    n521
  );


  buf
  g735
  (
    n688,
    n557
  );


  not
  g736
  (
    n728,
    n576
  );


  buf
  g737
  (
    n735,
    n579
  );


  buf
  g738
  (
    n610,
    n397
  );


  not
  g739
  (
    n771,
    n536
  );


  buf
  g740
  (
    n756,
    n548
  );


  not
  g741
  (
    n761,
    n476
  );


  buf
  g742
  (
    n614,
    n440
  );


  buf
  g743
  (
    n653,
    n380
  );


  not
  g744
  (
    n725,
    n561
  );


  buf
  g745
  (
    n791,
    n549
  );


  buf
  g746
  (
    n636,
    n495
  );


  not
  g747
  (
    KeyWire_0_39,
    n551
  );


  not
  g748
  (
    n731,
    n508
  );


  not
  g749
  (
    n709,
    n485
  );


  buf
  g750
  (
    n664,
    n535
  );


  buf
  g751
  (
    n634,
    n426
  );


  buf
  g752
  (
    n753,
    n402
  );


  not
  g753
  (
    n670,
    n503
  );


  not
  g754
  (
    n622,
    n567
  );


  buf
  g755
  (
    n713,
    n581
  );


  buf
  g756
  (
    n734,
    n403
  );


  not
  g757
  (
    n721,
    n390
  );


  not
  g758
  (
    n660,
    n445
  );


  not
  g759
  (
    n626,
    n574
  );


  buf
  g760
  (
    n638,
    n562
  );


  buf
  g761
  (
    n687,
    n492
  );


  buf
  g762
  (
    n737,
    n528
  );


  buf
  g763
  (
    n754,
    n419
  );


  not
  g764
  (
    n795,
    n511
  );


  buf
  g765
  (
    n611,
    n504
  );


  not
  g766
  (
    n703,
    n531
  );


  buf
  g767
  (
    n802,
    n525
  );


  buf
  g768
  (
    n666,
    n481
  );


  not
  g769
  (
    n676,
    n582
  );


  buf
  g770
  (
    n668,
    n478
  );


  buf
  g771
  (
    n649,
    n396
  );


  not
  g772
  (
    n698,
    n424
  );


  buf
  g773
  (
    n685,
    n457
  );


  buf
  g774
  (
    n777,
    n515
  );


  buf
  g775
  (
    n723,
    n506
  );


  not
  g776
  (
    n631,
    n473
  );


  buf
  g777
  (
    n783,
    n509
  );


  not
  g778
  (
    n708,
    n425
  );


  buf
  g779
  (
    n787,
    n460
  );


  buf
  g780
  (
    n607,
    n421
  );


  not
  g781
  (
    n749,
    n519
  );


  not
  g782
  (
    n711,
    n501
  );


  not
  g783
  (
    n780,
    n446
  );


  buf
  g784
  (
    n770,
    n578
  );


  buf
  g785
  (
    n800,
    n470
  );


  not
  g786
  (
    n758,
    n575
  );


  not
  g787
  (
    n781,
    n483
  );


  not
  g788
  (
    n629,
    n392
  );


  buf
  g789
  (
    n648,
    n456
  );


  not
  g790
  (
    n786,
    n405
  );


  buf
  g791
  (
    n684,
    n450
  );


  buf
  g792
  (
    n712,
    n559
  );


  buf
  g793
  (
    n620,
    n417
  );


  buf
  g794
  (
    n805,
    n441
  );


  buf
  g795
  (
    n901,
    n704
  );


  not
  g796
  (
    n886,
    n699
  );


  not
  g797
  (
    n973,
    n717
  );


  buf
  g798
  (
    n922,
    n663
  );


  not
  g799
  (
    n1010,
    n664
  );


  not
  g800
  (
    KeyWire_0_62,
    n696
  );


  buf
  g801
  (
    n979,
    n662
  );


  buf
  g802
  (
    n952,
    n660
  );


  not
  g803
  (
    n838,
    n690
  );


  not
  g804
  (
    n823,
    n726
  );


  buf
  g805
  (
    n921,
    n712
  );


  not
  g806
  (
    n891,
    n618
  );


  buf
  g807
  (
    n1045,
    n676
  );


  not
  g808
  (
    n948,
    n706
  );


  not
  g809
  (
    n1046,
    n716
  );


  not
  g810
  (
    n836,
    n613
  );


  buf
  g811
  (
    n830,
    n634
  );


  buf
  g812
  (
    n1023,
    n671
  );


  buf
  g813
  (
    n980,
    n700
  );


  not
  g814
  (
    n1002,
    n629
  );


  buf
  g815
  (
    n941,
    n711
  );


  buf
  g816
  (
    n824,
    n693
  );


  not
  g817
  (
    n983,
    n697
  );


  not
  g818
  (
    n970,
    n666
  );


  not
  g819
  (
    n914,
    n719
  );


  buf
  g820
  (
    n909,
    n642
  );


  not
  g821
  (
    n841,
    n617
  );


  not
  g822
  (
    n912,
    n616
  );


  buf
  g823
  (
    n868,
    n659
  );


  buf
  g824
  (
    n816,
    n626
  );


  buf
  g825
  (
    n1041,
    n623
  );


  not
  g826
  (
    n866,
    n642
  );


  not
  g827
  (
    n857,
    n670
  );


  not
  g828
  (
    n883,
    n678
  );


  buf
  g829
  (
    n907,
    n634
  );


  not
  g830
  (
    KeyWire_0_38,
    n663
  );


  buf
  g831
  (
    n1024,
    n633
  );


  not
  g832
  (
    n839,
    n665
  );


  not
  g833
  (
    n833,
    n622
  );


  not
  g834
  (
    n887,
    n679
  );


  buf
  g835
  (
    n937,
    n653
  );


  not
  g836
  (
    n933,
    n643
  );


  buf
  g837
  (
    KeyWire_0_30,
    n696
  );


  not
  g838
  (
    n964,
    n700
  );


  not
  g839
  (
    n1008,
    n698
  );


  buf
  g840
  (
    n852,
    n693
  );


  buf
  g841
  (
    n1015,
    n711
  );


  buf
  g842
  (
    n859,
    n660
  );


  buf
  g843
  (
    n1032,
    n710
  );


  buf
  g844
  (
    KeyWire_0_4,
    n633
  );


  buf
  g845
  (
    n998,
    n722
  );


  not
  g846
  (
    n855,
    n683
  );


  not
  g847
  (
    n1029,
    n718
  );


  buf
  g848
  (
    n1040,
    n614
  );


  not
  g849
  (
    n828,
    n643
  );


  buf
  g850
  (
    n1048,
    n616
  );


  not
  g851
  (
    n853,
    n645
  );


  buf
  g852
  (
    n1052,
    n691
  );


  buf
  g853
  (
    n894,
    n635
  );


  not
  g854
  (
    n858,
    n656
  );


  not
  g855
  (
    n847,
    n652
  );


  buf
  g856
  (
    n1014,
    n606
  );


  buf
  g857
  (
    n1026,
    n623
  );


  buf
  g858
  (
    n988,
    n635
  );


  not
  g859
  (
    n827,
    n640
  );


  not
  g860
  (
    n825,
    n714
  );


  not
  g861
  (
    n972,
    n617
  );


  buf
  g862
  (
    n959,
    n640
  );


  not
  g863
  (
    n873,
    n651
  );


  not
  g864
  (
    n1051,
    n608
  );


  not
  g865
  (
    n878,
    n615
  );


  buf
  g866
  (
    n896,
    n678
  );


  not
  g867
  (
    n867,
    n721
  );


  buf
  g868
  (
    n876,
    n612
  );


  not
  g869
  (
    n931,
    n689
  );


  not
  g870
  (
    n1013,
    n676
  );


  buf
  g871
  (
    n943,
    n610
  );


  buf
  g872
  (
    n1037,
    n679
  );


  not
  g873
  (
    n993,
    n675
  );


  buf
  g874
  (
    n1036,
    n720
  );


  buf
  g875
  (
    n946,
    n610
  );


  not
  g876
  (
    n955,
    n624
  );


  not
  g877
  (
    n906,
    n715
  );


  buf
  g878
  (
    n935,
    n637
  );


  not
  g879
  (
    n986,
    n647
  );


  buf
  g880
  (
    n1000,
    n649
  );


  not
  g881
  (
    n958,
    n722
  );


  not
  g882
  (
    n826,
    n621
  );


  not
  g883
  (
    n1031,
    n685
  );


  not
  g884
  (
    n938,
    n685
  );


  buf
  g885
  (
    n844,
    n674
  );


  buf
  g886
  (
    n978,
    n699
  );


  buf
  g887
  (
    KeyWire_0_22,
    n705
  );


  buf
  g888
  (
    n1009,
    n625
  );


  not
  g889
  (
    n999,
    n657
  );


  buf
  g890
  (
    n834,
    n692
  );


  buf
  g891
  (
    n1016,
    n719
  );


  not
  g892
  (
    n877,
    n631
  );


  buf
  g893
  (
    n969,
    n655
  );


  buf
  g894
  (
    n920,
    n713
  );


  buf
  g895
  (
    n888,
    n725
  );


  not
  g896
  (
    n814,
    n629
  );


  not
  g897
  (
    n872,
    n706
  );


  not
  g898
  (
    n1025,
    n647
  );


  not
  g899
  (
    n997,
    n686
  );


  not
  g900
  (
    n929,
    n701
  );


  buf
  g901
  (
    n916,
    n611
  );


  not
  g902
  (
    n930,
    n626
  );


  not
  g903
  (
    n1022,
    n701
  );


  buf
  g904
  (
    KeyWire_0_34,
    n684
  );


  buf
  g905
  (
    n842,
    n698
  );


  not
  g906
  (
    n945,
    n708
  );


  not
  g907
  (
    n904,
    n664
  );


  not
  g908
  (
    n865,
    n639
  );


  buf
  g909
  (
    n965,
    n639
  );


  not
  g910
  (
    KeyWire_0_43,
    n668
  );


  buf
  g911
  (
    KeyWire_0_5,
    n620
  );


  not
  g912
  (
    n991,
    n672
  );


  buf
  g913
  (
    n987,
    n638
  );


  buf
  g914
  (
    n854,
    n717
  );


  buf
  g915
  (
    n919,
    n630
  );


  not
  g916
  (
    n915,
    n695
  );


  not
  g917
  (
    n893,
    n654
  );


  not
  g918
  (
    n1005,
    n707
  );


  buf
  g919
  (
    n953,
    n723
  );


  buf
  g920
  (
    n940,
    n682
  );


  buf
  g921
  (
    n879,
    n705
  );


  buf
  g922
  (
    n954,
    n687
  );


  not
  g923
  (
    n951,
    n702
  );


  buf
  g924
  (
    n884,
    n692
  );


  buf
  g925
  (
    KeyWire_0_58,
    n707
  );


  buf
  g926
  (
    n899,
    n723
  );


  buf
  g927
  (
    n869,
    n627
  );


  not
  g928
  (
    n990,
    n624
  );


  not
  g929
  (
    n815,
    n720
  );


  buf
  g930
  (
    n950,
    n609
  );


  not
  g931
  (
    n881,
    n653
  );


  not
  g932
  (
    n928,
    n669
  );


  not
  g933
  (
    n864,
    n681
  );


  buf
  g934
  (
    n875,
    n704
  );


  not
  g935
  (
    n897,
    n674
  );


  buf
  g936
  (
    n977,
    n677
  );


  not
  g937
  (
    n923,
    n668
  );


  buf
  g938
  (
    n818,
    n721
  );


  buf
  g939
  (
    n863,
    n712
  );


  buf
  g940
  (
    n917,
    n667
  );


  not
  g941
  (
    n1047,
    n709
  );


  buf
  g942
  (
    n882,
    n652
  );


  not
  g943
  (
    n871,
    n619
  );


  buf
  g944
  (
    n851,
    n657
  );


  not
  g945
  (
    n944,
    n621
  );


  buf
  g946
  (
    KeyWire_0_27,
    n609
  );


  buf
  g947
  (
    n939,
    n641
  );


  not
  g948
  (
    n932,
    n645
  );


  not
  g949
  (
    n892,
    n658
  );


  not
  g950
  (
    n934,
    n646
  );


  buf
  g951
  (
    n981,
    n641
  );


  buf
  g952
  (
    n1006,
    n648
  );


  buf
  g953
  (
    n860,
    n708
  );


  not
  g954
  (
    n908,
    n688
  );


  buf
  g955
  (
    n862,
    n644
  );


  buf
  g956
  (
    n1003,
    n690
  );


  buf
  g957
  (
    n870,
    n632
  );


  not
  g958
  (
    n1033,
    n718
  );


  not
  g959
  (
    n1004,
    n694
  );


  not
  g960
  (
    n902,
    n619
  );


  not
  g961
  (
    n995,
    n710
  );


  not
  g962
  (
    n975,
    n684
  );


  not
  g963
  (
    n905,
    n662
  );


  not
  g964
  (
    n1007,
    n681
  );


  buf
  g965
  (
    n967,
    n628
  );


  buf
  g966
  (
    n968,
    n670
  );


  not
  g967
  (
    n982,
    n703
  );


  buf
  g968
  (
    n1012,
    n646
  );


  buf
  g969
  (
    n850,
    n671
  );


  buf
  g970
  (
    n1030,
    n611
  );


  not
  g971
  (
    n989,
    n702
  );


  not
  g972
  (
    n984,
    n644
  );


  buf
  g973
  (
    n837,
    n680
  );


  not
  g974
  (
    n996,
    n695
  );


  buf
  g975
  (
    n1019,
    n669
  );


  buf
  g976
  (
    n925,
    n632
  );


  buf
  g977
  (
    KeyWire_0_55,
    n694
  );


  buf
  g978
  (
    n832,
    n715
  );


  not
  g979
  (
    n942,
    n666
  );


  not
  g980
  (
    n910,
    n687
  );


  not
  g981
  (
    n926,
    n607
  );


  not
  g982
  (
    n1039,
    n677
  );


  buf
  g983
  (
    n1049,
    n655
  );


  buf
  g984
  (
    n889,
    n686
  );


  buf
  g985
  (
    n1042,
    n651
  );


  not
  g986
  (
    n949,
    n630
  );


  not
  g987
  (
    n1043,
    n667
  );


  buf
  g988
  (
    n961,
    n688
  );


  buf
  g989
  (
    n821,
    n713
  );


  buf
  g990
  (
    n957,
    n691
  );


  not
  g991
  (
    n890,
    n714
  );


  buf
  g992
  (
    n974,
    n672
  );


  buf
  g993
  (
    n903,
    n726
  );


  not
  g994
  (
    n885,
    n661
  );


  buf
  g995
  (
    n835,
    n661
  );


  not
  g996
  (
    n947,
    n659
  );


  not
  g997
  (
    n1011,
    n697
  );


  not
  g998
  (
    n1027,
    n703
  );


  buf
  g999
  (
    n817,
    n612
  );


  buf
  g1000
  (
    n1020,
    n656
  );


  not
  g1001
  (
    n971,
    n637
  );


  buf
  g1002
  (
    n843,
    n727
  );


  not
  g1003
  (
    n819,
    n682
  );


  buf
  g1004
  (
    n924,
    n625
  );


  not
  g1005
  (
    n1001,
    n618
  );


  not
  g1006
  (
    n1021,
    n673
  );


  not
  g1007
  (
    n1050,
    n613
  );


  buf
  g1008
  (
    n918,
    n614
  );


  not
  g1009
  (
    n911,
    n636
  );


  buf
  g1010
  (
    n985,
    n675
  );


  buf
  g1011
  (
    n1034,
    n654
  );


  not
  g1012
  (
    n1044,
    n724
  );


  not
  g1013
  (
    n1038,
    n638
  );


  buf
  g1014
  (
    KeyWire_0_50,
    n620
  );


  buf
  g1015
  (
    n966,
    n615
  );


  not
  g1016
  (
    n1035,
    n627
  );


  buf
  g1017
  (
    n1018,
    n650
  );


  buf
  g1018
  (
    n856,
    n649
  );


  not
  g1019
  (
    n992,
    n648
  );


  not
  g1020
  (
    n963,
    n716
  );


  not
  g1021
  (
    n840,
    n725
  );


  not
  g1022
  (
    n1053,
    n658
  );


  not
  g1023
  (
    n898,
    n683
  );


  buf
  g1024
  (
    n994,
    n650
  );


  buf
  g1025
  (
    n956,
    n709
  );


  buf
  g1026
  (
    n900,
    n724
  );


  not
  g1027
  (
    n829,
    n665
  );


  buf
  g1028
  (
    n831,
    n680
  );


  buf
  g1029
  (
    n936,
    n636
  );


  not
  g1030
  (
    n976,
    n689
  );


  not
  g1031
  (
    n960,
    n673
  );


  buf
  g1032
  (
    KeyWire_0_17,
    n631
  );


  not
  g1033
  (
    n927,
    n622
  );


  not
  g1034
  (
    n846,
    n628
  );


  not
  g1035
  (
    n1056,
    n821
  );


  buf
  g1036
  (
    n1054,
    n818
  );


  not
  g1037
  (
    n1060,
    n816
  );


  not
  g1038
  (
    n1059,
    n819
  );


  buf
  g1039
  (
    n1061,
    n817
  );


  not
  g1040
  (
    n1057,
    n820
  );


  buf
  g1041
  (
    KeyWire_0_53,
    n814
  );


  buf
  g1042
  (
    n1058,
    n815
  );


  not
  g1043
  (
    n1071,
    n837
  );


  not
  g1044
  (
    KeyWire_0_13,
    n841
  );


  nor
  g1045
  (
    n1063,
    n1060,
    n823
  );


  nand
  g1046
  (
    n1062,
    n1056,
    n827,
    n839,
    n836
  );


  xnor
  g1047
  (
    n1065,
    n835,
    n1061,
    n843,
    n833
  );


  nor
  g1048
  (
    n1066,
    n1058,
    n1060,
    n825,
    n840
  );


  nand
  g1049
  (
    n1070,
    n1059,
    n832,
    n831,
    n830
  );


  nor
  g1050
  (
    n1064,
    n834,
    n822,
    n824,
    n1054
  );


  nor
  g1051
  (
    n1067,
    n1057,
    n842,
    n829,
    n1061
  );


  xor
  g1052
  (
    n1068,
    n828,
    n1055,
    n838,
    n826
  );


  not
  g1053
  (
    n1074,
    n1066
  );


  buf
  g1054
  (
    n1072,
    n1063
  );


  buf
  g1055
  (
    n1075,
    n1065
  );


  buf
  g1056
  (
    n1076,
    n844
  );


  or
  g1057
  (
    n1073,
    n1064,
    n1062
  );


  buf
  g1058
  (
    n1079,
    n1073
  );


  buf
  g1059
  (
    n1083,
    n1073
  );


  not
  g1060
  (
    n1081,
    n1072
  );


  buf
  g1061
  (
    n1084,
    n1073
  );


  buf
  g1062
  (
    n1077,
    n1072
  );


  buf
  g1063
  (
    n1078,
    n1074
  );


  not
  g1064
  (
    KeyWire_0_29,
    n1073
  );


  not
  g1065
  (
    n1082,
    n1074
  );


  buf
  g1066
  (
    n1099,
    n1079
  );


  not
  g1067
  (
    n1100,
    n737
  );


  not
  g1068
  (
    n1091,
    n1078
  );


  not
  g1069
  (
    n1094,
    n1083
  );


  xor
  g1070
  (
    n1085,
    n734,
    n730,
    n1081,
    n739
  );


  nor
  g1071
  (
    n1087,
    n736,
    n739,
    n1078,
    n730
  );


  and
  g1072
  (
    n1093,
    n727,
    n1080,
    n733,
    n1078
  );


  xnor
  g1073
  (
    n1092,
    n736,
    n1081,
    n738,
    n1077
  );


  nor
  g1074
  (
    n1096,
    n735,
    n733,
    n737,
    n738
  );


  xor
  g1075
  (
    n1098,
    n1080,
    n735,
    n729,
    n1077
  );


  or
  g1076
  (
    n1097,
    n1079,
    n734,
    n732,
    n1077
  );


  nor
  g1077
  (
    n1088,
    n1080,
    n729,
    n1082,
    n728
  );


  nor
  g1078
  (
    n1086,
    n1082,
    n740,
    n731,
    n732
  );


  or
  g1079
  (
    n1089,
    n731,
    n728,
    n1078,
    n1082
  );


  and
  g1080
  (
    n1095,
    n1081,
    n1082,
    n1079,
    n1083
  );


  nor
  g1081
  (
    n1090,
    n1081,
    n1077,
    n1079,
    n1080
  );


  and
  g1082
  (
    n1110,
    n759,
    n761,
    n747,
    n756
  );


  xnor
  g1083
  (
    n1108,
    n754,
    n749,
    n757,
    n752
  );


  nor
  g1084
  (
    n1102,
    n742,
    n741,
    n740
  );


  or
  g1085
  (
    n1113,
    n745,
    n1100,
    n759,
    n1088
  );


  nor
  g1086
  (
    n1111,
    n1091,
    n763,
    n1085,
    n752
  );


  xnor
  g1087
  (
    n1103,
    n758,
    n745,
    n756,
    n1097
  );


  xnor
  g1088
  (
    n1116,
    n748,
    n755,
    n754,
    n743
  );


  or
  g1089
  (
    n1105,
    n1099,
    n762,
    n750,
    n1096
  );


  nand
  g1090
  (
    n1109,
    n1087,
    n764,
    n760,
    n755
  );


  nor
  g1091
  (
    n1101,
    n1095,
    n1089,
    n750,
    n746
  );


  xor
  g1092
  (
    n1106,
    n1092,
    n1093,
    n743,
    n1086
  );


  and
  g1093
  (
    n1115,
    n1094,
    n753,
    n1098,
    n751
  );


  nor
  g1094
  (
    n1107,
    n753,
    n747,
    n758,
    n748
  );


  nor
  g1095
  (
    n1104,
    n744,
    n746,
    n757,
    n1090
  );


  nand
  g1096
  (
    n1112,
    n751,
    n763,
    n760,
    n762
  );


  or
  g1097
  (
    n1114,
    n761,
    n742,
    n744,
    n749
  );


  or
  g1098
  (
    n1143,
    n858,
    n848,
    n1102,
    n922
  );


  or
  g1099
  (
    n1140,
    n871,
    n1106,
    n908,
    n911
  );


  nand
  g1100
  (
    n1129,
    n921,
    n906,
    n914,
    n923
  );


  or
  g1101
  (
    n1142,
    n846,
    n907,
    n857,
    n880
  );


  or
  g1102
  (
    n1123,
    n916,
    n1103,
    n1104,
    n1101
  );


  and
  g1103
  (
    n1119,
    n919,
    n851,
    n1105,
    n912
  );


  and
  g1104
  (
    n1131,
    n915,
    n878,
    n1106,
    n861
  );


  xor
  g1105
  (
    n1135,
    n866,
    n865,
    n1102,
    n1107
  );


  or
  g1106
  (
    n1136,
    n918,
    n876,
    n850,
    n924
  );


  or
  g1107
  (
    n1134,
    n909,
    n910,
    n1104,
    n1101
  );


  nand
  g1108
  (
    n1121,
    n874,
    n893,
    n856,
    n864
  );


  nand
  g1109
  (
    n1124,
    n868,
    n875,
    n1101,
    n899
  );


  nand
  g1110
  (
    n1125,
    n888,
    n882,
    n872,
    n847
  );


  or
  g1111
  (
    n1138,
    n883,
    n895,
    n877,
    n859
  );


  or
  g1112
  (
    n1122,
    n860,
    n1103,
    n900,
    n903
  );


  or
  g1113
  (
    KeyWire_0_20,
    n879,
    n863,
    n881,
    n892
  );


  nor
  g1114
  (
    n1120,
    n898,
    n1106,
    n1107,
    n1102
  );


  nand
  g1115
  (
    n1141,
    n884,
    n897,
    n1105,
    n867
  );


  or
  g1116
  (
    n1130,
    n904,
    n845,
    n1103,
    n925
  );


  and
  g1117
  (
    n1133,
    n849,
    n853,
    n917,
    n854
  );


  or
  g1118
  (
    n1132,
    n852,
    n887,
    n886,
    n890
  );


  xor
  g1119
  (
    n1128,
    n855,
    n870,
    n902,
    n1104
  );


  nor
  g1120
  (
    n1127,
    n889,
    n1102,
    n885,
    n1105
  );


  xnor
  g1121
  (
    n1118,
    n894,
    n920,
    n869,
    n1105
  );


  nand
  g1122
  (
    KeyWire_0_10,
    n1106,
    n913,
    n1103,
    n1107
  );


  nand
  g1123
  (
    n1117,
    n896,
    n891,
    n901,
    n862
  );


  xor
  g1124
  (
    n1137,
    n1101,
    n1104,
    n905,
    n873
  );


  buf
  g1125
  (
    n1150,
    n1120
  );


  buf
  g1126
  (
    KeyWire_0_40,
    n1123
  );


  not
  g1127
  (
    n1146,
    n1119
  );


  buf
  g1128
  (
    n1147,
    n1124
  );


  not
  g1129
  (
    n1149,
    n1125
  );


  buf
  g1130
  (
    n1145,
    n1121
  );


  not
  g1131
  (
    n1144,
    n1126
  );


  not
  g1132
  (
    n1148,
    n1122
  );


  and
  g1133
  (
    n1163,
    n1131,
    n958,
    n1149,
    n1069
  );


  and
  g1134
  (
    n1176,
    n952,
    n1149,
    n596,
    n1144
  );


  and
  g1135
  (
    n1172,
    n598,
    n1129,
    n938,
    n1074
  );


  nor
  g1136
  (
    n1179,
    n370,
    n929,
    n926,
    n589
  );


  or
  g1137
  (
    n1174,
    n1146,
    n951,
    n1145,
    n956
  );


  nor
  g1138
  (
    n1180,
    n1151,
    n934,
    n1150,
    n371
  );


  or
  g1139
  (
    n1158,
    n1127,
    n766,
    n1144,
    n1148
  );


  or
  g1140
  (
    n1164,
    n943,
    n1147,
    n936,
    n594
  );


  and
  g1141
  (
    n1153,
    n765,
    n1147,
    n604,
    n595
  );


  or
  g1142
  (
    KeyWire_0_61,
    n599,
    n602,
    n932,
    n764
  );


  nor
  g1143
  (
    n1161,
    n371,
    n369,
    n1146,
    n368
  );


  nand
  g1144
  (
    n1154,
    n368,
    n1068,
    n948,
    n370
  );


  xor
  g1145
  (
    n1159,
    n950,
    n368,
    n1128,
    n587
  );


  xor
  g1146
  (
    n1162,
    n1150,
    n1144,
    n930,
    n1075
  );


  nor
  g1147
  (
    n1168,
    n942,
    n941,
    n945,
    n766
  );


  and
  g1148
  (
    n1181,
    n1067,
    n605,
    n765,
    n588
  );


  or
  g1149
  (
    n1170,
    n1075,
    n1075,
    n1148,
    n369
  );


  and
  g1150
  (
    n1169,
    n946,
    n931,
    n947,
    n1147
  );


  or
  g1151
  (
    n1175,
    n939,
    n1076,
    n1145,
    n370
  );


  xnor
  g1152
  (
    n1173,
    n600,
    n1076,
    n597,
    n593
  );


  or
  g1153
  (
    n1178,
    n937,
    n767,
    n962,
    n1130
  );


  xor
  g1154
  (
    n1167,
    n370,
    n1148,
    n1074
  );


  or
  g1155
  (
    n1165,
    n1150,
    n1132,
    n1147,
    n1144
  );


  and
  g1156
  (
    n1160,
    n944,
    n1149,
    n591,
    n1071
  );


  nand
  g1157
  (
    n1157,
    n949,
    n368,
    n955,
    n960
  );


  and
  g1158
  (
    n1177,
    n957,
    n601,
    n940,
    n1151
  );


  nor
  g1159
  (
    n1183,
    n367,
    n590,
    n592,
    n961
  );


  xnor
  g1160
  (
    n1156,
    n1150,
    n1075,
    n1146,
    n369
  );


  and
  g1161
  (
    n1171,
    n1151,
    n1145,
    n959,
    n1070
  );


  and
  g1162
  (
    n1155,
    n1149,
    n933,
    n1145,
    n927
  );


  nand
  g1163
  (
    n1166,
    n928,
    n369,
    n954,
    n1146
  );


  xor
  g1164
  (
    n1152,
    n935,
    n603,
    n1151,
    n953
  );


  xor
  g1165
  (
    n1198,
    n779,
    n769,
    n790
  );


  nor
  g1166
  (
    n1184,
    n784,
    n1154,
    n1157,
    n787
  );


  and
  g1167
  (
    n1191,
    n785,
    n1156,
    n771,
    n1153
  );


  and
  g1168
  (
    n1188,
    n783,
    n790,
    n772,
    n788
  );


  xor
  g1169
  (
    n1185,
    n781,
    n1152,
    n782,
    n1154
  );


  xor
  g1170
  (
    n1197,
    n1153,
    n777,
    n781,
    n778
  );


  xnor
  g1171
  (
    n1195,
    n786,
    n768,
    n1156,
    n789
  );


  xnor
  g1172
  (
    n1189,
    n770,
    n776,
    n771,
    n786
  );


  xnor
  g1173
  (
    n1199,
    n776,
    n767,
    n783,
    n778
  );


  nor
  g1174
  (
    n1193,
    n784,
    n774,
    n791,
    n775
  );


  xor
  g1175
  (
    n1186,
    n1155,
    n772,
    n1158,
    n787
  );


  nor
  g1176
  (
    n1187,
    n777,
    n779,
    n780,
    n773
  );


  or
  g1177
  (
    n1196,
    n1157,
    n770,
    n1159,
    n773
  );


  or
  g1178
  (
    n1192,
    n789,
    n1152,
    n785,
    n1158
  );


  xnor
  g1179
  (
    n1194,
    n788,
    n774,
    n768,
    n775
  );


  xnor
  g1180
  (
    n1190,
    n1159,
    n780,
    n1155,
    n782
  );


  xnor
  g1181
  (
    n1211,
    n974,
    n985,
    n1196,
    n997
  );


  xnor
  g1182
  (
    n1208,
    n968,
    n969,
    n1195,
    n976
  );


  or
  g1183
  (
    n1206,
    n972,
    n995,
    n970,
    n983
  );


  nand
  g1184
  (
    n1201,
    n994,
    n986,
    n1001,
    n977
  );


  and
  g1185
  (
    n1212,
    n989,
    n1198,
    n990,
    n1192
  );


  or
  g1186
  (
    n1204,
    n980,
    n1000,
    n1188,
    n993
  );


  and
  g1187
  (
    n1209,
    n999,
    n1197,
    n965,
    n966
  );


  nor
  g1188
  (
    n1205,
    n987,
    n1003,
    n1002,
    n996
  );


  and
  g1189
  (
    n1213,
    n1191,
    n964,
    n998,
    n984
  );


  and
  g1190
  (
    n1203,
    n982,
    n1187,
    n992,
    n988
  );


  nand
  g1191
  (
    n1202,
    n967,
    n1199,
    n979,
    n1004
  );


  xor
  g1192
  (
    n1207,
    n1193,
    n1190,
    n971,
    n973
  );


  nand
  g1193
  (
    n1200,
    n975,
    n978,
    n981,
    n1189
  );


  or
  g1194
  (
    n1210,
    n1194,
    n1186,
    n991,
    n963
  );


  buf
  g1195
  (
    n1215,
    n1160
  );


  not
  g1196
  (
    n1217,
    n1211
  );


  xor
  g1197
  (
    n1214,
    n1210,
    n1160,
    n1212
  );


  xor
  g1198
  (
    n1216,
    n1213,
    n1161
  );


  not
  g1199
  (
    n1233,
    n792
  );


  buf
  g1200
  (
    n1222,
    n792
  );


  buf
  g1201
  (
    n1232,
    n1217
  );


  buf
  g1202
  (
    n1218,
    n1215
  );


  buf
  g1203
  (
    n1231,
    n1163
  );


  xor
  g1204
  (
    n1223,
    n1007,
    n1011,
    n1166,
    n1216
  );


  nor
  g1205
  (
    n1227,
    n1164,
    n1214,
    n1166,
    n1165
  );


  nor
  g1206
  (
    n1228,
    n1217,
    n1010,
    n793,
    n1163
  );


  nor
  g1207
  (
    n1219,
    n1012,
    n791,
    n1215,
    n1167
  );


  and
  g1208
  (
    n1221,
    n1006,
    n1215,
    n1216,
    n1217
  );


  xor
  g1209
  (
    n1224,
    n1164,
    n1005,
    n1214,
    n1015
  );


  xnor
  g1210
  (
    n1226,
    n1162,
    n1020,
    n1018,
    n1008
  );


  xor
  g1211
  (
    n1225,
    n1016,
    n371,
    n1013,
    n1014
  );


  xor
  g1212
  (
    n1220,
    n1165,
    n1019,
    n1021,
    n1216
  );


  or
  g1213
  (
    n1229,
    n1217,
    n1017,
    n1214
  );


  and
  g1214
  (
    n1230,
    n1216,
    n1215,
    n1009,
    n1162
  );


  nor
  g1215
  (
    n1235,
    n1218,
    n372,
    n376,
    n373
  );


  xor
  g1216
  (
    n1234,
    n1218,
    n1219,
    n373
  );


  and
  g1217
  (
    n1237,
    n1218,
    n1219,
    n374,
    n373
  );


  xnor
  g1218
  (
    n1240,
    n374,
    n372,
    n376,
    n375
  );


  nor
  g1219
  (
    n1238,
    n373,
    n375,
    n372
  );


  xor
  g1220
  (
    n1239,
    n371,
    n1218,
    n376,
    n375
  );


  or
  g1221
  (
    n1236,
    n374,
    n374,
    n375,
    n376
  );


  not
  g1222
  (
    n1244,
    n1237
  );


  buf
  g1223
  (
    n1246,
    n1239
  );


  not
  g1224
  (
    n1247,
    n1083
  );


  buf
  g1225
  (
    n1241,
    n1083
  );


  buf
  g1226
  (
    n1248,
    n1240
  );


  buf
  g1227
  (
    n1243,
    n377
  );


  and
  g1228
  (
    n1245,
    n1238,
    n377
  );


  nor
  g1229
  (
    n1242,
    n1235,
    n1236,
    n1240,
    n1234
  );


  nand
  g1230
  (
    KeyWire_0_37,
    n807,
    n807,
    n805,
    n1242
  );


  xnor
  g1231
  (
    n1258,
    n798,
    n1242,
    n1243,
    n802
  );


  and
  g1232
  (
    n1257,
    n806,
    n808,
    n799,
    n809
  );


  nand
  g1233
  (
    n1252,
    n803,
    n793,
    n809,
    n1243
  );


  xnor
  g1234
  (
    n1259,
    n795,
    n1242,
    n801,
    n804
  );


  and
  g1235
  (
    n1254,
    n794,
    n794,
    n803,
    n796
  );


  nand
  g1236
  (
    n1249,
    n806,
    n797,
    n1241,
    n1243
  );


  xnor
  g1237
  (
    n1255,
    n1241,
    n804,
    n799,
    n801
  );


  nor
  g1238
  (
    n1251,
    n800,
    n795,
    n802,
    n1242
  );


  xor
  g1239
  (
    n1256,
    n797,
    n798,
    n805,
    n800
  );


  nand
  g1240
  (
    n1253,
    n796,
    n808,
    n1241
  );


  or
  g1241
  (
    n1266,
    n1031,
    n1024,
    n1022,
    n1030
  );


  and
  g1242
  (
    n1264,
    n1030,
    n1028,
    n1032,
    n1256
  );


  xor
  g1243
  (
    n1262,
    n1034,
    n1031,
    n1252,
    n1026
  );


  nand
  g1244
  (
    n1267,
    n1259,
    n1027,
    n1254,
    n1032
  );


  xor
  g1245
  (
    n1263,
    n1026,
    n1025,
    n1253
  );


  nor
  g1246
  (
    n1260,
    n1258,
    n1029,
    n1028,
    n1024
  );


  and
  g1247
  (
    n1265,
    n1029,
    n1033,
    n1023
  );


  nor
  g1248
  (
    n1261,
    n1257,
    n1255,
    n1034,
    n1027
  );


  not
  g1249
  (
    n1269,
    n1260
  );


  buf
  g1250
  (
    n1270,
    n1260
  );


  not
  g1251
  (
    n1268,
    n1260
  );


  buf
  g1252
  (
    n1271,
    n1260
  );


  not
  g1253
  (
    n1274,
    n1261
  );


  buf
  g1254
  (
    n1273,
    n1261
  );


  not
  g1255
  (
    n1272,
    n1261
  );


  nand
  g1256
  (
    n1277,
    n1037,
    n1044,
    n810
  );


  xor
  g1257
  (
    KeyWire_0_8,
    n1271,
    n1274,
    n1039,
    n1041
  );


  nand
  g1258
  (
    n1285,
    n811,
    n1041,
    n1274,
    n1043
  );


  or
  g1259
  (
    n1278,
    n1047,
    n1272,
    n813,
    n1269
  );


  and
  g1260
  (
    n1282,
    n1046,
    n1046,
    n1038,
    n1270
  );


  nor
  g1261
  (
    n1279,
    n1037,
    n812,
    n1270,
    n1042
  );


  xnor
  g1262
  (
    n1280,
    n1042,
    n1045,
    n1273,
    n1048
  );


  or
  g1263
  (
    n1284,
    n1035,
    n1043,
    n813,
    n810
  );


  nor
  g1264
  (
    n1281,
    n1271,
    n1268,
    n1036,
    n1040
  );


  nor
  g1265
  (
    n1283,
    n1273,
    n1040,
    n1047,
    n1035
  );


  and
  g1266
  (
    n1276,
    n811,
    n812,
    n1036,
    n1039
  );


  or
  g1267
  (
    n1286,
    n1048,
    n1272,
    n1038,
    n1045
  );


  or
  g1268
  (
    n1294,
    n1275,
    n1179
  );


  or
  g1269
  (
    n1297,
    n1279,
    n1275,
    n1172,
    n1170
  );


  nor
  g1270
  (
    n1296,
    n1173,
    n1180,
    n1177,
    n1169
  );


  or
  g1271
  (
    n1295,
    n1174,
    n1276,
    n1278,
    n1173
  );


  nand
  g1272
  (
    n1289,
    n1178,
    n1177,
    n1277,
    n1278
  );


  or
  g1273
  (
    KeyWire_0_26,
    n1168,
    n1171,
    n1180,
    n1169
  );


  nand
  g1274
  (
    n1291,
    n1279,
    n1174,
    n1175,
    n1180
  );


  xnor
  g1275
  (
    n1290,
    n1167,
    n1277,
    n1171,
    n1276
  );


  or
  g1276
  (
    n1288,
    n1180,
    n1168,
    n1172,
    n1170
  );


  xnor
  g1277
  (
    n1293,
    n1176,
    n1179,
    n1178
  );


  nor
  g1278
  (
    n1287,
    n1280,
    n1178,
    n1176,
    n1175
  );


  buf
  g1279
  (
    n1299,
    n1288
  );


  buf
  g1280
  (
    n1301,
    n1288
  );


  buf
  g1281
  (
    n1298,
    n1287
  );


  not
  g1282
  (
    n1300,
    n1287
  );


  buf
  g1283
  (
    n1310,
    n1288
  );


  not
  g1284
  (
    n1309,
    n1247
  );


  not
  g1285
  (
    n1305,
    n1244
  );


  buf
  g1286
  (
    n1313,
    n1246
  );


  buf
  g1287
  (
    n1307,
    n1299
  );


  not
  g1288
  (
    n1311,
    n1298
  );


  xor
  g1289
  (
    n1315,
    n1288,
    n1246,
    n1248
  );


  xor
  g1290
  (
    n1312,
    n1246,
    n1300,
    n1244,
    n1248
  );


  xor
  g1291
  (
    n1304,
    n1244,
    n1300,
    n1301
  );


  or
  g1292
  (
    n1308,
    n1298,
    n1248,
    n1244,
    n1301
  );


  nand
  g1293
  (
    n1302,
    n1243,
    n1245,
    n1301
  );


  xnor
  g1294
  (
    n1306,
    n1246,
    n1245,
    n1247
  );


  xnor
  g1295
  (
    n1303,
    n1247,
    n1299
  );


  xnor
  g1296
  (
    KeyWire_0_48,
    n1245,
    n1245,
    n1049,
    n1300
  );


  not
  g1297
  (
    n1345,
    n1309
  );


  not
  g1298
  (
    KeyWire_0_31,
    n1291
  );


  not
  g1299
  (
    n1323,
    n1306
  );


  not
  g1300
  (
    n1344,
    n1306
  );


  buf
  g1301
  (
    n1356,
    n1314
  );


  buf
  g1302
  (
    n1362,
    n1310
  );


  not
  g1303
  (
    n1341,
    n1112
  );


  not
  g1304
  (
    KeyWire_0_47,
    n1314
  );


  buf
  g1305
  (
    n1343,
    n1293
  );


  not
  g1306
  (
    n1327,
    n1116
  );


  buf
  g1307
  (
    n1363,
    n1113
  );


  buf
  g1308
  (
    n1338,
    n1307
  );


  not
  g1309
  (
    n1336,
    n1181
  );


  not
  g1310
  (
    n1329,
    n1109
  );


  buf
  g1311
  (
    n1328,
    n1308
  );


  not
  g1312
  (
    n1352,
    n1115
  );


  buf
  g1313
  (
    n1349,
    n1111
  );


  not
  g1314
  (
    n1317,
    n1307
  );


  xnor
  g1315
  (
    n1325,
    n1110,
    n1296,
    n1292,
    n1306
  );


  xor
  g1316
  (
    n1359,
    n1116,
    n378,
    n1111,
    n1113
  );


  or
  g1317
  (
    n1334,
    n1109,
    n1289,
    n1313,
    n1295
  );


  nor
  g1318
  (
    n1321,
    n1050,
    n1311,
    n1297,
    n1295
  );


  or
  g1319
  (
    n1335,
    n1309,
    n1290,
    n1107,
    n1110
  );


  xnor
  g1320
  (
    n1330,
    n1312,
    n378,
    n1111,
    n1308
  );


  xnor
  g1321
  (
    n1360,
    n1293,
    n1112,
    n1290
  );


  or
  g1322
  (
    n1331,
    n1312,
    n1312,
    n1303,
    n1307
  );


  or
  g1323
  (
    n1326,
    n1112,
    n1309,
    n1108,
    n1053
  );


  xor
  g1324
  (
    n1358,
    n1302,
    n1294,
    n1114
  );


  xnor
  g1325
  (
    n1333,
    n1295,
    n1304,
    n1311,
    n1084
  );


  xor
  g1326
  (
    n1357,
    n1115,
    n1313,
    n1051,
    n1296
  );


  and
  g1327
  (
    n1337,
    n1312,
    n1302,
    n1305,
    n1115
  );


  xor
  g1328
  (
    n1316,
    n1315,
    n1306,
    n1293,
    n1289
  );


  nand
  g1329
  (
    n1339,
    n1290,
    n1297,
    n1294,
    n1315
  );


  nor
  g1330
  (
    n1348,
    n1052,
    n1303,
    n1108,
    n1115
  );


  or
  g1331
  (
    n1347,
    n1314,
    n1310,
    n1295,
    n1110
  );


  xnor
  g1332
  (
    n1324,
    n1114,
    n1296,
    n1313,
    n1310
  );


  xor
  g1333
  (
    n1346,
    n1111,
    n1051,
    n1309,
    n1292
  );


  or
  g1334
  (
    n1350,
    n1109,
    n1114,
    n1307,
    n1308
  );


  xor
  g1335
  (
    n1340,
    n1292,
    n1108,
    n1314,
    n1294
  );


  xnor
  g1336
  (
    n1353,
    n1181,
    n1315,
    n1313,
    n1110
  );


  nor
  g1337
  (
    n1320,
    n1293,
    n1291,
    n1109,
    n1049
  );


  xnor
  g1338
  (
    KeyWire_0_36,
    n1310,
    n1114,
    n1297,
    n1304
  );


  and
  g1339
  (
    n1361,
    n1084,
    n1116,
    n1296,
    n1311
  );


  xor
  g1340
  (
    n1318,
    n1052,
    n1311,
    n1305,
    n1084
  );


  or
  g1341
  (
    n1354,
    n1289,
    n1053,
    n1297,
    n1308
  );


  nor
  g1342
  (
    n1342,
    n1116,
    n1112,
    n1113,
    n1050
  );


  nor
  g1343
  (
    n1332,
    n1291,
    n1113,
    n1084,
    n1289
  );


  nand
  g1344
  (
    n1351,
    n1291,
    n1292,
    n1315,
    n1108
  );


  buf
  g1345
  (
    n1417,
    n1347
  );


  buf
  g1346
  (
    n1371,
    n1233
  );


  buf
  g1347
  (
    n1437,
    n1353
  );


  buf
  g1348
  (
    n1465,
    n1358
  );


  not
  g1349
  (
    n1445,
    n1285
  );


  not
  g1350
  (
    n1468,
    n1282
  );


  not
  g1351
  (
    n1373,
    n1223
  );


  not
  g1352
  (
    n1422,
    n1224
  );


  not
  g1353
  (
    n1493,
    n1356
  );


  buf
  g1354
  (
    n1530,
    n1333
  );


  buf
  g1355
  (
    n1535,
    n1355
  );


  not
  g1356
  (
    n1393,
    n1343
  );


  not
  g1357
  (
    n1416,
    n1228
  );


  not
  g1358
  (
    n1386,
    n1334
  );


  not
  g1359
  (
    n1555,
    n1324
  );


  buf
  g1360
  (
    n1449,
    n1262
  );


  not
  g1361
  (
    n1524,
    n1336
  );


  not
  g1362
  (
    n1486,
    n1341
  );


  buf
  g1363
  (
    n1447,
    n1348
  );


  buf
  g1364
  (
    n1474,
    n1222
  );


  not
  g1365
  (
    n1523,
    n1220
  );


  not
  g1366
  (
    n1375,
    n1359
  );


  not
  g1367
  (
    n1433,
    n1330
  );


  buf
  g1368
  (
    n1483,
    n1342
  );


  not
  g1369
  (
    n1406,
    n1183
  );


  buf
  g1370
  (
    n1476,
    n1332
  );


  buf
  g1371
  (
    n1459,
    n1339
  );


  not
  g1372
  (
    n1421,
    n1232
  );


  buf
  g1373
  (
    n1463,
    n1357
  );


  buf
  g1374
  (
    n1529,
    n1230
  );


  not
  g1375
  (
    n1439,
    n1350
  );


  not
  g1376
  (
    n1384,
    n1344
  );


  not
  g1377
  (
    n1527,
    n1265
  );


  not
  g1378
  (
    n1489,
    n1286
  );


  not
  g1379
  (
    n1400,
    n1349
  );


  not
  g1380
  (
    n1381,
    n1183
  );


  buf
  g1381
  (
    n1453,
    n1233
  );


  not
  g1382
  (
    n1541,
    n1226
  );


  not
  g1383
  (
    n1516,
    n1362
  );


  buf
  g1384
  (
    n1467,
    n1329
  );


  buf
  g1385
  (
    n1514,
    n1332
  );


  buf
  g1386
  (
    n1511,
    n1344
  );


  buf
  g1387
  (
    n1538,
    n1267
  );


  not
  g1388
  (
    n1394,
    n1352
  );


  buf
  g1389
  (
    n1518,
    n1229
  );


  buf
  g1390
  (
    n1390,
    n1331
  );


  not
  g1391
  (
    n1396,
    n1363
  );


  not
  g1392
  (
    n1427,
    n1353
  );


  buf
  g1393
  (
    n1423,
    n1350
  );


  not
  g1394
  (
    n1457,
    n1351
  );


  not
  g1395
  (
    n1547,
    n1232
  );


  not
  g1396
  (
    n1482,
    n1326
  );


  not
  g1397
  (
    n1448,
    n1225
  );


  not
  g1398
  (
    n1405,
    n1182
  );


  buf
  g1399
  (
    n1515,
    n1322
  );


  buf
  g1400
  (
    n1369,
    n1359
  );


  buf
  g1401
  (
    n1451,
    n1320
  );


  buf
  g1402
  (
    n1455,
    n1227
  );


  not
  g1403
  (
    n1548,
    n1318
  );


  not
  g1404
  (
    n1395,
    n1324
  );


  not
  g1405
  (
    KeyWire_0_14,
    n1137
  );


  buf
  g1406
  (
    n1495,
    n1324
  );


  not
  g1407
  (
    n1540,
    n1327
  );


  buf
  g1408
  (
    KeyWire_0_42,
    n1350
  );


  buf
  g1409
  (
    n1408,
    n1332
  );


  not
  g1410
  (
    n1522,
    n1354
  );


  not
  g1411
  (
    n1546,
    n1349
  );


  not
  g1412
  (
    n1380,
    n1330
  );


  buf
  g1413
  (
    n1365,
    n1134
  );


  not
  g1414
  (
    n1364,
    n1327
  );


  not
  g1415
  (
    n1436,
    n1232
  );


  not
  g1416
  (
    n1424,
    n1223
  );


  buf
  g1417
  (
    n1469,
    n1266
  );


  buf
  g1418
  (
    n1372,
    n1333
  );


  not
  g1419
  (
    n1413,
    n1326
  );


  buf
  g1420
  (
    n1415,
    n1356
  );


  not
  g1421
  (
    n1440,
    n1341
  );


  not
  g1422
  (
    n1426,
    n1319
  );


  buf
  g1423
  (
    n1434,
    n1282
  );


  buf
  g1424
  (
    n1501,
    n1136
  );


  buf
  g1425
  (
    n1487,
    n1321
  );


  buf
  g1426
  (
    n1500,
    n1283
  );


  buf
  g1427
  (
    n1401,
    n1319
  );


  not
  g1428
  (
    n1528,
    n1222
  );


  not
  g1429
  (
    n1484,
    n1338
  );


  buf
  g1430
  (
    n1499,
    n1340
  );


  buf
  g1431
  (
    n1450,
    n1331
  );


  not
  g1432
  (
    n1389,
    n1321
  );


  buf
  g1433
  (
    n1549,
    n1323
  );


  not
  g1434
  (
    KeyWire_0_60,
    n1329
  );


  not
  g1435
  (
    n1404,
    n1135
  );


  not
  g1436
  (
    n1477,
    n1342
  );


  not
  g1437
  (
    n1512,
    n1325
  );


  buf
  g1438
  (
    n1544,
    n1266
  );


  not
  g1439
  (
    n1480,
    n1338
  );


  buf
  g1440
  (
    n1475,
    n1334
  );


  not
  g1441
  (
    n1458,
    n1220
  );


  buf
  g1442
  (
    n1553,
    n1359
  );


  not
  g1443
  (
    n1551,
    n1340
  );


  not
  g1444
  (
    n1441,
    n1344
  );


  buf
  g1445
  (
    n1552,
    n1323
  );


  buf
  g1446
  (
    n1513,
    n1362
  );


  buf
  g1447
  (
    KeyWire_0_23,
    n1266
  );


  buf
  g1448
  (
    n1397,
    n1221
  );


  buf
  g1449
  (
    n1506,
    n1264
  );


  not
  g1450
  (
    n1526,
    n1228
  );


  buf
  g1451
  (
    n1517,
    n1142
  );


  not
  g1452
  (
    n1402,
    n1327
  );


  not
  g1453
  (
    n1509,
    n1322
  );


  not
  g1454
  (
    n1366,
    n1327
  );


  not
  g1455
  (
    n1479,
    n1330
  );


  buf
  g1456
  (
    n1391,
    n1349
  );


  not
  g1457
  (
    n1382,
    n1339
  );


  buf
  g1458
  (
    n1510,
    n1347
  );


  buf
  g1459
  (
    n1520,
    n1284
  );


  buf
  g1460
  (
    n1502,
    n1231
  );


  not
  g1461
  (
    n1503,
    n1233
  );


  buf
  g1462
  (
    n1473,
    n1262
  );


  not
  g1463
  (
    n1532,
    n1230
  );


  buf
  g1464
  (
    n1414,
    n1335
  );


  buf
  g1465
  (
    n1472,
    n1339
  );


  buf
  g1466
  (
    n1407,
    n378
  );


  not
  g1467
  (
    n1370,
    n1318
  );


  buf
  g1468
  (
    n1409,
    n1354
  );


  buf
  g1469
  (
    n1429,
    n1263
  );


  not
  g1470
  (
    n1462,
    n1345
  );


  not
  g1471
  (
    n1410,
    n1343
  );


  buf
  g1472
  (
    n1542,
    n1338
  );


  buf
  g1473
  (
    n1378,
    n1262
  );


  buf
  g1474
  (
    n1377,
    n1076
  );


  not
  g1475
  (
    n1545,
    n1335
  );


  not
  g1476
  (
    n1505,
    n1227
  );


  not
  g1477
  (
    n1508,
    n1317
  );


  buf
  g1478
  (
    n1443,
    n1325
  );


  not
  g1479
  (
    n1461,
    n1358
  );


  not
  g1480
  (
    n1418,
    n1266
  );


  not
  g1481
  (
    n1446,
    n1341
  );


  buf
  g1482
  (
    n1442,
    n1229
  );


  not
  g1483
  (
    n1411,
    n1320
  );


  not
  g1484
  (
    n1470,
    n1363
  );


  not
  g1485
  (
    n1398,
    n1355
  );


  not
  g1486
  (
    n1525,
    n1286
  );


  not
  g1487
  (
    n1497,
    n1267
  );


  buf
  g1488
  (
    n1403,
    n1318
  );


  not
  g1489
  (
    n1452,
    n1352
  );


  not
  g1490
  (
    n1456,
    n1320
  );


  buf
  g1491
  (
    n1464,
    n1325
  );


  buf
  g1492
  (
    n1534,
    n1267
  );


  buf
  g1493
  (
    n1444,
    n1228
  );


  not
  g1494
  (
    n1430,
    n1231
  );


  buf
  g1495
  (
    n1490,
    n1346
  );


  xor
  g1496
  (
    n1428,
    n1337,
    n1143,
    n1224
  );


  and
  g1497
  (
    n1419,
    n1359,
    n1340,
    n1221,
    n1337
  );


  xor
  g1498
  (
    n1478,
    n1356,
    n1345,
    n1316,
    n1224
  );


  xor
  g1499
  (
    n1521,
    n1231,
    n1264,
    n1138,
    n1183
  );


  xnor
  g1500
  (
    n1531,
    n1330,
    n1230,
    n1224,
    n1332
  );


  xnor
  g1501
  (
    n1536,
    n378,
    n1328,
    n1357,
    n1182
  );


  and
  g1502
  (
    n1387,
    n1347,
    n1358,
    n1348,
    n1344
  );


  xor
  g1503
  (
    n1460,
    n1317,
    n1362,
    n1324,
    n1319
  );


  xnor
  g1504
  (
    n1385,
    n1229,
    n1357,
    n1336,
    n1361
  );


  or
  g1505
  (
    KeyWire_0_11,
    n1329,
    n1323,
    n1346,
    n1348
  );


  or
  g1506
  (
    n1488,
    n1347,
    n1220,
    n1219,
    n1326
  );


  or
  g1507
  (
    n1537,
    n1338,
    n1319,
    n1263,
    n1182
  );


  or
  g1508
  (
    n1438,
    n1322,
    n1350,
    n1360,
    n1221
  );


  and
  g1509
  (
    n1368,
    n1230,
    n1345,
    n1363,
    n1286
  );


  and
  g1510
  (
    n1471,
    n1261,
    n1321,
    n1343,
    n1342
  );


  nand
  g1511
  (
    n1367,
    n1343,
    n1225,
    n1316,
    n1220
  );


  nor
  g1512
  (
    n1431,
    n1339,
    n1363,
    n1225,
    n1336
  );


  and
  g1513
  (
    n1496,
    n1357,
    n1329,
    n1326,
    n1334
  );


  nand
  g1514
  (
    n1507,
    n1349,
    n1286,
    n1264,
    n1328
  );


  or
  g1515
  (
    n1494,
    n1346,
    n1336,
    n1348,
    n1262
  );


  nand
  g1516
  (
    n1425,
    n1354,
    n1181,
    n1328,
    n1233
  );


  nand
  g1517
  (
    n1554,
    n1320,
    n1226,
    n1361,
    n1331
  );


  xor
  g1518
  (
    n1492,
    n1316,
    n1223,
    n1334,
    n1265
  );


  xnor
  g1519
  (
    n1485,
    n1361,
    n1141,
    n1227,
    n1140
  );


  nand
  g1520
  (
    n1519,
    n1356,
    n1182,
    n1264,
    n1318
  );


  or
  g1521
  (
    n1550,
    n1342,
    n1352,
    n1351,
    n1076
  );


  xnor
  g1522
  (
    n1533,
    n1360,
    n1265,
    n1317
  );


  nor
  g1523
  (
    n1498,
    n1337,
    n1285,
    n1283,
    n1335
  );


  and
  g1524
  (
    n1376,
    n1223,
    n1355,
    n1362,
    n1226
  );


  or
  g1525
  (
    n1491,
    n1355,
    n1183,
    n1227,
    n1280
  );


  nand
  g1526
  (
    n1454,
    n1263,
    n1139,
    n1267,
    n1322
  );


  or
  g1527
  (
    n1504,
    n1335,
    n1353,
    n1325,
    n1361
  );


  nor
  g1528
  (
    n1420,
    n1133,
    n1333,
    n1231,
    n1351
  );


  and
  g1529
  (
    n1435,
    n1265,
    n1263,
    n1341,
    n1181
  );


  or
  g1530
  (
    n1374,
    n1284,
    n1328,
    n1321,
    n1360
  );


  and
  g1531
  (
    n1392,
    n1354,
    n1226,
    n1337,
    n1229
  );


  nor
  g1532
  (
    n1383,
    n1222,
    n1353,
    n1345,
    n1225
  );


  or
  g1533
  (
    n1399,
    n1352,
    n1222,
    n1323,
    n1360
  );


  xor
  g1534
  (
    n1432,
    n1358,
    n1281,
    n1351,
    n1228
  );


  xnor
  g1535
  (
    n1388,
    n1316,
    n1340,
    n1221,
    n1232
  );


  nor
  g1536
  (
    n1379,
    n1346,
    n1331,
    n1333,
    n1281
  );


  not
  g1537
  (
    n1570,
    n1388
  );


  buf
  g1538
  (
    n1578,
    n1383
  );


  not
  g1539
  (
    n1559,
    n1376
  );


  not
  g1540
  (
    n1581,
    n1369
  );


  buf
  g1541
  (
    n1567,
    n1387
  );


  buf
  g1542
  (
    n1563,
    n1375
  );


  not
  g1543
  (
    n1576,
    n1368
  );


  not
  g1544
  (
    n1572,
    n1380
  );


  buf
  g1545
  (
    n1575,
    n1385
  );


  buf
  g1546
  (
    n1558,
    n1367
  );


  buf
  g1547
  (
    n1562,
    n1381
  );


  buf
  g1548
  (
    n1580,
    n1377
  );


  not
  g1549
  (
    n1566,
    n1374
  );


  buf
  g1550
  (
    n1574,
    n1378
  );


  buf
  g1551
  (
    n1569,
    n1373
  );


  buf
  g1552
  (
    n1579,
    n1371
  );


  not
  g1553
  (
    n1561,
    n1384
  );


  not
  g1554
  (
    n1577,
    n1370
  );


  not
  g1555
  (
    n1571,
    n1364
  );


  buf
  g1556
  (
    n1560,
    n1379
  );


  buf
  g1557
  (
    n1573,
    n1386
  );


  buf
  g1558
  (
    n1564,
    n1389
  );


  buf
  g1559
  (
    n1556,
    n1366
  );


  buf
  g1560
  (
    n1557,
    n1365
  );


  buf
  g1561
  (
    KeyWire_0_24,
    n1372
  );


  buf
  g1562
  (
    n1565,
    n1382
  );


  xor
  g1563
  (
    n1587,
    n1580,
    n1436,
    n1512,
    n1411
  );


  nand
  g1564
  (
    n1603,
    n1551,
    n1562,
    n1457,
    n1554
  );


  xnor
  g1565
  (
    n1636,
    n1548,
    n1556,
    n1569,
    n1463
  );


  or
  g1566
  (
    n1628,
    n1567,
    n1454,
    n1555,
    n1566
  );


  xnor
  g1567
  (
    n1635,
    n1475,
    n1444,
    n1563,
    n1572
  );


  nor
  g1568
  (
    n1616,
    n1465,
    n1443,
    n1490,
    n1557
  );


  xor
  g1569
  (
    n1597,
    n1502,
    n1568,
    n1408,
    n1496
  );


  and
  g1570
  (
    n1621,
    n1570,
    n1573,
    n1578,
    n1493
  );


  nand
  g1571
  (
    n1630,
    n1532,
    n1564,
    n1519,
    n1579
  );


  xnor
  g1572
  (
    n1589,
    n1570,
    n1425,
    n1545,
    n1553
  );


  nand
  g1573
  (
    n1639,
    n1451,
    n1553,
    n1421,
    n1453
  );


  and
  g1574
  (
    n1601,
    n1468,
    n1456,
    n1546,
    n1525
  );


  or
  g1575
  (
    n1612,
    n1581,
    n1471,
    n1445,
    n1488
  );


  xor
  g1576
  (
    n1638,
    n1554,
    n1497,
    n1409,
    n1460
  );


  nand
  g1577
  (
    n1586,
    n1571,
    n1573,
    n1510,
    n1434
  );


  or
  g1578
  (
    n1633,
    n1543,
    n1559,
    n1561,
    n1398
  );


  xnor
  g1579
  (
    n1609,
    n1489,
    n1413,
    n1580,
    n1576
  );


  nor
  g1580
  (
    n1615,
    n1418,
    n1564,
    n1415,
    n1539
  );


  nand
  g1581
  (
    n1640,
    n1528,
    n1544,
    n1547,
    n1426
  );


  xnor
  g1582
  (
    n1618,
    n1419,
    n1467,
    n1558,
    n1574
  );


  and
  g1583
  (
    n1596,
    n1535,
    n1478,
    n1499,
    n1412
  );


  xor
  g1584
  (
    n1637,
    n1414,
    n1550,
    n1508,
    n1404
  );


  or
  g1585
  (
    n1619,
    n1534,
    n1495,
    n1545,
    n1513
  );


  and
  g1586
  (
    n1641,
    n1579,
    n1532,
    n1410,
    n1565
  );


  and
  g1587
  (
    n1642,
    n1482,
    n1474,
    n1516,
    n1433
  );


  xor
  g1588
  (
    n1644,
    n1542,
    n1530,
    n1576,
    n1391
  );


  or
  g1589
  (
    KeyWire_0_52,
    n1473,
    n1432,
    n1548,
    n1539
  );


  nor
  g1590
  (
    KeyWire_0_33,
    n1530,
    n1536,
    n1578,
    n1438
  );


  nand
  g1591
  (
    n1591,
    n1403,
    n1561,
    n1483,
    n1515
  );


  xor
  g1592
  (
    n1629,
    n1555,
    n1427,
    n1533,
    n1578
  );


  and
  g1593
  (
    n1625,
    n1484,
    n1557,
    n1562,
    n1392
  );


  xor
  g1594
  (
    n1593,
    n1550,
    n1401,
    n1450,
    n1479
  );


  and
  g1595
  (
    n1631,
    n1581,
    n1544,
    n1514,
    n1429
  );


  xnor
  g1596
  (
    n1590,
    n1534,
    n1399,
    n1556,
    n1537
  );


  nor
  g1597
  (
    n1626,
    n1509,
    n1501,
    n1420,
    n1500
  );


  nand
  g1598
  (
    n1583,
    n1579,
    n1565,
    n1574,
    n1449
  );


  xor
  g1599
  (
    n1627,
    n1393,
    n1581,
    n1577,
    n1405
  );


  nor
  g1600
  (
    n1599,
    n1466,
    n1506,
    n1435,
    n1494
  );


  nand
  g1601
  (
    n1594,
    n1441,
    n1422,
    n1538,
    n1447
  );


  or
  g1602
  (
    n1614,
    n1567,
    n1535,
    n1558,
    n1523
  );


  xor
  g1603
  (
    n1632,
    n1452,
    n1396,
    n1529,
    n1520
  );


  xor
  g1604
  (
    n1645,
    n1575,
    n1462,
    n1480,
    n1448
  );


  xnor
  g1605
  (
    n1613,
    n1491,
    n1577,
    n1458,
    n1481
  );


  xor
  g1606
  (
    n1585,
    n1576,
    n1504,
    n1507,
    n1531
  );


  and
  g1607
  (
    n1608,
    n1543,
    n1430,
    n1390,
    n1547
  );


  xor
  g1608
  (
    n1622,
    n1579,
    n1549,
    n1472,
    n1439
  );


  xnor
  g1609
  (
    n1643,
    n1455,
    n1569,
    n1576,
    n1394
  );


  xnor
  g1610
  (
    n1600,
    n1503,
    n1533,
    n1470,
    n1538
  );


  xnor
  g1611
  (
    n1592,
    n1397,
    n1469,
    n1446,
    n1402
  );


  nand
  g1612
  (
    n1582,
    n1511,
    n1526,
    n1498,
    n1563
  );


  xor
  g1613
  (
    n1605,
    n1536,
    n1428,
    n1540,
    n1417
  );


  or
  g1614
  (
    n1584,
    n1560,
    n1486,
    n1546,
    n1522
  );


  nand
  g1615
  (
    n1620,
    n1581,
    n1572,
    n1459,
    n1549
  );


  nor
  g1616
  (
    n1606,
    n1537,
    n1518,
    n1406,
    n1531
  );


  or
  g1617
  (
    n1611,
    n1395,
    n1577,
    n1541,
    n1505
  );


  nor
  g1618
  (
    n1598,
    n1431,
    n1560,
    n1552
  );


  xor
  g1619
  (
    n1604,
    n1580,
    n1541,
    n1578,
    n1577
  );


  xnor
  g1620
  (
    n1588,
    n1485,
    n1477,
    n1416,
    n1580
  );


  xnor
  g1621
  (
    n1602,
    n1542,
    n1440,
    n1571,
    n1461
  );


  xor
  g1622
  (
    n1607,
    n1521,
    n1527,
    n1476,
    n1524
  );


  xnor
  g1623
  (
    n1624,
    n1575,
    n1551,
    n1566,
    n1540
  );


  and
  g1624
  (
    n1634,
    n1442,
    n1487,
    n1492,
    n1424
  );


  xor
  g1625
  (
    n1617,
    n1568,
    n1407,
    n1423,
    n1437
  );


  nor
  g1626
  (
    n1595,
    n1517,
    n1400,
    n1559,
    n1464
  );


  xor
  g1627
  (
    n1661,
    n1614,
    n1617,
    n1639,
    n1588
  );


  nand
  g1628
  (
    n1653,
    n1594,
    n1637,
    n1602,
    n1625
  );


  nand
  g1629
  (
    n1660,
    n1595,
    n1615,
    n1630,
    n1621
  );


  and
  g1630
  (
    n1649,
    n1631,
    n1636,
    n1638,
    n1592
  );


  and
  g1631
  (
    n1655,
    n1616,
    n1619,
    n1641,
    n1628
  );


  xnor
  g1632
  (
    n1650,
    n1585,
    n1644,
    n1607,
    n1597
  );


  nor
  g1633
  (
    n1647,
    n1642,
    n1583,
    n1582,
    n1584
  );


  nand
  g1634
  (
    n1656,
    n1622,
    n1598,
    n1593,
    n1609
  );


  nand
  g1635
  (
    n1659,
    n1608,
    n1620,
    n1590,
    n1618
  );


  xor
  g1636
  (
    n1657,
    n1627,
    n1610,
    n1586,
    n1601
  );


  nand
  g1637
  (
    n1658,
    n1604,
    n1603,
    n1613,
    n1612
  );


  xor
  g1638
  (
    n1646,
    n1640,
    n1599,
    n1634,
    n1606
  );


  or
  g1639
  (
    n1654,
    n1596,
    n1611,
    n1632,
    n1587
  );


  xnor
  g1640
  (
    n1652,
    n1591,
    n1626,
    n1589,
    n1645
  );


  nand
  g1641
  (
    n1651,
    n1623,
    n1635,
    n1643,
    n1629
  );


  nor
  g1642
  (
    n1648,
    n1605,
    n1600,
    n1624,
    n1633
  );


  nand
  g1643
  (
    n1665,
    n1652,
    n1651,
    n1648,
    n1653
  );


  xor
  g1644
  (
    n1663,
    n1657,
    n1650,
    n1646,
    n1649
  );


  xnor
  g1645
  (
    n1664,
    n1658,
    n1656,
    n1659,
    n1647
  );


  and
  g1646
  (
    n1662,
    n1655,
    n1661,
    n1654,
    n1660
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n673,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n313,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n467,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n746,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n895,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n820,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n516,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n717,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1275,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n751,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n1139,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1412,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n59,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1069,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1481,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n369,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n407,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1017,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n587,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n136,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1126,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n107,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n861,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n1543,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n1568,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n234,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1292,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1028,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n223,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1080,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n845,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1322,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n477,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n1623,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n822,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n339,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1355,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n1250,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n913,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n743,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n1151,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n207,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n1539,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n874,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n679,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n29,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n125,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n1319,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1314,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n594,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n848,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n354,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n1610,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1055,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n401,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n880,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n659,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n419,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n962,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n772,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n1466,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n1182,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n849,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n249,
    KeyNOTWire_0_63
  );


endmodule

