// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_202 written by SynthGen on 2021/04/05 11:23:24
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_202 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n659, n657, n632, n660, n627, n654, n644, n628,
 n634, n635, n646, n641, n648, n661, n652, n624,
 n906, n900, n896, n910, n983, n958, n1006, n973,
 n1017, n999, n976, n1011, n967, n1943, n2031, n2032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n659, n657, n632, n660, n627, n654, n644, n628,
 n634, n635, n646, n641, n648, n661, n652, n624,
 n906, n900, n896, n910, n983, n958, n1006, n973,
 n1017, n999, n976, n1011, n967, n1943, n2031, n2032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n625,
 n626, n629, n630, n631, n633, n636, n637, n638,
 n639, n640, n642, n643, n645, n647, n649, n650,
 n651, n653, n655, n656, n658, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n897,
 n898, n899, n901, n902, n903, n904, n905, n907,
 n908, n909, n911, n912, n913, n914, n915, n916,
 n917, n918, n919, n920, n921, n922, n923, n924,
 n925, n926, n927, n928, n929, n930, n931, n932,
 n933, n934, n935, n936, n937, n938, n939, n940,
 n941, n942, n943, n944, n945, n946, n947, n948,
 n949, n950, n951, n952, n953, n954, n955, n956,
 n957, n959, n960, n961, n962, n963, n964, n965,
 n966, n968, n969, n970, n971, n972, n974, n975,
 n977, n978, n979, n980, n981, n982, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n1000, n1001, n1002,
 n1003, n1004, n1005, n1007, n1008, n1009, n1010, n1012,
 n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021,
 n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
 n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
 n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
 n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
 n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
 n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
 n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
 n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
 n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
 n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
 n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
 n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
 n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
 n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
 n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
 n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
 n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
 n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
 n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
 n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
 n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
 n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
 n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
 n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
 n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
 n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
 n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
 n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
 n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
 n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
 n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
 n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
 n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
 n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
 n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
 n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
 n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
 n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
 n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
 n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
 n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
 n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
 n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
 n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
 n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
 n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
 n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
 n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
 n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
 n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
 n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
 n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
 n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
 n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
 n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
 n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
 n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
 n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
 n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
 n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
 n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
 n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
 n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
 n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
 n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
 n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
 n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
 n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
 n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
 n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
 n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
 n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
 n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
 n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
 n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
 n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
 n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
 n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
 n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
 n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
 n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
 n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
 n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
 n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
 n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
 n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
 n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
 n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
 n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
 n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
 n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
 n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
 n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
 n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
 n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
 n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
 n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
 n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
 n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
 n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
 n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
 n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
 n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
 n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
 n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
 n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
 n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
 n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
 n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
 n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
 n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
 n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
 n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
 n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
 n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
 n1942, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
 n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
 n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
 n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
 n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
 n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
 n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
 n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
 n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
 n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
 n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;

buf  g0 (n53, n26);
buf  g1 (n125, n9);
not  g2 (n127, n4);
not  g3 (n132, n6);
not  g4 (n99, n2);
not  g5 (n155, n14);
not  g6 (n74, n12);
not  g7 (n76, n13);
not  g8 (n55, n20);
buf  g9 (n157, n18);
not  g10 (n34, n11);
buf  g11 (n87, n21);
buf  g12 (n41, n10);
not  g13 (n129, n28);
buf  g14 (n50, n26);
buf  g15 (n150, n25);
buf  g16 (n82, n5);
buf  g17 (n63, n6);
not  g18 (n124, n6);
buf  g19 (n65, n18);
buf  g20 (n66, n15);
buf  g21 (n100, n4);
buf  g22 (n151, n24);
not  g23 (n89, n28);
not  g24 (n137, n25);
buf  g25 (n154, n1);
not  g26 (n88, n7);
not  g27 (n78, n30);
buf  g28 (n85, n25);
buf  g29 (n111, n32);
buf  g30 (n112, n3);
not  g31 (n62, n3);
buf  g32 (n57, n11);
buf  g33 (n49, n16);
not  g34 (n70, n32);
not  g35 (n114, n32);
buf  g36 (n119, n29);
buf  g37 (n71, n29);
not  g38 (n102, n18);
buf  g39 (n98, n32);
not  g40 (n68, n17);
not  g41 (n54, n19);
buf  g42 (n156, n25);
buf  g43 (n90, n21);
buf  g44 (n46, n23);
not  g45 (n149, n26);
buf  g46 (n110, n1);
not  g47 (n118, n27);
not  g48 (n38, n5);
not  g49 (n69, n22);
not  g50 (n103, n29);
not  g51 (n126, n14);
buf  g52 (n133, n8);
buf  g53 (n160, n29);
buf  g54 (n59, n31);
not  g55 (n152, n17);
not  g56 (n141, n6);
not  g57 (n113, n14);
buf  g58 (n44, n24);
buf  g59 (n61, n19);
buf  g60 (n117, n3);
not  g61 (n153, n12);
not  g62 (n92, n31);
not  g63 (n122, n4);
buf  g64 (n115, n10);
buf  g65 (n138, n2);
buf  g66 (n35, n11);
not  g67 (n95, n16);
not  g68 (n67, n7);
not  g69 (n86, n5);
not  g70 (n123, n22);
buf  g71 (n72, n24);
not  g72 (n77, n31);
not  g73 (n60, n28);
not  g74 (n33, n20);
not  g75 (n64, n21);
buf  g76 (n130, n10);
buf  g77 (n91, n22);
buf  g78 (n148, n11);
not  g79 (n145, n7);
not  g80 (n121, n23);
buf  g81 (n37, n17);
buf  g82 (n109, n9);
not  g83 (n84, n31);
not  g84 (n108, n15);
not  g85 (n51, n8);
not  g86 (n80, n9);
buf  g87 (n107, n30);
not  g88 (n75, n8);
buf  g89 (n131, n24);
buf  g90 (n42, n2);
not  g91 (n116, n2);
not  g92 (n93, n1);
buf  g93 (n73, n20);
not  g94 (n94, n17);
buf  g95 (n45, n13);
buf  g96 (n39, n18);
not  g97 (n139, n30);
buf  g98 (n147, n19);
not  g99 (n97, n9);
not  g100 (n40, n27);
buf  g101 (n136, n21);
buf  g102 (n144, n15);
buf  g103 (n58, n26);
buf  g104 (n36, n20);
not  g105 (n142, n27);
not  g106 (n48, n4);
not  g107 (n81, n14);
buf  g108 (n140, n13);
buf  g109 (n104, n23);
buf  g110 (n146, n15);
not  g111 (n135, n19);
buf  g112 (n158, n3);
buf  g113 (n83, n27);
not  g114 (n101, n16);
buf  g115 (n56, n23);
buf  g116 (n143, n1);
not  g117 (n105, n22);
buf  g118 (n52, n16);
buf  g119 (n128, n5);
not  g120 (n106, n8);
buf  g121 (n47, n7);
not  g122 (n79, n13);
not  g123 (n159, n28);
buf  g124 (n120, n10);
buf  g125 (n43, n12);
buf  g126 (n134, n12);
not  g127 (n96, n30);
not  g128 (n331, n33);
buf  g129 (n204, n48);
not  g130 (n203, n71);
buf  g131 (n293, n78);
not  g132 (n248, n59);
not  g133 (n229, n65);
buf  g134 (n241, n62);
not  g135 (n339, n56);
buf  g136 (n260, n51);
not  g137 (n325, n62);
not  g138 (n302, n76);
not  g139 (n333, n44);
not  g140 (n242, n58);
buf  g141 (n181, n68);
buf  g142 (n163, n65);
not  g143 (n244, n51);
not  g144 (n271, n55);
buf  g145 (n323, n64);
buf  g146 (n250, n72);
buf  g147 (n224, n67);
not  g148 (n329, n42);
not  g149 (n295, n42);
not  g150 (n274, n37);
not  g151 (n263, n45);
buf  g152 (n230, n64);
buf  g153 (n200, n48);
buf  g154 (n187, n77);
not  g155 (n313, n53);
buf  g156 (n310, n33);
buf  g157 (n175, n34);
not  g158 (n220, n78);
buf  g159 (n183, n76);
buf  g160 (n177, n58);
not  g161 (n174, n47);
buf  g162 (n179, n54);
not  g163 (n235, n44);
not  g164 (n164, n56);
not  g165 (n268, n35);
not  g166 (n321, n54);
not  g167 (n236, n70);
not  g168 (n275, n57);
buf  g169 (n217, n52);
not  g170 (n211, n35);
buf  g171 (n249, n46);
not  g172 (n286, n70);
buf  g173 (n305, n71);
buf  g174 (n343, n72);
not  g175 (n195, n57);
buf  g176 (n266, n40);
buf  g177 (n269, n43);
not  g178 (n334, n71);
not  g179 (n223, n79);
buf  g180 (n345, n45);
not  g181 (n228, n52);
not  g182 (n327, n33);
buf  g183 (n283, n40);
buf  g184 (n280, n57);
buf  g185 (n189, n61);
not  g186 (n287, n63);
not  g187 (n185, n46);
not  g188 (n259, n74);
buf  g189 (n320, n61);
not  g190 (n208, n38);
not  g191 (n328, n47);
not  g192 (n316, n48);
buf  g193 (n319, n60);
buf  g194 (n344, n61);
not  g195 (n304, n45);
not  g196 (n289, n71);
buf  g197 (n272, n33);
buf  g198 (n258, n49);
buf  g199 (n337, n73);
buf  g200 (n335, n59);
not  g201 (n265, n67);
not  g202 (n308, n68);
buf  g203 (n225, n58);
buf  g204 (n199, n69);
buf  g205 (n178, n66);
not  g206 (n276, n38);
not  g207 (n300, n76);
not  g208 (n197, n78);
buf  g209 (n284, n56);
buf  g210 (n218, n41);
not  g211 (n166, n41);
not  g212 (n253, n50);
buf  g213 (n309, n69);
buf  g214 (n307, n35);
not  g215 (n221, n78);
buf  g216 (n246, n39);
buf  g217 (n296, n61);
not  g218 (n173, n79);
buf  g219 (n194, n52);
not  g220 (n182, n60);
not  g221 (n215, n59);
not  g222 (n167, n50);
not  g223 (n170, n34);
buf  g224 (n162, n49);
not  g225 (n226, n62);
not  g226 (n292, n55);
not  g227 (n330, n65);
not  g228 (n238, n55);
buf  g229 (n227, n40);
not  g230 (n172, n63);
not  g231 (n188, n75);
not  g232 (n257, n56);
not  g233 (n267, n39);
not  g234 (n186, n34);
buf  g235 (n326, n77);
buf  g236 (n212, n44);
not  g237 (n322, n36);
not  g238 (n243, n70);
not  g239 (n306, n69);
not  g240 (n240, n73);
not  g241 (n340, n55);
not  g242 (n288, n53);
buf  g243 (n234, n34);
buf  g244 (n324, n51);
not  g245 (n303, n67);
not  g246 (n279, n36);
not  g247 (n256, n70);
buf  g248 (n202, n59);
buf  g249 (n201, n65);
buf  g250 (n315, n63);
buf  g251 (n252, n60);
buf  g252 (n233, n52);
buf  g253 (n314, n60);
not  g254 (n318, n74);
buf  g255 (n277, n41);
buf  g256 (n176, n64);
not  g257 (n262, n66);
not  g258 (n180, n42);
buf  g259 (n206, n43);
buf  g260 (n161, n73);
not  g261 (n285, n77);
buf  g262 (n346, n38);
not  g263 (n297, n73);
buf  g264 (n261, n66);
buf  g265 (n245, n46);
buf  g266 (n222, n68);
buf  g267 (n198, n44);
not  g268 (n281, n62);
buf  g269 (n301, n75);
not  g270 (n171, n42);
not  g271 (n291, n38);
not  g272 (n273, n37);
not  g273 (n254, n36);
buf  g274 (n332, n47);
not  g275 (n169, n35);
not  g276 (n278, n43);
not  g277 (n270, n39);
buf  g278 (n191, n47);
buf  g279 (n264, n72);
not  g280 (n210, n39);
buf  g281 (n338, n37);
not  g282 (n192, n66);
not  g283 (n255, n58);
not  g284 (n282, n57);
not  g285 (n232, n77);
buf  g286 (n290, n63);
buf  g287 (n251, n67);
buf  g288 (n209, n41);
buf  g289 (n207, n53);
not  g290 (n237, n50);
not  g291 (n205, n51);
not  g292 (n165, n54);
not  g293 (n216, n74);
buf  g294 (n219, n43);
buf  g295 (n342, n69);
not  g296 (n168, n45);
not  g297 (n213, n75);
not  g298 (n193, n76);
buf  g299 (n214, n64);
buf  g300 (n184, n53);
buf  g301 (n190, n50);
not  g302 (n311, n40);
buf  g303 (n299, n54);
buf  g304 (n298, n72);
not  g305 (n196, n49);
not  g306 (n341, n37);
buf  g307 (n336, n46);
not  g308 (n294, n75);
not  g309 (n231, n74);
buf  g310 (n317, n49);
not  g311 (n239, n48);
not  g312 (n312, n68);
buf  g313 (n247, n36);
not  g314 (n608, n211);
buf  g315 (n442, n287);
not  g316 (n582, n124);
buf  g317 (n418, n103);
not  g318 (n507, n154);
buf  g319 (n531, n270);
buf  g320 (n443, n129);
buf  g321 (n530, n142);
buf  g322 (n532, n130);
not  g323 (n552, n279);
buf  g324 (n491, n290);
buf  g325 (n524, n136);
not  g326 (n371, n257);
not  g327 (n470, n88);
buf  g328 (n449, n208);
buf  g329 (n489, n90);
buf  g330 (n368, n125);
not  g331 (n607, n189);
buf  g332 (n559, n256);
not  g333 (n444, n288);
buf  g334 (n410, n115);
buf  g335 (n372, n258);
buf  g336 (n569, n180);
not  g337 (n541, n254);
buf  g338 (n590, n114);
buf  g339 (n595, n247);
not  g340 (n415, n240);
buf  g341 (n610, n295);
not  g342 (n562, n236);
buf  g343 (n563, n95);
buf  g344 (n367, n195);
not  g345 (n550, n274);
not  g346 (n479, n203);
buf  g347 (n589, n126);
buf  g348 (n515, n282);
not  g349 (n476, n159);
not  g350 (n574, n143);
buf  g351 (n370, n241);
not  g352 (n396, n98);
buf  g353 (n452, n289);
not  g354 (n510, n288);
not  g355 (n435, n110);
buf  g356 (n437, n211);
not  g357 (n616, n93);
buf  g358 (n394, n80);
buf  g359 (n596, n131);
buf  g360 (n555, n210);
buf  g361 (n518, n183);
not  g362 (n487, n243);
not  g363 (n619, n141);
not  g364 (n440, n265);
not  g365 (n480, n141);
not  g366 (n409, n93);
buf  g367 (n420, n254);
buf  g368 (n473, n253);
not  g369 (n511, n127);
not  g370 (n427, n230);
not  g371 (n355, n136);
buf  g372 (n502, n258);
not  g373 (n430, n202);
buf  g374 (n587, n92);
buf  g375 (n349, n89);
buf  g376 (n542, n213);
buf  g377 (n615, n284);
not  g378 (n408, n221);
buf  g379 (n392, n91);
buf  g380 (n465, n121);
not  g381 (n428, n218);
buf  g382 (n389, n251);
buf  g383 (n477, n289);
not  g384 (n348, n96);
buf  g385 (n434, n155);
buf  g386 (n528, n101);
not  g387 (n436, n138);
buf  g388 (n441, n99);
buf  g389 (n475, n218);
not  g390 (n454, n286);
not  g391 (n356, n280);
buf  g392 (n488, n184);
buf  g393 (n404, n149);
buf  g394 (n463, n186);
not  g395 (n591, n89);
buf  g396 (n469, n272);
buf  g397 (n593, n281);
buf  g398 (n503, n132);
not  g399 (n419, n139);
not  g400 (n519, n81);
buf  g401 (n433, n235);
buf  g402 (n594, n231);
buf  g403 (n579, n156);
buf  g404 (n352, n256);
buf  g405 (n377, n263);
not  g406 (n557, n275);
buf  g407 (n583, n115);
not  g408 (n597, n235);
buf  g409 (n405, n120);
buf  g410 (n584, n188);
not  g411 (n588, n81);
not  g412 (n570, n117);
not  g413 (n585, n205);
not  g414 (n421, n110);
not  g415 (n361, n118);
buf  g416 (n453, n265);
not  g417 (n397, n200);
not  g418 (n412, n80);
buf  g419 (n496, n106);
not  g420 (n575, n145);
buf  g421 (n380, n279);
buf  g422 (n606, n118);
not  g423 (n544, n130);
buf  g424 (n572, n281);
not  g425 (n536, n223);
not  g426 (n383, n276);
buf  g427 (n365, n251);
buf  g428 (n450, n139);
not  g429 (n603, n105);
buf  g430 (n534, n107);
not  g431 (n364, n205);
not  g432 (n484, n114);
not  g433 (n467, n113);
buf  g434 (n546, n113);
not  g435 (n540, n148);
not  g436 (n390, n90);
buf  g437 (n611, n246);
not  g438 (n612, n273);
buf  g439 (n353, n143);
buf  g440 (n400, n107);
buf  g441 (n369, n252);
not  g442 (n567, n156);
buf  g443 (n483, n144);
not  g444 (n513, n285);
buf  g445 (n547, n158);
not  g446 (n388, n101);
not  g447 (n517, n130);
not  g448 (n432, n137);
not  g449 (n514, n236);
buf  g450 (n375, n247);
not  g451 (n374, n92);
buf  g452 (n499, n244);
buf  g453 (n581, n84);
buf  g454 (n521, n144);
buf  g455 (n558, n245);
not  g456 (n359, n98);
buf  g457 (n573, n108);
not  g458 (n598, n146);
buf  g459 (n568, n85);
buf  g460 (n527, n154);
not  g461 (n577, n269);
not  g462 (n347, n229);
buf  g463 (n382, n145);
not  g464 (n482, n257);
buf  g465 (n578, n290);
buf  g466 (n429, n134);
not  g467 (n402, n263);
buf  g468 (n509, n246);
buf  g469 (n414, n130);
not  g470 (n481, n87);
not  g471 (n423, n133);
not  g472 (n447, n234);
buf  g473 (n529, n91);
nor  g474 (n554, n292, n101, n90, n100);
nor  g475 (n592, n296, n114, n177, n145);
or   g476 (n399, n97, n277, n106, n185);
nor  g477 (n537, n141, n198, n95, n127);
xnor g478 (n535, n261, n110, n138, n226);
nand g479 (n501, n224, n151, n79, n96);
xnor g480 (n354, n135, n132, n262, n198);
and  g481 (n495, n121, n247, n81, n240);
or   g482 (n520, n87, n181, n185, n115);
xnor g483 (n360, n282, n229, n102, n139);
xor  g484 (n468, n90, n155, n183, n113);
or   g485 (n600, n102, n293, n233, n210);
nor  g486 (n466, n135, n125, n249, n284);
nand g487 (n508, n122, n137, n230, n81);
and  g488 (n526, n270, n106, n107, n248);
nor  g489 (n464, n228, n83, n151, n179);
nor  g490 (n556, n212, n114, n136, n242);
xor  g491 (n472, n148, n227, n184, n214);
nor  g492 (n564, n112, n140, n157, n142);
xor  g493 (n366, n116, n287, n283);
nand g494 (n500, n267, n111, n287, n192);
xor  g495 (n586, n154, n194, n193, n273);
nor  g496 (n460, n104, n201, n278, n217);
xnor g497 (n560, n233, n275, n142, n190);
xor  g498 (n358, n268, n272, n278, n106);
and  g499 (n457, n224, n103, n291, n134);
xnor g500 (n553, n294, n79, n128, n134);
xor  g501 (n576, n182, n158, n115);
nor  g502 (n492, n140, n132, n295, n197);
nand g503 (n494, n137, n225, n126, n279);
xor  g504 (n566, n97, n89, n104, n290);
nand g505 (n406, n104, n112, n249, n262);
nand g506 (n545, n82, n244, n151, n105);
nand g507 (n571, n84, n269, n128, n131);
xor  g508 (n373, n255, n199, n98, n249);
xor  g509 (n613, n241, n264, n232, n121);
nor  g510 (n471, n294, n296, n276, n128);
or   g511 (n490, n269, n293, n239, n83);
nand g512 (n522, n237, n251, n207, n186);
xor  g513 (n416, n255, n213, n120, n248);
xnor g514 (n381, n153, n191, n223, n96);
xor  g515 (n474, n239, n286, n266, n117);
xor  g516 (n618, n148, n103, n88, n86);
nand g517 (n533, n109, n84, n267, n129);
and  g518 (n512, n149, n126, n87, n138);
nand g519 (n425, n209, n85, n242, n132);
nor  g520 (n411, n111, n271, n144, n252);
nand g521 (n395, n291, n285, n284, n146);
xnor g522 (n431, n120, n189, n277, n85);
nand g523 (n580, n121, n82, n216, n125);
nand g524 (n561, n260, n119, n195, n110);
xor  g525 (n357, n83, n138, n266, n259);
nand g526 (n378, n82, n94, n101, n149);
xor  g527 (n549, n98, n212, n99, n147);
xor  g528 (n505, n86, n262, n133, n144);
xnor g529 (n525, n158, n246, n257, n86);
nor  g530 (n363, n153, n146, n143, n271);
xor  g531 (n422, n91, n105, n120, n243);
xnor g532 (n461, n152, n260, n116, n202);
or   g533 (n504, n252, n122, n295, n245);
or   g534 (n403, n253, n95, n187, n125);
and  g535 (n451, n150, n143, n153, n95);
xnor g536 (n448, n155, n237, n219, n197);
and  g537 (n386, n228, n196, n234, n84);
or   g538 (n497, n127, n219, n190, n118);
xnor g539 (n376, n275, n258, n221, n268);
xnor g540 (n506, n192, n127, n118, n199);
nand g541 (n362, n274, n281, n261, n100);
nand g542 (n614, n194, n292, n265, n150);
or   g543 (n523, n232, n153, n93, n274);
or   g544 (n458, n113, n244, n157, n250);
nor  g545 (n393, n214, n286, n222, n282);
and  g546 (n485, n159, n137, n294, n278);
or   g547 (n401, n80, n141, n108, n260);
and  g548 (n350, n225, n270, n83, n112);
and  g549 (n417, n204, n291, n253, n261);
nand g550 (n424, n220, n243, n119, n104);
xnor g551 (n538, n111, n117, n92, n241);
nand g552 (n379, n135, n196, n248, n102);
xnor g553 (n462, n146, n94, n119);
nor  g554 (n455, n123, n182, n107, n108);
xnor g555 (n609, n93, n250, n157, n124);
xor  g556 (n565, n123, n191, n254, n82);
xnor g557 (n548, n216, n272, n129, n147);
nand g558 (n602, n208, n289, n207, n89);
and  g559 (n617, n85, n135, n99, n86);
nand g560 (n498, n222, n88, n215, n80);
and  g561 (n516, n259, n264, n126, n200);
nor  g562 (n426, n152, n97, n123, n117);
nand g563 (n439, n148, n103, n187, n131);
and  g564 (n445, n156, n288, n109, n87);
or   g565 (n385, n250, n122, n152, n131);
xor  g566 (n486, n255, n268, n112, n285);
xor  g567 (n478, n109, n193, n116, n215);
or   g568 (n446, n124, n178, n140, n271);
xnor g569 (n459, n155, n150, n283);
nand g570 (n413, n119, n129, n242, n256);
xnor g571 (n438, n152, n123, n111, n133);
xnor g572 (n391, n267, n217, n201, n276);
nand g573 (n351, n293, n128, n91, n97);
nand g574 (n456, n188, n100, n149, n151);
xor  g575 (n604, n292, n245, n147, n263);
xnor g576 (n543, n159, n238, n259, n204);
nand g577 (n387, n116, n99, n96, n266);
nor  g578 (n384, n100, n134, n209, n122);
nand g579 (n407, n139, n136, n92, n105);
and  g580 (n601, n140, n206, n157, n264);
and  g581 (n605, n226, n206, n156, n142);
and  g582 (n493, n227, n109, n159, n154);
and  g583 (n398, n238, n94, n133, n88);
xor  g584 (n599, n203, n277, n124, n273);
nor  g585 (n551, n231, n102, n220, n145);
nand g586 (n539, n147, n280, n108);
not  g587 (n655, n361);
buf  g588 (n654, n355);
buf  g589 (n624, n383);
buf  g590 (n659, n362);
buf  g591 (n652, n360);
buf  g592 (n642, n376);
not  g593 (n648, n379);
not  g594 (n622, n375);
buf  g595 (n658, n365);
buf  g596 (n638, n351);
buf  g597 (n626, n353);
not  g598 (n651, n349);
buf  g599 (n627, n386);
not  g600 (n643, n369);
not  g601 (n660, n374);
not  g602 (n625, n370);
buf  g603 (n641, n371);
buf  g604 (n623, n388);
not  g605 (n632, n350);
not  g606 (n650, n373);
buf  g607 (n637, n359);
buf  g608 (n636, n378);
not  g609 (n628, n368);
buf  g610 (n646, n348);
buf  g611 (n649, n372);
buf  g612 (n657, n347);
not  g613 (n656, n367);
buf  g614 (n620, n354);
not  g615 (n633, n352);
not  g616 (n639, n387);
not  g617 (n647, n358);
not  g618 (n644, n363);
buf  g619 (n640, n377);
buf  g620 (n629, n382);
not  g621 (n631, n357);
not  g622 (n661, n385);
buf  g623 (n634, n366);
buf  g624 (n645, n364);
not  g625 (n653, n356);
buf  g626 (n621, n384);
not  g627 (n630, n380);
not  g628 (n635, n381);
buf  g629 (n727, n620);
not  g630 (n761, n649);
buf  g631 (n704, n487);
not  g632 (n746, n412);
not  g633 (n747, n482);
buf  g634 (n705, n460);
not  g635 (n680, n479);
not  g636 (n763, n654);
not  g637 (n670, n623);
buf  g638 (n716, n631);
not  g639 (n718, n406);
buf  g640 (n675, n629);
not  g641 (n767, n428);
buf  g642 (n698, n659);
not  g643 (n699, n494);
buf  g644 (n734, n391);
buf  g645 (n684, n394);
not  g646 (n742, n500);
buf  g647 (n754, n627);
buf  g648 (n773, n503);
buf  g649 (n781, n431);
buf  g650 (n772, n493);
not  g651 (n725, n621);
not  g652 (n715, n648);
not  g653 (n723, n644);
buf  g654 (n768, n450);
not  g655 (n749, n441);
buf  g656 (n710, n625);
not  g657 (n757, n397);
not  g658 (n735, n474);
buf  g659 (n674, n415);
not  g660 (n721, n644);
not  g661 (n711, n443);
not  g662 (n738, n659);
buf  g663 (n726, n484);
not  g664 (n744, n650);
not  g665 (n697, n422);
buf  g666 (n766, n449);
buf  g667 (n717, n437);
not  g668 (n682, n480);
buf  g669 (n770, n398);
not  g670 (n759, n399);
not  g671 (n708, n409);
buf  g672 (n732, n429);
buf  g673 (n664, n447);
buf  g674 (n758, n489);
buf  g675 (n774, n632);
not  g676 (n776, n462);
buf  g677 (n692, n456);
buf  g678 (n671, n496);
not  g679 (n683, n639);
buf  g680 (n756, n435);
not  g681 (n709, n625);
not  g682 (n729, n626);
buf  g683 (n700, n490);
buf  g684 (n688, n628);
buf  g685 (n740, n469);
buf  g686 (n753, n621);
not  g687 (n663, n622);
not  g688 (n779, n402);
or   g689 (n672, n476, n470, n643);
xor  g690 (n771, n632, n466, n644);
nor  g691 (n764, n463, n433, n650);
xor  g692 (n669, n446, n423, n646);
or   g693 (n695, n646, n629, n438);
or   g694 (n681, n504, n392, n657);
xor  g695 (n712, n645, n624, n486);
xnor g696 (n687, n408, n637, n471);
and  g697 (n706, n419, n414, n626);
nor  g698 (n666, n396, n622, n635);
or   g699 (n728, n620, n652, n418);
or   g700 (n714, n654, n401, n393);
nand g701 (n755, n641, n630, n404);
nand g702 (n769, n426, n461, n637);
nor  g703 (n679, n472, n389, n459);
xnor g704 (n775, n651, n631, n465);
or   g705 (n686, n656, n458, n395);
or   g706 (n696, n636, n626, n468);
xor  g707 (n777, n647, n634, n633);
xnor g708 (n713, n658, n507, n457);
and  g709 (n737, n648, n656, n453);
xor  g710 (n724, n467, n652, n628);
nor  g711 (n668, n646, n623, n491);
xor  g712 (n707, n464, n439, n645);
nand g713 (n741, n630, n651, n637);
and  g714 (n739, n432, n657, n643);
nand g715 (n662, n647, n400, n653);
nor  g716 (n752, n481, n417, n508);
nor  g717 (n743, n655, n636, n640);
or   g718 (n733, n483, n451, n440);
and  g719 (n691, n407, n639, n649);
xnor g720 (n690, n623, n624, n657);
xor  g721 (n720, n658, n448, n444);
and  g722 (n677, n621, n454, n434);
nand g723 (n676, n655, n497, n654);
nor  g724 (n736, n648, n642, n629);
or   g725 (n778, n625, n405, n638);
nor  g726 (n762, n410, n477, n424);
and  g727 (n731, n633, n420, n442);
and  g728 (n667, n638, n620, n632);
xor  g729 (n748, n653, n641, n634);
xnor g730 (n678, n622, n488, n635);
nand g731 (n685, n498, n416, n390);
xnor g732 (n780, n492, n642, n403);
nand g733 (n722, n653, n647, n505);
nor  g734 (n689, n645, n495, n485);
nand g735 (n765, n652, n436, n627);
or   g736 (n760, n455, n445, n649);
nor  g737 (n719, n640, n633, n473);
nor  g738 (n701, n427, n475, n478);
nand g739 (n702, n628, n636, n655);
xnor g740 (n673, n630, n640, n425);
or   g741 (n751, n650, n421, n639);
and  g742 (n750, n635, n501, n430);
xor  g743 (n745, n411, n499, n656);
nor  g744 (n693, n643, n634, n642);
nor  g745 (n730, n506, n624, n641);
xor  g746 (n665, n452, n627, n651);
and  g747 (n694, n631, n502, n413);
xor  g748 (n703, n658, n659, n638);
xor  g749 (n790, n330, n304, n311, n329);
xnor g750 (n810, n312, n300, n338, n662);
or   g751 (n800, n336, n297, n680, n314);
nor  g752 (n793, n303, n346, n695, n333);
xor  g753 (n795, n298, n330, n343, n306);
xnor g754 (n802, n337, n686, n314, n318);
and  g755 (n785, n696, n336, n666, n327);
xnor g756 (n799, n302, n309, n300, n310);
xor  g757 (n809, n298, n328, n675, n324);
nand g758 (n801, n704, n320, n344, n331);
nor  g759 (n798, n682, n338, n331, n707);
nor  g760 (n797, n308, n683, n681, n708);
xor  g761 (n794, n312, n303, n302, n335);
nand g762 (n829, n697, n318, n671, n304);
xor  g763 (n821, n312, n345, n700, n324);
nor  g764 (n787, n332, n307, n667, n509);
or   g765 (n811, n325, n332, n692, n330);
xnor g766 (n828, n301, n344, n314, n322);
xor  g767 (n816, n313, n301, n337, n706);
nand g768 (n815, n321, n690, n342, n323);
xnor g769 (n813, n339, n332, n321, n305);
nor  g770 (n817, n670, n337, n676, n694);
xor  g771 (n792, n328, n334, n319, n299);
xor  g772 (n806, n340, n344, n674, n326);
xnor g773 (n827, n313, n687, n688, n705);
or   g774 (n805, n308, n709, n341, n342);
xor  g775 (n822, n307, n320, n685, n298);
nand g776 (n788, n322, n340, n343, n335);
or   g777 (n826, n663, n678, n300, n323);
xnor g778 (n789, n335, n345, n317, n339);
xnor g779 (n808, n664, n311, n702, n333);
xor  g780 (n786, n334, n315, n309);
or   g781 (n823, n693, n306, n329);
xnor g782 (n819, n310, n684, n304, n673);
nand g783 (n820, n308, n669, n323, n336);
xnor g784 (n830, n331, n299, n339, n703);
and  g785 (n783, n672, n319, n305, n689);
or   g786 (n796, n297, n317, n303, n333);
xor  g787 (n824, n668, n321, n309, n318);
xnor g788 (n807, n325, n305, n334, n701);
or   g789 (n818, n345, n691, n324, n341);
xor  g790 (n803, n327, n297, n307, n302);
or   g791 (n825, n329, n342, n665, n677);
and  g792 (n784, n698, n296, n340, n320);
xnor g793 (n831, n316, n328, n299, n338);
and  g794 (n782, n311, n327, n326, n317);
xnor g795 (n814, n301, n315, n319, n343);
or   g796 (n791, n710, n326, n322, n341);
xor  g797 (n804, n313, n310, n316);
nand g798 (n812, n711, n699, n679, n325);
buf  g799 (n842, n565);
buf  g800 (n888, n796);
buf  g801 (n878, n795);
buf  g802 (n889, n602);
not  g803 (n844, n782);
buf  g804 (n859, n566);
buf  g805 (n854, n786);
not  g806 (n874, n790);
buf  g807 (n846, n608);
buf  g808 (n840, n797);
buf  g809 (n834, n559);
not  g810 (n865, n586);
buf  g811 (n864, n580);
not  g812 (n881, n596);
buf  g813 (n845, n795);
not  g814 (n867, n712);
buf  g815 (n858, n526);
not  g816 (n838, n792);
buf  g817 (n860, n796);
not  g818 (n849, n521);
not  g819 (n879, n594);
buf  g820 (n850, n532);
not  g821 (n877, n784);
not  g822 (n856, n572);
not  g823 (n873, n550);
and  g824 (n866, n564, n569, n796);
xnor g825 (n851, n796, n605, n552, n535);
and  g826 (n841, n563, n786, n588, n790);
xnor g827 (n876, n787, n795, n528, n589);
xor  g828 (n884, n593, n579, n542, n567);
and  g829 (n862, n603, n585, n788, n793);
and  g830 (n872, n571, n544, n789, n520);
xnor g831 (n855, n561, n714, n797, n514);
xor  g832 (n843, n530, n546, n788, n573);
or   g833 (n871, n533, n537, n536, n551);
and  g834 (n869, n787, n793, n590, n513);
xnor g835 (n880, n539, n578, n785, n555);
and  g836 (n832, n789, n568, n548, n538);
and  g837 (n870, n785, n782, n597, n613);
and  g838 (n863, n790, n784, n609, n793);
or   g839 (n891, n788, n547, n560, n529);
xnor g840 (n882, n599, n791, n519, n581);
xnor g841 (n883, n793, n527, n786, n787);
nor  g842 (n885, n554, n788, n545, n595);
xnor g843 (n837, n574, n516, n524, n610);
xor  g844 (n835, n517, n510, n525, n607);
or   g845 (n875, n562, n791, n518, n556);
nand g846 (n861, n511, n540, n785, n794);
and  g847 (n853, n794, n790, n543, n591);
and  g848 (n857, n587, n592, n515, n582);
nor  g849 (n890, n792, n612, n782, n797);
and  g850 (n852, n601, n606, n557, n783);
xnor g851 (n886, n534, n604, n783, n576);
or   g852 (n892, n789, n792, n512, n577);
or   g853 (n868, n784, n523, n522, n787);
xor  g854 (n847, n575, n795, n786, n553);
nand g855 (n839, n794, n598, n570, n558);
xor  g856 (n848, n600, n791, n531, n789);
xor  g857 (n836, n783, n611, n797, n583);
nand g858 (n833, n584, n792, n549, n791);
nor  g859 (n887, n713, n541, n794, n785);
xor  g860 (n910, n834, n835, n732, n740);
xnor g861 (n899, n738, n717, n834, n833);
or   g862 (n902, n724, n798, n718);
or   g863 (n903, n832, n738, n727, n835);
or   g864 (n894, n723, n737, n739, n832);
or   g865 (n895, n736, n660, n728, n835);
and  g866 (n896, n725, n735, n833, n726);
or   g867 (n893, n834, n743, n798);
or   g868 (n909, n736, n660, n728);
and  g869 (n900, n740, n661, n833);
and  g870 (n908, n722, n734, n661, n833);
and  g871 (n904, n743, n836, n733, n742);
nand g872 (n898, n715, n744, n732, n836);
or   g873 (n897, n737, n741, n729, n739);
nand g874 (n901, n729, n836, n730, n742);
xnor g875 (n912, n741, n744, n731, n727);
or   g876 (n906, n836, n837, n735, n730);
nor  g877 (n905, n835, n733, n834, n720);
nand g878 (n907, n721, n731, n660, n832);
nand g879 (n911, n716, n734, n719, n661);
buf  g880 (n916, n747);
not  g881 (n915, n905);
not  g882 (n919, n900);
buf  g883 (n913, n897);
and  g884 (n914, n901, n899, n748, n749);
and  g885 (n921, n751, n745, n746, n747);
and  g886 (n917, n751, n745, n898, n750);
xor  g887 (n918, n749, n752, n903, n750);
or   g888 (n920, n746, n904, n748, n902);
xor  g889 (n957, n814, n815, n813, n810);
nor  g890 (n955, n918, n818, n914, n804);
nand g891 (n922, n804, n913, n917, n817);
or   g892 (n951, n810, n817, n913, n921);
nor  g893 (n949, n811, n815, n810, n916);
nor  g894 (n952, n814, n916, n808, n801);
nor  g895 (n931, n914, n811, n802, n803);
nand g896 (n932, n801, n824, n805, n806);
nor  g897 (n943, n824, n819, n812, n822);
or   g898 (n937, n802, n807, n819, n808);
nor  g899 (n946, n800, n816, n913, n814);
nand g900 (n942, n801, n811, n816, n920);
or   g901 (n936, n814, n805, n813, n810);
nand g902 (n940, n920, n803, n915, n806);
and  g903 (n956, n818, n807, n808, n800);
and  g904 (n941, n799, n812, n820, n813);
nor  g905 (n935, n809, n917, n916, n821);
and  g906 (n938, n920, n915, n799, n919);
and  g907 (n925, n809, n918, n823, n807);
xor  g908 (n948, n823, n802, n822);
or   g909 (n939, n805, n812, n915, n809);
nand g910 (n929, n815, n919, n820);
nand g911 (n944, n813, n917, n799, n811);
xor  g912 (n954, n825, n818, n918, n914);
nor  g913 (n923, n917, n801, n804, n803);
and  g914 (n924, n800, n918, n819, n820);
or   g915 (n930, n800, n752, n817, n921);
nor  g916 (n945, n753, n821, n914);
and  g917 (n950, n805, n817, n815, n823);
or   g918 (n953, n915, n816, n920, n913);
nand g919 (n926, n816, n821, n753, n812);
nand g920 (n927, n806, n808, n818, n804);
and  g921 (n947, n803, n921, n807, n809);
xor  g922 (n928, n820, n921, n806, n802);
nand g923 (n933, n919, n823, n824, n822);
and  g924 (n934, n824, n819, n916, n799);
and  g925 (n1014, n876, n843, n869, n928);
xnor g926 (n1003, n839, n856, n875, n867);
xnor g927 (n981, n850, n841, n937, n938);
and  g928 (n983, n848, n875, n863, n844);
xor  g929 (n1011, n853, n949, n889, n944);
xnor g930 (n1001, n838, n888, n883, n940);
or   g931 (n1017, n863, n948, n945, n886);
or   g932 (n1026, n842, n941, n888, n868);
or   g933 (n993, n936, n855, n878);
xnor g934 (n986, n861, n932, n930, n945);
xnor g935 (n1009, n866, n841, n862, n846);
and  g936 (n994, n859, n885, n875, n851);
xnor g937 (n1004, n870, n869, n857, n860);
nand g938 (n1024, n878, n841, n890, n845);
xnor g939 (n965, n862, n931, n847, n876);
and  g940 (n1025, n879, n855, n876, n926);
or   g941 (n1028, n843, n943, n935, n874);
xor  g942 (n977, n852, n838, n879, n864);
xor  g943 (n1005, n853, n856, n930, n852);
nor  g944 (n968, n924, n838, n883, n881);
nand g945 (n1000, n859, n861, n937, n865);
nand g946 (n1021, n874, n840, n842, n947);
nor  g947 (n961, n849, n928, n861, n883);
nor  g948 (n974, n890, n875, n862, n837);
xor  g949 (n1030, n924, n889, n943, n860);
nor  g950 (n1012, n856, n881, n939, n864);
nand g951 (n997, n932, n938, n891, n863);
xor  g952 (n978, n855, n845, n851, n868);
and  g953 (n976, n935, n840, n939, n877);
nor  g954 (n991, n871, n888, n950, n857);
xnor g955 (n1020, n882, n847, n858, n870);
xnor g956 (n1018, n884, n859, n891, n882);
xnor g957 (n989, n949, n844, n866, n838);
nand g958 (n980, n890, n945, n948, n942);
and  g959 (n988, n869, n922, n848, n843);
and  g960 (n975, n873, n840, n870, n889);
nor  g961 (n1002, n880, n881, n940, n841);
nand g962 (n1019, n871, n858, n865, n849);
xnor g963 (n996, n844, n852, n944, n949);
and  g964 (n1007, n942, n874, n950, n868);
xor  g965 (n966, n837, n864, n839, n871);
or   g966 (n979, n943, n863, n941, n946);
or   g967 (n1015, n873, n845, n851, n860);
nor  g968 (n1022, n947, n868, n933, n941);
xnor g969 (n969, n869, n940, n938, n854);
or   g970 (n973, n936, n880, n864, n850);
xor  g971 (n1029, n887, n926, n853, n867);
nor  g972 (n971, n891, n888, n925, n877);
xor  g973 (n1023, n882, n848, n887, n854);
and  g974 (n1006, n839, n946, n850, n934);
and  g975 (n1008, n847, n872, n923, n874);
and  g976 (n982, n950, n933, n891, n844);
xnor g977 (n963, n854, n878, n853, n846);
nor  g978 (n972, n872, n854, n849, n846);
xor  g979 (n958, n877, n879, n866, n843);
nor  g980 (n1027, n884, n885, n927, n939);
nor  g981 (n959, n871, n858, n840, n872);
xnor g982 (n970, n946, n847, n887, n883);
or   g983 (n990, n886, n884, n934, n859);
xnor g984 (n998, n865, n885, n837, n882);
nand g985 (n1013, n923, n873, n852, n944);
xnor g986 (n1016, n866, n925, n842, n942);
or   g987 (n992, n880, n947, n929, n879);
xnor g988 (n987, n862, n922, n881, n858);
and  g989 (n999, n860, n884, n846, n867);
xor  g990 (n984, n929, n927, n880, n887);
xor  g991 (n967, n845, n885, n861, n850);
xor  g992 (n964, n876, n878, n877, n870);
nor  g993 (n960, n857, n839, n886);
xor  g994 (n985, n856, n848, n889, n842);
and  g995 (n1010, n948, n873, n872, n931);
or   g996 (n995, n849, n851, n936, n867);
xnor g997 (n962, n890, n857, n937, n865);
not  g998 (n1077, n974);
buf  g999 (n1065, n759);
not  g1000 (n1034, n984);
buf  g1001 (n1060, n911);
buf  g1002 (n1080, n757);
buf  g1003 (n1085, n827);
not  g1004 (n1037, n828);
buf  g1005 (n1051, n1011);
not  g1006 (n1071, n754);
not  g1007 (n1032, n908);
buf  g1008 (n1056, n1016);
not  g1009 (n1086, n975);
buf  g1010 (n1061, n971);
not  g1011 (n1041, n754);
not  g1012 (n1053, n1020);
not  g1013 (n1031, n967);
not  g1014 (n1042, n826);
not  g1015 (n1048, n825);
buf  g1016 (n1045, n829);
not  g1017 (n1093, n907);
buf  g1018 (n1057, n1010);
buf  g1019 (n1070, n758);
not  g1020 (n1054, n1001);
not  g1021 (n1064, n755);
buf  g1022 (n1069, n1026);
buf  g1023 (n1036, n761);
not  g1024 (n1047, n828);
not  g1025 (n1076, n764);
not  g1026 (n1067, n764);
buf  g1027 (n1079, n827);
not  g1028 (n1058, n997);
buf  g1029 (n1068, n1014);
buf  g1030 (n1039, n983);
not  g1031 (n1043, n757);
buf  g1032 (n1081, n988);
buf  g1033 (n1038, n826);
buf  g1034 (n1084, n1012);
buf  g1035 (n1050, n1007);
buf  g1036 (n1062, n980);
buf  g1037 (n1040, n1019);
not  g1038 (n1083, n995);
not  g1039 (n1066, n979);
buf  g1040 (n1052, n770);
buf  g1041 (n1033, n825);
xor  g1042 (n1078, n999, n973, n1009, n978);
and  g1043 (n1082, n756, n986, n758, n1022);
nor  g1044 (n1046, n1015, n976, n910, n1027);
xor  g1045 (n1049, n765, n756, n1017, n991);
or   g1046 (n1075, n968, n1003, n759, n760);
nand g1047 (n1094, n990, n989, n1000, n987);
xor  g1048 (n1055, n765, n763, n1004);
nand g1049 (n1072, n972, n827, n767, n906);
or   g1050 (n1035, n1029, n985, n969, n826);
or   g1051 (n1091, n767, n1030, n829, n768);
and  g1052 (n1044, n1021, n826, n829, n977);
nand g1053 (n1074, n1024, n1028, n1002, n909);
xnor g1054 (n1063, n1006, n770, n828, n825);
nand g1055 (n1059, n998, n762, n1023, n994);
xor  g1056 (n1092, n1018, n830, n1005, n827);
nand g1057 (n1089, n993, n996, n755, n981);
and  g1058 (n1087, n766, n769, n762);
and  g1059 (n1090, n761, n1025, n766, n828);
or   g1060 (n1073, n1008, n768, n760, n982);
nor  g1061 (n1088, n829, n992, n1013, n970);
not  g1062 (n1159, n1052);
not  g1063 (n1133, n1082);
buf  g1064 (n1191, n1090);
not  g1065 (n1342, n1046);
not  g1066 (n1151, n1039);
buf  g1067 (n1155, n1040);
not  g1068 (n1265, n1056);
buf  g1069 (n1317, n1075);
buf  g1070 (n1282, n1032);
buf  g1071 (n1242, n1093);
buf  g1072 (n1225, n1042);
not  g1073 (n1222, n1054);
buf  g1074 (n1332, n1035);
buf  g1075 (n1219, n1061);
buf  g1076 (n1289, n1044);
buf  g1077 (n1240, n1070);
not  g1078 (n1212, n1055);
buf  g1079 (n1156, n1034);
buf  g1080 (n1308, n1043);
not  g1081 (n1194, n1078);
not  g1082 (n1261, n1092);
buf  g1083 (n1182, n1065);
buf  g1084 (n1276, n1038);
not  g1085 (n1290, n1032);
buf  g1086 (n1127, n1038);
not  g1087 (n1295, n1089);
not  g1088 (n1142, n1061);
not  g1089 (n1246, n1091);
not  g1090 (n1239, n1087);
not  g1091 (n1196, n1043);
buf  g1092 (n1237, n1037);
not  g1093 (n1220, n1079);
not  g1094 (n1108, n1058);
not  g1095 (n1329, n1063);
buf  g1096 (n1326, n1031);
buf  g1097 (n1097, n1033);
buf  g1098 (n1341, n1043);
not  g1099 (n1331, n1069);
not  g1100 (n1128, n1076);
buf  g1101 (n1300, n1073);
not  g1102 (n1333, n1059);
not  g1103 (n1328, n1058);
buf  g1104 (n1105, n1094);
not  g1105 (n1173, n1064);
not  g1106 (n1218, n1040);
not  g1107 (n1186, n1081);
not  g1108 (n1302, n1077);
buf  g1109 (n1248, n1055);
not  g1110 (n1176, n1071);
not  g1111 (n1233, n1071);
not  g1112 (n1313, n1084);
buf  g1113 (n1161, n1093);
buf  g1114 (n1198, n1059);
not  g1115 (n1221, n1072);
buf  g1116 (n1320, n1056);
not  g1117 (n1287, n1068);
not  g1118 (n1310, n1050);
not  g1119 (n1203, n1045);
not  g1120 (n1213, n1082);
buf  g1121 (n1335, n1078);
buf  g1122 (n1103, n1052);
not  g1123 (n1149, n1042);
buf  g1124 (n1279, n1083);
buf  g1125 (n1228, n1059);
not  g1126 (n1192, n1082);
buf  g1127 (n1293, n1052);
not  g1128 (n1263, n1085);
not  g1129 (n1267, n1033);
buf  g1130 (n1119, n1085);
buf  g1131 (n1280, n1055);
not  g1132 (n1325, n1031);
buf  g1133 (n1136, n1035);
not  g1134 (n1181, n1049);
buf  g1135 (n1347, n1080);
buf  g1136 (n1299, n1085);
buf  g1137 (n1231, n1063);
not  g1138 (n1109, n1033);
not  g1139 (n1318, n1083);
buf  g1140 (n1346, n1092);
buf  g1141 (n1315, n1037);
buf  g1142 (n1134, n1046);
not  g1143 (n1122, n1060);
buf  g1144 (n1324, n1066);
buf  g1145 (n1146, n1053);
not  g1146 (n1141, n1041);
not  g1147 (n1338, n1048);
not  g1148 (n1202, n1057);
buf  g1149 (n1226, n1048);
not  g1150 (n1157, n1047);
buf  g1151 (n1185, n1068);
buf  g1152 (n1135, n1075);
not  g1153 (n1168, n1094);
not  g1154 (n1232, n1077);
not  g1155 (n1345, n1033);
not  g1156 (n1166, n1054);
not  g1157 (n1316, n1069);
not  g1158 (n1207, n1072);
not  g1159 (n1111, n1051);
buf  g1160 (n1211, n1092);
not  g1161 (n1188, n1064);
buf  g1162 (n1130, n1066);
not  g1163 (n1340, n1057);
not  g1164 (n1336, n1062);
not  g1165 (n1292, n1083);
buf  g1166 (n1165, n1080);
not  g1167 (n1264, n1088);
buf  g1168 (n1337, n1046);
buf  g1169 (n1210, n1046);
not  g1170 (n1247, n1091);
buf  g1171 (n1120, n1053);
not  g1172 (n1230, n1060);
buf  g1173 (n1095, n1076);
buf  g1174 (n1216, n1045);
not  g1175 (n1286, n1038);
not  g1176 (n1164, n1066);
not  g1177 (n1116, n1047);
not  g1178 (n1102, n1073);
not  g1179 (n1277, n1043);
not  g1180 (n1307, n1076);
buf  g1181 (n1137, n772);
not  g1182 (n1256, n1060);
not  g1183 (n1229, n1066);
not  g1184 (n1174, n1089);
not  g1185 (n1281, n1077);
not  g1186 (n1139, n1051);
buf  g1187 (n1348, n1078);
not  g1188 (n1140, n1058);
not  g1189 (n1170, n771);
not  g1190 (n1169, n1044);
buf  g1191 (n1209, n773);
buf  g1192 (n1180, n1090);
not  g1193 (n1143, n1062);
buf  g1194 (n1273, n1087);
not  g1195 (n1104, n1034);
not  g1196 (n1150, n1090);
not  g1197 (n1124, n1047);
buf  g1198 (n1309, n1091);
buf  g1199 (n1254, n1031);
not  g1200 (n1262, n1038);
not  g1201 (n1189, n773);
not  g1202 (n1350, n1070);
not  g1203 (n1339, n1067);
not  g1204 (n1271, n1058);
not  g1205 (n1251, n1049);
not  g1206 (n1301, n1075);
buf  g1207 (n1270, n1037);
buf  g1208 (n1100, n1051);
not  g1209 (n1125, n1067);
buf  g1210 (n1201, n1032);
not  g1211 (n1115, n1071);
not  g1212 (n1129, n1065);
buf  g1213 (n1330, n1072);
not  g1214 (n1311, n1088);
not  g1215 (n1208, n1067);
not  g1216 (n1183, n1086);
buf  g1217 (n1154, n1085);
buf  g1218 (n1096, n1065);
not  g1219 (n1344, n1049);
not  g1220 (n1145, n1048);
not  g1221 (n1117, n1082);
buf  g1222 (n1190, n1078);
not  g1223 (n1195, n1089);
not  g1224 (n1243, n1031);
not  g1225 (n1227, n1088);
not  g1226 (n1314, n1064);
buf  g1227 (n1234, n1086);
buf  g1228 (n1241, n1090);
buf  g1229 (n1312, n1041);
buf  g1230 (n1187, n1039);
buf  g1231 (n1238, n1091);
not  g1232 (n1178, n1079);
not  g1233 (n1193, n1055);
not  g1234 (n1250, n1084);
not  g1235 (n1235, n1056);
buf  g1236 (n1138, n1086);
buf  g1237 (n1275, n1070);
buf  g1238 (n1285, n1048);
not  g1239 (n1304, n1047);
buf  g1240 (n1306, n1087);
buf  g1241 (n1321, n1049);
not  g1242 (n1132, n1077);
not  g1243 (n1205, n1062);
buf  g1244 (n1147, n1079);
buf  g1245 (n1148, n1041);
not  g1246 (n1126, n1036);
not  g1247 (n1249, n1069);
buf  g1248 (n1131, n1044);
not  g1249 (n1305, n1041);
not  g1250 (n1172, n1074);
not  g1251 (n1274, n1054);
buf  g1252 (n1123, n1042);
not  g1253 (n1294, n1074);
not  g1254 (n1245, n1074);
buf  g1255 (n1199, n772);
not  g1256 (n1278, n1045);
buf  g1257 (n1303, n1040);
buf  g1258 (n1197, n1072);
not  g1259 (n1260, n1081);
buf  g1260 (n1291, n1042);
buf  g1261 (n1283, n1084);
not  g1262 (n1171, n1057);
buf  g1263 (n1252, n1032);
buf  g1264 (n1175, n1035);
not  g1265 (n1215, n1065);
buf  g1266 (n1284, n1064);
buf  g1267 (n1322, n1073);
buf  g1268 (n1223, n1057);
not  g1269 (n1114, n1040);
buf  g1270 (n1259, n1081);
buf  g1271 (n1244, n1053);
buf  g1272 (n1163, n1089);
buf  g1273 (n1152, n1039);
buf  g1274 (n1269, n1054);
not  g1275 (n1113, n1059);
not  g1276 (n1121, n1079);
not  g1277 (n1144, n1074);
buf  g1278 (n1217, n1087);
not  g1279 (n1153, n1050);
not  g1280 (n1343, n1063);
not  g1281 (n1204, n1053);
not  g1282 (n1258, n1037);
buf  g1283 (n1349, n1067);
not  g1284 (n1298, n1070);
not  g1285 (n1160, n1051);
not  g1286 (n1272, n1062);
not  g1287 (n1098, n1092);
not  g1288 (n1253, n1084);
buf  g1289 (n1323, n1036);
buf  g1290 (n1200, n1044);
buf  g1291 (n1099, n1039);
buf  g1292 (n1106, n1083);
buf  g1293 (n1334, n1061);
not  g1294 (n1112, n1050);
not  g1295 (n1297, n1036);
not  g1296 (n1319, n1045);
buf  g1297 (n1206, n1088);
not  g1298 (n1266, n1094);
not  g1299 (n1101, n1034);
not  g1300 (n1296, n1036);
buf  g1301 (n1327, n1069);
buf  g1302 (n1167, n1063);
not  g1303 (n1257, n1093);
buf  g1304 (n1236, n1073);
buf  g1305 (n1177, n1035);
not  g1306 (n1214, n1052);
buf  g1307 (n1118, n1061);
buf  g1308 (n1179, n1093);
not  g1309 (n1162, n1086);
not  g1310 (n1107, n1068);
not  g1311 (n1268, n1080);
buf  g1312 (n1255, n771);
buf  g1313 (n1288, n1050);
not  g1314 (n1110, n1080);
not  g1315 (n1158, n1075);
or   g1316 (n1224, n1068, n1094, n1060, n1034);
and  g1317 (n1184, n1076, n1056, n1071, n1081);
not  g1318 (n1364, n1141);
not  g1319 (n1396, n1161);
buf  g1320 (n1354, n1136);
not  g1321 (n1612, n1124);
buf  g1322 (n1504, n1130);
buf  g1323 (n1374, n1120);
buf  g1324 (n1419, n1113);
not  g1325 (n1573, n1150);
not  g1326 (n1484, n1115);
buf  g1327 (n1506, n1170);
buf  g1328 (n1556, n1102);
buf  g1329 (n1530, n1147);
buf  g1330 (n1498, n1146);
not  g1331 (n1388, n1098);
not  g1332 (n1561, n780);
buf  g1333 (n1464, n1118);
not  g1334 (n1439, n1102);
not  g1335 (n1480, n346);
not  g1336 (n1550, n1102);
buf  g1337 (n1647, n1114);
buf  g1338 (n1355, n1160);
buf  g1339 (n1602, n1131);
not  g1340 (n1361, n1108);
not  g1341 (n1427, n1161);
buf  g1342 (n1594, n1170);
buf  g1343 (n1524, n1144);
buf  g1344 (n1485, n1112);
not  g1345 (n1539, n1158);
buf  g1346 (n1406, n1111);
not  g1347 (n1589, n1095);
buf  g1348 (n1366, n617);
buf  g1349 (n1644, n1166);
not  g1350 (n1353, n1165);
buf  g1351 (n1554, n778);
buf  g1352 (n1389, n1139);
not  g1353 (n1508, n1109);
buf  g1354 (n1569, n1095);
not  g1355 (n1648, n1148);
buf  g1356 (n1462, n1125);
not  g1357 (n1395, n1114);
not  g1358 (n1566, n1145);
not  g1359 (n1571, n778);
not  g1360 (n1581, n1111);
buf  g1361 (n1629, n1169);
buf  g1362 (n1563, n953);
not  g1363 (n1449, n1162);
buf  g1364 (n1471, n781);
buf  g1365 (n1616, n1141);
not  g1366 (n1555, n1128);
buf  g1367 (n1436, n1107);
buf  g1368 (n1620, n1166);
not  g1369 (n1630, n775);
buf  g1370 (n1520, n1132);
not  g1371 (n1523, n1099);
not  g1372 (n1625, n956);
not  g1373 (n1450, n1162);
buf  g1374 (n1398, n1135);
not  g1375 (n1510, n160);
not  g1376 (n1577, n1103);
not  g1377 (n1372, n1152);
not  g1378 (n1392, n1139);
buf  g1379 (n1433, n1149);
not  g1380 (n1386, n1128);
not  g1381 (n1548, n892);
not  g1382 (n1601, n1147);
not  g1383 (n1591, n1098);
buf  g1384 (n1631, n1115);
not  g1385 (n1410, n1121);
buf  g1386 (n1380, n952);
not  g1387 (n1624, n1103);
not  g1388 (n1603, n1156);
not  g1389 (n1460, n1097);
not  g1390 (n1444, n1157);
not  g1391 (n1515, n1142);
not  g1392 (n1635, n1127);
buf  g1393 (n1422, n1142);
buf  g1394 (n1512, n1153);
buf  g1395 (n1509, n346);
buf  g1396 (n1617, n1111);
not  g1397 (n1399, n1167);
not  g1398 (n1584, n1105);
buf  g1399 (n1579, n830);
not  g1400 (n1356, n1134);
not  g1401 (n1409, n1144);
buf  g1402 (n1588, n1101);
not  g1403 (n1543, n1116);
not  g1404 (n1496, n1129);
buf  g1405 (n1455, n1119);
buf  g1406 (n1442, n1106);
not  g1407 (n1487, n779);
not  g1408 (n1475, n1146);
buf  g1409 (n1611, n1126);
not  g1410 (n1465, n1100);
buf  g1411 (n1572, n1096);
not  g1412 (n1453, n1130);
buf  g1413 (n1382, n1152);
buf  g1414 (n1413, n1134);
not  g1415 (n1549, n957);
buf  g1416 (n1521, n1145);
buf  g1417 (n1459, n1124);
buf  g1418 (n1478, n1114);
buf  g1419 (n1593, n1133);
buf  g1420 (n1514, n1110);
not  g1421 (n1637, n774);
not  g1422 (n1638, n1155);
buf  g1423 (n1477, n1122);
buf  g1424 (n1619, n1171);
not  g1425 (n1608, n1099);
buf  g1426 (n1476, n1138);
not  g1427 (n1610, n1169);
not  g1428 (n1446, n1153);
not  g1429 (n1456, n1096);
buf  g1430 (n1488, n780);
buf  g1431 (n1605, n1118);
buf  g1432 (n1431, n1122);
buf  g1433 (n1373, n954);
not  g1434 (n1614, n1159);
not  g1435 (n1551, n1112);
buf  g1436 (n1536, n1109);
buf  g1437 (n1621, n953);
not  g1438 (n1385, n1109);
not  g1439 (n1502, n1158);
not  g1440 (n1447, n1136);
not  g1441 (n1408, n1119);
not  g1442 (n1639, n1154);
not  g1443 (n1371, n1095);
buf  g1444 (n1495, n1152);
not  g1445 (n1578, n1134);
buf  g1446 (n1636, n1166);
buf  g1447 (n1559, n1123);
not  g1448 (n1404, n1137);
not  g1449 (n1434, n831);
buf  g1450 (n1576, n1143);
not  g1451 (n1424, n1134);
not  g1452 (n1586, n1109);
not  g1453 (n1393, n1141);
buf  g1454 (n1599, n1135);
buf  g1455 (n1640, n1124);
buf  g1456 (n1469, n1149);
not  g1457 (n1390, n956);
buf  g1458 (n1547, n1129);
not  g1459 (n1405, n1116);
not  g1460 (n1360, n1151);
buf  g1461 (n1545, n615);
not  g1462 (n1500, n1120);
not  g1463 (n1486, n1126);
buf  g1464 (n1416, n1128);
not  g1465 (n1527, n1147);
not  g1466 (n1560, n1133);
buf  g1467 (n1468, n1107);
buf  g1468 (n1583, n1107);
buf  g1469 (n1622, n1138);
buf  g1470 (n1582, n1150);
buf  g1471 (n1600, n1143);
not  g1472 (n1466, n1097);
not  g1473 (n1497, n1161);
not  g1474 (n1597, n1123);
buf  g1475 (n1632, n1115);
not  g1476 (n1362, n1112);
not  g1477 (n1457, n830);
not  g1478 (n1649, n1152);
not  g1479 (n1526, n955);
buf  g1480 (n1452, n1106);
not  g1481 (n1542, n831);
not  g1482 (n1378, n1099);
not  g1483 (n1580, n951);
buf  g1484 (n1558, n1097);
buf  g1485 (n1428, n775);
not  g1486 (n1618, n892);
buf  g1487 (n1592, n1117);
buf  g1488 (n1623, n831);
buf  g1489 (n1463, n1167);
buf  g1490 (n1546, n1115);
buf  g1491 (n1585, n1104);
not  g1492 (n1552, n1124);
buf  g1493 (n1414, n1164);
not  g1494 (n1626, n952);
buf  g1495 (n1567, n1140);
not  g1496 (n1606, n1116);
buf  g1497 (n1633, n1139);
not  g1498 (n1493, n1153);
not  g1499 (n1651, n1117);
not  g1500 (n1489, n1125);
not  g1501 (n1383, n1129);
not  g1502 (n1642, n1159);
buf  g1503 (n1634, n779);
not  g1504 (n1517, n1169);
buf  g1505 (n1426, n1100);
buf  g1506 (n1369, n1105);
not  g1507 (n1575, n1122);
buf  g1508 (n1375, n1143);
not  g1509 (n1490, n1149);
not  g1510 (n1458, n1113);
buf  g1511 (n1531, n1126);
buf  g1512 (n1607, n1120);
not  g1513 (n1430, n831);
buf  g1514 (n1363, n1138);
not  g1515 (n1604, n1137);
buf  g1516 (n1441, n912);
not  g1517 (n1370, n1106);
not  g1518 (n1401, n1098);
buf  g1519 (n1454, n1104);
buf  g1520 (n1381, n1169);
buf  g1521 (n1533, n1118);
buf  g1522 (n1544, n1153);
not  g1523 (n1568, n1127);
not  g1524 (n1535, n1095);
not  g1525 (n1359, n1157);
buf  g1526 (n1519, n1143);
not  g1527 (n1423, n1114);
not  g1528 (n1513, n776);
not  g1529 (n1445, n776);
buf  g1530 (n1596, n1163);
not  g1531 (n1472, n1110);
buf  g1532 (n1397, n1103);
not  g1533 (n1411, n1146);
not  g1534 (n1451, n1096);
buf  g1535 (n1562, n1140);
not  g1536 (n1412, n1160);
buf  g1537 (n1609, n1107);
buf  g1538 (n1570, n1163);
not  g1539 (n1420, n1130);
not  g1540 (n1473, n1167);
buf  g1541 (n1587, n1139);
not  g1542 (n1627, n1121);
not  g1543 (n1357, n1113);
buf  g1544 (n1507, n1145);
not  g1545 (n1650, n1106);
buf  g1546 (n1491, n1168);
buf  g1547 (n1481, n1142);
buf  g1548 (n1499, n1155);
not  g1549 (n1503, n1161);
buf  g1550 (n1553, n1164);
not  g1551 (n1516, n1148);
not  g1552 (n1641, n1150);
not  g1553 (n1501, n1160);
buf  g1554 (n1407, n1170);
buf  g1555 (n1628, n1159);
buf  g1556 (n1438, n1151);
not  g1557 (n1479, n957);
buf  g1558 (n1421, n1151);
buf  g1559 (n1432, n955);
buf  g1560 (n1541, n1168);
not  g1561 (n1402, n1164);
buf  g1562 (n1394, n953);
not  g1563 (n1425, n1096);
buf  g1564 (n1352, n1150);
buf  g1565 (n1525, n1110);
not  g1566 (n1522, n1119);
not  g1567 (n1391, n1140);
not  g1568 (n1595, n1102);
buf  g1569 (n1467, n1156);
not  g1570 (n1415, n1108);
not  g1571 (n1376, n1101);
not  g1572 (n1492, n951);
buf  g1573 (n1400, n614);
buf  g1574 (n1351, n1101);
buf  g1575 (n1435, n1126);
not  g1576 (n1537, n1117);
not  g1577 (n1557, n1125);
not  g1578 (n1574, n957);
buf  g1579 (n1528, n777);
buf  g1580 (n1448, n1171);
buf  g1581 (n1494, n1112);
buf  g1582 (n1565, n1113);
buf  g1583 (n1532, n1132);
not  g1584 (n1598, n1154);
not  g1585 (n1368, n1123);
not  g1586 (n1482, n1119);
not  g1587 (n1538, n777);
buf  g1588 (n1646, n954);
buf  g1589 (n1615, n1117);
not  g1590 (n1518, n1155);
not  g1591 (n1417, n1111);
not  g1592 (n1358, n1157);
buf  g1593 (n1483, n951);
not  g1594 (n1429, n1118);
not  g1595 (n1377, n1105);
not  g1596 (n1403, n1158);
buf  g1597 (n1474, n781);
and  g1598 (n1387, n1159, n1146, n1141, n1156);
xor  g1599 (n1564, n1167, n1137, n774, n1136);
nand g1600 (n1365, n1144, n1142, n1132, n1136);
or   g1601 (n1461, n1147, n1156, n1154, n1101);
xnor g1602 (n1645, n1149, n1105, n1168, n1125);
nand g1603 (n1384, n830, n1138, n1104);
nor  g1604 (n1440, n1165, n1144, n1155, n1170);
nor  g1605 (n1529, n160, n1110, n1120, n616);
and  g1606 (n1418, n1158, n1133, n952, n160);
and  g1607 (n1643, n1166, n1151, n1145, n892);
nand g1608 (n1443, n1129, n1133, n1116, n1098);
xor  g1609 (n1470, n1121, n1165, n1099, n1127);
or   g1610 (n1379, n1122, n1100, n1128, n1160);
nand g1611 (n1590, n1154, n1137, n1127, n1097);
nand g1612 (n1367, n1108, n1135, n1164, n1148);
or   g1613 (n1540, n1163, n954, n1131, n1108);
and  g1614 (n1613, n1123, n1162, n1100);
xnor g1615 (n1511, n1130, n1168, n955, n1131);
or   g1616 (n1534, n892, n1135, n1132, n1148);
or   g1617 (n1437, n1103, n1131, n1163, n1140);
or   g1618 (n1505, n1121, n956, n1157, n1165);
or   g1619 (n1713, n1627, n1176);
xor  g1620 (n1834, n1253, n1295);
xnor g1621 (n1889, n1367, n1288);
xor  g1622 (n1811, n1625, n1631);
nand g1623 (n1692, n1271, n1293);
xnor g1624 (n1867, n1191, n1382, n1206, n1230);
or   g1625 (n1727, n1181, n1270, n1391, n1298);
xnor g1626 (n1810, n1257, n1502, n1493, n1411);
nand g1627 (n1804, n1468, n1338, n1210, n1319);
nand g1628 (n1896, n1218, n1465, n1268, n1301);
xor  g1629 (n1933, n1360, n1430, n1262, n1288);
or   g1630 (n1908, n1602, n1451, n1224, n1646);
nand g1631 (n1919, n1222, n1533, n1318, n1254);
xnor g1632 (n1738, n1315, n1459, n1252, n1225);
and  g1633 (n1931, n1347, n1349, n1199, n1598);
or   g1634 (n1895, n1205, n1179, n1245, n1256);
nor  g1635 (n1735, n1259, n1422, n1549, n1236);
and  g1636 (n1687, n1223, n1348, n1618, n1631);
nor  g1637 (n1877, n1575, n1364, n1570, n1198);
nand g1638 (n1654, n1535, n1487, n1264, n1247);
xnor g1639 (n1802, n1175, n1629, n1610, n1222);
nand g1640 (n1677, n1241, n1246, n1392, n1435);
xnor g1641 (n1803, n1607, n1331, n1208, n1268);
or   g1642 (n1756, n1340, n1621, n1179, n1221);
or   g1643 (n1824, n1322, n1196, n1265, n1243);
or   g1644 (n1830, n1240, n1599, n1538, n1302);
xor  g1645 (n1904, n1269, n1286, n1339, n1501);
and  g1646 (n1717, n1174, n1643, n1226, n1349);
and  g1647 (n1697, n1284, n1321, n1238, n1455);
or   g1648 (n1890, n1280, n1304, n1426, n1516);
or   g1649 (n1920, n1563, n1243, n1526, n1447);
or   g1650 (n1917, n1190, n1283, n1212, n1220);
nand g1651 (n1840, n1186, n1216, n1200, n1287);
xor  g1652 (n1750, n1587, n1618, n1349, n1201);
xnor g1653 (n1854, n1223, n1216, n1233, n1291);
or   g1654 (n1884, n1542, n1202, n1309, n1299);
nand g1655 (n1859, n1325, n1542, n1581, n1571);
and  g1656 (n1792, n1284, n1587, n1252, n1576);
or   g1657 (n1669, n1197, n1579, n1286, n1211);
xor  g1658 (n1716, n1292, n1244, n1424, n1180);
and  g1659 (n1746, n1554, n1449, n1358, n1472);
and  g1660 (n1674, n1547, n1417, n1176, n1216);
nand g1661 (n1764, n1420, n1198, n1208, n1621);
or   g1662 (n1790, n1644, n1228, n1195, n1186);
nor  g1663 (n1652, n1205, n1540, n1597, n1337);
or   g1664 (n1894, n1323, n1215, n1399, n1303);
or   g1665 (n1762, n1185, n1578, n1627, n1194);
nor  g1666 (n1852, n1346, n1637, n1340, n1603);
or   g1667 (n1843, n1187, n1567, n1223, n1552);
xor  g1668 (n1748, n1329, n1240, n1540, n1312);
xor  g1669 (n1733, n1456, n1172, n1419, n1193);
nor  g1670 (n1671, n1546, n1461, n1616, n1593);
xnor g1671 (n1696, n1274, n1580, n1638, n1334);
xor  g1672 (n1845, n1291, n1494, n1277, n1350);
and  g1673 (n1729, n1479, n1406, n1269, n1612);
and  g1674 (n1875, n1189, n1341, n1371, n1323);
xor  g1675 (n1722, n1234, n1286, n1275, n1529);
nand g1676 (n1685, n1250, n1278, n1336, n1171);
nand g1677 (n1797, n1513, n1553, n1259, n1243);
nor  g1678 (n1848, n1197, n1244, n1189, n1332);
xor  g1679 (n1666, n1236, n1244, n1217, n1546);
xor  g1680 (n1712, n1298, n1605, n1445, n1242);
nand g1681 (n1778, n1248, n1569, n1317, n1288);
and  g1682 (n1771, n1277, n1550, n1649, n1283);
nand g1683 (n1751, n1650, n1336, n1267, n1186);
nand g1684 (n1715, n1192, n1335, n1207, n1251);
xor  g1685 (n1846, n1279, n1324, n1243, n1647);
xor  g1686 (n1780, n1213, n1639, n1568, n1188);
nor  g1687 (n1873, n1385, n1577, n1551, n1314);
or   g1688 (n1839, n1281, n1262, n1195, n1218);
xnor g1689 (n1885, n1555, n1208, n1440, n1596);
nand g1690 (n1740, n1266, n1238, n1172, n1633);
and  g1691 (n1849, n1598, n1390, n1608, n1318);
xnor g1692 (n1863, n1315, n1327, n1640, n1184);
or   g1693 (n1928, n1294, n1590, n1272, n1350);
xor  g1694 (n1711, n1594, n1299, n1312, n1211);
nor  g1695 (n1822, n1297, n1444, n1527, n1254);
nand g1696 (n1864, n1251, n1230, n1550, n1192);
nand g1697 (n1660, n1345, n1326, n1321, n1193);
xor  g1698 (n1903, n1596, n1376, n1290, n1626);
or   g1699 (n1847, n1384, n1204, n1221, n1295);
or   g1700 (n1878, n1226, n1477, n1267, n1316);
and  g1701 (n1888, n1344, n1614, n1443, n1327);
xor  g1702 (n1892, n1231, n1327, n1250, n1308);
or   g1703 (n1857, n1279, n1271, n1562, n1346);
xnor g1704 (n1865, n1612, n1434, n1256, n1309);
nand g1705 (n1719, n1316, n1475, n1600, n1223);
nand g1706 (n1680, n1191, n1531, n1270, n1374);
nor  g1707 (n1815, n1273, n1244, n1327, n1340);
and  g1708 (n1708, n1232, n1474, n1320, n1263);
nor  g1709 (n1765, n1261, n1204, n1218, n1642);
xor  g1710 (n1667, n1259, n1563, n1219, n1568);
nor  g1711 (n1682, n1348, n1330, n1416, n1202);
xnor g1712 (n1714, n1350, n1308, n1270, n1423);
nand g1713 (n1786, n1274, n1305, n1566, n1574);
nor  g1714 (n1883, n1203, n1383, n1496, n1249);
xor  g1715 (n1731, n1481, n1213, n1573, n1337);
or   g1716 (n1862, n1307, n1395, n1324, n1293);
nand g1717 (n1791, n1614, n1208, n1242, n1448);
xnor g1718 (n1684, n1258, n1336, n1279);
nand g1719 (n1755, n1381, n1316, n1620, n1184);
and  g1720 (n1800, n1324, n1201, n1256, n1304);
and  g1721 (n1930, n1281, n1649, n1225, n1490);
xor  g1722 (n1835, n1190, n1300, n1272, n1641);
nor  g1723 (n1679, n1585, n1397, n1173, n1204);
or   g1724 (n1906, n1495, n1403, n1373, n1177);
nand g1725 (n1709, n1595, n1549, n1305, n1319);
nor  g1726 (n1912, n1182, n1646, n1305, n1272);
xnor g1727 (n1837, n1273, n1184, n1354, n1398);
and  g1728 (n1747, n1560, n1233, n1275, n1438);
and  g1729 (n1730, n1175, n1615, n1588, n1604);
nor  g1730 (n1785, n1431, n1293, n1264, n1269);
xor  g1731 (n1703, n1258, n1331, n1302, n1328);
nand g1732 (n1720, n1582, n1262, n1242, n1349);
nand g1733 (n1818, n1339, n1561, n1484, n1464);
nor  g1734 (n1869, n1321, n1263, n1343, n1375);
nand g1735 (n1916, n1193, n1648, n1285, n1278);
nand g1736 (n1825, n1589, n1310, n1368, n1630);
xor  g1737 (n1882, n1571, n1184, n1418, n1644);
xor  g1738 (n1900, n1210, n1269, n1557, n1548);
xor  g1739 (n1808, n1648, n1203, n1266, n1335);
nor  g1740 (n1773, n1207, n1307, n1603, n1215);
or   g1741 (n1768, n1638, n1251, n1510, n1558);
and  g1742 (n1793, n1466, n1282, n1637, n1225);
and  g1743 (n1898, n1341, n1362, n1264, n1179);
and  g1744 (n1718, n1345, n1452, n1237, n1255);
and  g1745 (n1861, n1228, n1304, n1326, n1314);
nand g1746 (n1876, n1592, n1252, n1273, n1209);
and  g1747 (n1723, n1213, n1635, n1338, n1551);
nor  g1748 (n1787, n1567, n1640, n1219, n1522);
or   g1749 (n1705, n1559, n1387, n1181, n1604);
xnor g1750 (n1925, n1343, n1232, n1306, n1497);
xnor g1751 (n1910, n1583, n1185, n1203, n1409);
xor  g1752 (n1659, n1572, n1485, n1258, n1247);
xnor g1753 (n1907, n1289, n1199, n1508, n1365);
nand g1754 (n1820, n1293, n1601, n1191, n1338);
or   g1755 (n1686, n1177, n1189, n1498, n1295);
xor  g1756 (n1655, n1183, n1471, n1347, n1322);
and  g1757 (n1743, n1565, n1235, n1492, n1347);
or   g1758 (n1668, n1334, n1476, n1308, n1339);
nand g1759 (n1741, n1237, n1330, n1311, n1187);
or   g1760 (n1770, n1228, n1297, n1341, n1266);
xnor g1761 (n1656, n1400, n1217, n1333, n1436);
nor  g1762 (n1812, n1279, n1276, n1318, n1410);
or   g1763 (n1763, n1249, n1317, n1286, n1222);
and  g1764 (n1827, n1333, n1335, n1172, n1599);
nor  g1765 (n1689, n1199, n1623, n1363, n1389);
or   g1766 (n1658, n1331, n1408, n1200, n1544);
nor  g1767 (n1798, n1194, n1241, n1582, n1313);
xnor g1768 (n1683, n1482, n1624, n1275, n1346);
or   g1769 (n1886, n1241, n1266, n1180, n1556);
nor  g1770 (n1922, n1632, n1307, n1246, n1296);
nor  g1771 (n1758, n1523, n1317, n1331, n1290);
xnor g1772 (n1657, n1359, n1181, n1229, n1205);
nor  g1773 (n1879, n1611, n1287, n1235, n1366);
xor  g1774 (n1901, n1232, n1314, n1521, n1317);
nor  g1775 (n1871, n1532, n1350, n1272, n1217);
and  g1776 (n1672, n1344, n1217, n1234, n1320);
nor  g1777 (n1844, n1348, n1173, n1589, n1342);
and  g1778 (n1831, n1287, n1200, n1203, n1558);
nor  g1779 (n1914, n1229, n1388, n1597, n1301);
xor  g1780 (n1734, n1310, n1326, n1281, n1210);
nand g1781 (n1935, n1469, n1480, n1488, n1261);
nor  g1782 (n1742, n1348, n1285, n1559, n1183);
nor  g1783 (n1860, n1230, n1178, n1507, n1292);
or   g1784 (n1784, n1536, n1248, n1219, n1294);
xor  g1785 (n1782, n1214, n1277, n1564, n1478);
nor  g1786 (n1868, n1220, n1378, n1177, n1641);
nor  g1787 (n1813, n1594, n1188, n1216, n1517);
nor  g1788 (n1921, n1226, n1427, n1187, n1602);
and  g1789 (n1927, n1341, n1302, n1609, n1323);
or   g1790 (n1829, n1311, n1425, n1306, n1209);
or   g1791 (n1700, n1324, n1463, n1591, n1296);
xor  g1792 (n1691, n1231, n1547, n1428, n1180);
and  g1793 (n1681, n1450, n1271, n1414, n1247);
or   g1794 (n1752, n1514, n1569, n1626, n1625);
nor  g1795 (n1833, n1633, n1229, n1233, n1239);
xnor g1796 (n1779, n1642, n1322, n1467, n1185);
or   g1797 (n1745, n1259, n1290, n1257, n1305);
nor  g1798 (n1766, n1647, n1178, n1212, n1191);
xnor g1799 (n1856, n1607, n1619, n1329, n1309);
and  g1800 (n1832, n1292, n1613, n1310, n1294);
xor  g1801 (n1805, n1611, n1296, n1544, n1421);
nand g1802 (n1781, n1282, n1628, n1296, n1268);
or   g1803 (n1725, n1289, n1302, n1572, n1337);
xor  g1804 (n1902, n1263, n1325, n1393, n1312);
and  g1805 (n1721, n1189, n1174, n1240, n1630);
and  g1806 (n1788, n1528, n1209, n1271, n1330);
or   g1807 (n1934, n1173, n1511, n1340, n1457);
xor  g1808 (n1851, n1345, n1210, n1462, n1316);
nand g1809 (n1688, n1181, n1273, n1323, n1311);
and  g1810 (n1929, n1636, n1377, n1584, n1174);
xor  g1811 (n1694, n1545, n1192, n1294, n1329);
and  g1812 (n1704, n1446, n1261, n1247, n1215);
and  g1813 (n1838, n1303, n1556, n1206, n1442);
xnor g1814 (n1905, n1239, n1407, n1255, n1454);
xnor g1815 (n1662, n1283, n1277, n1352, n1193);
or   g1816 (n1663, n1206, n1634, n1519, n1175);
and  g1817 (n1855, n1298, n1342, n1228, n1226);
and  g1818 (n1707, n1332, n1282, n1328, n1234);
nand g1819 (n1913, n1285, n1543, n1227, n1574);
or   g1820 (n1665, n1288, n1345, n1315, n1576);
or   g1821 (n1932, n1192, n1586, n1332, n1608);
nand g1822 (n1728, n1473, n1562, n1251, n1301);
xnor g1823 (n1874, n1224, n1617, n1307, n1212);
xnor g1824 (n1673, n1372, n1312, n1541, n1622);
nand g1825 (n1821, n1301, n1380, n1588, n1254);
nor  g1826 (n1783, n1263, n1636, n1617, n1579);
and  g1827 (n1816, n1541, n1214, n1554, n1275);
xor  g1828 (n1866, n1174, n1276, n1248, n1214);
nor  g1829 (n1695, n1319, n1289, n1237, n1429);
and  g1830 (n1795, n1278, n1353, n1202, n1267);
nand g1831 (n1767, n1321, n1236, n1235, n1592);
xor  g1832 (n1858, n1234, n1342, n1356, n1183);
and  g1833 (n1776, n1308, n1245, n1261, n1609);
or   g1834 (n1826, n1314, n1176, n1242, n1441);
nor  g1835 (n1853, n1322, n1270, n1333, n1291);
nor  g1836 (n1698, n1326, n1555, n1188, n1186);
xnor g1837 (n1870, n1415, n1282, n1343, n1591);
and  g1838 (n1749, n1311, n1204, n1328, n1402);
xnor g1839 (n1807, n1530, n1586, n1584, n1320);
xor  g1840 (n1926, n1183, n1396, n1284, n1583);
nor  g1841 (n1724, n1566, n1218, n1267, n1553);
and  g1842 (n1678, n1632, n1460, n1255, n1347);
and  g1843 (n1923, n1231, n1194, n1458, n1483);
or   g1844 (n1732, n1197, n1287, n1285, n1280);
nor  g1845 (n1911, n1334, n1361, n1173, n1209);
and  g1846 (n1760, n1178, n1564, n1334, n1593);
xnor g1847 (n1675, n1211, n1239, n1254, n1175);
xor  g1848 (n1676, n1578, n1299, n1229, n1620);
xor  g1849 (n1769, n1306, n1539, n1297, n1240);
and  g1850 (n1872, n1249, n1236, n1338, n1300);
nand g1851 (n1841, n1265, n1643, n1355, n1320);
or   g1852 (n1737, n1503, n1188, n1238, n1537);
nor  g1853 (n1836, n1245, n1344, n1227, n1525);
and  g1854 (n1772, n1211, n1573, n1585, n1187);
nand g1855 (n1744, n1257, n1199, n1258, n1313);
nor  g1856 (n1909, n1190, n1299, n1575, n1265);
xor  g1857 (n1789, n1303, n1198, n1520, n1628);
or   g1858 (n1736, n1278, n1605, n1329, n1212);
xnor g1859 (n1842, n1198, n1412, n1600, n1645);
and  g1860 (n1661, n1227, n1518, n1225, n1500);
and  g1861 (n1881, n1274, n1313, n1509, n1610);
nor  g1862 (n1775, n1201, n1230, n1196, n1231);
or   g1863 (n1828, n1232, n1241, n1202, n1570);
and  g1864 (n1774, n1245, n1595, n1257, n1601);
or   g1865 (n1806, n1280, n1437, n1577, n1224);
or   g1866 (n1936, n1539, n1176, n1504, n1246);
and  g1867 (n1761, n1512, n1250, n1506, n1260);
xor  g1868 (n1701, n1171, n1295, n1239, n1623);
nor  g1869 (n1915, n1561, n1253, n1335, n1246);
nor  g1870 (n1702, n1224, n1557, n1179, n1325);
or   g1871 (n1880, n1180, n1276, n1260, n1250);
nor  g1872 (n1817, n1178, n1325, n1433, n1639);
nor  g1873 (n1693, n1580, n1337, n1306, n1260);
nor  g1874 (n1670, n1268, n1543, n1291, n1284);
and  g1875 (n1850, n1214, n1297, n1303, n1545);
xor  g1876 (n1819, n1613, n1206, n1255, n1221);
and  g1877 (n1706, n1194, n1343, n1252, n1264);
xnor g1878 (n1897, n1524, n1262, n1439, n1565);
or   g1879 (n1653, n1195, n1237, n1344, n1339);
xor  g1880 (n1664, n1207, n1342, n1309, n1394);
or   g1881 (n1814, n1629, n1196, n1197, n1499);
nand g1882 (n1893, n1298, n1182, n1470, n1190);
nand g1883 (n1726, n1238, n1634, n1207, n1172);
and  g1884 (n1809, n1379, n1606, n1233, n1276);
xnor g1885 (n1891, n1635, n1369, n1205, n1215);
xor  g1886 (n1823, n1235, n1219, n1315, n1292);
or   g1887 (n1924, n1248, n1453, n1328, n1182);
or   g1888 (n1699, n1290, n1220, n1357, n1274);
and  g1889 (n1799, n1489, n1622, n1249, n1201);
and  g1890 (n1794, n1505, n1318, n1491, n1624);
xnor g1891 (n1899, n1280, n1289, n1581, n1300);
nand g1892 (n1757, n1548, n1222, n1386, n1606);
nor  g1893 (n1759, n1413, n1552, n1330, n1283);
and  g1894 (n1777, n1220, n1310, n1370, n1650);
xnor g1895 (n1754, n1332, n1560, n1195, n1304);
or   g1896 (n1753, n1182, n1486, n1227, n1196);
xor  g1897 (n1796, n1313, n1534, n1432, n1200);
or   g1898 (n1710, n1319, n1256, n1615, n1619);
nor  g1899 (n1739, n1300, n1281, n1405, n1590);
nand g1900 (n1887, n1213, n1221, n1253);
and  g1901 (n1801, n1333, n1265, n1346, n1401);
xnor g1902 (n1918, n1351, n1185, n1616, n1515);
xnor g1903 (n1690, n1177, n1404, n1260, n1645);
xor  g1904 (n1964, n1733, n1767, n1745, n1699);
xnor g1905 (n1968, n1654, n1709, n1764, n1723);
and  g1906 (n1966, n1737, n1781, n1683, n1710);
and  g1907 (n1942, n1729, n1681, n1760, n1782);
nor  g1908 (n1953, n1720, n1742, n1675, n1778);
xnor g1909 (n1944, n1722, n1713, n1670, n1653);
nand g1910 (n1957, n1665, n1652, n1669, n1712);
or   g1911 (n1946, n1695, n1735, n1739, n1765);
xor  g1912 (n1940, n1685, n1711, n1730, n1783);
xnor g1913 (n1938, n1751, n1750, n1721, n1775);
nand g1914 (n1962, n1757, n1756, n1655, n1771);
or   g1915 (n1937, n1668, n1719, n1731, n1659);
or   g1916 (n1941, n1700, n1740, n1662, n1776);
xor  g1917 (n1963, n1738, n1785, n1706, n1688);
xnor g1918 (n1952, n1703, n1770, n1747, n1746);
or   g1919 (n1956, n1741, n1761, n1656, n1680);
or   g1920 (n1961, n1671, n1718, n1690, n1724);
nor  g1921 (n1950, n1697, n1743, n1715, n1777);
and  g1922 (n1943, n1678, n1784, n1780, n1657);
or   g1923 (n1949, n1734, n1772, n1755, n1663);
nor  g1924 (n1959, n1661, n1726, n1707, n1768);
nand g1925 (n1970, n1701, n1677, n1727, n1651);
xor  g1926 (n1955, n1679, n1673, n1774, n1704);
xor  g1927 (n1969, n1779, n1666, n1694, n1664);
and  g1928 (n1958, n1773, n1651, n1660, n1732);
nand g1929 (n1951, n1762, n1754, n1748, n1687);
xnor g1930 (n1954, n1708, n1672, n1716, n1702);
or   g1931 (n1948, n1692, n1684, n1758, n1693);
nand g1932 (n1960, n1698, n1689, n1725, n1686);
or   g1933 (n1965, n1763, n1691, n1696, n1759);
or   g1934 (n1939, n1717, n1752, n1769, n1766);
xor  g1935 (n1945, n1753, n1658, n1705, n1676);
nand g1936 (n1947, n1714, n1744, n1667, n1682);
nor  g1937 (n1967, n1728, n1736, n1749, n1674);
xnor g1938 (n1996, n1852, n1835, n1955, n1957);
or   g1939 (n1985, n1942, n1854, n1954, n1822);
or   g1940 (n2003, n1941, n1867, n1958, n1952);
nand g1941 (n1991, n1799, n1792, n1877, n1851);
xor  g1942 (n1993, n1949, n1808, n1811, n1848);
or   g1943 (n1982, n1853, n1857, n1875, n1850);
xor  g1944 (n1987, n1815, n1810, n1796, n1879);
xnor g1945 (n2002, n1951, n1790, n1863, n1964);
nor  g1946 (n1981, n1832, n1880, n1940, n1946);
nand g1947 (n1983, n1819, n1787, n1884, n1836);
and  g1948 (n1995, n1807, n1806, n1801, n1814);
and  g1949 (n1992, n1948, n1834, n1859, n1849);
xnor g1950 (n1976, n1829, n1959, n1786, n1858);
nand g1951 (n1998, n1825, n1864, n1874, n1789);
nand g1952 (n1988, n1800, n1883, n1813, n1860);
and  g1953 (n1979, n1969, n1960, n1947, n1847);
nor  g1954 (n1971, n1966, n1837, n1950, n1818);
xor  g1955 (n1984, n1841, n1826, n1868, n1838);
nor  g1956 (n2000, n1961, n1816, n1823, n1827);
xor  g1957 (n1990, n1794, n1791, n1965, n1809);
nand g1958 (n1980, n1881, n1956, n1812, n1803);
or   g1959 (n1975, n1871, n1817, n1830, n1970);
nor  g1960 (n1973, n1831, n1967, n1802, n1963);
xnor g1961 (n1974, n1804, n1872, n1788, n1828);
xor  g1962 (n1994, n1855, n1845, n1962, n1844);
xor  g1963 (n2001, n1882, n1842, n1856, n1938);
nand g1964 (n1972, n1870, n1878, n1833, n1839);
xnor g1965 (n1989, n1861, n1869, n1876, n1873);
xnor g1966 (n1986, n1866, n1805, n1824, n1843);
and  g1967 (n1997, n1795, n1953, n1865, n1846);
nand g1968 (n1978, n1793, n1820, n1840, n1821);
nand g1969 (n1977, n1943, n1798, n1944, n1862);
or   g1970 (n1999, n1968, n1945, n1797, n1939);
nand g1971 (n2008, n1975, n1901, n1924, n1909);
xnor g1972 (n2010, n1918, n1903, n1934, n1893);
or   g1973 (n2014, n1887, n1917, n1907, n1888);
nand g1974 (n2004, n1892, n1915, n1910, n1889);
or   g1975 (n2021, n1902, n1891, n1971, n1912);
and  g1976 (n2020, n1894, n618, n1983, n1990);
xor  g1977 (n2018, n1988, n1906, n1992, n1899);
and  g1978 (n2016, n1980, n1987, n1885, n1935);
xnor g1979 (n2006, n1977, n1925, n1900, n1922);
xnor g1980 (n2005, n1886, n1931, n1897, n1981);
xor  g1981 (n2013, n1929, n1890, n1979, n1923);
nor  g1982 (n2022, n1927, n1898, n1986, n1933);
or   g1983 (n2009, n1913, n1908, n1905, n1982);
nor  g1984 (n2019, n1991, n1973, n1930, n1920);
nor  g1985 (n2015, n1921, n1984, n1926, n1896);
and  g1986 (n2011, n1972, n1928, n1914, n1989);
nand g1987 (n2017, n1936, n1895, n1976, n1916);
nor  g1988 (n2012, n1985, n619, n1978, n1919);
xor  g1989 (n2007, n1911, n1932, n1904, n1974);
nand g1990 (n2028, n2002, n2015, n2003, n1997);
nor  g1991 (n2027, n1994, n1998, n2001, n2014);
nor  g1992 (n2030, n2022, n1995, n2004, n1993);
nand g1993 (n2023, n2013, n2012, n2008, n2020);
nor  g1994 (n2029, n2000, n2006, n2017, n2011);
and  g1995 (n2025, n2021, n2019, n2003, n2010);
nor  g1996 (n2024, n160, n2007, n1996, n2016);
xnor g1997 (n2026, n2009, n2005, n1999, n2018);
or   g1998 (n2032, n2025, n2026, n2023, n2029);
nor  g1999 (n2031, n2027, n2030, n2024, n2028);
endmodule
