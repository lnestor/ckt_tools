// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_325 written by SynthGen on 2021/04/05 11:24:15
module Stat_3000_325( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n2378, n2382, n2380, n2368, n2373, n2369, n2376, n2377,
 n2370, n2911, n2910, n2913, n2900, n2898, n2919, n2917,
 n2916, n2920, n3019, n3025, n3021, n3032, n3027, n3031,
 n3023, n3030, n3024, n3028, n3020, n3026, n3022, n3029);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n2378, n2382, n2380, n2368, n2373, n2369, n2376, n2377,
 n2370, n2911, n2910, n2913, n2900, n2898, n2919, n2917,
 n2916, n2920, n3019, n3025, n3021, n3032, n3027, n3031,
 n3023, n3030, n3024, n3028, n3020, n3026, n3022, n3029;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
 n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
 n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
 n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
 n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
 n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
 n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
 n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
 n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
 n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
 n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
 n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
 n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
 n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
 n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
 n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
 n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
 n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
 n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
 n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
 n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
 n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
 n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
 n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
 n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
 n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
 n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
 n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
 n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
 n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
 n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
 n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
 n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
 n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
 n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
 n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
 n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
 n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
 n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
 n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
 n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
 n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
 n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
 n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
 n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
 n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
 n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
 n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
 n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
 n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
 n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
 n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
 n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
 n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
 n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
 n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
 n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
 n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
 n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
 n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
 n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
 n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
 n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
 n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
 n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
 n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
 n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
 n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
 n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
 n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
 n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
 n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
 n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
 n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
 n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
 n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
 n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
 n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
 n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
 n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
 n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
 n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
 n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
 n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
 n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
 n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
 n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
 n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
 n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
 n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
 n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
 n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
 n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
 n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
 n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
 n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
 n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
 n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
 n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
 n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
 n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
 n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
 n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
 n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2371,
 n2372, n2374, n2375, n2379, n2381, n2383, n2384, n2385,
 n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
 n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
 n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
 n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
 n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
 n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
 n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
 n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
 n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
 n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
 n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
 n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
 n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
 n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
 n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
 n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
 n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
 n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
 n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
 n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
 n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
 n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
 n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
 n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
 n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
 n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
 n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
 n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
 n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
 n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
 n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
 n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
 n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
 n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
 n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
 n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
 n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
 n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
 n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
 n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
 n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
 n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
 n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
 n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
 n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
 n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
 n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
 n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
 n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
 n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
 n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
 n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
 n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
 n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
 n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
 n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
 n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
 n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
 n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
 n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
 n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
 n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
 n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
 n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
 n2899, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
 n2908, n2909, n2912, n2914, n2915, n2918, n2921, n2922,
 n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
 n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
 n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
 n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
 n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
 n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
 n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
 n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
 n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
 n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
 n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
 n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018;

buf  g0 (n145, n31);
buf  g1 (n68, n26);
buf  g2 (n46, n31);
not  g3 (n75, n13);
buf  g4 (n82, n17);
not  g5 (n152, n6);
not  g6 (n102, n13);
buf  g7 (n131, n15);
not  g8 (n122, n8);
not  g9 (n98, n9);
not  g10 (n115, n18);
not  g11 (n101, n32);
not  g12 (n69, n14);
buf  g13 (n76, n12);
not  g14 (n83, n30);
buf  g15 (n62, n28);
buf  g16 (n133, n2);
buf  g17 (n81, n6);
not  g18 (n34, n13);
buf  g19 (n151, n7);
buf  g20 (n70, n31);
not  g21 (n125, n15);
buf  g22 (n106, n30);
buf  g23 (n91, n11);
not  g24 (n121, n26);
buf  g25 (n45, n16);
buf  g26 (n35, n3);
buf  g27 (n112, n8);
not  g28 (n144, n25);
buf  g29 (n108, n21);
buf  g30 (n130, n31);
buf  g31 (n137, n17);
not  g32 (n139, n14);
not  g33 (n52, n24);
not  g34 (n65, n16);
buf  g35 (n113, n20);
buf  g36 (n66, n5);
not  g37 (n103, n1);
buf  g38 (n126, n10);
buf  g39 (n146, n17);
buf  g40 (n120, n5);
buf  g41 (n92, n2);
buf  g42 (n150, n25);
buf  g43 (n127, n5);
buf  g44 (n73, n10);
not  g45 (n42, n2);
buf  g46 (n50, n8);
buf  g47 (n107, n7);
not  g48 (n94, n10);
not  g49 (n156, n30);
not  g50 (n36, n1);
buf  g51 (n147, n29);
buf  g52 (n118, n27);
buf  g53 (n44, n24);
not  g54 (n128, n7);
not  g55 (n78, n21);
not  g56 (n55, n29);
buf  g57 (n64, n28);
not  g58 (n37, n18);
not  g59 (n141, n12);
not  g60 (n40, n1);
buf  g61 (n67, n23);
not  g62 (n63, n16);
not  g63 (n97, n29);
not  g64 (n155, n27);
buf  g65 (n109, n4);
not  g66 (n119, n4);
not  g67 (n104, n23);
buf  g68 (n149, n2);
buf  g69 (n41, n3);
buf  g70 (n56, n22);
not  g71 (n90, n18);
buf  g72 (n79, n28);
not  g73 (n116, n12);
buf  g74 (n142, n19);
buf  g75 (n88, n19);
not  g76 (n105, n27);
not  g77 (n38, n26);
buf  g78 (n51, n24);
buf  g79 (n77, n27);
not  g80 (n153, n30);
not  g81 (n71, n15);
not  g82 (n84, n23);
buf  g83 (n96, n28);
not  g84 (n53, n18);
buf  g85 (n110, n4);
not  g86 (n117, n5);
buf  g87 (n72, n14);
not  g88 (n136, n21);
buf  g89 (n159, n12);
not  g90 (n148, n9);
not  g91 (n138, n6);
not  g92 (n123, n20);
buf  g93 (n160, n17);
buf  g94 (n140, n20);
not  g95 (n47, n13);
buf  g96 (n54, n6);
buf  g97 (n80, n11);
not  g98 (n129, n25);
not  g99 (n135, n19);
not  g100 (n124, n14);
buf  g101 (n99, n25);
not  g102 (n59, n22);
buf  g103 (n57, n32);
buf  g104 (n134, n19);
not  g105 (n154, n3);
not  g106 (n61, n11);
buf  g107 (n143, n4);
not  g108 (n89, n9);
buf  g109 (n157, n11);
not  g110 (n87, n20);
not  g111 (n111, n23);
buf  g112 (n100, n10);
not  g113 (n85, n32);
buf  g114 (n48, n32);
not  g115 (n49, n7);
not  g116 (n43, n8);
buf  g117 (n95, n22);
buf  g118 (n39, n24);
buf  g119 (n74, n1);
buf  g120 (n132, n15);
buf  g121 (n114, n16);
not  g122 (n158, n21);
buf  g123 (n60, n26);
buf  g124 (n58, n9);
buf  g125 (n93, n22);
not  g126 (n33, n3);
not  g127 (n86, n29);
buf  g128 (n256, n82);
buf  g129 (n432, n56);
not  g130 (n670, n82);
not  g131 (n490, n91);
not  g132 (n411, n148);
not  g133 (n352, n44);
not  g134 (n186, n117);
buf  g135 (n239, n148);
buf  g136 (n348, n149);
buf  g137 (n660, n109);
not  g138 (n513, n76);
not  g139 (n259, n33);
buf  g140 (n629, n126);
not  g141 (n580, n92);
buf  g142 (n632, n116);
not  g143 (n219, n107);
not  g144 (n622, n64);
buf  g145 (n515, n51);
not  g146 (n511, n54);
not  g147 (n551, n66);
buf  g148 (n644, n93);
buf  g149 (n625, n119);
buf  g150 (n571, n38);
not  g151 (n476, n43);
not  g152 (n667, n145);
not  g153 (n270, n119);
buf  g154 (n479, n134);
buf  g155 (n509, n57);
not  g156 (n520, n126);
buf  g157 (n474, n106);
buf  g158 (n415, n140);
buf  g159 (n426, n109);
not  g160 (n453, n158);
buf  g161 (n313, n157);
not  g162 (n535, n50);
not  g163 (n569, n60);
buf  g164 (n231, n47);
not  g165 (n375, n156);
buf  g166 (n350, n130);
not  g167 (n640, n90);
not  g168 (n209, n106);
buf  g169 (n316, n83);
buf  g170 (n454, n47);
buf  g171 (n654, n84);
not  g172 (n178, n103);
buf  g173 (n423, n127);
buf  g174 (n251, n111);
not  g175 (n198, n60);
buf  g176 (n579, n74);
buf  g177 (n643, n93);
not  g178 (n393, n115);
buf  g179 (n366, n98);
buf  g180 (n635, n97);
buf  g181 (n430, n80);
buf  g182 (n340, n147);
buf  g183 (n594, n37);
not  g184 (n387, n84);
not  g185 (n621, n108);
buf  g186 (n176, n103);
buf  g187 (n463, n43);
buf  g188 (n312, n145);
buf  g189 (n344, n138);
buf  g190 (n524, n133);
not  g191 (n433, n33);
not  g192 (n531, n80);
buf  g193 (n372, n88);
not  g194 (n488, n57);
not  g195 (n402, n151);
not  g196 (n438, n117);
buf  g197 (n308, n89);
buf  g198 (n404, n114);
not  g199 (n582, n78);
buf  g200 (n599, n144);
not  g201 (n380, n78);
not  g202 (n195, n150);
buf  g203 (n280, n124);
not  g204 (n518, n39);
buf  g205 (n498, n36);
not  g206 (n578, n112);
not  g207 (n321, n107);
buf  g208 (n371, n84);
not  g209 (n555, n113);
not  g210 (n369, n72);
buf  g211 (n653, n159);
buf  g212 (n566, n113);
buf  g213 (n462, n138);
not  g214 (n317, n55);
not  g215 (n403, n86);
buf  g216 (n249, n129);
not  g217 (n365, n136);
not  g218 (n549, n33);
not  g219 (n218, n143);
buf  g220 (n530, n118);
not  g221 (n457, n120);
not  g222 (n536, n56);
not  g223 (n391, n48);
buf  g224 (n424, n128);
not  g225 (n318, n69);
not  g226 (n492, n61);
not  g227 (n258, n95);
buf  g228 (n480, n114);
not  g229 (n341, n79);
not  g230 (n425, n124);
buf  g231 (n382, n44);
not  g232 (n330, n87);
buf  g233 (n367, n67);
not  g234 (n436, n96);
buf  g235 (n327, n69);
buf  g236 (n494, n138);
not  g237 (n624, n151);
buf  g238 (n534, n131);
not  g239 (n449, n124);
buf  g240 (n378, n67);
buf  g241 (n326, n67);
buf  g242 (n664, n150);
buf  g243 (n416, n122);
not  g244 (n191, n47);
not  g245 (n421, n107);
buf  g246 (n274, n158);
not  g247 (n538, n35);
buf  g248 (n671, n91);
buf  g249 (n276, n153);
buf  g250 (n273, n97);
not  g251 (n557, n154);
buf  g252 (n361, n48);
buf  g253 (n605, n86);
not  g254 (n460, n42);
buf  g255 (n215, n90);
buf  g256 (n461, n92);
buf  g257 (n305, n158);
not  g258 (n633, n132);
buf  g259 (n362, n133);
not  g260 (n172, n160);
buf  g261 (n514, n141);
not  g262 (n564, n156);
not  g263 (n657, n58);
not  g264 (n478, n141);
not  g265 (n440, n58);
not  g266 (n510, n84);
not  g267 (n619, n105);
buf  g268 (n439, n147);
buf  g269 (n207, n52);
not  g270 (n336, n72);
buf  g271 (n243, n155);
not  g272 (n523, n85);
buf  g273 (n290, n34);
buf  g274 (n627, n74);
buf  g275 (n618, n126);
buf  g276 (n663, n53);
not  g277 (n615, n45);
not  g278 (n441, n130);
buf  g279 (n354, n90);
buf  g280 (n601, n144);
not  g281 (n346, n89);
buf  g282 (n634, n35);
buf  g283 (n617, n45);
buf  g284 (n289, n147);
buf  g285 (n166, n155);
not  g286 (n396, n143);
buf  g287 (n641, n142);
buf  g288 (n495, n77);
not  g289 (n174, n145);
buf  g290 (n194, n38);
buf  g291 (n427, n59);
not  g292 (n613, n58);
not  g293 (n279, n110);
buf  g294 (n253, n74);
not  g295 (n659, n64);
buf  g296 (n585, n109);
buf  g297 (n163, n99);
not  g298 (n187, n68);
buf  g299 (n537, n70);
not  g300 (n282, n129);
not  g301 (n482, n129);
buf  g302 (n521, n130);
not  g303 (n502, n71);
not  g304 (n431, n152);
buf  g305 (n568, n88);
buf  g306 (n591, n76);
not  g307 (n244, n60);
buf  g308 (n169, n133);
buf  g309 (n237, n151);
buf  g310 (n604, n104);
buf  g311 (n196, n56);
not  g312 (n584, n52);
not  g313 (n185, n140);
not  g314 (n516, n153);
not  g315 (n303, n108);
not  g316 (n260, n65);
not  g317 (n419, n51);
buf  g318 (n264, n149);
buf  g319 (n322, n103);
buf  g320 (n558, n55);
buf  g321 (n268, n150);
not  g322 (n299, n33);
buf  g323 (n379, n104);
buf  g324 (n473, n100);
not  g325 (n293, n153);
not  g326 (n493, n72);
not  g327 (n503, n152);
buf  g328 (n413, n104);
buf  g329 (n467, n120);
not  g330 (n227, n113);
buf  g331 (n333, n82);
not  g332 (n220, n128);
not  g333 (n489, n134);
buf  g334 (n499, n49);
buf  g335 (n595, n34);
not  g336 (n188, n154);
buf  g337 (n554, n57);
not  g338 (n637, n114);
not  g339 (n353, n76);
buf  g340 (n301, n146);
buf  g341 (n228, n148);
buf  g342 (n281, n41);
not  g343 (n234, n158);
buf  g344 (n505, n124);
not  g345 (n283, n42);
not  g346 (n526, n53);
not  g347 (n587, n127);
not  g348 (n325, n116);
buf  g349 (n307, n72);
not  g350 (n294, n123);
buf  g351 (n500, n41);
buf  g352 (n265, n115);
buf  g353 (n358, n66);
not  g354 (n414, n105);
not  g355 (n338, n46);
buf  g356 (n261, n41);
not  g357 (n355, n87);
buf  g358 (n608, n46);
buf  g359 (n252, n108);
buf  g360 (n412, n68);
not  g361 (n173, n49);
buf  g362 (n248, n155);
not  g363 (n668, n92);
buf  g364 (n610, n143);
not  g365 (n484, n125);
not  g366 (n315, n135);
buf  g367 (n590, n69);
not  g368 (n374, n92);
not  g369 (n639, n86);
not  g370 (n363, n98);
buf  g371 (n184, n136);
buf  g372 (n394, n132);
buf  g373 (n197, n117);
not  g374 (n602, n112);
not  g375 (n177, n54);
not  g376 (n203, n51);
buf  g377 (n247, n63);
not  g378 (n581, n96);
not  g379 (n335, n122);
buf  g380 (n567, n83);
not  g381 (n202, n102);
not  g382 (n669, n100);
not  g383 (n300, n63);
buf  g384 (n550, n85);
buf  g385 (n288, n100);
buf  g386 (n451, n132);
buf  g387 (n342, n147);
not  g388 (n399, n81);
buf  g389 (n540, n141);
not  g390 (n420, n35);
not  g391 (n501, n59);
buf  g392 (n319, n106);
not  g393 (n470, n146);
buf  g394 (n222, n101);
not  g395 (n349, n97);
buf  g396 (n496, n94);
not  g397 (n193, n71);
buf  g398 (n631, n47);
not  g399 (n388, n137);
buf  g400 (n250, n98);
buf  g401 (n309, n101);
not  g402 (n200, n75);
not  g403 (n213, n115);
not  g404 (n477, n160);
not  g405 (n628, n110);
not  g406 (n269, n64);
not  g407 (n435, n94);
not  g408 (n405, n42);
not  g409 (n389, n148);
not  g410 (n409, n36);
buf  g411 (n295, n74);
buf  g412 (n182, n136);
buf  g413 (n612, n133);
buf  g414 (n606, n79);
not  g415 (n533, n37);
not  g416 (n609, n112);
buf  g417 (n271, n130);
not  g418 (n277, n44);
buf  g419 (n257, n123);
not  g420 (n392, n52);
not  g421 (n230, n34);
buf  g422 (n211, n153);
not  g423 (n407, n40);
not  g424 (n339, n55);
buf  g425 (n646, n103);
buf  g426 (n208, n116);
not  g427 (n543, n146);
buf  g428 (n360, n70);
not  g429 (n395, n127);
not  g430 (n444, n125);
buf  g431 (n385, n62);
buf  g432 (n161, n68);
buf  g433 (n486, n119);
not  g434 (n577, n157);
buf  g435 (n661, n146);
not  g436 (n542, n93);
buf  g437 (n614, n135);
buf  g438 (n255, n41);
buf  g439 (n508, n78);
buf  g440 (n216, n118);
buf  g441 (n242, n106);
not  g442 (n466, n121);
buf  g443 (n226, n66);
not  g444 (n655, n61);
buf  g445 (n442, n49);
buf  g446 (n232, n51);
not  g447 (n171, n111);
not  g448 (n570, n43);
not  g449 (n240, n62);
buf  g450 (n650, n88);
not  g451 (n469, n94);
not  g452 (n267, n96);
buf  g453 (n235, n121);
buf  g454 (n323, n81);
not  g455 (n410, n48);
buf  g456 (n170, n137);
not  g457 (n417, n55);
not  g458 (n575, n102);
not  g459 (n456, n126);
not  g460 (n556, n77);
not  g461 (n464, n61);
not  g462 (n468, n136);
buf  g463 (n397, n77);
not  g464 (n636, n69);
buf  g465 (n665, n44);
buf  g466 (n381, n81);
not  g467 (n221, n144);
not  g468 (n297, n118);
not  g469 (n507, n68);
buf  g470 (n370, n36);
not  g471 (n386, n73);
buf  g472 (n656, n77);
buf  g473 (n544, n75);
buf  g474 (n310, n101);
not  g475 (n304, n135);
not  g476 (n201, n91);
buf  g477 (n649, n99);
buf  g478 (n376, n58);
not  g479 (n561, n53);
buf  g480 (n314, n65);
buf  g481 (n332, n56);
buf  g482 (n210, n98);
not  g483 (n246, n111);
buf  g484 (n373, n121);
not  g485 (n547, n73);
buf  g486 (n337, n83);
not  g487 (n334, n140);
buf  g488 (n351, n36);
not  g489 (n406, n134);
buf  g490 (n532, n114);
not  g491 (n164, n159);
buf  g492 (n574, n139);
not  g493 (n598, n159);
not  g494 (n320, n122);
not  g495 (n162, n73);
buf  g496 (n206, n118);
buf  g497 (n546, n80);
buf  g498 (n287, n54);
not  g499 (n552, n149);
buf  g500 (n192, n79);
buf  g501 (n623, n137);
not  g502 (n658, n88);
buf  g503 (n642, n139);
buf  g504 (n465, n86);
buf  g505 (n285, n50);
not  g506 (n238, n94);
not  g507 (n539, n128);
buf  g508 (n607, n105);
buf  g509 (n217, n60);
not  g510 (n278, n150);
buf  g511 (n357, n157);
buf  g512 (n573, n63);
buf  g513 (n225, n123);
buf  g514 (n179, n93);
not  g515 (n229, n97);
buf  g516 (n548, n156);
buf  g517 (n576, n39);
not  g518 (n529, n121);
buf  g519 (n491, n157);
buf  g520 (n377, n37);
buf  g521 (n541, n45);
not  g522 (n284, n64);
not  g523 (n626, n62);
buf  g524 (n400, n129);
not  g525 (n306, n65);
not  g526 (n204, n145);
buf  g527 (n214, n131);
buf  g528 (n560, n120);
buf  g529 (n302, n70);
not  g530 (n190, n139);
not  g531 (n181, n111);
buf  g532 (n364, n100);
not  g533 (n506, n101);
buf  g534 (n630, n57);
buf  g535 (n286, n70);
not  g536 (n448, n91);
buf  g537 (n383, n154);
not  g538 (n458, n138);
buf  g539 (n522, n85);
not  g540 (n616, n120);
buf  g541 (n328, n142);
buf  g542 (n565, n35);
buf  g543 (n620, n65);
buf  g544 (n408, n144);
not  g545 (n292, n116);
buf  g546 (n167, n95);
not  g547 (n600, n53);
buf  g548 (n545, n39);
not  g549 (n638, n90);
buf  g550 (n189, n154);
not  g551 (n443, n119);
not  g552 (n311, n104);
not  g553 (n647, n75);
not  g554 (n603, n128);
buf  g555 (n611, n155);
not  g556 (n418, n152);
buf  g557 (n553, n46);
not  g558 (n459, n34);
buf  g559 (n175, n45);
buf  g560 (n672, n149);
buf  g561 (n483, n73);
buf  g562 (n666, n95);
buf  g563 (n296, n95);
buf  g564 (n272, n125);
not  g565 (n471, n63);
not  g566 (n455, n54);
not  g567 (n662, n80);
not  g568 (n597, n40);
buf  g569 (n384, n102);
buf  g570 (n429, n112);
buf  g571 (n572, n143);
buf  g572 (n398, n48);
not  g573 (n475, n107);
buf  g574 (n651, n131);
not  g575 (n437, n96);
buf  g576 (n596, n50);
not  g577 (n528, n52);
not  g578 (n517, n50);
not  g579 (n434, n87);
not  g580 (n359, n139);
buf  g581 (n446, n127);
buf  g582 (n262, n42);
buf  g583 (n487, n79);
not  g584 (n212, n82);
not  g585 (n593, n123);
buf  g586 (n266, n137);
buf  g587 (n481, n78);
buf  g588 (n275, n142);
buf  g589 (n329, n66);
not  g590 (n245, n141);
buf  g591 (n504, n159);
not  g592 (n445, n75);
not  g593 (n485, n115);
buf  g594 (n298, n59);
buf  g595 (n497, n89);
buf  g596 (n428, n110);
buf  g597 (n241, n46);
buf  g598 (n347, n117);
buf  g599 (n324, n89);
not  g600 (n559, n131);
not  g601 (n401, n38);
buf  g602 (n452, n40);
not  g603 (n254, n105);
not  g604 (n525, n49);
not  g605 (n356, n71);
buf  g606 (n331, n99);
buf  g607 (n645, n125);
not  g608 (n562, n160);
buf  g609 (n563, n110);
not  g610 (n199, n156);
buf  g611 (n343, n113);
buf  g612 (n233, n61);
not  g613 (n224, n108);
buf  g614 (n472, n83);
not  g615 (n447, n140);
not  g616 (n512, n62);
not  g617 (n168, n81);
buf  g618 (n183, n99);
not  g619 (n236, n71);
not  g620 (n588, n102);
buf  g621 (n205, n76);
buf  g622 (n527, n135);
not  g623 (n592, n134);
not  g624 (n165, n132);
buf  g625 (n519, n85);
not  g626 (n368, n142);
buf  g627 (n589, n122);
not  g628 (n223, n37);
not  g629 (n390, n38);
not  g630 (n422, n87);
buf  g631 (n450, n109);
buf  g632 (n345, n160);
buf  g633 (n263, n59);
buf  g634 (n652, n152);
buf  g635 (n583, n39);
buf  g636 (n291, n43);
not  g637 (n586, n40);
buf  g638 (n180, n67);
buf  g639 (n648, n151);
not  g640 (n1176, n200);
not  g641 (n1404, n427);
buf  g642 (n815, n560);
buf  g643 (n863, n327);
not  g644 (n1984, n514);
buf  g645 (n1926, n490);
not  g646 (n992, n639);
not  g647 (n1976, n192);
not  g648 (n1393, n633);
buf  g649 (n1119, n379);
buf  g650 (n1184, n342);
buf  g651 (n1385, n271);
buf  g652 (n1298, n197);
not  g653 (n1880, n353);
buf  g654 (n1470, n524);
not  g655 (n1153, n235);
buf  g656 (n1566, n333);
buf  g657 (n779, n545);
not  g658 (n1143, n407);
not  g659 (n1797, n212);
not  g660 (n740, n392);
buf  g661 (n861, n493);
buf  g662 (n1693, n303);
not  g663 (n1979, n425);
buf  g664 (n816, n468);
not  g665 (n1239, n405);
not  g666 (n1414, n619);
buf  g667 (n1685, n552);
not  g668 (n1730, n649);
buf  g669 (n1937, n349);
buf  g670 (n1401, n513);
buf  g671 (n806, n415);
not  g672 (n1758, n567);
buf  g673 (n1552, n550);
not  g674 (n1073, n288);
not  g675 (n1275, n658);
buf  g676 (n1613, n315);
not  g677 (n978, n195);
not  g678 (n719, n515);
buf  g679 (n731, n364);
not  g680 (n1063, n290);
buf  g681 (n1811, n354);
buf  g682 (n1016, n615);
buf  g683 (n772, n223);
not  g684 (n1326, n381);
buf  g685 (n998, n365);
not  g686 (n682, n340);
not  g687 (n790, n498);
not  g688 (n1112, n293);
buf  g689 (n696, n544);
not  g690 (n1828, n578);
not  g691 (n1860, n609);
buf  g692 (n1410, n426);
not  g693 (n1780, n610);
buf  g694 (n1922, n325);
not  g695 (n683, n428);
not  g696 (n1429, n518);
not  g697 (n1158, n367);
not  g698 (n1936, n255);
buf  g699 (n1686, n372);
not  g700 (n1731, n478);
buf  g701 (n1286, n261);
buf  g702 (n1966, n333);
buf  g703 (n1457, n472);
buf  g704 (n1005, n287);
buf  g705 (n1174, n474);
not  g706 (n1588, n421);
not  g707 (n1062, n234);
not  g708 (n1565, n240);
not  g709 (n780, n312);
not  g710 (n1909, n624);
buf  g711 (n1647, n443);
buf  g712 (n1316, n324);
not  g713 (n1015, n279);
buf  g714 (n1083, n443);
buf  g715 (n1992, n430);
buf  g716 (n1202, n323);
not  g717 (n982, n538);
buf  g718 (n1204, n445);
buf  g719 (n1628, n191);
not  g720 (n1026, n176);
buf  g721 (n883, n418);
not  g722 (n1609, n474);
buf  g723 (n846, n518);
buf  g724 (n929, n297);
buf  g725 (n1506, n347);
not  g726 (n1141, n568);
not  g727 (n1216, n621);
buf  g728 (n898, n189);
buf  g729 (n1952, n341);
not  g730 (n1471, n546);
buf  g731 (n1230, n640);
buf  g732 (n753, n177);
buf  g733 (n1807, n177);
buf  g734 (n1453, n627);
buf  g735 (n1490, n585);
not  g736 (n1717, n183);
not  g737 (n1111, n237);
not  g738 (n1580, n281);
not  g739 (n1514, n401);
not  g740 (n768, n533);
buf  g741 (n766, n626);
not  g742 (n937, n276);
not  g743 (n1182, n181);
buf  g744 (n1343, n360);
buf  g745 (n1048, n525);
not  g746 (n1555, n345);
not  g747 (n1113, n201);
not  g748 (n1077, n660);
not  g749 (n938, n194);
buf  g750 (n1712, n661);
buf  g751 (n1739, n227);
not  g752 (n1528, n273);
buf  g753 (n1480, n452);
buf  g754 (n1545, n437);
not  g755 (n1496, n532);
buf  g756 (n755, n482);
not  g757 (n1579, n668);
buf  g758 (n1257, n393);
buf  g759 (n1368, n484);
not  g760 (n1150, n367);
not  g761 (n1249, n312);
buf  g762 (n1959, n579);
buf  g763 (n1595, n224);
not  g764 (n1208, n581);
buf  g765 (n1439, n438);
not  g766 (n1715, n243);
not  g767 (n1713, n246);
not  g768 (n1869, n569);
not  g769 (n830, n318);
not  g770 (n1200, n417);
not  g771 (n1965, n245);
buf  g772 (n1370, n439);
not  g773 (n1803, n294);
buf  g774 (n1955, n665);
not  g775 (n1582, n220);
buf  g776 (n1229, n524);
not  g777 (n1755, n391);
not  g778 (n824, n458);
buf  g779 (n1052, n599);
buf  g780 (n1638, n659);
buf  g781 (n1667, n666);
buf  g782 (n1584, n286);
buf  g783 (n904, n229);
buf  g784 (n912, n640);
not  g785 (n1919, n486);
buf  g786 (n1900, n192);
not  g787 (n1219, n366);
not  g788 (n1155, n528);
not  g789 (n1818, n665);
not  g790 (n1525, n667);
not  g791 (n769, n371);
buf  g792 (n1866, n582);
not  g793 (n1165, n565);
buf  g794 (n729, n350);
not  g795 (n1978, n231);
not  g796 (n1245, n269);
not  g797 (n1315, n278);
not  g798 (n1804, n645);
buf  g799 (n1655, n344);
not  g800 (n1627, n169);
buf  g801 (n758, n432);
buf  g802 (n1235, n444);
buf  g803 (n765, n312);
not  g804 (n954, n319);
not  g805 (n745, n473);
not  g806 (n925, n413);
not  g807 (n1832, n436);
not  g808 (n744, n454);
buf  g809 (n1574, n174);
buf  g810 (n1222, n614);
not  g811 (n1935, n547);
buf  g812 (n1932, n171);
buf  g813 (n1640, n307);
buf  g814 (n1199, n343);
not  g815 (n997, n351);
not  g816 (n1433, n638);
not  g817 (n1908, n376);
not  g818 (n920, n341);
buf  g819 (n1762, n617);
buf  g820 (n1633, n515);
not  g821 (n1277, n556);
not  g822 (n673, n308);
buf  g823 (n1511, n510);
not  g824 (n1617, n195);
not  g825 (n1741, n406);
buf  g826 (n985, n250);
not  g827 (n1639, n316);
not  g828 (n1341, n305);
not  g829 (n736, n667);
not  g830 (n1331, n357);
buf  g831 (n1768, n522);
buf  g832 (n1029, n479);
buf  g833 (n1195, n586);
buf  g834 (n864, n386);
buf  g835 (n1918, n343);
buf  g836 (n1875, n601);
not  g837 (n1134, n600);
buf  g838 (n1972, n461);
buf  g839 (n1748, n391);
not  g840 (n1040, n669);
buf  g841 (n1554, n431);
not  g842 (n807, n164);
not  g843 (n1534, n566);
buf  g844 (n1347, n246);
buf  g845 (n770, n567);
not  g846 (n852, n376);
not  g847 (n1250, n650);
buf  g848 (n777, n648);
not  g849 (n1697, n324);
not  g850 (n1749, n384);
not  g851 (n1201, n522);
buf  g852 (n1775, n478);
buf  g853 (n1690, n377);
buf  g854 (n1577, n592);
buf  g855 (n1017, n388);
buf  g856 (n1102, n353);
not  g857 (n1785, n185);
not  g858 (n1898, n498);
buf  g859 (n1567, n279);
buf  g860 (n1232, n327);
not  g861 (n1968, n664);
buf  g862 (n1967, n242);
buf  g863 (n838, n189);
not  g864 (n1809, n564);
not  g865 (n1246, n644);
not  g866 (n1927, n495);
not  g867 (n814, n475);
buf  g868 (n1161, n326);
buf  g869 (n1197, n219);
not  g870 (n1355, n603);
not  g871 (n1556, n516);
not  g872 (n1413, n310);
buf  g873 (n1561, n268);
not  g874 (n1665, n230);
not  g875 (n1289, n289);
buf  g876 (n1242, n263);
not  g877 (n968, n343);
not  g878 (n1663, n359);
buf  g879 (n1189, n238);
not  g880 (n709, n330);
not  g881 (n1318, n226);
buf  g882 (n1151, n354);
buf  g883 (n1144, n335);
buf  g884 (n1808, n446);
not  g885 (n1795, n199);
not  g886 (n1600, n395);
buf  g887 (n1290, n262);
not  g888 (n1362, n577);
not  g889 (n928, n175);
not  g890 (n720, n493);
buf  g891 (n1962, n399);
buf  g892 (n718, n629);
buf  g893 (n1352, n274);
not  g894 (n1886, n507);
not  g895 (n1622, n510);
not  g896 (n1604, n609);
not  g897 (n1537, n338);
not  g898 (n1256, n642);
buf  g899 (n1445, n539);
not  g900 (n1503, n535);
not  g901 (n1078, n466);
not  g902 (n1397, n326);
buf  g903 (n1312, n427);
not  g904 (n1253, n547);
not  g905 (n1894, n472);
buf  g906 (n1774, n494);
buf  g907 (n1380, n169);
buf  g908 (n1434, n285);
not  g909 (n805, n641);
buf  g910 (n1706, n240);
not  g911 (n1532, n366);
buf  g912 (n952, n635);
not  g913 (n1501, n637);
not  g914 (n1076, n486);
buf  g915 (n702, n589);
not  g916 (n1887, n371);
not  g917 (n1864, n488);
not  g918 (n1363, n522);
not  g919 (n784, n208);
not  g920 (n1897, n416);
buf  g921 (n1314, n496);
buf  g922 (n1190, n221);
not  g923 (n886, n537);
buf  g924 (n873, n642);
buf  g925 (n730, n421);
buf  g926 (n927, n546);
buf  g927 (n1881, n548);
buf  g928 (n1116, n508);
not  g929 (n1754, n493);
not  g930 (n1572, n172);
buf  g931 (n1440, n575);
buf  g932 (n1702, n235);
not  g933 (n1548, n629);
not  g934 (n717, n659);
not  g935 (n1065, n598);
buf  g936 (n847, n638);
buf  g937 (n713, n435);
buf  g938 (n1039, n272);
not  g939 (n1133, n477);
not  g940 (n836, n167);
not  g941 (n1024, n259);
buf  g942 (n988, n215);
not  g943 (n686, n464);
not  g944 (n1895, n672);
not  g945 (n1814, n227);
not  g946 (n1110, n184);
not  g947 (n1943, n242);
not  g948 (n697, n444);
not  g949 (n1276, n264);
buf  g950 (n1179, n355);
buf  g951 (n823, n208);
not  g952 (n1090, n660);
buf  g953 (n1193, n453);
not  g954 (n1166, n540);
buf  g955 (n1435, n601);
not  g956 (n1261, n596);
buf  g957 (n1294, n557);
not  g958 (n1226, n417);
not  g959 (n800, n222);
not  g960 (n1046, n505);
buf  g961 (n939, n475);
not  g962 (n1304, n292);
not  g963 (n1645, n583);
buf  g964 (n1420, n383);
not  g965 (n1280, n637);
buf  g966 (n1870, n571);
not  g967 (n1425, n423);
buf  g968 (n1441, n643);
buf  g969 (n843, n181);
not  g970 (n1668, n276);
buf  g971 (n1837, n588);
buf  g972 (n1949, n187);
buf  g973 (n712, n521);
buf  g974 (n1842, n558);
buf  g975 (n1549, n416);
buf  g976 (n1454, n429);
buf  g977 (n727, n257);
not  g978 (n1779, n444);
not  g979 (n909, n523);
not  g980 (n828, n450);
not  g981 (n1862, n492);
buf  g982 (n906, n516);
buf  g983 (n1101, n226);
not  g984 (n1971, n577);
not  g985 (n953, n433);
buf  g986 (n716, n314);
buf  g987 (n1474, n491);
buf  g988 (n1516, n355);
buf  g989 (n1293, n485);
not  g990 (n1233, n671);
not  g991 (n1497, n639);
buf  g992 (n1356, n567);
buf  g993 (n1183, n313);
not  g994 (n1231, n339);
not  g995 (n809, n446);
not  g996 (n1732, n347);
not  g997 (n1542, n241);
not  g998 (n1846, n190);
not  g999 (n1092, n294);
buf  g1000 (n885, n365);
buf  g1001 (n1263, n336);
buf  g1002 (n1626, n354);
not  g1003 (n1834, n216);
not  g1004 (n797, n194);
buf  g1005 (n1657, n543);
not  g1006 (n1989, n448);
buf  g1007 (n1623, n606);
buf  g1008 (n1904, n536);
not  g1009 (n1742, n429);
not  g1010 (n796, n190);
not  g1011 (n1265, n514);
buf  g1012 (n1191, n208);
buf  g1013 (n1325, n192);
not  g1014 (n1529, n652);
not  g1015 (n1852, n238);
buf  g1016 (n1391, n400);
buf  g1017 (n1213, n547);
not  g1018 (n1423, n559);
buf  g1019 (n711, n563);
not  g1020 (n774, n582);
buf  g1021 (n1011, n278);
buf  g1022 (n1666, n363);
buf  g1023 (n1344, n311);
buf  g1024 (n1139, n223);
buf  g1025 (n1057, n521);
not  g1026 (n1699, n605);
buf  g1027 (n1095, n392);
not  g1028 (n943, n583);
not  g1029 (n1778, n212);
not  g1030 (n866, n166);
not  g1031 (n812, n531);
buf  g1032 (n1675, n203);
buf  g1033 (n1430, n237);
not  g1034 (n1196, n292);
buf  g1035 (n1032, n396);
buf  g1036 (n1964, n590);
not  g1037 (n1008, n203);
not  g1038 (n1513, n480);
not  g1039 (n1939, n266);
buf  g1040 (n1763, n621);
not  g1041 (n1418, n470);
not  g1042 (n1462, n570);
not  g1043 (n1973, n375);
not  g1044 (n1218, n398);
not  g1045 (n1386, n382);
buf  g1046 (n1969, n300);
buf  g1047 (n1912, n414);
buf  g1048 (n1892, n243);
buf  g1049 (n1099, n362);
buf  g1050 (n1185, n578);
buf  g1051 (n1075, n263);
not  g1052 (n1759, n545);
buf  g1053 (n808, n583);
buf  g1054 (n701, n594);
not  g1055 (n1338, n662);
not  g1056 (n1890, n556);
buf  g1057 (n1871, n655);
not  g1058 (n1392, n441);
buf  g1059 (n1688, n648);
not  g1060 (n793, n407);
buf  g1061 (n1268, n657);
not  g1062 (n1771, n212);
not  g1063 (n1096, n294);
not  g1064 (n1540, n644);
buf  g1065 (n1181, n626);
buf  g1066 (n1982, n364);
buf  g1067 (n1586, n284);
buf  g1068 (n1776, n388);
not  g1069 (n1827, n379);
buf  g1070 (n1980, n352);
buf  g1071 (n829, n342);
not  g1072 (n1054, n313);
buf  g1073 (n1535, n653);
buf  g1074 (n1933, n467);
not  g1075 (n1320, n201);
not  g1076 (n1074, n595);
not  g1077 (n786, n180);
buf  g1078 (n1679, n334);
buf  g1079 (n1883, n278);
buf  g1080 (n1030, n618);
buf  g1081 (n1168, n597);
not  g1082 (n921, n187);
buf  g1083 (n1615, n323);
not  g1084 (n1327, n634);
not  g1085 (n1526, n429);
buf  g1086 (n1473, n198);
not  g1087 (n1757, n395);
not  g1088 (n1172, n597);
not  g1089 (n1995, n337);
buf  g1090 (n1192, n304);
not  g1091 (n1616, n451);
buf  g1092 (n983, n502);
not  g1093 (n1491, n521);
not  g1094 (n1854, n613);
buf  g1095 (n1359, n196);
buf  g1096 (n826, n244);
not  g1097 (n1996, n504);
buf  g1098 (n1390, n666);
not  g1099 (n1488, n461);
not  g1100 (n1210, n189);
buf  g1101 (n1993, n371);
buf  g1102 (n1212, n517);
buf  g1103 (n675, n198);
buf  g1104 (n1700, n613);
not  g1105 (n947, n220);
not  g1106 (n1387, n562);
buf  g1107 (n1823, n480);
not  g1108 (n1123, n466);
not  g1109 (n1942, n193);
buf  g1110 (n1861, n185);
buf  g1111 (n1751, n286);
not  g1112 (n778, n611);
not  g1113 (n1389, n585);
not  g1114 (n1375, n410);
buf  g1115 (n1381, n334);
not  g1116 (n1388, n308);
not  g1117 (n1303, n364);
buf  g1118 (n1028, n230);
buf  g1119 (n1125, n333);
buf  g1120 (n869, n465);
buf  g1121 (n989, n240);
buf  g1122 (n1041, n348);
not  g1123 (n1658, n224);
not  g1124 (n703, n233);
not  g1125 (n1371, n164);
buf  g1126 (n1591, n301);
not  g1127 (n1209, n242);
buf  g1128 (n1681, n552);
buf  g1129 (n1906, n266);
buf  g1130 (n1902, n619);
buf  g1131 (n750, n319);
not  g1132 (n773, n602);
not  g1133 (n1521, n368);
buf  g1134 (n1499, n604);
not  g1135 (n1136, n179);
not  g1136 (n919, n501);
buf  g1137 (n962, n528);
not  g1138 (n822, n325);
not  g1139 (n1510, n612);
buf  g1140 (n1308, n455);
not  g1141 (n708, n320);
not  g1142 (n1374, n490);
buf  g1143 (n1899, n657);
not  g1144 (n1769, n442);
buf  g1145 (n676, n374);
not  g1146 (n738, n439);
not  g1147 (n781, n640);
buf  g1148 (n1800, n527);
buf  g1149 (n1531, n178);
buf  g1150 (n1406, n241);
not  g1151 (n1081, n499);
not  g1152 (n1324, n627);
not  g1153 (n1448, n324);
buf  g1154 (n1879, n300);
buf  g1155 (n1476, n547);
not  g1156 (n1252, n236);
not  g1157 (n1940, n472);
not  g1158 (n1402, n529);
not  g1159 (n922, n570);
buf  g1160 (n1653, n383);
not  g1161 (n1928, n270);
buf  g1162 (n1475, n385);
not  g1163 (n990, n519);
buf  g1164 (n694, n447);
buf  g1165 (n1154, n195);
not  g1166 (n677, n380);
not  g1167 (n915, n211);
not  g1168 (n1925, n614);
not  g1169 (n1705, n540);
not  g1170 (n879, n650);
buf  g1171 (n1121, n477);
buf  g1172 (n1664, n244);
buf  g1173 (n1722, n434);
not  g1174 (n1247, n357);
buf  g1175 (n839, n369);
buf  g1176 (n1127, n182);
not  g1177 (n986, n363);
buf  g1178 (n1203, n308);
not  g1179 (n1954, n302);
not  g1180 (n840, n573);
buf  g1181 (n1849, n634);
not  g1182 (n1422, n436);
buf  g1183 (n1281, n530);
not  g1184 (n1553, n622);
not  g1185 (n1103, n524);
buf  g1186 (n963, n636);
buf  g1187 (n959, n239);
not  g1188 (n1288, n586);
buf  g1189 (n1601, n642);
not  g1190 (n1287, n468);
buf  g1191 (n1848, n204);
not  g1192 (n1427, n633);
buf  g1193 (n1736, n572);
not  g1194 (n723, n574);
not  g1195 (n741, n259);
not  g1196 (n1794, n469);
buf  g1197 (n1305, n647);
not  g1198 (n1876, n389);
buf  g1199 (n1021, n380);
not  g1200 (n1369, n621);
buf  g1201 (n1207, n422);
buf  g1202 (n1505, n550);
not  g1203 (n1033, n180);
not  g1204 (n1098, n633);
not  g1205 (n1042, n659);
not  g1206 (n896, n351);
buf  g1207 (n882, n614);
not  g1208 (n1527, n263);
buf  g1209 (n1224, n513);
buf  g1210 (n692, n413);
not  g1211 (n1117, n649);
buf  g1212 (n1292, n494);
buf  g1213 (n1610, n376);
not  g1214 (n1711, n452);
not  g1215 (n1129, n189);
not  g1216 (n958, n503);
not  g1217 (n1345, n529);
not  g1218 (n913, n512);
buf  g1219 (n1585, n304);
buf  g1220 (n1157, n355);
buf  g1221 (n1752, n519);
buf  g1222 (n1118, n205);
not  g1223 (n1421, n630);
buf  g1224 (n1524, n268);
not  g1225 (n1563, n553);
not  g1226 (n1632, n610);
not  g1227 (n1456, n378);
not  g1228 (n795, n307);
not  g1229 (n930, n222);
not  g1230 (n1047, n575);
not  g1231 (n995, n467);
not  g1232 (n1882, n609);
buf  g1233 (n724, n232);
not  g1234 (n1784, n638);
buf  g1235 (n757, n213);
buf  g1236 (n1598, n413);
not  g1237 (n1272, n216);
not  g1238 (n1772, n352);
buf  g1239 (n1990, n657);
not  g1240 (n1307, n188);
not  g1241 (n1167, n512);
buf  g1242 (n818, n459);
buf  g1243 (n1648, n344);
not  g1244 (n1336, n213);
not  g1245 (n1999, n167);
not  g1246 (n1614, n345);
buf  g1247 (n1630, n254);
not  g1248 (n698, n287);
not  g1249 (n813, n615);
not  g1250 (n1659, n435);
buf  g1251 (n1517, n262);
not  g1252 (n1455, n411);
not  g1253 (n1677, n183);
not  g1254 (n1850, n247);
not  g1255 (n1502, n642);
buf  g1256 (n941, n252);
buf  g1257 (n1350, n311);
buf  g1258 (n1970, n398);
buf  g1259 (n1340, n587);
not  g1260 (n1003, n269);
buf  g1261 (n1160, n450);
not  g1262 (n1379, n217);
buf  g1263 (n1518, n290);
buf  g1264 (n832, n481);
not  g1265 (n1093, n281);
buf  g1266 (n1634, n517);
buf  g1267 (n934, n191);
buf  g1268 (n1255, n395);
buf  g1269 (n1091, n561);
buf  g1270 (n1793, n402);
buf  g1271 (n1512, n541);
buf  g1272 (n1006, n325);
not  g1273 (n1469, n329);
buf  g1274 (n1236, n631);
buf  g1275 (n1671, n538);
buf  g1276 (n1539, n620);
buf  g1277 (n1500, n436);
buf  g1278 (n821, n356);
buf  g1279 (n1351, n247);
not  g1280 (n783, n636);
not  g1281 (n1788, n289);
buf  g1282 (n944, n481);
not  g1283 (n1743, n180);
buf  g1284 (n1703, n168);
buf  g1285 (n1237, n485);
buf  g1286 (n946, n496);
buf  g1287 (n1284, n644);
buf  g1288 (n1443, n581);
not  g1289 (n1045, n482);
buf  g1290 (n970, n617);
not  g1291 (n1452, n249);
buf  g1292 (n1104, n631);
buf  g1293 (n900, n639);
buf  g1294 (n693, n284);
not  g1295 (n1559, n240);
buf  g1296 (n865, n417);
not  g1297 (n1468, n556);
buf  g1298 (n833, n283);
buf  g1299 (n1729, n628);
buf  g1300 (n1447, n305);
not  g1301 (n1296, n473);
buf  g1302 (n1383, n163);
buf  g1303 (n1910, n439);
buf  g1304 (n1641, n234);
buf  g1305 (n1661, n496);
buf  g1306 (n1704, n241);
not  g1307 (n1198, n344);
buf  g1308 (n1587, n389);
buf  g1309 (n1815, n428);
buf  g1310 (n1631, n570);
buf  g1311 (n1486, n163);
not  g1312 (n1960, n405);
buf  g1313 (n700, n664);
not  g1314 (n848, n161);
not  g1315 (n887, n574);
not  g1316 (n1789, n661);
not  g1317 (n1411, n288);
not  g1318 (n1988, n654);
not  g1319 (n1373, n300);
not  g1320 (n1007, n211);
buf  g1321 (n1206, n289);
buf  g1322 (n993, n316);
buf  g1323 (n1805, n558);
not  g1324 (n880, n441);
buf  g1325 (n1520, n486);
not  g1326 (n1737, n562);
not  g1327 (n1415, n201);
buf  g1328 (n1000, n271);
buf  g1329 (n1796, n464);
buf  g1330 (n1863, n213);
not  g1331 (n1132, n440);
not  g1332 (n1825, n668);
not  g1333 (n969, n440);
buf  g1334 (n893, n346);
buf  g1335 (n1025, n490);
buf  g1336 (n1728, n603);
buf  g1337 (n899, n500);
not  g1338 (n908, n591);
buf  g1339 (n845, n379);
buf  g1340 (n1084, n373);
not  g1341 (n960, n309);
not  g1342 (n1100, n384);
buf  g1343 (n1405, n381);
buf  g1344 (n1164, n272);
buf  g1345 (n984, n225);
not  g1346 (n1560, n345);
not  g1347 (n1186, n489);
buf  g1348 (n1509, n250);
buf  g1349 (n1187, n663);
buf  g1350 (n1901, n271);
not  g1351 (n1654, n514);
not  g1352 (n1673, n306);
not  g1353 (n1258, n278);
not  g1354 (n1558, n267);
buf  g1355 (n1254, n317);
buf  g1356 (n1546, n596);
buf  g1357 (n1896, n626);
not  g1358 (n1056, n374);
buf  g1359 (n1958, n535);
not  g1360 (n1330, n497);
buf  g1361 (n895, n569);
not  g1362 (n1377, n199);
not  g1363 (n1914, n338);
buf  g1364 (n1485, n581);
buf  g1365 (n1777, n470);
buf  g1366 (n881, n532);
not  g1367 (n728, n382);
buf  g1368 (n1396, n380);
not  g1369 (n1472, n275);
buf  g1370 (n1354, n510);
not  g1371 (n1142, n492);
buf  g1372 (n810, n432);
not  g1373 (n1953, n511);
not  g1374 (n782, n473);
not  g1375 (n1251, n497);
buf  g1376 (n994, n402);
not  g1377 (n1279, n187);
buf  g1378 (n1066, n625);
not  g1379 (n1605, n448);
buf  g1380 (n1266, n590);
buf  g1381 (n877, n270);
not  g1382 (n1740, n258);
not  g1383 (n1050, n531);
not  g1384 (n974, n314);
buf  g1385 (n1813, n624);
not  g1386 (n1214, n424);
buf  g1387 (n945, n453);
not  g1388 (n911, n668);
buf  g1389 (n975, n264);
not  g1390 (n1306, n162);
not  g1391 (n981, n233);
not  g1392 (n820, n595);
buf  g1393 (n1140, n332);
buf  g1394 (n1603, n487);
buf  g1395 (n1676, n612);
buf  g1396 (n1241, n579);
buf  g1397 (n825, n600);
buf  g1398 (n1467, n392);
buf  g1399 (n1297, n237);
buf  g1400 (n1934, n568);
buf  g1401 (n1035, n286);
buf  g1402 (n1707, n214);
buf  g1403 (n1735, n353);
not  g1404 (n1660, n236);
not  g1405 (n979, n424);
buf  g1406 (n1211, n212);
not  g1407 (n1494, n599);
not  g1408 (n964, n651);
not  g1409 (n1431, n576);
not  g1410 (n1987, n250);
not  g1411 (n1002, n193);
not  g1412 (n1820, n313);
buf  g1413 (n1856, n300);
not  g1414 (n1541, n404);
not  g1415 (n1444, n317);
buf  g1416 (n759, n484);
buf  g1417 (n1915, n402);
not  g1418 (n1309, n396);
buf  g1419 (n1571, n614);
not  g1420 (n1997, n180);
buf  g1421 (n949, n623);
not  g1422 (n1781, n353);
buf  g1423 (n976, n587);
not  g1424 (n1812, n166);
buf  g1425 (n1608, n309);
buf  g1426 (n1851, n622);
not  g1427 (n1822, n368);
buf  g1428 (n888, n582);
not  g1429 (n1624, n235);
buf  g1430 (n1903, n639);
buf  g1431 (n739, n304);
not  g1432 (n1115, n261);
buf  g1433 (n1547, n514);
not  g1434 (n1152, n611);
not  g1435 (n1365, n454);
buf  g1436 (n1612, n308);
not  g1437 (n1259, n528);
not  g1438 (n1097, n480);
not  g1439 (n767, n328);
buf  g1440 (n1865, n296);
not  g1441 (n1124, n350);
buf  g1442 (n1037, n340);
buf  g1443 (n1924, n419);
not  g1444 (n1360, n210);
buf  g1445 (n1720, n579);
buf  g1446 (n722, n296);
buf  g1447 (n1721, n322);
not  g1448 (n1551, n432);
buf  g1449 (n1859, n217);
buf  g1450 (n1438, n310);
buf  g1451 (n1416, n627);
not  g1452 (n674, n358);
not  g1453 (n1599, n468);
buf  g1454 (n1597, n391);
buf  g1455 (n932, n424);
not  g1456 (n1782, n457);
not  g1457 (n1868, n242);
not  g1458 (n801, n401);
not  g1459 (n1376, n422);
buf  g1460 (n714, n628);
buf  g1461 (n1051, n476);
buf  g1462 (n1043, n281);
buf  g1463 (n1508, n197);
not  g1464 (n1515, n291);
buf  g1465 (n1493, n162);
not  g1466 (n1946, n563);
not  g1467 (n841, n657);
buf  g1468 (n1642, n495);
not  g1469 (n1044, n394);
not  g1470 (n1923, n589);
not  g1471 (n1727, n216);
buf  g1472 (n1747, n176);
not  g1473 (n1145, n172);
buf  g1474 (n1719, n663);
buf  g1475 (n1346, n594);
buf  g1476 (n1372, n592);
buf  g1477 (n1921, n217);
buf  g1478 (n1714, n660);
buf  g1479 (n1643, n463);
buf  g1480 (n1107, n669);
buf  g1481 (n1361, n569);
buf  g1482 (n1977, n272);
buf  g1483 (n1644, n362);
not  g1484 (n1929, n209);
buf  g1485 (n894, n369);
not  g1486 (n1507, n497);
not  g1487 (n1985, n560);
not  g1488 (n1170, n447);
buf  g1489 (n751, n615);
buf  g1490 (n1328, n401);
buf  g1491 (n1282, n501);
not  g1492 (n844, n233);
not  g1493 (n1020, n541);
not  g1494 (n725, n591);
buf  g1495 (n1426, n254);
buf  g1496 (n1543, n295);
buf  g1497 (n1138, n576);
not  g1498 (n870, n264);
buf  g1499 (n878, n426);
not  g1500 (n1710, n602);
buf  g1501 (n884, n331);
buf  g1502 (n1244, n531);
buf  g1503 (n1135, n275);
not  g1504 (n907, n203);
buf  g1505 (n1761, n449);
not  g1506 (n684, n447);
buf  g1507 (n966, n265);
buf  g1508 (n1635, n370);
not  g1509 (n1482, n341);
buf  g1510 (n1269, n554);
buf  g1511 (n991, n541);
buf  g1512 (n1273, n246);
buf  g1513 (n1357, n530);
buf  g1514 (n1650, n383);
not  g1515 (n1055, n285);
buf  g1516 (n1082, n291);
buf  g1517 (n1678, n448);
not  g1518 (n1223, n256);
buf  g1519 (n1698, n455);
buf  g1520 (n853, n327);
buf  g1521 (n1951, n672);
buf  g1522 (n1399, n257);
not  g1523 (n1228, n564);
not  g1524 (n1023, n609);
not  g1525 (n1072, n198);
buf  g1526 (n1461, n254);
not  g1527 (n1106, n437);
buf  g1528 (n1773, n533);
buf  g1529 (n903, n631);
not  g1530 (n789, n425);
not  g1531 (n1873, n245);
buf  g1532 (n1120, n482);
not  g1533 (n1465, n290);
not  g1534 (n1948, n223);
buf  g1535 (n1691, n573);
not  g1536 (n1329, n494);
not  g1537 (n1672, n188);
buf  g1538 (n1175, n268);
buf  g1539 (n871, n478);
buf  g1540 (n1696, n585);
not  g1541 (n737, n542);
buf  g1542 (n1756, n530);
buf  g1543 (n890, n652);
not  g1544 (n1689, n650);
buf  g1545 (n1913, n541);
buf  g1546 (n1845, n367);
buf  g1547 (n923, n409);
buf  g1548 (n706, n235);
buf  g1549 (n763, n662);
buf  g1550 (n856, n578);
not  g1551 (n897, n538);
not  g1552 (n1619, n231);
not  g1553 (n874, n218);
buf  g1554 (n1802, n534);
not  g1555 (n1844, n269);
buf  g1556 (n854, n375);
not  g1557 (n1417, n506);
buf  g1558 (n1260, n500);
buf  g1559 (n746, n516);
buf  g1560 (n1839, n372);
not  g1561 (n1149, n227);
not  g1562 (n1086, n205);
not  g1563 (n948, n611);
buf  g1564 (n1602, n182);
buf  g1565 (n1994, n196);
buf  g1566 (n688, n457);
buf  g1567 (n1409, n270);
not  g1568 (n977, n239);
buf  g1569 (n1446, n229);
not  g1570 (n1424, n454);
not  g1571 (n1683, n655);
buf  g1572 (n967, n312);
not  g1573 (n916, n323);
not  g1574 (n1504, n184);
not  g1575 (n1333, n163);
not  g1576 (n1726, n168);
not  g1577 (n1162, n292);
buf  g1578 (n1695, n265);
not  g1579 (n1367, n299);
not  g1580 (n1734, n605);
buf  g1581 (n1838, n324);
buf  g1582 (n1147, n218);
buf  g1583 (n1583, n319);
not  g1584 (n1459, n204);
buf  g1585 (n1058, n326);
buf  g1586 (n1339, n515);
buf  g1587 (n1264, n279);
buf  g1588 (n942, n588);
buf  g1589 (n1105, n641);
not  g1590 (n1238, n403);
buf  g1591 (n1094, n350);
buf  g1592 (n1156, n309);
buf  g1593 (n1637, n636);
not  g1594 (n1829, n626);
buf  g1595 (n1464, n305);
not  g1596 (n1412, n302);
buf  g1597 (n1460, n625);
not  g1598 (n867, n162);
buf  g1599 (n1300, n338);
buf  g1600 (n752, n340);
buf  g1601 (n1744, n407);
not  g1602 (n1877, n582);
not  g1603 (n1271, n503);
buf  g1604 (n732, n164);
not  g1605 (n935, n252);
not  g1606 (n1220, n612);
not  g1607 (n1606, n605);
buf  g1608 (n1891, n630);
buf  g1609 (n1819, n564);
not  g1610 (n1986, n277);
not  g1611 (n1087, n311);
buf  g1612 (n872, n417);
not  g1613 (n695, n386);
not  g1614 (n2000, n201);
buf  g1615 (n1944, n178);
not  g1616 (n1646, n375);
buf  g1617 (n1975, n631);
buf  g1618 (n1855, n643);
buf  g1619 (n1384, n209);
buf  g1620 (n1578, n384);
not  g1621 (n955, n648);
not  g1622 (n1395, n248);
not  g1623 (n1745, n231);
buf  g1624 (n1088, n651);
buf  g1625 (n756, n346);
buf  g1626 (n680, n460);
not  g1627 (n1394, n198);
buf  g1628 (n1569, n260);
buf  g1629 (n743, n222);
not  g1630 (n1070, n190);
not  g1631 (n1419, n237);
buf  g1632 (n1835, n372);
buf  g1633 (n1544, n273);
not  g1634 (n1436, n285);
not  g1635 (n1334, n421);
not  g1636 (n1941, n281);
not  g1637 (n1798, n204);
buf  g1638 (n1027, n643);
not  g1639 (n819, n211);
buf  g1640 (n1701, n258);
buf  g1641 (n1278, n430);
not  g1642 (n1843, n534);
buf  g1643 (n1137, n606);
buf  g1644 (n835, n218);
buf  g1645 (n1285, n339);
buf  g1646 (n858, n571);
not  g1647 (n1570, n228);
not  g1648 (n1492, n410);
not  g1649 (n1061, n187);
buf  g1650 (n1981, n311);
buf  g1651 (n1169, n419);
buf  g1652 (n1188, n348);
not  g1653 (n681, n591);
not  g1654 (n1108, n210);
not  g1655 (n1458, n628);
buf  g1656 (n1621, n347);
not  g1657 (n1576, n590);
not  g1658 (n1225, n214);
buf  g1659 (n1765, n429);
buf  g1660 (n1905, n430);
buf  g1661 (n1787, n670);
buf  g1662 (n1594, n595);
buf  g1663 (n1487, n328);
buf  g1664 (n699, n310);
not  g1665 (n1911, n470);
buf  g1666 (n1466, n390);
not  g1667 (n1122, n581);
buf  g1668 (n936, n671);
buf  g1669 (n1568, n418);
not  g1670 (n687, n375);
not  g1671 (n1335, n408);
buf  g1672 (n726, n434);
buf  g1673 (n957, n169);
not  g1674 (n1295, n185);
not  g1675 (n794, n289);
not  g1676 (n1723, n633);
buf  g1677 (n1301, n330);
not  g1678 (n1267, n399);
buf  g1679 (n1611, n364);
buf  g1680 (n834, n299);
not  g1681 (n799, n443);
buf  g1682 (n1767, n182);
buf  g1683 (n851, n267);
buf  g1684 (n1071, n291);
not  g1685 (n1945, n506);
buf  g1686 (n860, n555);
not  g1687 (n1983, n331);
not  g1688 (n1684, n456);
not  g1689 (n827, n170);
not  g1690 (n1291, n634);
not  g1691 (n1366, n174);
buf  g1692 (n1857, n239);
buf  g1693 (n901, n288);
buf  g1694 (n1930, n350);
not  g1695 (n1792, n499);
not  g1696 (n761, n527);
not  g1697 (n1833, n654);
buf  g1698 (n1816, n266);
buf  g1699 (n940, n662);
not  g1700 (n748, n443);
not  g1701 (n1299, n632);
not  g1702 (n1831, n584);
buf  g1703 (n1428, n363);
not  g1704 (n1770, n553);
not  g1705 (n1853, n327);
not  g1706 (n1878, n473);
not  g1707 (n762, n320);
not  g1708 (n1562, n282);
not  g1709 (n1080, n165);
buf  g1710 (n690, n592);
not  g1711 (n791, n195);
not  g1712 (n1173, n359);
buf  g1713 (n811, n544);
not  g1714 (n1353, n580);
buf  g1715 (n1783, n267);
not  g1716 (n1109, n428);
not  g1717 (n1656, n387);
not  g1718 (n910, n249);
not  g1719 (n972, n433);
not  g1720 (n917, n179);
not  g1721 (n1538, n362);
not  g1722 (n837, n578);
not  g1723 (n1938, n322);
not  g1724 (n747, n173);
not  g1725 (n862, n348);
not  g1726 (n831, n458);
buf  g1727 (n1649, n607);
nor  g1728 (n1974, n502, n272, n549, n260);
or   g1729 (n1991, n348, n610, n347, n199);
nand g1730 (n1437, n178, n166, n462, n501);
nand g1731 (n1750, n575, n539, n221, n532);
xor  g1732 (n1262, n262, n460, n492, n555);
or   g1733 (n1519, n523, n339, n209, n170);
xor  g1734 (n1718, n220, n387, n496, n161);
xnor g1735 (n792, n206, n526, n607, n481);
xnor g1736 (n1407, n604, n276, n295, n256);
nor  g1737 (n1342, n407, n385, n231, n232);
and  g1738 (n754, n592, n662, n465, n559);
nand g1739 (n1089, n552, n637, n392, n440);
and  g1740 (n1575, n511, n249, n420, n170);
nor  g1741 (n1248, n608, n301, n510, n455);
nor  g1742 (n1114, n248, n393, n530, n238);
or   g1743 (n1550, n406, n546, n503, n397);
nor  g1744 (n1957, n388, n318, n361, n335);
nand g1745 (n996, n415, n332, n296, n236);
nor  g1746 (n1917, n169, n665, n294, n413);
nand g1747 (n971, n397, n425, n203, n529);
or   g1748 (n1378, n275, n194, n207, n619);
xnor g1749 (n1564, n544, n481, n603, n445);
nor  g1750 (n1893, n545, n596, n411, n464);
xnor g1751 (n1670, n570, n498, n620, n322);
nor  g1752 (n850, n228, n388, n518, n572);
nand g1753 (n1130, n184, n219, n583, n525);
nand g1754 (n1038, n499, n576, n171, n366);
nand g1755 (n1836, n332, n527, n529, n600);
xnor g1756 (n1725, n467, n361, n504, n229);
xor  g1757 (n1830, n168, n221, n433, n625);
or   g1758 (n1947, n587, n342, n457, n435);
nor  g1759 (n1310, n507, n175, n427, n655);
nor  g1760 (n1012, n505, n399, n185, n322);
xor  g1761 (n1205, n399, n397, n484, n230);
xor  g1762 (n1592, n197, n319, n563, n498);
or   g1763 (n1956, n276, n453, n284, n602);
xor  g1764 (n787, n508, n623, n334, n666);
or   g1765 (n710, n359, n584, n450, n419);
xnor g1766 (n1709, n605, n317, n379, n420);
xor  g1767 (n891, n670, n540, n207, n446);
xnor g1768 (n734, n173, n367, n409, n495);
and  g1769 (n924, n296, n374, n440, n172);
nor  g1770 (n1884, n297, n414, n663, n500);
xor  g1771 (n1432, n425, n370, n565, n505);
xor  g1772 (n1221, n580, n329, n504, n389);
nand g1773 (n691, n337, n415, n298, n273);
xor  g1774 (n1589, n251, n448, n479, n546);
nor  g1775 (n1013, n243, n365, n215, n666);
xor  g1776 (n859, n561, n222, n589, n632);
xnor g1777 (n1961, n655, n554, n645, n204);
nor  g1778 (n1620, n434, n178, n535, n219);
nand g1779 (n1692, n539, n526, n303, n493);
nand g1780 (n1180, n619, n622, n403, n554);
xnor g1781 (n956, n587, n298, n458, n543);
xor  g1782 (n1067, n612, n205, n384, n402);
and  g1783 (n1662, n604, n640, n598, n186);
xor  g1784 (n1004, n335, n561, n259, n302);
nor  g1785 (n973, n426, n329, n331, n667);
xnor g1786 (n1031, n523, n622, n543, n351);
xnor g1787 (n1014, n247, n641, n526, n572);
nor  g1788 (n1313, n310, n551, n394, n236);
nand g1789 (n1636, n661, n279, n531, n568);
xnor g1790 (n679, n556, n566, n396, n403);
and  g1791 (n876, n553, n361, n220, n210);
xnor g1792 (n1888, n274, n172, n618, n254);
nand g1793 (n1059, n433, n257, n580, n230);
nand g1794 (n1009, n193, n637, n406, n206);
or   g1795 (n1593, n408, n550, n634, n186);
or   g1796 (n1724, n458, n393, n179, n555);
nand g1797 (n1817, n580, n591, n313, n215);
nand g1798 (n1069, n671, n437, n295, n438);
xor  g1799 (n1786, n460, n405, n656, n306);
xnor g1800 (n689, n224, n461, n306, n246);
or   g1801 (n1858, n618, n549, n227, n190);
xor  g1802 (n1669, n283, n537, n207);
xor  g1803 (n705, n566, n442, n293, n600);
xor  g1804 (n842, n256, n482, n334, n536);
nand g1805 (n1680, n476, n576, n165, n466);
xor  g1806 (n817, n651, n439, n470, n594);
xor  g1807 (n1178, n584, n446, n283, n321);
xnor g1808 (n1270, n360, n377, n459, n176);
or   g1809 (n1449, n275, n357, n534, n646);
xnor g1810 (n1746, n287, n485, n618, n286);
nand g1811 (n1018, n672, n593, n638, n174);
xor  g1812 (n1146, n226, n613, n495, n608);
or   g1813 (n931, n647, n549, n335, n670);
nand g1814 (n1400, n257, n464, n508, n586);
or   g1815 (n1053, n535, n412, n536, n423);
and  g1816 (n1217, n517, n542, n390);
nor  g1817 (n1931, n537, n356, n177, n368);
and  g1818 (n1916, n277, n492, n652, n604);
nor  g1819 (n855, n648, n280, n574, n476);
and  g1820 (n1322, n370, n513, n654, n349);
and  g1821 (n678, n465, n330, n217, n199);
nand g1822 (n1302, n450, n228, n411, n297);
xor  g1823 (n933, n163, n422, n431, n330);
xnor g1824 (n1651, n501, n186, n332, n249);
nand g1825 (n1049, n660, n562, n669, n234);
nand g1826 (n914, n208, n462, n321, n641);
xnor g1827 (n1824, n442, n268, n560, n455);
xor  g1828 (n1001, n293, n255, n459, n196);
xnor g1829 (n1477, n161, n386, n669, n548);
and  g1830 (n1806, n404, n563, n461, n451);
and  g1831 (n1311, n337, n259, n194, n406);
xor  g1832 (n1708, n162, n206, n434, n460);
nand g1833 (n980, n671, n369, n261, n616);
xor  g1834 (n760, n518, n188, n277, n653);
and  g1835 (n1791, n486, n282, n562, n166);
xnor g1836 (n1872, n396, n416, n474, n266);
or   g1837 (n1687, n372, n658, n176, n352);
xor  g1838 (n1674, n390, n488, n377, n632);
or   g1839 (n1319, n523, n467, n412, n445);
nand g1840 (n1126, n616, n505, n298, n282);
and  g1841 (n889, n416, n504, n665, n508);
and  g1842 (n1733, n649, n472, n421, n401);
nor  g1843 (n803, n260, n437, n559, n607);
or   g1844 (n1581, n378, n265, n170, n572);
nand g1845 (n788, n382, n385, n218, n599);
nand g1846 (n987, n221, n398, n451, n186);
nor  g1847 (n1874, n354, n225, n290, n567);
and  g1848 (n1766, n224, n635, n646, n373);
nand g1849 (n902, n588, n277, n410, n331);
nand g1850 (n1533, n298, n397, n320, n550);
nor  g1851 (n1194, n664, n463, n394, n175);
and  g1852 (n733, n621, n661, n342, n520);
or   g1853 (n1403, n668, n423, n321, n623);
nor  g1854 (n704, n597, n366, n326, n381);
or   g1855 (n1068, n422, n239, n644, n491);
xnor g1856 (n1498, n202, n478, n381, n232);
or   g1857 (n1801, n555, n428, n271, n409);
or   g1858 (n721, n551, n566, n475, n558);
xnor g1859 (n1867, n297, n574, n256, n414);
nand g1860 (n1128, n554, n252, n349, n647);
nand g1861 (n1716, n656, n525, n577, n430);
nor  g1862 (n1629, n251, n636, n306, n479);
xor  g1863 (n1522, n394, n643, n445, n483);
nor  g1864 (n775, n302, n280, n573, n362);
xnor g1865 (n918, n469, n435, n509, n427);
nand g1866 (n1625, n645, n511, n497, n182);
nor  g1867 (n749, n253, n571, n575, n532);
nand g1868 (n1148, n244, n359, n258, n403);
nand g1869 (n905, n515, n377, n274, n408);
and  g1870 (n950, n241, n293, n376, n593);
xnor g1871 (n1799, n309, n316, n395, n594);
nand g1872 (n1950, n232, n597, n315, n601);
or   g1873 (n1234, n557, n352, n373, n449);
xnor g1874 (n1885, n568, n551, n654, n561);
nand g1875 (n892, n282, n526, n491, n598);
and  g1876 (n1481, n596, n483, n646, n509);
xnor g1877 (n1323, n436, n480, n632, n285);
nand g1878 (n1159, n611, n357, n420, n658);
and  g1879 (n1321, n499, n627, n456, n652);
xor  g1880 (n1826, n630, n565, n338, n244);
nor  g1881 (n1847, n452, n412, n489, n483);
nand g1882 (n735, n540, n284, n371, n610);
and  g1883 (n1450, n645, n595, n409, n485);
xnor g1884 (n1998, n321, n400, n441, n248);
xnor g1885 (n1907, n184, n307, n462, n512);
or   g1886 (n1483, n370, n305, n343, n280);
and  g1887 (n1060, n404, n488, n656, n629);
nand g1888 (n1694, n183, n603, n528, n346);
xor  g1889 (n1442, n415, n465, n459, n456);
xnor g1890 (n1274, n502, n382, n635, n387);
xor  g1891 (n1364, n196, n663, n165, n288);
and  g1892 (n1790, n351, n542, n431, n585);
nand g1893 (n1652, n527, n432, n164, n368);
or   g1894 (n1463, n533, n200, n522, n267);
xnor g1895 (n1215, n650, n213, n349, n524);
or   g1896 (n1760, n295, n491, n463, n608);
nor  g1897 (n1573, n511, n355, n360, n356);
or   g1898 (n1889, n400, n520, n173);
nand g1899 (n1019, n234, n602, n325, n536);
xor  g1900 (n1840, n553, n588, n336, n539);
and  g1901 (n849, n616, n412, n405, n538);
or   g1902 (n1036, n209, n624, n314, n258);
nor  g1903 (n804, n599, n253, n548, n171);
xor  g1904 (n1382, n264, n374, n517, n358);
xnor g1905 (n1240, n646, n476, n358, n345);
or   g1906 (n1478, n216, n269, n346, n487);
nand g1907 (n1618, n393, n564, n586, n579);
or   g1908 (n1495, n251, n391, n263, n494);
and  g1909 (n1034, n542, n453, n344, n551);
nor  g1910 (n1530, n361, n653, n516, n670);
nor  g1911 (n776, n214, n247, n571, n474);
or   g1912 (n1358, n360, n183, n506, n489);
nor  g1913 (n1596, n487, n408, n543, n462);
or   g1914 (n1963, n552, n202, n457, n307);
nand g1915 (n1022, n513, n291, n617, n506);
or   g1916 (n1177, n451, n387, n651, n223);
nor  g1917 (n1920, n378, n449, n426, n500);
and  g1918 (n999, n253, n616, n419, n383);
xor  g1919 (n1171, n454, n165, n193, n336);
xor  g1920 (n1227, n573, n507, n483, n469);
nor  g1921 (n771, n479, n245, n211, n191);
nor  g1922 (n868, n569, n519, n548, n468);
nor  g1923 (n1607, n340, n615, n456, n226);
nand g1924 (n1557, n205, n503, n317, n590);
and  g1925 (n961, n647, n206, n509, n385);
nand g1926 (n802, n488, n620, n265, n420);
and  g1927 (n1317, n664, n248, n635, n507);
or   g1928 (n857, n620, n471, n606, n534);
nor  g1929 (n965, n229, n303, n519, n260);
xor  g1930 (n1283, n521, n438, n171, n386);
or   g1931 (n1489, n659, n520, n270, n175);
nand g1932 (n1753, n252, n557, n658, n283);
or   g1933 (n875, n484, n245, n363, n444);
nand g1934 (n685, n287, n341, n181);
and  g1935 (n1821, n623, n607, n490, n250);
xnor g1936 (n951, n452, n601, n471, n442);
xnor g1937 (n1010, n255, n512, n398, n207);
nor  g1938 (n1332, n509, n656, n316, n471);
or   g1939 (n1536, n544, n299, n502, n200);
nand g1940 (n1764, n463, n447, n233, n625);
and  g1941 (n785, n261, n215, n304, n558);
nor  g1942 (n1243, n173, n225, n423, n200);
and  g1943 (n1810, n167, n301, n253, n559);
and  g1944 (n1451, n210, n469, n549, n323);
xor  g1945 (n926, n214, n318, n410, n219);
xor  g1946 (n1085, n653, n202, n174, n339);
and  g1947 (n1349, n630, n400, n179, n560);
nor  g1948 (n742, n336, n565, n533, n613);
nand g1949 (n1348, n365, n161, n477, n577);
nand g1950 (n1131, n584, n466, n489, n333);
and  g1951 (n707, n329, n628, n251, n243);
or   g1952 (n1064, n369, n262, n431, n280);
or   g1953 (n1682, n274, n192, n667, n188);
nor  g1954 (n1479, n167, n414, n477, n373);
or   g1955 (n798, n545, n608, n487, n589);
or   g1956 (n1523, n177, n328, n303, n438);
xor  g1957 (n1337, n411, n273, n337, n299);
and  g1958 (n1590, n593, n191, n315, n471);
xnor g1959 (n1738, n168, n301, n525, n197);
xnor g1960 (n764, n557, n228, n672, n649);
and  g1961 (n715, n593, n418, n617, n424);
nor  g1962 (n1408, n441, n378, n598, n358);
and  g1963 (n1079, n380, n314, n320, n418);
nand g1964 (n1484, n449, n255, n292, n225);
xor  g1965 (n1163, n404, n629, n238, n202);
and  g1966 (n1398, n315, n356, n606, n389);
and  g1967 (n1841, n475, n624, n328, n318);
xnor g1968 (n2044, n1209, n1572, n798, n1827);
and  g1969 (n2266, n1478, n1670, n825, n1539);
xnor g1970 (n2204, n1179, n1413, n995, n1464);
and  g1971 (n2029, n1503, n1565, n1567, n1162);
xor  g1972 (n2146, n1453, n1178, n1534, n1759);
xor  g1973 (n2123, n1530, n1546, n1094, n960);
xor  g1974 (n2034, n1270, n1438, n852, n943);
or   g1975 (n2223, n1292, n1786, n1247, n894);
or   g1976 (n2275, n836, n1961, n1314, n922);
or   g1977 (n2111, n1678, n992, n1493, n1665);
and  g1978 (n2103, n720, n1580, n1281, n1624);
or   g1979 (n2096, n1316, n1367, n858, n763);
and  g1980 (n2133, n1684, n1122, n1851, n1638);
nand g1981 (n2109, n1930, n1435, n1452, n1389);
nor  g1982 (n2256, n1507, n1707, n1123, n832);
or   g1983 (n2060, n1520, n1241, n1431, n1234);
or   g1984 (n2011, n1529, n1189, n1448, n1661);
xnor g1985 (n2216, n1754, n1199, n780, n953);
nor  g1986 (n2043, n849, n988, n1644, n1811);
xnor g1987 (n2086, n1005, n1817, n1057, n1602);
xor  g1988 (n2083, n1333, n1498, n865, n848);
nor  g1989 (n2226, n1901, n913, n1866, n1802);
nand g1990 (n2173, n991, n1111, n1711, n869);
nand g1991 (n2062, n1884, n1249, n944, n711);
and  g1992 (n2009, n1744, n1355, n1252, n1518);
nor  g1993 (n2042, n808, n1007, n1588, n1922);
and  g1994 (n2280, n1144, n1070, n1014, n1445);
xnor g1995 (n2220, n1324, n722, n1377, n1597);
nor  g1996 (n2193, n678, n1479, n1980, n1578);
and  g1997 (n2001, n1084, n1075, n1832, n1044);
xor  g1998 (n2228, n904, n1061, n1841, n1584);
xor  g1999 (n2162, n1698, n1917, n1517, n1787);
xnor g2000 (n2245, n1660, n1618, n1939, n1606);
nand g2001 (n2047, n1623, n876, n679, n1043);
xor  g2002 (n2237, n1193, n1248, n1040, n1873);
xor  g2003 (n2107, n1317, n1766, n1024, n774);
xor  g2004 (n2231, n854, n1370, n1978, n1336);
or   g2005 (n2268, n693, n1009, n1482, n1257);
xor  g2006 (n2023, n1164, n1916, n1476, n857);
nand g2007 (n2196, n835, n1018, n952, n1169);
nor  g2008 (n2113, n896, n1612, n1437, n1207);
xnor g2009 (n2142, n860, n1251, n1592, n1815);
xnor g2010 (n2312, n1415, n695, n1049, n961);
or   g2011 (n2063, n1835, n1447, n1614, n1474);
and  g2012 (n2329, n1158, n1829, n1900, n1228);
nand g2013 (n2313, n1533, n1635, n1284, n1214);
xnor g2014 (n2024, n885, n1959, n1451, n844);
xnor g2015 (n2296, n775, n866, n1219, n1163);
and  g2016 (n2189, n1538, n1659, n1000, n1818);
xnor g2017 (n2278, n1762, n1103, n814, n874);
and  g2018 (n2203, n1718, n1704, n989, n909);
or   g2019 (n2325, n704, n1908, n1372, n1975);
nand g2020 (n2240, n1771, n1120, n1840, n1570);
and  g2021 (n2045, n1646, n1082, n1450, n1677);
xor  g2022 (n2246, n700, n1921, n889, n1626);
nor  g2023 (n2031, n1760, n1573, n1710, n1366);
nor  g2024 (n2112, n1957, n1351, n1414, n958);
nor  g2025 (n2059, n939, n1194, n873, n915);
nand g2026 (n2138, n779, n727, n1204, n691);
or   g2027 (n2163, n681, n1941, n1583, n1537);
and  g2028 (n2014, n1839, n1637, n914, n1467);
and  g2029 (n2208, n1170, n1505, n1246, n1739);
and  g2030 (n2099, n1442, n1275, n893, n1266);
xnor g2031 (n2254, n1868, n1903, n1410, n937);
and  g2032 (n2180, n999, n1232, n1566, n1872);
and  g2033 (n2169, n1979, n1460, n1912, n1823);
nor  g2034 (n2274, n1937, n1862, n755, n1616);
nand g2035 (n2010, n1642, n1980, n1885, n1932);
or   g2036 (n2117, n1403, n956, n1106, n1648);
xnor g2037 (n2186, n1243, n1747, n1544, n1589);
nor  g2038 (n2127, n1608, n1807, n1871, n778);
xnor g2039 (n2027, n717, n1918, n1600, n701);
or   g2040 (n2057, n1320, n1831, n1462, n987);
or   g2041 (n2079, n1968, n767, n1850, n1655);
xor  g2042 (n2287, n1259, n1830, n1076, n1238);
nor  g2043 (n2035, n1757, n1188, n1065, n1221);
and  g2044 (n2140, n1004, n1748, n1949, n694);
xnor g2045 (n2055, n1662, n1774, n1631, n1001);
xor  g2046 (n2253, n1198, n1563, n1615, n1386);
nor  g2047 (n2302, n804, n1339, n1310, n965);
and  g2048 (n2230, n1195, n724, n930, n1081);
or   g2049 (n2082, n829, n903, n1318, n1233);
or   g2050 (n2007, n1155, n1323, n1935, n1115);
xnor g2051 (n2137, n1595, n1374, n846, n1861);
nor  g2052 (n2078, n737, n839, n1629, n1156);
and  g2053 (n2039, n1343, n1093, n813, n1109);
xor  g2054 (n2324, n1303, n1789, n1781, n1449);
xor  g2055 (n2006, n1132, n1373, n1965, n1387);
and  g2056 (n2319, n1694, n1581, n1315, n1041);
and  g2057 (n2234, n1847, n1056, n1060, n697);
xnor g2058 (n2104, n1913, n1879, n782, n1621);
nor  g2059 (n2143, n729, n1290, n1867, n1279);
nor  g2060 (n2328, n1693, n702, n1311, n1302);
xnor g2061 (n2244, n1053, n1039, n1376, n1636);
nor  g2062 (n2210, n747, n1669, n789, n982);
or   g2063 (n2314, n673, n1446, n1828, n1177);
nand g2064 (n2155, n713, n1149, n1721, n892);
or   g2065 (n2227, n1124, n1102, n1304, n1184);
xor  g2066 (n2281, n900, n1746, n1726, n1473);
nor  g2067 (n2272, n745, n1887, n1794, n902);
nand g2068 (n2264, n1671, n1855, n1480, n945);
xnor g2069 (n2070, n1955, n1231, n1481, n1441);
nor  g2070 (n2145, n1205, n794, n1015, n993);
nand g2071 (n2288, n833, n1118, n1213, n783);
and  g2072 (n2327, n1526, n1135, n1687, n1017);
and  g2073 (n2238, n1689, n1673, n1619, n1100);
and  g2074 (n2050, n1151, n879, n1816, n1808);
and  g2075 (n2105, n887, n1695, n1947, n1716);
xnor g2076 (n2075, n770, n1008, n827, n1819);
and  g2077 (n2202, n1294, n1427, n932, n1598);
nor  g2078 (n2051, n872, n1653, n1335, n683);
xor  g2079 (n2167, n877, n1552, n979, n1751);
nand g2080 (n2191, n1550, n1960, n1641, n1825);
nand g2081 (n2307, n1690, n1369, n1019, n751);
nor  g2082 (n2211, n1273, n1803, n1714, n1593);
nor  g2083 (n2236, n1574, n1215, n1489, n1801);
nand g2084 (n2129, n1944, n1782, n1559, n1838);
and  g2085 (n2094, n1525, n1657, n1679, n743);
nor  g2086 (n2091, n1392, n1891, n1634, n1826);
nor  g2087 (n2168, n1731, n740, n1737, n1658);
and  g2088 (n2089, n764, n1845, n1216, n963);
nor  g2089 (n2232, n1161, n1116, n1003, n1535);
and  g2090 (n2217, n1364, n1806, n1870, n1211);
or   g2091 (n2072, n1883, n1080, n1237, n812);
nor  g2092 (n2040, n1540, n1286, n1730, n1399);
nor  g2093 (n2156, n1814, n1033, n820, n1013);
nand g2094 (n2290, n1532, n799, n1006, n1777);
xnor g2095 (n2219, n1134, n1967, n1599, n976);
or   g2096 (n2157, n1601, n870, n1962, n969);
nor  g2097 (n2150, n1688, n1280, n924, n862);
xor  g2098 (n2225, n1190, n1976, n1911, n1795);
nor  g2099 (n2069, n1647, n1604, n1088, n1072);
and  g2100 (n2110, n689, n710, n1531, n1129);
and  g2101 (n2025, n1021, n921, n905, n1051);
xor  g2102 (n2098, n1380, n1296, n1098, n1105);
nand g2103 (n2126, n971, n1728, n1383, n1743);
or   g2104 (n2071, n1812, n749, n1749, n756);
xor  g2105 (n2002, n1035, n1756, n954, n1542);
nor  g2106 (n2174, n1332, n821, n1338, n1236);
xnor g2107 (n2182, n1331, n1894, n1632, n1078);
xor  g2108 (n2222, n1528, n1143, n1192, n935);
xor  g2109 (n2299, n1675, n1723, n803, n1267);
xor  g2110 (n2181, n1220, n1888, n1471, n883);
nor  g2111 (n2068, n941, n1416, n1404, n1208);
nor  g2112 (n2291, n1804, n986, n1863, n1287);
nand g2113 (n2198, n781, n1548, n1262, n1980);
or   g2114 (n2255, n1150, n1258, n1717, n769);
nand g2115 (n2165, n1643, n951, n1755, n1650);
xor  g2116 (n2056, n1740, n1180, n1274, n1649);
nand g2117 (n2304, n1627, n705, n1224, n1764);
or   g2118 (n2317, n746, n1406, n984, n1036);
xnor g2119 (n2295, n1893, n1363, n1842, n738);
and  g2120 (n2183, n1068, n1767, n1395, n1114);
xor  g2121 (n2205, n1240, n1409, n1099, n1904);
or   g2122 (n2085, n1761, n1854, n1981, n1126);
xor  g2123 (n2012, n907, n851, n1725, n1974);
or   g2124 (n2251, n1864, n807, n1433, n977);
nor  g2125 (n2270, n970, n706, n1268, n739);
nor  g2126 (n2252, n1313, n1073, n1133, n1899);
nand g2127 (n2124, n882, n1172, n1645, n1485);
or   g2128 (n2207, n1843, n1973, n1742, n785);
or   g2129 (n2073, n1769, n1472, n1463, n1852);
xor  g2130 (n2139, n1562, n981, n997, n1860);
and  g2131 (n2215, n1720, n819, n1536, n1368);
or   g2132 (n2195, n933, n1419, n1349, n1074);
or   g2133 (n2233, n806, n1651, n1500, n842);
nand g2134 (n2271, n1085, n1022, n791, n1859);
xor  g2135 (n2257, n1605, n1326, n1587, n1128);
xor  g2136 (n2077, n853, n1800, n1964, n1953);
nand g2137 (n2032, n1420, n1308, n1954, n1483);
xor  g2138 (n2022, n1052, n1895, n897, n1793);
xnor g2139 (n2214, n1226, n1067, n1722, n910);
xnor g2140 (n2286, n890, n1966, n1175, n1622);
or   g2141 (n2316, n1182, n1491, n1681, n1344);
xnor g2142 (n2020, n1365, n823, n957, n831);
nand g2143 (n2200, n1950, n974, n1522, n1502);
xnor g2144 (n2037, n1579, n1173, n1187, n1138);
or   g2145 (n2017, n1271, n1285, n966, n1712);
xnor g2146 (n2178, n1112, n736, n888, n899);
nand g2147 (n2164, n837, n809, n1853, n1735);
nor  g2148 (n2283, n1582, n838, n1347, n1924);
or   g2149 (n2321, n1300, n1734, n1168, n801);
xor  g2150 (n2260, n1719, n765, n1822, n761);
and  g2151 (n2176, n934, n855, n1920, n1063);
and  g2152 (n2041, n949, n1979, n1560, n843);
and  g2153 (n2248, n1079, n1557, n692, n677);
xor  g2154 (n2090, n1683, n817, n1486, n891);
or   g2155 (n2267, n690, n1283, n919, n1200);
nand g2156 (n2289, n1506, n1443, n1496, n1145);
and  g2157 (n2005, n723, n1301, n1524, n1527);
xnor g2158 (n2261, n1288, n1110, n1071, n712);
nor  g2159 (n2128, n1979, n675, n1512, n1424);
xor  g2160 (n2159, n867, n1104, n850, n1325);
nand g2161 (n2201, n1571, n1197, n1701, n1312);
xnor g2162 (n2221, n1554, n1946, n1685, n1352);
or   g2163 (n2134, n1309, n841, n1772, n1466);
nand g2164 (n2301, n1152, n926, n1709, n967);
and  g2165 (n2116, n1390, n1136, n1405, n1391);
nand g2166 (n2015, n1328, n1425, n1378, n1291);
xor  g2167 (n2004, n1833, n1508, n1576, n916);
xor  g2168 (n2106, n1858, n1628, n1551, n1773);
nor  g2169 (n2131, n1421, n1484, n901, n1456);
xor  g2170 (n2065, n1558, n1255, n1130, n1715);
and  g2171 (n2054, n1032, n1875, n1012, n1590);
nor  g2172 (n2269, n1620, n962, n797, n1222);
nand g2173 (n2262, n1069, n1191, n787, n1147);
nor  g2174 (n2118, n884, n1201, n1203, n748);
xor  g2175 (n2019, n918, n906, n1890, n1159);
or   g2176 (n2120, n1045, n776, n777, n1881);
nand g2177 (n2038, n1330, n1971, n1350, n1160);
xor  g2178 (n2209, n1613, n1357, n1936, n1514);
nand g2179 (n2213, n1568, n950, n1091, n676);
nor  g2180 (n2311, n1821, n1768, n1097, n1384);
and  g2181 (n2152, n753, n815, n1305, n1837);
and  g2182 (n2309, n696, n1824, n1820, n1210);
and  g2183 (n2276, n699, n1692, n948, n1902);
nor  g2184 (n2258, n1107, n1663, n1030, n1470);
xnor g2185 (n2076, n680, n1411, n955, n1555);
nand g2186 (n2166, n1519, n1412, n1938, n1245);
xnor g2187 (n2095, n1277, n1633, n1849, n1250);
or   g2188 (n2305, n1142, n714, n1148, n1702);
nand g2189 (n2016, n1298, n1515, n1477, n1680);
xnor g2190 (n2293, n750, n1440, n1418, n1603);
or   g2191 (n2100, n1121, n1023, n1549, n1092);
nand g2192 (n2320, n1906, n1058, n1927, n1055);
nor  g2193 (n2241, n1289, n1732, n1956, n990);
and  g2194 (n2066, n733, n1455, n1223, n875);
xor  g2195 (n2292, n1886, n1066, n1086, n1029);
xor  g2196 (n2303, n1738, n959, n1137, n1796);
nand g2197 (n2101, n1329, n1117, n1458, n1423);
and  g2198 (n2087, n886, n1108, n1494, n1062);
nor  g2199 (n2048, n1297, n1083, n1654, n1753);
xor  g2200 (n2185, n1909, n1388, n1230, n1358);
nor  g2201 (n2018, n1054, n1541, n1846, n1729);
and  g2202 (n2141, n1708, n1877, n1026, n1575);
or   g2203 (n2080, n1356, n1461, n1907, n826);
xnor g2204 (n2074, n792, n830, n1171, n1706);
and  g2205 (n2323, n1218, n1269, n726, n1596);
nand g2206 (n2279, n674, n1703, n1434, n1011);
and  g2207 (n2160, n762, n1361, n1556, n793);
and  g2208 (n2218, n1242, n1244, n1475, n911);
and  g2209 (n2277, n1783, n1394, n1027, n1282);
xnor g2210 (n2239, n752, n1454, n1400, n1038);
xnor g2211 (n2148, n1235, n1096, n1016, n1432);
nand g2212 (n2121, n1487, n1047, n1790, n947);
or   g2213 (n2058, n732, n1031, n1969, n1865);
xnor g2214 (n2310, n1509, n1342, n1928, n1700);
xor  g2215 (n2297, n928, n1492, n1345, n861);
or   g2216 (n2318, n1141, n1140, n1457, n1696);
nor  g2217 (n2028, n1942, n1724, n1625, n1183);
xor  g2218 (n2053, n1272, n920, n734, n925);
and  g2219 (n2224, n1146, n1025, n1630, n1306);
and  g2220 (n2194, n824, n1260, n1253, n1382);
nand g2221 (n2308, n1553, n1157, n1951, n1354);
xor  g2222 (n2114, n1153, n929, n728, n1341);
and  g2223 (n2179, n1254, n1741, n721, n796);
xor  g2224 (n2115, n766, n1577, n1119, n685);
or   g2225 (n2153, n1504, n1664, n1101, n1265);
xnor g2226 (n2026, n1915, n708, n816, n1892);
xnor g2227 (n2263, n1809, n759, n978, n828);
or   g2228 (n2013, n946, n1176, n1276, n709);
nand g2229 (n2197, n1836, n834, n682, n1439);
nor  g2230 (n2250, n1674, n1792, n1799, n725);
nand g2231 (n2284, n1561, n1417, n1206, n985);
nor  g2232 (n2132, n1334, n1385, n1952, n1977);
xnor g2233 (n2172, n686, n1958, n1095, n1307);
and  g2234 (n2188, n1293, n1401, n760, n1779);
xnor g2235 (n2125, n1186, n908, n1666, n1497);
nand g2236 (n2190, n917, n1020, n859, n1727);
or   g2237 (n2322, n730, n938, n703, n1940);
or   g2238 (n2298, n1778, n1090, n1691, n1407);
nand g2239 (n2235, n1943, n1784, n1926, n1002);
or   g2240 (n2170, n927, n931, n1791, n1776);
xor  g2241 (n2171, n840, n912, n880, n1933);
xnor g2242 (n2064, n1174, n1640, n744, n1857);
or   g2243 (n2184, n1980, n1087, n1181, n1459);
xor  g2244 (n2247, n1844, n1125, n1880, n1263);
nor  g2245 (n2052, n1131, n1426, n1089, n1750);
xor  g2246 (n2084, n972, n1611, n1225, n1428);
and  g2247 (n2243, n1037, n1185, n898, n1963);
and  g2248 (n2021, n1765, n1878, n1758, n1511);
xor  g2249 (n2144, n847, n998, n1705, n1166);
or   g2250 (n2061, n1501, n1770, n1656, n895);
xnor g2251 (n2265, n1429, n1034, n1934, n1353);
and  g2252 (n2242, n1914, n1697, n1585, n1212);
nor  g2253 (n2326, n1510, n784, n715, n1543);
xnor g2254 (n2097, n758, n1848, n1699, n1397);
or   g2255 (n2212, n964, n1064, n771, n1436);
nand g2256 (n2136, n735, n800, n1780, n1594);
nand g2257 (n2003, n1227, n1929, n1586, n1805);
or   g2258 (n2033, n1396, n1381, n786, n881);
xnor g2259 (n2300, n1813, n1889, n802, n1925);
nand g2260 (n2030, n1046, n994, n1010, n1444);
and  g2261 (n2081, n1970, n996, n1468, n878);
nand g2262 (n2008, n1547, n1322, n741, n1229);
nand g2263 (n2315, n716, n772, n1059, n1874);
or   g2264 (n2036, n845, n1337, n1202, n1763);
xor  g2265 (n2119, n1856, n1910, n871, n973);
nor  g2266 (n2206, n707, n1798, n1785, n810);
nand g2267 (n2147, n1617, n1398, n788, n698);
nand g2268 (n2049, n1256, n805, n1490, n936);
and  g2269 (n2175, n1261, n1672, n1028, n1465);
and  g2270 (n2154, n1713, n1499, n1050, n1408);
and  g2271 (n2092, n1591, n1834, n757, n1360);
xnor g2272 (n2199, n1521, n1048, n684, n942);
or   g2273 (n2192, n1327, n1513, n1686, n811);
xnor g2274 (n2135, n1775, n1676, n1402, n868);
xnor g2275 (n2273, n1264, n795, n923, n1393);
xnor g2276 (n2102, n1609, n1898, n719, n1897);
nor  g2277 (n2282, n968, n1165, n1869, n1810);
nor  g2278 (n2088, n1167, n1077, n1422, n1564);
xor  g2279 (n2294, n1154, n1196, n1797, n1488);
and  g2280 (n2149, n1545, n1295, n1340, n1348);
xnor g2281 (n2187, n1876, n1919, n1569, n1375);
and  g2282 (n2130, n940, n1359, n742, n1745);
or   g2283 (n2108, n1923, n1981, n1607, n983);
and  g2284 (n2259, n731, n1042, n1319, n1239);
or   g2285 (n2177, n1752, n856, n1127, n1321);
nand g2286 (n2229, n864, n687, n1788, n1217);
xnor g2287 (n2249, n1278, n1882, n980, n1652);
nor  g2288 (n2306, n768, n1733, n688, n1736);
nor  g2289 (n2161, n1945, n1668, n863, n818);
nor  g2290 (n2046, n1495, n1948, n773, n1371);
nor  g2291 (n2067, n1523, n1905, n1516, n1299);
nand g2292 (n2158, n1362, n1931, n790, n1972);
and  g2293 (n2122, n822, n975, n1430, n1346);
or   g2294 (n2285, n1979, n1113, n1379, n1896);
xnor g2295 (n2093, n1139, n718, n1682, n1469);
nor  g2296 (n2151, n1639, n1610, n1667, n754);
nor  g2297 (n2347, n2029, n2064, n2061, n2007);
and  g2298 (n2331, n2020, n2042, n2001, n2024);
xnor g2299 (n2342, n2002, n2019, n2047, n2023);
and  g2300 (n2340, n2062, n2026, n2022, n2015);
nand g2301 (n2345, n2030, n2006, n2065, n2021);
nor  g2302 (n2339, n2027, n2033, n2014, n2057);
xor  g2303 (n2337, n2036, n2011, n2005, n2016);
xor  g2304 (n2334, n2025, n2009, n2017, n2041);
nor  g2305 (n2333, n2028, n2039, n2051, n2068);
nor  g2306 (n2330, n2004, n2060, n2066, n2071);
and  g2307 (n2332, n2059, n2018, n2037, n2013);
and  g2308 (n2343, n2040, n2045, n2046, n2058);
xor  g2309 (n2344, n2048, n2053, n2070, n2034);
and  g2310 (n2346, n2049, n2044, n2031, n2055);
or   g2311 (n2336, n2056, n2050, n2063, n2038);
xnor g2312 (n2335, n2069, n2072, n2067, n2054);
or   g2313 (n2341, n2032, n2010, n2008, n2003);
nor  g2314 (n2338, n2035, n2012, n2052, n2043);
buf  g2315 (n2357, n2339);
buf  g2316 (n2362, n2334);
buf  g2317 (n2351, n2337);
not  g2318 (n2353, n2341);
buf  g2319 (n2356, n2338);
buf  g2320 (n2354, n2345);
not  g2321 (n2364, n2333);
not  g2322 (n2363, n2336);
buf  g2323 (n2352, n2331);
not  g2324 (n2359, n2346);
buf  g2325 (n2355, n2342);
buf  g2326 (n2360, n2330);
not  g2327 (n2361, n2340);
buf  g2328 (n2348, n2332);
buf  g2329 (n2358, n2344);
buf  g2330 (n2350, n2335);
buf  g2331 (n2349, n2343);
nand g2332 (n2365, n2354, n2361, n2349);
nor  g2333 (n2367, n2357, n2349, n2363);
xor  g2334 (n2377, n2359, n2352, n2361, n2364);
xor  g2335 (n2383, n1982, n1982, n2361, n2353);
xor  g2336 (n2380, n2350, n1982, n2360, n2357);
xor  g2337 (n2378, n2348, n2358, n2350, n2354);
and  g2338 (n2371, n2360, n2351, n2355, n2357);
and  g2339 (n2373, n2355, n1981, n2363, n2360);
xnor g2340 (n2374, n2358, n2351, n2357, n2364);
nand g2341 (n2375, n2351, n2359, n2362);
and  g2342 (n2366, n2350, n1981, n2348, n2356);
xnor g2343 (n2369, n2364, n2352, n2354);
nand g2344 (n2382, n2353, n2356, n2355);
and  g2345 (n2372, n2361, n2363, n2355, n2348);
or   g2346 (n2381, n2350, n2358, n2349);
or   g2347 (n2370, n2358, n2364, n2352, n2360);
or   g2348 (n2376, n1982, n2348, n2351, n2362);
nand g2349 (n2379, n2363, n2356, n2353);
and  g2350 (n2368, n2354, n2359, n2362);
nand g2351 (n2391, n2080, n2091, n2076, n2374);
nor  g2352 (n2385, n2382, n2082, n2093, n2381);
and  g2353 (n2393, n2073, n2078, n2090, n2086);
xor  g2354 (n2384, n2378, n2095, n2097, n2099);
nor  g2355 (n2390, n2101, n2075, n2085, n2077);
and  g2356 (n2392, n2081, n2379, n2098, n2088);
and  g2357 (n2387, n2074, n2377, n2380, n2100);
xor  g2358 (n2386, n2087, n2084, n2094, n2092);
or   g2359 (n2389, n2375, n2089, n2083, n2079);
or   g2360 (n2388, n2102, n2096, n2383, n2376);
not  g2361 (n2395, n2386);
buf  g2362 (n2396, n2387);
or   g2363 (n2394, n2385, n2388, n2389, n2384);
and  g2364 (n2397, n2395, n2394, n2396);
nand g2365 (n2399, n2104, n2107, n2105, n2106);
xor  g2366 (n2398, n2397, n2397, n2108, n2103);
or   g2367 (n2400, n2109, n2398);
nor  g2368 (n2401, n2400, n2113, n2110, n2118);
xnor g2369 (n2404, n2115, n2112, n2111, n2400);
xor  g2370 (n2403, n2121, n2400, n2116, n2120);
nand g2371 (n2402, n2119, n2114, n2117, n2400);
buf  g2372 (n2406, n2402);
not  g2373 (n2408, n2403);
not  g2374 (n2410, n2401);
not  g2375 (n2405, n2403);
buf  g2376 (n2411, n2404);
buf  g2377 (n2407, n2404);
buf  g2378 (n2412, n2404);
buf  g2379 (n2409, n2404);
not  g2380 (n2419, n2405);
not  g2381 (n2414, n2409);
not  g2382 (n2436, n2410);
not  g2383 (n2431, n2406);
not  g2384 (n2415, n2390);
buf  g2385 (n2432, n2407);
buf  g2386 (n2428, n2407);
not  g2387 (n2437, n2409);
buf  g2388 (n2427, n2399);
not  g2389 (n2439, n2412);
not  g2390 (n2425, n2407);
buf  g2391 (n2423, n2406);
not  g2392 (n2435, n2407);
buf  g2393 (n2421, n2391);
not  g2394 (n2417, n2411);
buf  g2395 (n2416, n2405);
not  g2396 (n2440, n2398);
not  g2397 (n2420, n2409);
not  g2398 (n2434, n2412);
not  g2399 (n2426, n2406);
buf  g2400 (n2430, n2405);
buf  g2401 (n2413, n2411);
buf  g2402 (n2438, n2408);
nand g2403 (n2418, n2410, n2398);
or   g2404 (n2433, n2408, n2391, n2406, n2410);
nand g2405 (n2424, n2408, n2391, n2392);
nand g2406 (n2422, n2410, n2408, n2412);
xnor g2407 (n2429, n2405, n2411, n2409);
buf  g2408 (n2481, n2435);
buf  g2409 (n2480, n2125);
buf  g2410 (n2493, n2439);
not  g2411 (n2447, n2414);
buf  g2412 (n2497, n2426);
buf  g2413 (n2474, n2419);
buf  g2414 (n2518, n2421);
buf  g2415 (n2517, n2422);
buf  g2416 (n2472, n2433);
not  g2417 (n2492, n2413);
buf  g2418 (n2543, n2432);
not  g2419 (n2441, n2436);
buf  g2420 (n2530, n2433);
not  g2421 (n2473, n2424);
not  g2422 (n2531, n2426);
not  g2423 (n2506, n2424);
buf  g2424 (n2535, n2431);
buf  g2425 (n2479, n2438);
buf  g2426 (n2522, n2439);
not  g2427 (n2507, n2440);
not  g2428 (n2508, n2418);
not  g2429 (n2446, n2428);
not  g2430 (n2483, n2422);
buf  g2431 (n2548, n2123);
buf  g2432 (n2490, n2424);
buf  g2433 (n2444, n2437);
not  g2434 (n2516, n2427);
buf  g2435 (n2505, n2416);
not  g2436 (n2503, n2415);
not  g2437 (n2460, n2440);
buf  g2438 (n2526, n2429);
not  g2439 (n2527, n2425);
not  g2440 (n2540, n2429);
not  g2441 (n2450, n2435);
buf  g2442 (n2538, n2392);
not  g2443 (n2524, n2431);
not  g2444 (n2521, n2435);
buf  g2445 (n2495, n2427);
buf  g2446 (n2512, n2416);
buf  g2447 (n2510, n2432);
buf  g2448 (n2455, n2430);
buf  g2449 (n2536, n2431);
not  g2450 (n2457, n2393);
buf  g2451 (n2443, n2124);
buf  g2452 (n2477, n2424);
not  g2453 (n2542, n2423);
not  g2454 (n2486, n2416);
not  g2455 (n2546, n2438);
not  g2456 (n2551, n2428);
not  g2457 (n2476, n2126);
buf  g2458 (n2514, n2393);
not  g2459 (n2488, n2415);
not  g2460 (n2501, n2435);
buf  g2461 (n2547, n2414);
buf  g2462 (n2498, n2431);
buf  g2463 (n2494, n2427);
buf  g2464 (n2537, n2135);
not  g2465 (n2484, n2134);
buf  g2466 (n2504, n2439);
not  g2467 (n2520, n2437);
buf  g2468 (n2502, n2413);
not  g2469 (n2519, n2422);
not  g2470 (n2545, n2426);
not  g2471 (n2452, n2432);
not  g2472 (n2552, n2393);
buf  g2473 (n2467, n2392);
buf  g2474 (n2549, n2392);
buf  g2475 (n2513, n2421);
buf  g2476 (n2499, n2415);
buf  g2477 (n2482, n2122);
not  g2478 (n2449, n2418);
buf  g2479 (n2509, n2430);
not  g2480 (n2534, n2438);
not  g2481 (n2464, n2127);
buf  g2482 (n2475, n2416);
not  g2483 (n2462, n2423);
buf  g2484 (n2539, n2429);
buf  g2485 (n2525, n2434);
not  g2486 (n2456, n2128);
not  g2487 (n2541, n2137);
not  g2488 (n2478, n2417);
buf  g2489 (n2511, n2413);
buf  g2490 (n2469, n2138);
buf  g2491 (n2468, n2419);
not  g2492 (n2515, n2422);
not  g2493 (n2459, n2430);
not  g2494 (n2465, n2417);
buf  g2495 (n2487, n2434);
buf  g2496 (n2550, n2428);
not  g2497 (n2448, n2425);
buf  g2498 (n2442, n2437);
not  g2499 (n2529, n2419);
not  g2500 (n2451, n2429);
not  g2501 (n2485, n2136);
buf  g2502 (n2453, n2420);
buf  g2503 (n2533, n2421);
not  g2504 (n2496, n2420);
buf  g2505 (n2470, n2433);
buf  g2506 (n2445, n2129);
not  g2507 (n2466, n2420);
buf  g2508 (n2471, n2133);
not  g2509 (n2458, n2425);
buf  g2510 (n2461, n2434);
buf  g2511 (n2489, n2436);
nand g2512 (n2532, n2413, n2439, n2428, n2414);
xnor g2513 (n2500, n2426, n2436, n2440, n2415);
nor  g2514 (n2544, n2418, n2433, n2434, n2130);
nand g2515 (n2523, n2418, n2423, n2437, n2432);
nand g2516 (n2491, n2417, n2393, n2440, n2438);
or   g2517 (n2463, n2436, n2420, n2430, n2423);
xor  g2518 (n2454, n2417, n2414, n2427, n2425);
and  g2519 (n2528, n2419, n2131, n2421, n2132);
nand g2520 (n2560, n2483, n2454, n2459, n2481);
and  g2521 (n2566, n2484, n2462, n2492, n2447);
xor  g2522 (n2555, n2139, n2451, n2491, n2478);
or   g2523 (n2564, n2472, n2479, n2453, n2445);
xor  g2524 (n2557, n2450, n2482, n2455, n2465);
xor  g2525 (n2554, n2458, n2456, n2446, n2477);
nor  g2526 (n2558, n2489, n2448, n2441, n2449);
nor  g2527 (n2563, n2485, n2490, n2488, n2140);
nor  g2528 (n2561, n2468, n2467, n2463, n2487);
xor  g2529 (n2562, n2141, n2443, n2470, n2475);
nand g2530 (n2556, n2480, n2452, n2457, n2474);
nor  g2531 (n2565, n2469, n2444, n2476, n2442);
nand g2532 (n2559, n2493, n2473, n2464, n2460);
or   g2533 (n2553, n2461, n2466, n2486, n2471);
or   g2534 (n2568, n2146, n2553, n2144);
or   g2535 (n2569, n2555, n2143, n2556);
or   g2536 (n2567, n2142, n2145, n2147, n2554);
not  g2537 (n2575, n2568);
not  g2538 (n2576, n2153);
not  g2539 (n2571, n2148);
not  g2540 (n2570, n2569);
not  g2541 (n2572, n2154);
xor  g2542 (n2574, n2569, n2568);
and  g2543 (n2577, n2149, n2569, n2152, n2150);
or   g2544 (n2573, n2568, n2567, n2151, n2155);
buf  g2545 (n2594, n2522);
buf  g2546 (n2581, n2571);
buf  g2547 (n2593, n2531);
not  g2548 (n2588, n2572);
not  g2549 (n2609, n2507);
not  g2550 (n2608, n2573);
buf  g2551 (n2585, n2539);
buf  g2552 (n2579, n2542);
buf  g2553 (n2590, n2512);
buf  g2554 (n2606, n2499);
buf  g2555 (n2600, n2545);
buf  g2556 (n2592, n2495);
buf  g2557 (n2582, n2504);
xnor g2558 (n2589, n2570, n2572);
nand g2559 (n2595, n2547, n2508, n2510, n2156);
and  g2560 (n2602, n2527, n2540, n2544, n2529);
or   g2561 (n2586, n2538, n2574, n2530, n2575);
nand g2562 (n2584, n2571, n2546, n2535, n2518);
or   g2563 (n2587, n2505, n2571, n2576, n2528);
nand g2564 (n2601, n2496, n2494, n2525, n2533);
xnor g2565 (n2597, n2575, n2541, n2506, n2577);
xnor g2566 (n2605, n2570, n2576, n2517, n2501);
xor  g2567 (n2607, n2577, n2576, n2574);
nand g2568 (n2583, n2524, n2577, n2570, n2498);
xor  g2569 (n2596, n2534, n2570, n2521, n2537);
or   g2570 (n2603, n2519, n2526, n2575, n2516);
and  g2571 (n2598, n2509, n2520, n2577, n2497);
xor  g2572 (n2578, n2511, n2572, n2575, n2573);
xnor g2573 (n2599, n2543, n2576, n2536, n2572);
nor  g2574 (n2580, n2513, n2532, n2573, n2515);
or   g2575 (n2604, n2502, n2523, n2571, n2573);
xor  g2576 (n2591, n2574, n2500, n2503, n2514);
not  g2577 (n2613, n2599);
buf  g2578 (n2644, n2601);
buf  g2579 (n2611, n2589);
not  g2580 (n2629, n2583);
not  g2581 (n2618, n2583);
buf  g2582 (n2630, n2560);
buf  g2583 (n2627, n2590);
buf  g2584 (n2615, n2584);
buf  g2585 (n2631, n2399);
buf  g2586 (n2647, n2559);
buf  g2587 (n2621, n2563);
not  g2588 (n2637, n2592);
not  g2589 (n2658, n2562);
buf  g2590 (n2617, n2599);
not  g2591 (n2641, n2588);
buf  g2592 (n2620, n2564);
buf  g2593 (n2640, n2605);
or   g2594 (n2638, n2599, n2582, n2587, n2564);
nor  g2595 (n2628, n2605, n2607, n2609, n2601);
xnor g2596 (n2636, n2583, n2580, n2603, n2591);
xor  g2597 (n2653, n2579, n2597, n2590, n2588);
xor  g2598 (n2633, n2562, n2563, n2604, n2583);
xor  g2599 (n2650, n2593, n2592, n2582, n2608);
xnor g2600 (n2625, n2596, n2607, n2580, n2565);
nor  g2601 (n2632, n2606, n2595, n2157, n2581);
or   g2602 (n2643, n2582, n2399, n2609, n2590);
nand g2603 (n2649, n2578, n2586, n2600, n2609);
xor  g2604 (n2623, n2580, n2598, n2589, n2594);
xor  g2605 (n2610, n2588, n2601, n2562, n2580);
and  g2606 (n2642, n2594, n2594, n2586, n2585);
nand g2607 (n2635, n2585, n2588, n2598, n2591);
xor  g2608 (n2646, n2600, n2605, n2596);
xnor g2609 (n2659, n2581, n2603, n2584, n2604);
or   g2610 (n2624, n2606, n2579, n2561, n2600);
nor  g2611 (n2634, n2599, n2602, n2579, n2587);
xor  g2612 (n2660, n2584, n2593, n2587, n2591);
nand g2613 (n2616, n2585, n2585, n2587, n2607);
nor  g2614 (n2622, n2606, n2595, n2608, n2563);
xnor g2615 (n2626, n2602, n2597, n2578);
nand g2616 (n2645, n2581, n2564, n2609, n2565);
nor  g2617 (n2612, n2592, n2564, n2602, n2595);
xnor g2618 (n2652, n2582, n2600, n2603, n2563);
xnor g2619 (n2619, n2596, n2598, n2581, n2595);
xor  g2620 (n2651, n2603, n2604, n2606, n2586);
and  g2621 (n2614, n2592, n2601, n2565, n2589);
xor  g2622 (n2657, n2607, n2562, n2561, n2591);
or   g2623 (n2655, n2584, n2590, n2604, n2598);
nor  g2624 (n2654, n2558, n2594, n2608, n2579);
nor  g2625 (n2648, n2586, n2578, n2605, n2557);
xnor g2626 (n2639, n2399, n2589, n2593, n2602);
xnor g2627 (n2656, n2597, n2608, n2578, n2593);
not  g2628 (n2666, n2613);
buf  g2629 (n2664, n2620);
buf  g2630 (n2673, n2160);
not  g2631 (n2668, n2619);
not  g2632 (n2669, n2612);
buf  g2633 (n2662, n2610);
buf  g2634 (n2663, n2615);
not  g2635 (n2672, n2622);
buf  g2636 (n2665, n2616);
not  g2637 (n2670, n2614);
nand g2638 (n2661, n2159, n2618);
nor  g2639 (n2667, n2611, n2621);
xnor g2640 (n2671, n2158, n2617);
xor  g2641 (n2683, n2662, n2667);
and  g2642 (n2678, n2661, n2551);
or   g2643 (n2686, n2161, n2664);
nand g2644 (n2675, n2672, n2550);
xnor g2645 (n2684, n2549, n2673);
xor  g2646 (n2682, n2164, n2668);
xor  g2647 (n2680, n2672, n2669);
or   g2648 (n2677, n2162, n2165);
xor  g2649 (n2685, n2673, n2671);
and  g2650 (n2681, n2663, n2548);
xor  g2651 (n2687, n2665, n2670);
xor  g2652 (n2679, n2163, n2672);
nand g2653 (n2674, n2666, n2673);
xor  g2654 (n2676, n2672, n2673);
not  g2655 (n2728, n2683);
not  g2656 (n2727, n2682);
not  g2657 (n2708, n2679);
buf  g2658 (n2734, n2685);
buf  g2659 (n2721, n2676);
not  g2660 (n2711, n2681);
buf  g2661 (n2720, n2675);
not  g2662 (n2692, n2687);
not  g2663 (n2690, n2684);
buf  g2664 (n2696, n2679);
buf  g2665 (n2706, n2680);
buf  g2666 (n2715, n2683);
not  g2667 (n2737, n2681);
buf  g2668 (n2731, n2674);
buf  g2669 (n2729, n2166);
buf  g2670 (n2716, n2681);
not  g2671 (n2693, n2687);
buf  g2672 (n2701, n2167);
buf  g2673 (n2697, n2173);
not  g2674 (n2733, n2686);
not  g2675 (n2712, n2675);
not  g2676 (n2695, n2678);
not  g2677 (n2714, n2679);
not  g2678 (n2699, n2685);
buf  g2679 (n2704, n2684);
buf  g2680 (n2724, n2680);
not  g2681 (n2691, n2687);
not  g2682 (n2698, n2684);
not  g2683 (n2688, n2680);
buf  g2684 (n2707, n2675);
buf  g2685 (n2694, n2677);
not  g2686 (n2705, n2685);
not  g2687 (n2742, n2677);
buf  g2688 (n2703, n2676);
not  g2689 (n2740, n2678);
not  g2690 (n2725, n2686);
buf  g2691 (n2689, n2686);
buf  g2692 (n2726, n2679);
buf  g2693 (n2730, n2687);
not  g2694 (n2722, n2683);
not  g2695 (n2735, n2168);
not  g2696 (n2717, n2682);
not  g2697 (n2738, n2682);
buf  g2698 (n2743, n2170);
buf  g2699 (n2719, n2677);
buf  g2700 (n2718, n2686);
not  g2701 (n2713, n2674);
not  g2702 (n2741, n2683);
and  g2703 (n2700, n2680, n2682);
xnor g2704 (n2709, n2677, n2681);
and  g2705 (n2702, n2171, n2169);
not  g2706 (n2736, n2676);
and  g2707 (n2723, n2685, n2675);
buf  g2708 (n2739, n2678);
xnor g2709 (n2732, n2684, n2172);
buf  g2710 (n2710, n2674);
not  g2711 (n2764, n2688);
not  g2712 (n2851, n2712);
not  g2713 (n2834, n2723);
buf  g2714 (n2887, n2637);
not  g2715 (n2759, n2702);
buf  g2716 (n2778, n2728);
buf  g2717 (n2844, n2702);
not  g2718 (n2782, n2645);
not  g2719 (n2817, n2638);
not  g2720 (n2772, n2700);
not  g2721 (n2805, n2695);
buf  g2722 (n2830, n2716);
not  g2723 (n2761, n2731);
not  g2724 (n2824, n2715);
buf  g2725 (n2754, n2742);
not  g2726 (n2857, n2741);
not  g2727 (n2791, n2706);
buf  g2728 (n2871, n2566);
buf  g2729 (n2746, n2711);
buf  g2730 (n2836, n2705);
buf  g2731 (n2813, n2702);
not  g2732 (n2804, n2725);
not  g2733 (n2823, n2629);
buf  g2734 (n2802, n2735);
buf  g2735 (n2783, n2727);
not  g2736 (n2766, n2722);
not  g2737 (n2765, n2728);
not  g2738 (n2849, n2723);
not  g2739 (n2771, n2727);
buf  g2740 (n2841, n2691);
buf  g2741 (n2884, n2732);
not  g2742 (n2889, n2741);
buf  g2743 (n2758, n2690);
buf  g2744 (n2837, n2734);
buf  g2745 (n2864, n2566);
not  g2746 (n2763, n2701);
buf  g2747 (n2770, n2719);
not  g2748 (n2838, n2656);
not  g2749 (n2752, n2730);
buf  g2750 (n2774, n2659);
not  g2751 (n2788, n2690);
not  g2752 (n2888, n2636);
not  g2753 (n2881, n2729);
not  g2754 (n2747, n2728);
buf  g2755 (n2876, n2727);
buf  g2756 (n2756, n2738);
not  g2757 (n2828, n2704);
not  g2758 (n2869, n2706);
not  g2759 (n2861, n2711);
buf  g2760 (n2868, n2650);
not  g2761 (n2814, n2703);
buf  g2762 (n2874, n2689);
buf  g2763 (n2879, n2647);
not  g2764 (n2822, n2688);
not  g2765 (n2781, n2689);
not  g2766 (n2762, n2729);
buf  g2767 (n2862, n2700);
buf  g2768 (n2832, n2729);
buf  g2769 (n2749, n2632);
not  g2770 (n2840, n2565);
buf  g2771 (n2767, n2552);
not  g2772 (n2855, n2691);
not  g2773 (n2893, n2721);
buf  g2774 (n2894, n2717);
buf  g2775 (n2751, n2737);
not  g2776 (n2847, n2743);
not  g2777 (n2794, n2711);
buf  g2778 (n2867, n2700);
not  g2779 (n2860, n2732);
buf  g2780 (n2773, n2698);
buf  g2781 (n2819, n2692);
not  g2782 (n2806, n2735);
not  g2783 (n2843, n2634);
not  g2784 (n2835, n2698);
buf  g2785 (n2827, n2660);
not  g2786 (n2809, n2714);
buf  g2787 (n2786, n2700);
buf  g2788 (n2748, n2693);
not  g2789 (n2811, n2736);
not  g2790 (n2775, n2706);
buf  g2791 (n2839, n2716);
not  g2792 (n2883, n2720);
not  g2793 (n2768, n2737);
buf  g2794 (n2865, n2717);
buf  g2795 (n2833, n2694);
buf  g2796 (n2852, n2719);
not  g2797 (n2755, n2696);
buf  g2798 (n2878, n2704);
buf  g2799 (n2780, n2566);
buf  g2800 (n2793, n2623);
buf  g2801 (n2820, n2646);
buf  g2802 (n2826, n2731);
not  g2803 (n2753, n2639);
buf  g2804 (n2760, n2739);
buf  g2805 (n2800, n2710);
not  g2806 (n2891, n2704);
buf  g2807 (n2831, n2703);
buf  g2808 (n2792, n2698);
not  g2809 (n2784, n2724);
not  g2810 (n2799, n2698);
not  g2811 (n2872, n2720);
buf  g2812 (n2882, n2714);
not  g2813 (n2776, n2740);
buf  g2814 (n2850, n2699);
buf  g2815 (n2829, n2649);
buf  g2816 (n2892, n2712);
not  g2817 (n2870, n2734);
buf  g2818 (n2807, n2635);
not  g2819 (n2842, n2718);
not  g2820 (n2816, n2640);
buf  g2821 (n2797, n2725);
buf  g2822 (n2810, n2710);
xnor g2823 (n2873, n2703, n2738, n2690, n2655);
and  g2824 (n2777, n2658, n2708, n2709, n2705);
xor  g2825 (n2863, n2694, n2722, n2741, n2734);
xor  g2826 (n2750, n2688, n2708, n2709, n2696);
nand g2827 (n2880, n2712, n2552, n2716, n2730);
nand g2828 (n2859, n2696, n2713, n2627, n2697);
nand g2829 (n2779, n2733, n2726, n2718, n2732);
nor  g2830 (n2812, n2657, n2693, n2688, n2692);
and  g2831 (n2856, n2714, n2699, n2707, n2715);
xor  g2832 (n2825, n2692, n2713, n2707, n2721);
nor  g2833 (n2798, n2652, n2569, n2743, n2552);
nand g2834 (n2818, n2701, n2653, n2694, n2709);
nor  g2835 (n2808, n2651, n2728, n2734, n2732);
nand g2836 (n2866, n2701, n2743, n2735, n2736);
and  g2837 (n2885, n2723, n2648, n2696, n2740);
or   g2838 (n2803, n2708, n2624, n2736, n2722);
or   g2839 (n2875, n2722, n2730, n2713, n2729);
xnor g2840 (n2787, n2705, n2695, n2737, n2726);
nand g2841 (n2854, n2711, n2642, n2717, n2630);
xnor g2842 (n2848, n2739, n2697, n2735, n2716);
and  g2843 (n2757, n2720, n2697, n2693, n2730);
and  g2844 (n2845, n2644, n2739, n2738, n2702);
nor  g2845 (n2815, n2713, n2733, n2741, n2689);
nand g2846 (n2769, n2731, n2714, n2631, n2717);
xor  g2847 (n2853, n2694, n2742, n2733, n2727);
nor  g2848 (n2744, n2692, n2690, n2695, n2719);
and  g2849 (n2789, n2740, n2709, n2721, n2724);
xor  g2850 (n2895, n2715, n2552, n2725, n2718);
xor  g2851 (n2796, n2689, n2710, n2726, n2699);
or   g2852 (n2890, n2710, n2707, n2721, n2715);
xor  g2853 (n2745, n2705, n2708, n2703, n2626);
or   g2854 (n2846, n2731, n2743, n2740, n2701);
nor  g2855 (n2821, n2693, n2654, n2733, n2704);
nor  g2856 (n2886, n2641, n2697, n2742, n2633);
and  g2857 (n2790, n2739, n2725, n2724, n2723);
nor  g2858 (n2785, n2706, n2742, n2738, n2566);
and  g2859 (n2795, n2718, n2691, n2720);
nand g2860 (n2858, n2719, n2628, n2643, n2707);
nand g2861 (n2801, n2625, n2724, n2726, n2712);
nor  g2862 (n2877, n2695, n2736, n2699, n2737);
xnor g2863 (n2898, n2746, n2819, n2818, n2798);
xor  g2864 (n2915, n2781, n2786, n2750, n2782);
nor  g2865 (n2914, n2745, n2788, n2822, n2777);
nand g2866 (n2902, n2762, n2772, n2806, n2793);
xnor g2867 (n2901, n2814, n2770, n2800, n2773);
or   g2868 (n2899, n2792, n2771, n2754, n2790);
xor  g2869 (n2904, n2823, n2811, n2763, n2757);
xnor g2870 (n2909, n2752, n2753, n2787, n2774);
xor  g2871 (n2897, n2797, n2810, n2760, n2795);
nor  g2872 (n2896, n2769, n2799, n2807, n2789);
and  g2873 (n2913, n2756, n2776, n2748, n2803);
or   g2874 (n2905, n2751, n2749, n2809, n2780);
xnor g2875 (n2906, n2805, n2785, n2813, n2775);
and  g2876 (n2912, n2755, n2779, n2784, n2778);
nor  g2877 (n2908, n2768, n2820, n2759, n2821);
xnor g2878 (n2911, n2744, n2804, n2802, n2783);
xnor g2879 (n2903, n2791, n2767, n2801, n2816);
and  g2880 (n2910, n2764, n2808, n2812, n2761);
and  g2881 (n2900, n2758, n2817, n2815, n2766);
xnor g2882 (n2907, n2747, n2796, n2765, n2794);
and  g2883 (n2919, n2903, n2837, n2831, n2832);
and  g2884 (n2920, n2905, n2904, n2825, n2827);
or   g2885 (n2917, n2907, n2826, n2901, n2902);
or   g2886 (n2916, n2838, n2834, n2908, n2833);
xnor g2887 (n2921, n2824, n2828, n2835, n2829);
xnor g2888 (n2918, n2174, n2906, n2836, n2830);
and  g2889 (n2922, n2839, n2921, n1983);
xnor g2890 (n2923, n2920, n2840, n1983);
xor  g2891 (n2925, n2851, n2847, n2864, n2862);
or   g2892 (n2929, n2922, n2857, n2843, n2841);
nand g2893 (n2930, n2858, n2922, n2852, n2923);
xor  g2894 (n2926, n2923, n2861, n2856, n2849);
nor  g2895 (n2931, n2855, n2860, n2845, n2844);
or   g2896 (n2924, n2923, n2853, n2863, n2854);
nor  g2897 (n2927, n2848, n2923, n2850, n2922);
xor  g2898 (n2928, n2859, n2922, n2842, n2846);
nand g2899 (n2957, n1989, n1985, n2929, n2925);
xor  g2900 (n2948, n1995, n1985, n2883, n2881);
xnor g2901 (n2961, n1997, n1986, n1988, n2912);
nor  g2902 (n2955, n2000, n2911, n2865, n1991);
xor  g2903 (n2934, n2925, n2926, n2931, n2882);
nor  g2904 (n2946, n2000, n1991, n1994);
nand g2905 (n2940, n2930, n1990, n2876, n2871);
and  g2906 (n2942, n2928, n1987, n1995);
and  g2907 (n2937, n2877, n2873, n2927, n1992);
xnor g2908 (n2951, n1984, n1989, n1992, n2926);
nor  g2909 (n2943, n1997, n1987, n1990, n1985);
xnor g2910 (n2947, n2347, n1993, n1992, n1998);
and  g2911 (n2932, n1991, n1993, n2925, n2927);
nor  g2912 (n2960, n2927, n1994, n1998, n2930);
xor  g2913 (n2941, n1984, n1989, n1993, n2910);
or   g2914 (n2949, n1988, n1984, n2929, n2931);
nor  g2915 (n2958, n2924, n1997, n1987, n2928);
nor  g2916 (n2938, n1999, n2929, n2928, n1996);
xor  g2917 (n2933, n2926, n1994, n2874, n2879);
xnor g2918 (n2959, n2924, n2872, n2915, n2000);
xor  g2919 (n2935, n1996, n2927, n2931, n2926);
or   g2920 (n2962, n1993, n2867, n1988, n2930);
nor  g2921 (n2956, n1984, n2913, n2884, n1989);
xnor g2922 (n2953, n1999, n1990, n1985, n1995);
xor  g2923 (n2954, n2924, n1999, n2914, n1986);
nand g2924 (n2952, n1997, n2925, n1986, n1995);
and  g2925 (n2950, n2000, n2880, n1996);
or   g2926 (n2945, n2878, n2924, n2866, n1986);
and  g2927 (n2936, n2875, n2869, n1998, n1999);
or   g2928 (n2944, n1992, n2870, n2868, n1998);
and  g2929 (n2963, n2929, n2931, n1994, n2928);
xnor g2930 (n2939, n2909, n1988, n1990, n2930);
or   g2931 (n3012, n2275, n2183, n2962, n2251);
xnor g2932 (n3002, n2310, n2254, n2293, n2276);
nor  g2933 (n2984, n2221, n2230, n2959, n2323);
xor  g2934 (n2975, n2253, n2280, n2288, n2933);
nor  g2935 (n2973, n2937, n2281, n2886, n2952);
nand g2936 (n2992, n2242, n2302, n2278, n2296);
xnor g2937 (n3018, n2944, n2316, n2939, n2958);
nand g2938 (n3011, n2189, n2191, n2244, n2201);
xor  g2939 (n2972, n2279, n2954, n2177, n2292);
nor  g2940 (n3007, n2215, n2206, n2962, n2955);
nor  g2941 (n2969, n2325, n2208, n2198, n2960);
nor  g2942 (n3010, n2247, n2252, n2181, n2263);
and  g2943 (n2985, n2284, n2321, n2236, n2320);
or   g2944 (n2996, n2237, n2312, n2243, n2235);
or   g2945 (n2967, n2226, n2283, n2958, n2943);
nor  g2946 (n2974, n2257, n2959, n2285, n2274);
or   g2947 (n3000, n2264, n2234, n2892, n2239);
and  g2948 (n3016, n2179, n2241, n2948, n2960);
xor  g2949 (n3004, n2887, n2211, n2245, n2219);
nor  g2950 (n3003, n2314, n2178, n2962, n2318);
nor  g2951 (n3009, n2938, n2963, n2240, n2893);
and  g2952 (n2994, n2246, n2956, n2295, n2216);
xor  g2953 (n2990, n2960, n2936, n2207, n2260);
xor  g2954 (n3005, n2959, n2304, n2270, n2228);
nor  g2955 (n3014, n2193, n2209, n2214, n2203);
nand g2956 (n3015, n2290, n2286, n2180, n2955);
xnor g2957 (n2971, n2266, n2959, n2250, n2961);
nand g2958 (n2999, n2949, n2950, n2328, n2192);
nor  g2959 (n2965, n2894, n2233, n2309, n2273);
xnor g2960 (n2980, n2197, n2232, n2282, n2324);
or   g2961 (n3008, n2962, n2935, n2188, n2213);
nor  g2962 (n2970, n2297, n2956, n2305, n2255);
nand g2963 (n2979, n2291, n2248, n2176, n2259);
xnor g2964 (n2989, n2961, n2277, n2289, n2322);
xnor g2965 (n3017, n2225, n2319, n2963, n2265);
or   g2966 (n2988, n2195, n2185, n2238, n2190);
and  g2967 (n2991, n2287, n2957, n2329, n2941);
xnor g2968 (n2976, n2262, n2961, n2947, n2218);
xor  g2969 (n2966, n2315, n2303, n2890, n2249);
nand g2970 (n2987, n2217, n2220, n2256, n2223);
or   g2971 (n3006, n2963, n2300, n2888, n2307);
or   g2972 (n2993, n2268, n2940, n2301, n2958);
nand g2973 (n3001, n2308, n2224, n2945, n2184);
and  g2974 (n2964, n2175, n2326, n2210, n2942);
and  g2975 (n2995, n2196, n2957, n2199, n2311);
xor  g2976 (n2977, n2951, n2891, n2212, n2960);
and  g2977 (n2983, n2261, n2327, n2231, n2889);
and  g2978 (n3013, n2957, n2186, n2205, n2299);
xor  g2979 (n2982, n2271, n2182, n2200, n2272);
xnor g2980 (n2968, n2953, n2958, n2267, n2229);
nand g2981 (n2978, n2187, n2294, n2932, n2946);
and  g2982 (n2998, n2269, n2306, n2317, n2227);
or   g2983 (n2997, n2202, n2298, n2934, n2204);
nand g2984 (n2981, n2961, n2222, n2313, n2194);
or   g2985 (n2986, n2885, n2957, n2258, n2963);
nand g2986 (n3026, n2964, n3018, n2984, n2999);
xor  g2987 (n3027, n2995, n2988, n2980, n2971);
or   g2988 (n3030, n3013, n3015, n2990, n2974);
nand g2989 (n3029, n3007, n2977, n2972, n2976);
nor  g2990 (n3020, n2983, n3012, n2996, n2985);
and  g2991 (n3032, n3017, n3005, n3009, n2994);
nand g2992 (n3025, n2993, n2969, n2965, n3002);
nand g2993 (n3031, n2968, n3003, n2986, n2998);
xnor g2994 (n3028, n2987, n3011, n3014, n2982);
xor  g2995 (n3019, n3001, n3000, n2979, n3010);
xor  g2996 (n3024, n2991, n2975, n3008, n2970);
xnor g2997 (n3022, n3016, n2966, n2997, n2992);
or   g2998 (n3021, n2895, n3006, n2989, n2973);
nor  g2999 (n3023, n3004, n2981, n2978, n2967);
endmodule
