

module Stat_403_1822
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n193,
  n210,
  n211,
  n204,
  n189,
  n202,
  n212,
  n364,
  n368,
  n367,
  n371,
  n372,
  n377,
  n375,
  n418,
  n421,
  n417,
  n419,
  n422,
  n420
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n193;output n210;output n211;output n204;output n189;output n202;output n212;output n364;output n368;output n367;output n371;output n372;output n377;output n375;output n418;output n421;output n417;output n419;output n422;output n420;
  wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n190;wire n191;wire n192;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n203;wire n205;wire n206;wire n207;wire n208;wire n209;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n365;wire n366;wire n369;wire n370;wire n373;wire n374;wire n376;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;

  buf
  g0
  (
    n39,
    n12
  );


  not
  g1
  (
    n94,
    n1
  );


  buf
  g2
  (
    n32,
    n17
  );


  buf
  g3
  (
    n73,
    n8
  );


  buf
  g4
  (
    n78,
    n3
  );


  buf
  g5
  (
    n22,
    n19
  );


  not
  g6
  (
    n59,
    n1
  );


  buf
  g7
  (
    n27,
    n11
  );


  not
  g8
  (
    n89,
    n18
  );


  not
  g9
  (
    n40,
    n14
  );


  buf
  g10
  (
    n20,
    n18
  );


  buf
  g11
  (
    n74,
    n9
  );


  buf
  g12
  (
    n82,
    n5
  );


  not
  g13
  (
    n63,
    n8
  );


  buf
  g14
  (
    n42,
    n9
  );


  not
  g15
  (
    n43,
    n17
  );


  buf
  g16
  (
    n80,
    n10
  );


  not
  g17
  (
    n35,
    n2
  );


  buf
  g18
  (
    KeyWire_0_5,
    n10
  );


  not
  g19
  (
    n56,
    n8
  );


  buf
  g20
  (
    n50,
    n3
  );


  not
  g21
  (
    n70,
    n5
  );


  buf
  g22
  (
    n44,
    n16
  );


  buf
  g23
  (
    n68,
    n6
  );


  not
  g24
  (
    n81,
    n4
  );


  not
  g25
  (
    n41,
    n9
  );


  not
  g26
  (
    n26,
    n2
  );


  buf
  g27
  (
    n53,
    n13
  );


  buf
  g28
  (
    n29,
    n5
  );


  buf
  g29
  (
    n88,
    n16
  );


  not
  g30
  (
    n38,
    n18
  );


  buf
  g31
  (
    n51,
    n3
  );


  not
  g32
  (
    n46,
    n18
  );


  not
  g33
  (
    n90,
    n13
  );


  buf
  g34
  (
    n49,
    n1
  );


  not
  g35
  (
    n25,
    n8
  );


  not
  g36
  (
    n31,
    n9
  );


  not
  g37
  (
    n34,
    n5
  );


  not
  g38
  (
    n58,
    n3
  );


  buf
  g39
  (
    n71,
    n13
  );


  not
  g40
  (
    n37,
    n7
  );


  not
  g41
  (
    n47,
    n13
  );


  buf
  g42
  (
    n93,
    n19
  );


  buf
  g43
  (
    n86,
    n2
  );


  not
  g44
  (
    n91,
    n6
  );


  buf
  g45
  (
    n45,
    n12
  );


  buf
  g46
  (
    n55,
    n17
  );


  buf
  g47
  (
    n61,
    n11
  );


  buf
  g48
  (
    n33,
    n14
  );


  buf
  g49
  (
    n83,
    n17
  );


  not
  g50
  (
    n79,
    n1
  );


  not
  g51
  (
    n24,
    n10
  );


  buf
  g52
  (
    n87,
    n11
  );


  not
  g53
  (
    n62,
    n16
  );


  buf
  g54
  (
    n77,
    n12
  );


  not
  g55
  (
    n69,
    n7
  );


  not
  g56
  (
    n92,
    n15
  );


  buf
  g57
  (
    n60,
    n7
  );


  buf
  g58
  (
    n28,
    n10
  );


  buf
  g59
  (
    n76,
    n15
  );


  buf
  g60
  (
    KeyWire_0_12,
    n16
  );


  buf
  g61
  (
    n84,
    n2
  );


  buf
  g62
  (
    n95,
    n19
  );


  buf
  g63
  (
    KeyWire_0_13,
    n6
  );


  not
  g64
  (
    n30,
    n14
  );


  not
  g65
  (
    n64,
    n4
  );


  not
  g66
  (
    n23,
    n11
  );


  not
  g67
  (
    n72,
    n4
  );


  not
  g68
  (
    n36,
    n15
  );


  buf
  g69
  (
    n54,
    n12
  );


  not
  g70
  (
    n48,
    n14
  );


  not
  g71
  (
    n85,
    n4
  );


  not
  g72
  (
    n52,
    n15
  );


  not
  g73
  (
    n75,
    n19
  );


  buf
  g74
  (
    n57,
    n6
  );


  buf
  g75
  (
    n66,
    n7
  );


  not
  g76
  (
    n115,
    n36
  );


  buf
  g77
  (
    n124,
    n47
  );


  not
  g78
  (
    n156,
    n37
  );


  buf
  g79
  (
    n123,
    n37
  );


  buf
  g80
  (
    n152,
    n57
  );


  buf
  g81
  (
    n168,
    n57
  );


  buf
  g82
  (
    n153,
    n54
  );


  not
  g83
  (
    n137,
    n33
  );


  buf
  g84
  (
    n159,
    n30
  );


  not
  g85
  (
    n132,
    n34
  );


  not
  g86
  (
    n136,
    n53
  );


  not
  g87
  (
    n148,
    n33
  );


  buf
  g88
  (
    n135,
    n29
  );


  buf
  g89
  (
    n130,
    n23
  );


  not
  g90
  (
    n160,
    n39
  );


  buf
  g91
  (
    n141,
    n26
  );


  buf
  g92
  (
    n133,
    n53
  );


  buf
  g93
  (
    n112,
    n34
  );


  buf
  g94
  (
    KeyWire_0_7,
    n47
  );


  buf
  g95
  (
    n107,
    n21
  );


  not
  g96
  (
    n151,
    n41
  );


  not
  g97
  (
    n171,
    n40
  );


  buf
  g98
  (
    n158,
    n45
  );


  buf
  g99
  (
    n169,
    n52
  );


  buf
  g100
  (
    n176,
    n50
  );


  buf
  g101
  (
    n125,
    n30
  );


  not
  g102
  (
    n108,
    n59
  );


  buf
  g103
  (
    n175,
    n44
  );


  buf
  g104
  (
    n119,
    n43
  );


  not
  g105
  (
    n116,
    n46
  );


  not
  g106
  (
    n161,
    n26
  );


  buf
  g107
  (
    n157,
    n51
  );


  not
  g108
  (
    n105,
    n42
  );


  buf
  g109
  (
    n163,
    n48
  );


  not
  g110
  (
    n99,
    n22
  );


  buf
  g111
  (
    n179,
    n60
  );


  buf
  g112
  (
    n117,
    n49
  );


  buf
  g113
  (
    n178,
    n50
  );


  not
  g114
  (
    n102,
    n49
  );


  buf
  g115
  (
    n131,
    n51
  );


  buf
  g116
  (
    n182,
    n36
  );


  buf
  g117
  (
    n165,
    n27
  );


  not
  g118
  (
    n166,
    n30
  );


  buf
  g119
  (
    n167,
    n24
  );


  buf
  g120
  (
    n113,
    n55
  );


  buf
  g121
  (
    n188,
    n50
  );


  buf
  g122
  (
    n172,
    n61
  );


  buf
  g123
  (
    n177,
    n42
  );


  buf
  g124
  (
    n147,
    n58
  );


  not
  g125
  (
    n185,
    n48
  );


  not
  g126
  (
    KeyWire_0_0,
    n27
  );


  buf
  g127
  (
    n111,
    n41
  );


  not
  g128
  (
    n122,
    n60
  );


  buf
  g129
  (
    n164,
    n60
  );


  not
  g130
  (
    n120,
    n29
  );


  not
  g131
  (
    n101,
    n60
  );


  buf
  g132
  (
    n104,
    n31
  );


  not
  g133
  (
    KeyWire_0_4,
    n57
  );


  not
  g134
  (
    n110,
    n61
  );


  buf
  g135
  (
    n106,
    n59
  );


  buf
  g136
  (
    n126,
    n43
  );


  buf
  g137
  (
    n128,
    n53
  );


  not
  g138
  (
    n121,
    n35
  );


  buf
  g139
  (
    n154,
    n35
  );


  buf
  g140
  (
    n114,
    n20
  );


  not
  g141
  (
    n187,
    n52
  );


  buf
  g142
  (
    n96,
    n44
  );


  buf
  g143
  (
    n186,
    n38
  );


  not
  g144
  (
    n146,
    n56
  );


  not
  g145
  (
    n180,
    n51
  );


  not
  g146
  (
    n155,
    n28
  );


  not
  g147
  (
    n144,
    n55
  );


  nor
  g148
  (
    n134,
    n42,
    n61
  );


  nor
  g149
  (
    n162,
    n25,
    n46,
    n40,
    n50
  );


  xnor
  g150
  (
    n97,
    n48,
    n58,
    n40,
    n56
  );


  xor
  g151
  (
    n183,
    n28,
    n28,
    n38,
    n55
  );


  nor
  g152
  (
    n143,
    n36,
    n49,
    n35,
    n37
  );


  nand
  g153
  (
    n139,
    n56,
    n54,
    n27,
    n55
  );


  xor
  g154
  (
    n184,
    n52,
    n53,
    n32,
    n58
  );


  nor
  g155
  (
    n140,
    n47,
    n34,
    n32,
    n46
  );


  xnor
  g156
  (
    n109,
    n52,
    n56,
    n22,
    n45
  );


  nor
  g157
  (
    n127,
    n33,
    n54,
    n42,
    n59
  );


  nand
  g158
  (
    n150,
    n41,
    n21,
    n59,
    n40
  );


  xnor
  g159
  (
    n142,
    n28,
    n47,
    n48,
    n41
  );


  xnor
  g160
  (
    n149,
    n38,
    n32,
    n25,
    n61
  );


  xor
  g161
  (
    n173,
    n44,
    n43,
    n58,
    n31
  );


  xnor
  g162
  (
    n138,
    n31,
    n39,
    n45,
    n57
  );


  xnor
  g163
  (
    n118,
    n45,
    n32,
    n30,
    n37
  );


  nor
  g164
  (
    n103,
    n23,
    n24,
    n20,
    n44
  );


  nor
  g165
  (
    n129,
    n31,
    n38,
    n34,
    n46
  );


  xor
  g166
  (
    n100,
    n49,
    n35,
    n33,
    n51
  );


  nand
  g167
  (
    n174,
    n29,
    n29,
    n39,
    n36
  );


  or
  g168
  (
    n170,
    n43,
    n54,
    n27,
    n39
  );


  xor
  g169
  (
    n191,
    n75,
    n100,
    n64,
    n70
  );


  xnor
  g170
  (
    n204,
    n63,
    n125,
    n71,
    n97
  );


  nand
  g171
  (
    n199,
    n104,
    n72,
    n98,
    n74
  );


  xnor
  g172
  (
    n196,
    n101,
    n111,
    n115,
    n76
  );


  and
  g173
  (
    n189,
    n65,
    n124,
    n106,
    n129
  );


  and
  g174
  (
    n203,
    n65,
    n77,
    n74
  );


  xor
  g175
  (
    n208,
    n96,
    n126,
    n120,
    n122
  );


  xor
  g176
  (
    n192,
    n68,
    n119,
    n65,
    n113
  );


  xor
  g177
  (
    n190,
    n70,
    n99,
    n67
  );


  nand
  g178
  (
    n197,
    n76,
    n71,
    n77,
    n107
  );


  nor
  g179
  (
    n205,
    n127,
    n62,
    n68,
    n66
  );


  nor
  g180
  (
    n201,
    n65,
    n62,
    n73,
    n117
  );


  or
  g181
  (
    n206,
    n76,
    n69,
    n123,
    n71
  );


  and
  g182
  (
    n207,
    n67,
    n75,
    n118,
    n108
  );


  nand
  g183
  (
    n210,
    n69,
    n72,
    n64,
    n78
  );


  nor
  g184
  (
    n194,
    n73,
    n73,
    n63,
    n75
  );


  or
  g185
  (
    n211,
    n128,
    n63,
    n72,
    n110
  );


  and
  g186
  (
    n200,
    n72,
    n74,
    n64,
    n69
  );


  nand
  g187
  (
    n195,
    n105,
    n66,
    n77,
    n62
  );


  and
  g188
  (
    n213,
    n70,
    n74,
    n68,
    n62
  );


  and
  g189
  (
    n202,
    n102,
    n112,
    n121,
    n66
  );


  and
  g190
  (
    n193,
    n116,
    n109,
    n63,
    n66
  );


  or
  g191
  (
    n209,
    n114,
    n68,
    n78,
    n73
  );


  nor
  g192
  (
    n198,
    n64,
    n70,
    n69,
    n76
  );


  xnor
  g193
  (
    n212,
    n67,
    n71,
    n103,
    n75
  );


  buf
  g194
  (
    n223,
    n205
  );


  buf
  g195
  (
    n225,
    n197
  );


  not
  g196
  (
    n219,
    n145
  );


  buf
  g197
  (
    n221,
    n137
  );


  not
  g198
  (
    n217,
    n138
  );


  buf
  g199
  (
    n214,
    n135
  );


  xor
  g200
  (
    n220,
    n131,
    n196
  );


  xnor
  g201
  (
    n215,
    n207,
    n136,
    n201,
    n130
  );


  and
  g202
  (
    n222,
    n202,
    n140,
    n198,
    n203
  );


  and
  g203
  (
    n224,
    n142,
    n139,
    n133,
    n200
  );


  xor
  g204
  (
    n216,
    n144,
    n143,
    n199,
    n206
  );


  nand
  g205
  (
    n218,
    n204,
    n141,
    n132,
    n134
  );


  buf
  g206
  (
    n246,
    n220
  );


  not
  g207
  (
    KeyWire_0_6,
    n214
  );


  buf
  g208
  (
    n242,
    n217
  );


  buf
  g209
  (
    n241,
    n225
  );


  not
  g210
  (
    n227,
    n210
  );


  not
  g211
  (
    n226,
    n225
  );


  buf
  g212
  (
    KeyWire_0_2,
    n221
  );


  buf
  g213
  (
    n236,
    n218
  );


  not
  g214
  (
    n235,
    n223
  );


  buf
  g215
  (
    n231,
    n215
  );


  buf
  g216
  (
    n234,
    n224
  );


  buf
  g217
  (
    n239,
    n222
  );


  buf
  g218
  (
    n228,
    n224
  );


  not
  g219
  (
    KeyWire_0_1,
    n222
  );


  buf
  g220
  (
    n233,
    n221
  );


  buf
  g221
  (
    n247,
    n208
  );


  not
  g222
  (
    n245,
    n216
  );


  not
  g223
  (
    n244,
    n219
  );


  buf
  g224
  (
    n237,
    n220
  );


  buf
  g225
  (
    n238,
    n216
  );


  buf
  g226
  (
    n230,
    n223
  );


  xor
  g227
  (
    n229,
    n217,
    n218,
    n209,
    n219
  );


  not
  g228
  (
    n250,
    n230
  );


  not
  g229
  (
    n255,
    n232
  );


  buf
  g230
  (
    n254,
    n227
  );


  buf
  g231
  (
    n253,
    n226
  );


  not
  g232
  (
    n265,
    n229
  );


  buf
  g233
  (
    n258,
    n229
  );


  buf
  g234
  (
    n249,
    n232
  );


  buf
  g235
  (
    KeyWire_0_10,
    n233
  );


  buf
  g236
  (
    n259,
    n230
  );


  buf
  g237
  (
    n263,
    n232
  );


  not
  g238
  (
    KeyWire_0_8,
    n231
  );


  buf
  g239
  (
    n264,
    n232
  );


  not
  g240
  (
    n266,
    n228
  );


  not
  g241
  (
    n251,
    n231
  );


  buf
  g242
  (
    n252,
    n231
  );


  buf
  g243
  (
    n261,
    n226
  );


  not
  g244
  (
    n262,
    n228
  );


  buf
  g245
  (
    n248,
    n231
  );


  not
  g246
  (
    n257,
    n227
  );


  and
  g247
  (
    n291,
    n149,
    n147,
    n234,
    n253
  );


  nor
  g248
  (
    KeyWire_0_11,
    n166,
    n235,
    n236,
    n168
  );


  nor
  g249
  (
    n279,
    n255,
    n252,
    n153,
    n233
  );


  nand
  g250
  (
    n270,
    n241,
    n243,
    n239,
    n257
  );


  nor
  g251
  (
    n277,
    n160,
    n241,
    n249
  );


  xnor
  g252
  (
    n286,
    n256,
    n254,
    n179,
    n173
  );


  nand
  g253
  (
    n290,
    n250,
    n248,
    n253,
    n239
  );


  xor
  g254
  (
    n268,
    n243,
    n237,
    n250,
    n236
  );


  nand
  g255
  (
    n281,
    n167,
    n238,
    n161,
    n239
  );


  nand
  g256
  (
    n282,
    n242,
    n242,
    n234,
    n238
  );


  xor
  g257
  (
    n267,
    n235,
    n233,
    n163,
    n236
  );


  or
  g258
  (
    n271,
    n169,
    n237,
    n248,
    n254
  );


  xnor
  g259
  (
    n292,
    n146,
    n256,
    n251,
    n158
  );


  nand
  g260
  (
    n273,
    n157,
    n174,
    n243,
    n162
  );


  xnor
  g261
  (
    n284,
    n171,
    n176,
    n155,
    n256
  );


  xor
  g262
  (
    n278,
    n257,
    n152,
    n175,
    n178
  );


  xnor
  g263
  (
    n272,
    n254,
    n256,
    n177,
    n255
  );


  nor
  g264
  (
    n283,
    n255,
    n252,
    n240,
    n235
  );


  and
  g265
  (
    n269,
    n239,
    n151,
    n236,
    n165
  );


  or
  g266
  (
    n276,
    n159,
    n251,
    n164,
    n255
  );


  or
  g267
  (
    n280,
    n243,
    n238,
    n249,
    n241
  );


  xnor
  g268
  (
    n275,
    n235,
    n242,
    n233,
    n150
  );


  nor
  g269
  (
    n288,
    n240,
    n170,
    n172,
    n238
  );


  nor
  g270
  (
    n285,
    n234,
    n242,
    n240,
    n254
  );


  xnor
  g271
  (
    n289,
    n237,
    n154,
    n257,
    n240
  );


  nand
  g272
  (
    n287,
    n156,
    n237,
    n148,
    n234
  );


  or
  g273
  (
    n295,
    n257,
    n269,
    n270,
    n259
  );


  nor
  g274
  (
    n296,
    n268,
    n260,
    n258
  );


  or
  g275
  (
    n293,
    n259,
    n274,
    n272,
    n271
  );


  or
  g276
  (
    n297,
    n267,
    n258,
    n273
  );


  nor
  g277
  (
    n294,
    n260,
    n259
  );


  buf
  g278
  (
    n304,
    n294
  );


  not
  g279
  (
    n308,
    n297
  );


  buf
  g280
  (
    n309,
    n297
  );


  not
  g281
  (
    n311,
    n275
  );


  not
  g282
  (
    n301,
    n295
  );


  not
  g283
  (
    n310,
    n295
  );


  not
  g284
  (
    n307,
    n296
  );


  not
  g285
  (
    n305,
    n294
  );


  not
  g286
  (
    KeyWire_0_15,
    n295
  );


  not
  g287
  (
    n303,
    n293
  );


  buf
  g288
  (
    n298,
    n278
  );


  buf
  g289
  (
    n306,
    n296
  );


  buf
  g290
  (
    n313,
    n297
  );


  buf
  g291
  (
    n312,
    n296
  );


  and
  g292
  (
    n299,
    n276,
    n277
  );


  or
  g293
  (
    n302,
    n293,
    n295,
    n296,
    n297
  );


  not
  g294
  (
    n315,
    n78
  );


  xnor
  g295
  (
    n321,
    n284,
    n245
  );


  xor
  g296
  (
    n330,
    n300,
    n313,
    n80,
    n247
  );


  nor
  g297
  (
    n331,
    n244,
    n310,
    n213,
    n312
  );


  xor
  g298
  (
    n326,
    n244,
    n78,
    n79,
    n311
  );


  and
  g299
  (
    n328,
    n301,
    n290,
    n313,
    n79
  );


  or
  g300
  (
    n316,
    n279,
    n286,
    n312,
    n280
  );


  xnor
  g301
  (
    n332,
    n245,
    n212,
    n303,
    n310
  );


  and
  g302
  (
    n325,
    n246,
    n82,
    n81,
    n307
  );


  nor
  g303
  (
    n323,
    n285,
    n82,
    n81,
    n80
  );


  nand
  g304
  (
    n314,
    n247,
    n298,
    n306,
    n309
  );


  or
  g305
  (
    KeyWire_0_9,
    n79,
    n302,
    n247,
    n82
  );


  xor
  g306
  (
    n322,
    n311,
    n246,
    n289,
    n79
  );


  xor
  g307
  (
    n317,
    n245,
    n83,
    n246,
    n288
  );


  or
  g308
  (
    n320,
    n304,
    n281,
    n287,
    n80
  );


  nor
  g309
  (
    n324,
    n244,
    n308,
    n246,
    n291
  );


  nand
  g310
  (
    n318,
    n80,
    n211,
    n83,
    n282
  );


  and
  g311
  (
    n327,
    n299,
    n81,
    n247,
    n244
  );


  nor
  g312
  (
    n319,
    n305,
    n82,
    n81,
    n283
  );


  not
  g313
  (
    n347,
    n315
  );


  buf
  g314
  (
    n339,
    n318
  );


  not
  g315
  (
    n344,
    n318
  );


  not
  g316
  (
    n337,
    n317
  );


  not
  g317
  (
    n350,
    n322
  );


  buf
  g318
  (
    n340,
    n314
  );


  buf
  g319
  (
    n351,
    n316
  );


  buf
  g320
  (
    n349,
    n319
  );


  buf
  g321
  (
    n341,
    n321
  );


  buf
  g322
  (
    n345,
    n322
  );


  not
  g323
  (
    n346,
    n322
  );


  buf
  g324
  (
    n333,
    n315
  );


  buf
  g325
  (
    n342,
    n319
  );


  buf
  g326
  (
    KeyWire_0_14,
    n314
  );


  not
  g327
  (
    n335,
    n316
  );


  not
  g328
  (
    n338,
    n320
  );


  buf
  g329
  (
    n348,
    n322
  );


  not
  g330
  (
    n336,
    n320
  );


  not
  g331
  (
    n334,
    n321
  );


  not
  g332
  (
    n343,
    n317
  );


  and
  g333
  (
    n355,
    n335,
    n333,
    n326,
    n327
  );


  and
  g334
  (
    n353,
    n327,
    n328,
    n324,
    n323
  );


  xnor
  g335
  (
    n359,
    n335,
    n328,
    n334,
    n329
  );


  or
  g336
  (
    n354,
    n328,
    n323,
    n327,
    n326
  );


  and
  g337
  (
    n361,
    n336,
    n324,
    n325
  );


  xor
  g338
  (
    n357,
    n326,
    n333,
    n334,
    n328
  );


  or
  g339
  (
    n356,
    n329,
    n323,
    n324,
    n335
  );


  and
  g340
  (
    n360,
    n324,
    n327,
    n325,
    n336
  );


  xor
  g341
  (
    n358,
    n325,
    n335,
    n323,
    n326
  );


  or
  g342
  (
    n368,
    n342,
    n341,
    n356,
    n338
  );


  nor
  g343
  (
    n365,
    n353,
    n360,
    n342,
    n341
  );


  nand
  g344
  (
    n370,
    n337,
    n337,
    n343,
    n342
  );


  xor
  g345
  (
    n366,
    n343,
    n340
  );


  nand
  g346
  (
    n369,
    n337,
    n339,
    n338
  );


  and
  g347
  (
    n371,
    n336,
    n339,
    n337
  );


  and
  g348
  (
    n364,
    n359,
    n343,
    n358,
    n342
  );


  xor
  g349
  (
    n367,
    n355,
    n338,
    n361
  );


  xor
  g350
  (
    n363,
    n338,
    n340,
    n354,
    n357
  );


  nor
  g351
  (
    n362,
    n336,
    n341,
    n343
  );


  nor
  g352
  (
    n375,
    n85,
    n85,
    n369,
    n368
  );


  nand
  g353
  (
    n372,
    n83,
    n85,
    n87
  );


  xor
  g354
  (
    n376,
    n86,
    n84
  );


  nor
  g355
  (
    n377,
    n87,
    n86,
    n371,
    n370
  );


  and
  g356
  (
    n373,
    n84,
    n366,
    n367,
    n83
  );


  xnor
  g357
  (
    n374,
    n292,
    n85,
    n86
  );


  nand
  g358
  (
    n380,
    n188,
    n185,
    n182,
    n183
  );


  xor
  g359
  (
    n378,
    n186,
    n184,
    n375,
    n180
  );


  nand
  g360
  (
    n379,
    n376,
    n187,
    n181,
    n377
  );


  or
  g361
  (
    n381,
    n352,
    n379,
    n347,
    n345
  );


  xnor
  g362
  (
    n383,
    n352,
    n345,
    n348,
    n349
  );


  and
  g363
  (
    n390,
    n349,
    n345,
    n380,
    n379
  );


  or
  g364
  (
    n391,
    n379,
    n347,
    n380,
    n378
  );


  and
  g365
  (
    n389,
    n346,
    n352,
    n351,
    n344
  );


  xnor
  g366
  (
    n392,
    n379,
    n346,
    n378
  );


  xnor
  g367
  (
    n387,
    n378,
    n380,
    n346,
    n350
  );


  xor
  g368
  (
    KeyWire_0_3,
    n344,
    n349,
    n351,
    n348
  );


  or
  g369
  (
    n382,
    n345,
    n378,
    n344,
    n349
  );


  and
  g370
  (
    n388,
    n380,
    n350,
    n351
  );


  nand
  g371
  (
    n384,
    n348,
    n344,
    n347,
    n351
  );


  xnor
  g372
  (
    n385,
    n348,
    n350,
    n352,
    n347
  );


  xnor
  g373
  (
    n399,
    n263,
    n332,
    n89,
    n95
  );


  nand
  g374
  (
    n414,
    n91,
    n332,
    n264,
    n94
  );


  nor
  g375
  (
    n406,
    n266,
    n262,
    n261,
    n391
  );


  xnor
  g376
  (
    n410,
    n91,
    n386,
    n388,
    n93
  );


  xor
  g377
  (
    n396,
    n264,
    n330,
    n261,
    n93
  );


  or
  g378
  (
    n405,
    n389,
    n382,
    n262,
    n386
  );


  nor
  g379
  (
    n401,
    n93,
    n88,
    n94,
    n95
  );


  nor
  g380
  (
    n395,
    n383,
    n92,
    n331,
    n94
  );


  nor
  g381
  (
    n400,
    n260,
    n266,
    n88,
    n92
  );


  and
  g382
  (
    n394,
    n382,
    n90,
    n264,
    n332
  );


  and
  g383
  (
    n415,
    n389,
    n265,
    n261,
    n387
  );


  xor
  g384
  (
    n407,
    n330,
    n88,
    n263
  );


  xnor
  g385
  (
    n403,
    n266,
    n90,
    n390,
    n392
  );


  nor
  g386
  (
    n398,
    n329,
    n89,
    n90,
    n261
  );


  nor
  g387
  (
    n393,
    n332,
    n387,
    n263,
    n91
  );


  or
  g388
  (
    n397,
    n265,
    n330,
    n331,
    n390
  );


  and
  g389
  (
    n408,
    n95,
    n392,
    n92,
    n89
  );


  xor
  g390
  (
    n402,
    n263,
    n331,
    n262,
    n384
  );


  xor
  g391
  (
    n413,
    n381,
    n329,
    n331,
    n262
  );


  xor
  g392
  (
    n409,
    n385,
    n95,
    n90,
    n89
  );


  xnor
  g393
  (
    n411,
    n265,
    n381,
    n385,
    n94
  );


  nand
  g394
  (
    n416,
    n383,
    n391,
    n92,
    n265
  );


  and
  g395
  (
    n412,
    n330,
    n87,
    n266,
    n91
  );


  xor
  g396
  (
    n404,
    n93,
    n264,
    n388,
    n384
  );


  and
  g397
  (
    n420,
    n412,
    n400,
    n398,
    n413
  );


  nand
  g398
  (
    n421,
    n405,
    n415,
    n397,
    n409
  );


  nor
  g399
  (
    n419,
    n403,
    n393,
    n408,
    n411
  );


  xnor
  g400
  (
    n418,
    n396,
    n406,
    n401,
    n416
  );


  and
  g401
  (
    n422,
    n414,
    n394,
    n399,
    n402
  );


  and
  g402
  (
    n417,
    n407,
    n410,
    n404,
    n395
  );


  xor
  KeyGate_0_0
  (
    n98,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n243,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n240,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n386,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n145,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n67,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n232,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n181,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n256,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n329,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n260,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n274,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n65,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n21,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n352,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n300,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


