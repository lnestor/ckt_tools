

module Stat_1619_32_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n1525,
  n1539,
  n1537,
  n1538,
  n1610,
  n1619,
  n1620,
  n1612,
  n1611,
  n1614,
  n1628,
  n1637,
  n1632,
  n1643,
  n1634,
  n1630,
  n1636,
  n1642,
  n1635,
  n1638,
  n1640,
  n1639,
  n1641,
  n1631,
  n1629,
  n1651,
  n1650,
  n1653,
  n1649,
  n1658,
  n1654,
  n1657,
  n1652,
  n1655,
  n1656
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1525;output n1539;output n1537;output n1538;output n1610;output n1619;output n1620;output n1612;output n1611;output n1614;output n1628;output n1637;output n1632;output n1643;output n1634;output n1630;output n1636;output n1642;output n1635;output n1638;output n1640;output n1639;output n1641;output n1631;output n1629;output n1651;output n1650;output n1653;output n1649;output n1658;output n1654;output n1657;output n1652;output n1655;output n1656;
  wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1613;wire n1615;wire n1616;wire n1617;wire n1618;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1633;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n47,
    n32
  );


  not
  g1
  (
    n45,
    n16
  );


  not
  g2
  (
    n168,
    n4
  );


  buf
  g3
  (
    n143,
    n31
  );


  not
  g4
  (
    n161,
    n31
  );


  buf
  g5
  (
    n80,
    n31
  );


  not
  g6
  (
    n84,
    n13
  );


  buf
  g7
  (
    n60,
    n5
  );


  buf
  g8
  (
    n171,
    n35
  );


  buf
  g9
  (
    n91,
    n6
  );


  buf
  g10
  (
    n89,
    n36
  );


  not
  g11
  (
    n131,
    n2
  );


  buf
  g12
  (
    n147,
    n12
  );


  not
  g13
  (
    n132,
    n30
  );


  not
  g14
  (
    KeyWire_0_0,
    n22
  );


  not
  g15
  (
    n102,
    n27
  );


  not
  g16
  (
    n148,
    n13
  );


  buf
  g17
  (
    n93,
    n18
  );


  not
  g18
  (
    n74,
    n14
  );


  not
  g19
  (
    n153,
    n10
  );


  buf
  g20
  (
    n55,
    n12
  );


  not
  g21
  (
    n160,
    n7
  );


  not
  g22
  (
    n77,
    n37
  );


  buf
  g23
  (
    n92,
    n29
  );


  buf
  g24
  (
    n70,
    n8
  );


  buf
  g25
  (
    n69,
    n21
  );


  buf
  g26
  (
    n157,
    n5
  );


  buf
  g27
  (
    n62,
    n15
  );


  buf
  g28
  (
    n56,
    n28
  );


  buf
  g29
  (
    n122,
    n27
  );


  buf
  g30
  (
    n75,
    n14
  );


  not
  g31
  (
    n96,
    n15
  );


  not
  g32
  (
    n126,
    n20
  );


  buf
  g33
  (
    n94,
    n24
  );


  buf
  g34
  (
    n169,
    n27
  );


  buf
  g35
  (
    n152,
    n25
  );


  not
  g36
  (
    n53,
    n26
  );


  not
  g37
  (
    n124,
    n29
  );


  not
  g38
  (
    n127,
    n19
  );


  buf
  g39
  (
    n177,
    n33
  );


  not
  g40
  (
    n142,
    n20
  );


  buf
  g41
  (
    n64,
    n8
  );


  not
  g42
  (
    n82,
    n24
  );


  buf
  g43
  (
    n117,
    n28
  );


  buf
  g44
  (
    n111,
    n33
  );


  not
  g45
  (
    n166,
    n31
  );


  not
  g46
  (
    n167,
    n32
  );


  buf
  g47
  (
    n46,
    n11
  );


  not
  g48
  (
    n158,
    n13
  );


  not
  g49
  (
    n65,
    n23
  );


  not
  g50
  (
    n57,
    n17
  );


  not
  g51
  (
    n43,
    n26
  );


  buf
  g52
  (
    n134,
    n7
  );


  not
  g53
  (
    n83,
    n30
  );


  buf
  g54
  (
    n86,
    n4
  );


  buf
  g55
  (
    n49,
    n36
  );


  buf
  g56
  (
    n130,
    n16
  );


  not
  g57
  (
    n100,
    n34
  );


  not
  g58
  (
    n144,
    n23
  );


  buf
  g59
  (
    n163,
    n35
  );


  not
  g60
  (
    n165,
    n6
  );


  not
  g61
  (
    n72,
    n19
  );


  buf
  g62
  (
    n50,
    n18
  );


  buf
  g63
  (
    n121,
    n10
  );


  not
  g64
  (
    n112,
    n14
  );


  buf
  g65
  (
    n155,
    n20
  );


  not
  g66
  (
    n42,
    n25
  );


  buf
  g67
  (
    n170,
    n33
  );


  buf
  g68
  (
    n78,
    n7
  );


  buf
  g69
  (
    n99,
    n23
  );


  not
  g70
  (
    n120,
    n9
  );


  buf
  g71
  (
    n145,
    n9
  );


  not
  g72
  (
    n61,
    n22
  );


  buf
  g73
  (
    n41,
    n10
  );


  not
  g74
  (
    n175,
    n4
  );


  not
  g75
  (
    n71,
    n37
  );


  buf
  g76
  (
    n51,
    n8
  );


  not
  g77
  (
    n151,
    n12
  );


  not
  g78
  (
    n140,
    n15
  );


  not
  g79
  (
    n159,
    n28
  );


  not
  g80
  (
    n137,
    n19
  );


  not
  g81
  (
    n114,
    n5
  );


  not
  g82
  (
    n81,
    n28
  );


  not
  g83
  (
    n44,
    n16
  );


  buf
  g84
  (
    n150,
    n15
  );


  buf
  g85
  (
    n59,
    n26
  );


  buf
  g86
  (
    n164,
    n35
  );


  buf
  g87
  (
    n101,
    n25
  );


  buf
  g88
  (
    n156,
    n23
  );


  not
  g89
  (
    n136,
    n17
  );


  buf
  g90
  (
    n76,
    n21
  );


  buf
  g91
  (
    n67,
    n14
  );


  not
  g92
  (
    n129,
    n19
  );


  buf
  g93
  (
    n107,
    n32
  );


  not
  g94
  (
    n146,
    n8
  );


  buf
  g95
  (
    n118,
    n36
  );


  buf
  g96
  (
    n97,
    n5
  );


  not
  g97
  (
    n104,
    n11
  );


  buf
  g98
  (
    n48,
    n32
  );


  buf
  g99
  (
    n162,
    n33
  );


  not
  g100
  (
    n110,
    n3
  );


  buf
  g101
  (
    n172,
    n17
  );


  buf
  g102
  (
    n154,
    n27
  );


  not
  g103
  (
    n68,
    n24
  );


  not
  g104
  (
    n52,
    n13
  );


  buf
  g105
  (
    n103,
    n34
  );


  buf
  g106
  (
    n40,
    n34
  );


  not
  g107
  (
    n58,
    n16
  );


  buf
  g108
  (
    n79,
    n34
  );


  buf
  g109
  (
    n125,
    n21
  );


  buf
  g110
  (
    n135,
    n9
  );


  buf
  g111
  (
    n173,
    n7
  );


  not
  g112
  (
    n63,
    n22
  );


  not
  g113
  (
    n133,
    n37
  );


  not
  g114
  (
    KeyWire_0_18,
    n20
  );


  buf
  g115
  (
    n115,
    n21
  );


  buf
  g116
  (
    n54,
    n18
  );


  not
  g117
  (
    n106,
    n6
  );


  buf
  g118
  (
    n119,
    n11
  );


  not
  g119
  (
    n88,
    n29
  );


  not
  g120
  (
    n128,
    n12
  );


  not
  g121
  (
    n108,
    n30
  );


  not
  g122
  (
    n149,
    n11
  );


  not
  g123
  (
    n105,
    n4
  );


  not
  g124
  (
    n116,
    n17
  );


  buf
  g125
  (
    n123,
    n22
  );


  buf
  g126
  (
    n139,
    n10
  );


  buf
  g127
  (
    KeyWire_0_9,
    n6
  );


  buf
  g128
  (
    n138,
    n1
  );


  not
  g129
  (
    n98,
    n24
  );


  not
  g130
  (
    n73,
    n29
  );


  not
  g131
  (
    n109,
    n25
  );


  buf
  g132
  (
    n87,
    n26
  );


  not
  g133
  (
    n66,
    n36
  );


  not
  g134
  (
    n113,
    n35
  );


  not
  g135
  (
    n95,
    n9
  );


  not
  g136
  (
    n176,
    n30
  );


  not
  g137
  (
    n85,
    n18
  );


  buf
  g138
  (
    n396,
    n148
  );


  buf
  g139
  (
    n392,
    n58
  );


  buf
  g140
  (
    n362,
    n120
  );


  not
  g141
  (
    n370,
    n135
  );


  buf
  g142
  (
    n301,
    n92
  );


  not
  g143
  (
    n277,
    n46
  );


  buf
  g144
  (
    n343,
    n94
  );


  buf
  g145
  (
    n389,
    n149
  );


  not
  g146
  (
    n286,
    n49
  );


  not
  g147
  (
    n347,
    n156
  );


  buf
  g148
  (
    n247,
    n48
  );


  buf
  g149
  (
    n278,
    n95
  );


  buf
  g150
  (
    n195,
    n42
  );


  buf
  g151
  (
    n365,
    n159
  );


  buf
  g152
  (
    n284,
    n122
  );


  not
  g153
  (
    n314,
    n164
  );


  buf
  g154
  (
    n271,
    n74
  );


  not
  g155
  (
    n291,
    n160
  );


  not
  g156
  (
    n242,
    n91
  );


  not
  g157
  (
    n225,
    n163
  );


  buf
  g158
  (
    n191,
    n136
  );


  buf
  g159
  (
    n305,
    n142
  );


  buf
  g160
  (
    n182,
    n133
  );


  not
  g161
  (
    n267,
    n169
  );


  not
  g162
  (
    n212,
    n158
  );


  not
  g163
  (
    n299,
    n172
  );


  not
  g164
  (
    n334,
    n170
  );


  not
  g165
  (
    n315,
    n153
  );


  buf
  g166
  (
    n394,
    n128
  );


  not
  g167
  (
    n214,
    n173
  );


  not
  g168
  (
    n356,
    n96
  );


  buf
  g169
  (
    n261,
    n146
  );


  not
  g170
  (
    n378,
    n154
  );


  not
  g171
  (
    n197,
    n61
  );


  not
  g172
  (
    n223,
    n72
  );


  not
  g173
  (
    n241,
    n68
  );


  not
  g174
  (
    n181,
    n139
  );


  not
  g175
  (
    n338,
    n93
  );


  buf
  g176
  (
    n279,
    n137
  );


  not
  g177
  (
    n254,
    n117
  );


  not
  g178
  (
    n335,
    n100
  );


  buf
  g179
  (
    n388,
    n162
  );


  buf
  g180
  (
    n207,
    n173
  );


  buf
  g181
  (
    n228,
    n81
  );


  not
  g182
  (
    n302,
    n112
  );


  buf
  g183
  (
    n262,
    n157
  );


  not
  g184
  (
    n339,
    n102
  );


  buf
  g185
  (
    n382,
    n90
  );


  not
  g186
  (
    n189,
    n89
  );


  buf
  g187
  (
    n219,
    n43
  );


  buf
  g188
  (
    n344,
    n173
  );


  buf
  g189
  (
    n321,
    n153
  );


  not
  g190
  (
    n239,
    n111
  );


  buf
  g191
  (
    n198,
    n131
  );


  buf
  g192
  (
    n329,
    n40
  );


  buf
  g193
  (
    n345,
    n163
  );


  buf
  g194
  (
    n250,
    n41
  );


  buf
  g195
  (
    n381,
    n126
  );


  not
  g196
  (
    n213,
    n54
  );


  buf
  g197
  (
    n310,
    n162
  );


  not
  g198
  (
    n357,
    n156
  );


  not
  g199
  (
    n243,
    n147
  );


  buf
  g200
  (
    n322,
    n110
  );


  buf
  g201
  (
    n319,
    n80
  );


  not
  g202
  (
    n235,
    n51
  );


  buf
  g203
  (
    n289,
    n108
  );


  buf
  g204
  (
    n324,
    n151
  );


  not
  g205
  (
    n386,
    n154
  );


  not
  g206
  (
    n205,
    n158
  );


  not
  g207
  (
    n202,
    n87
  );


  not
  g208
  (
    n393,
    n167
  );


  buf
  g209
  (
    n367,
    n151
  );


  not
  g210
  (
    n185,
    n167
  );


  not
  g211
  (
    n255,
    n168
  );


  not
  g212
  (
    n265,
    n144
  );


  buf
  g213
  (
    n385,
    n171
  );


  not
  g214
  (
    n320,
    n162
  );


  buf
  g215
  (
    n318,
    n116
  );


  not
  g216
  (
    n337,
    n73
  );


  not
  g217
  (
    n366,
    n157
  );


  buf
  g218
  (
    n309,
    n164
  );


  buf
  g219
  (
    n358,
    n147
  );


  not
  g220
  (
    n364,
    n154
  );


  not
  g221
  (
    n273,
    n159
  );


  buf
  g222
  (
    n300,
    n129
  );


  not
  g223
  (
    n375,
    n150
  );


  buf
  g224
  (
    n374,
    n145
  );


  not
  g225
  (
    n192,
    n99
  );


  buf
  g226
  (
    n208,
    n146
  );


  not
  g227
  (
    n257,
    n121
  );


  buf
  g228
  (
    n281,
    n148
  );


  buf
  g229
  (
    n333,
    n169
  );


  not
  g230
  (
    n361,
    n155
  );


  not
  g231
  (
    n326,
    n167
  );


  not
  g232
  (
    n221,
    n84
  );


  buf
  g233
  (
    n179,
    n155
  );


  buf
  g234
  (
    n360,
    n70
  );


  buf
  g235
  (
    n316,
    n134
  );


  not
  g236
  (
    n246,
    n162
  );


  not
  g237
  (
    n293,
    n165
  );


  buf
  g238
  (
    n288,
    n153
  );


  buf
  g239
  (
    n311,
    n124
  );


  not
  g240
  (
    n351,
    n149
  );


  buf
  g241
  (
    n236,
    n138
  );


  buf
  g242
  (
    n353,
    n152
  );


  buf
  g243
  (
    n234,
    n165
  );


  not
  g244
  (
    n264,
    n161
  );


  not
  g245
  (
    n204,
    n170
  );


  buf
  g246
  (
    n184,
    n82
  );


  not
  g247
  (
    n331,
    n119
  );


  not
  g248
  (
    n325,
    n159
  );


  not
  g249
  (
    n290,
    n168
  );


  not
  g250
  (
    n248,
    n167
  );


  buf
  g251
  (
    n283,
    n160
  );


  buf
  g252
  (
    n256,
    n149
  );


  buf
  g253
  (
    n298,
    n63
  );


  not
  g254
  (
    n317,
    n169
  );


  not
  g255
  (
    n187,
    n163
  );


  buf
  g256
  (
    n194,
    n85
  );


  buf
  g257
  (
    n216,
    n141
  );


  not
  g258
  (
    n210,
    n64
  );


  not
  g259
  (
    n354,
    n148
  );


  buf
  g260
  (
    n297,
    n165
  );


  buf
  g261
  (
    n183,
    n79
  );


  buf
  g262
  (
    n359,
    n107
  );


  not
  g263
  (
    n259,
    n168
  );


  not
  g264
  (
    n231,
    n161
  );


  buf
  g265
  (
    n227,
    n161
  );


  not
  g266
  (
    n268,
    n114
  );


  buf
  g267
  (
    n330,
    n171
  );


  buf
  g268
  (
    n276,
    n154
  );


  buf
  g269
  (
    n395,
    n166
  );


  not
  g270
  (
    n270,
    n113
  );


  buf
  g271
  (
    n296,
    n150
  );


  buf
  g272
  (
    n178,
    n161
  );


  buf
  g273
  (
    n391,
    n148
  );


  buf
  g274
  (
    n253,
    n145
  );


  not
  g275
  (
    n229,
    n171
  );


  buf
  g276
  (
    n368,
    n140
  );


  buf
  g277
  (
    n222,
    n147
  );


  buf
  g278
  (
    n346,
    n150
  );


  not
  g279
  (
    n280,
    n130
  );


  buf
  g280
  (
    n232,
    n155
  );


  not
  g281
  (
    n252,
    n76
  );


  not
  g282
  (
    n312,
    n160
  );


  not
  g283
  (
    n215,
    n147
  );


  buf
  g284
  (
    n307,
    n101
  );


  not
  g285
  (
    n237,
    n86
  );


  not
  g286
  (
    n352,
    n103
  );


  not
  g287
  (
    n275,
    n105
  );


  not
  g288
  (
    n327,
    n127
  );


  not
  g289
  (
    n211,
    n78
  );


  buf
  g290
  (
    n199,
    n71
  );


  not
  g291
  (
    n372,
    n67
  );


  buf
  g292
  (
    n387,
    n160
  );


  not
  g293
  (
    n295,
    n125
  );


  buf
  g294
  (
    n383,
    n146
  );


  buf
  g295
  (
    n218,
    n146
  );


  buf
  g296
  (
    n379,
    n166
  );


  not
  g297
  (
    n233,
    n97
  );


  buf
  g298
  (
    n282,
    n171
  );


  buf
  g299
  (
    n292,
    n173
  );


  buf
  g300
  (
    n203,
    n45
  );


  buf
  g301
  (
    n209,
    n83
  );


  buf
  g302
  (
    n188,
    n59
  );


  not
  g303
  (
    n244,
    n98
  );


  buf
  g304
  (
    n220,
    n152
  );


  not
  g305
  (
    n313,
    n55
  );


  buf
  g306
  (
    n274,
    n169
  );


  not
  g307
  (
    n303,
    n44
  );


  not
  g308
  (
    n190,
    n164
  );


  not
  g309
  (
    n251,
    n123
  );


  not
  g310
  (
    n272,
    n168
  );


  not
  g311
  (
    KeyWire_0_3,
    n164
  );


  not
  g312
  (
    n240,
    n56
  );


  buf
  g313
  (
    n348,
    n66
  );


  buf
  g314
  (
    n230,
    n143
  );


  not
  g315
  (
    n224,
    n149
  );


  buf
  g316
  (
    n308,
    n115
  );


  buf
  g317
  (
    n371,
    n172
  );


  not
  g318
  (
    n390,
    n104
  );


  not
  g319
  (
    n269,
    n65
  );


  buf
  g320
  (
    n200,
    n69
  );


  not
  g321
  (
    n186,
    n62
  );


  buf
  g322
  (
    n397,
    n109
  );


  not
  g323
  (
    n376,
    n75
  );


  buf
  g324
  (
    n332,
    n52
  );


  not
  g325
  (
    n323,
    n155
  );


  buf
  g326
  (
    n369,
    n174
  );


  not
  g327
  (
    n355,
    n88
  );


  buf
  g328
  (
    n380,
    n158
  );


  buf
  g329
  (
    n263,
    n172
  );


  not
  g330
  (
    n363,
    n170
  );


  buf
  g331
  (
    n180,
    n158
  );


  buf
  g332
  (
    n238,
    n163
  );


  buf
  g333
  (
    n193,
    n157
  );


  buf
  g334
  (
    n306,
    n153
  );


  not
  g335
  (
    n350,
    n132
  );


  not
  g336
  (
    n206,
    n166
  );


  not
  g337
  (
    n266,
    n156
  );


  not
  g338
  (
    n196,
    n166
  );


  buf
  g339
  (
    n341,
    n165
  );


  buf
  g340
  (
    n294,
    n150
  );


  buf
  g341
  (
    n249,
    n57
  );


  not
  g342
  (
    n342,
    n152
  );


  not
  g343
  (
    n260,
    n118
  );


  buf
  g344
  (
    n336,
    n152
  );


  buf
  g345
  (
    n226,
    n172
  );


  buf
  g346
  (
    KeyWire_0_13,
    n159
  );


  buf
  g347
  (
    n258,
    n47
  );


  buf
  g348
  (
    n377,
    n106
  );


  not
  g349
  (
    n245,
    n151
  );


  buf
  g350
  (
    n287,
    n151
  );


  buf
  g351
  (
    n304,
    n156
  );


  buf
  g352
  (
    n384,
    n157
  );


  not
  g353
  (
    n340,
    n50
  );


  not
  g354
  (
    n217,
    n77
  );


  buf
  g355
  (
    n201,
    n53
  );


  buf
  g356
  (
    n373,
    n60
  );


  not
  g357
  (
    n285,
    n170
  );


  not
  g358
  (
    n715,
    n301
  );


  buf
  g359
  (
    n779,
    n193
  );


  not
  g360
  (
    n590,
    n263
  );


  buf
  g361
  (
    n667,
    n292
  );


  not
  g362
  (
    n569,
    n197
  );


  not
  g363
  (
    n625,
    n349
  );


  buf
  g364
  (
    n520,
    n350
  );


  not
  g365
  (
    n553,
    n271
  );


  buf
  g366
  (
    n435,
    n296
  );


  not
  g367
  (
    n506,
    n192
  );


  not
  g368
  (
    n444,
    n298
  );


  not
  g369
  (
    n863,
    n265
  );


  buf
  g370
  (
    n813,
    n386
  );


  not
  g371
  (
    n727,
    n312
  );


  buf
  g372
  (
    n1041,
    n315
  );


  buf
  g373
  (
    n414,
    n192
  );


  not
  g374
  (
    n424,
    n392
  );


  buf
  g375
  (
    n833,
    n184
  );


  not
  g376
  (
    n891,
    n259
  );


  not
  g377
  (
    n769,
    n297
  );


  not
  g378
  (
    n649,
    n364
  );


  buf
  g379
  (
    n743,
    n367
  );


  not
  g380
  (
    n449,
    n179
  );


  not
  g381
  (
    n431,
    n211
  );


  buf
  g382
  (
    n1042,
    n239
  );


  buf
  g383
  (
    n636,
    n390
  );


  buf
  g384
  (
    n1027,
    n260
  );


  buf
  g385
  (
    n918,
    n183
  );


  not
  g386
  (
    n934,
    n248
  );


  buf
  g387
  (
    n1014,
    n178
  );


  buf
  g388
  (
    n1015,
    n256
  );


  not
  g389
  (
    n429,
    n202
  );


  buf
  g390
  (
    n648,
    n302
  );


  buf
  g391
  (
    n706,
    n352
  );


  buf
  g392
  (
    n895,
    n367
  );


  not
  g393
  (
    n1021,
    n257
  );


  not
  g394
  (
    n577,
    n243
  );


  not
  g395
  (
    n407,
    n306
  );


  buf
  g396
  (
    n1005,
    n316
  );


  buf
  g397
  (
    n929,
    n254
  );


  not
  g398
  (
    n794,
    n277
  );


  not
  g399
  (
    n678,
    n284
  );


  buf
  g400
  (
    n995,
    n327
  );


  buf
  g401
  (
    n511,
    n238
  );


  not
  g402
  (
    KeyWire_0_30,
    n335
  );


  not
  g403
  (
    n997,
    n254
  );


  not
  g404
  (
    n627,
    n391
  );


  not
  g405
  (
    n544,
    n306
  );


  not
  g406
  (
    n482,
    n243
  );


  buf
  g407
  (
    n527,
    n207
  );


  buf
  g408
  (
    n723,
    n197
  );


  buf
  g409
  (
    n475,
    n264
  );


  buf
  g410
  (
    n879,
    n389
  );


  buf
  g411
  (
    n717,
    n206
  );


  buf
  g412
  (
    n748,
    n246
  );


  not
  g413
  (
    n543,
    n263
  );


  not
  g414
  (
    n848,
    n217
  );


  buf
  g415
  (
    n865,
    n396
  );


  not
  g416
  (
    n498,
    n295
  );


  not
  g417
  (
    n658,
    n231
  );


  buf
  g418
  (
    n812,
    n212
  );


  not
  g419
  (
    n936,
    n227
  );


  not
  g420
  (
    n808,
    n305
  );


  buf
  g421
  (
    n824,
    n252
  );


  not
  g422
  (
    n840,
    n251
  );


  buf
  g423
  (
    n857,
    n178
  );


  buf
  g424
  (
    n476,
    n341
  );


  buf
  g425
  (
    n460,
    n205
  );


  buf
  g426
  (
    n613,
    n308
  );


  not
  g427
  (
    n508,
    n279
  );


  not
  g428
  (
    n841,
    n383
  );


  not
  g429
  (
    n835,
    n319
  );


  not
  g430
  (
    n777,
    n310
  );


  buf
  g431
  (
    n898,
    n268
  );


  not
  g432
  (
    n878,
    n397
  );


  buf
  g433
  (
    n797,
    n383
  );


  buf
  g434
  (
    n581,
    n283
  );


  buf
  g435
  (
    n599,
    n229
  );


  not
  g436
  (
    n602,
    n330
  );


  buf
  g437
  (
    n849,
    n367
  );


  not
  g438
  (
    n593,
    n267
  );


  buf
  g439
  (
    n826,
    n228
  );


  buf
  g440
  (
    n643,
    n240
  );


  not
  g441
  (
    n908,
    n247
  );


  not
  g442
  (
    n564,
    n256
  );


  buf
  g443
  (
    n888,
    n250
  );


  not
  g444
  (
    n696,
    n219
  );


  buf
  g445
  (
    n802,
    n319
  );


  not
  g446
  (
    n418,
    n393
  );


  buf
  g447
  (
    n950,
    n353
  );


  not
  g448
  (
    n796,
    n234
  );


  not
  g449
  (
    n529,
    n315
  );


  not
  g450
  (
    n585,
    n391
  );


  not
  g451
  (
    n647,
    n392
  );


  not
  g452
  (
    n746,
    n373
  );


  not
  g453
  (
    n709,
    n237
  );


  buf
  g454
  (
    n839,
    n273
  );


  buf
  g455
  (
    n832,
    n378
  );


  not
  g456
  (
    n959,
    n269
  );


  not
  g457
  (
    n881,
    n238
  );


  not
  g458
  (
    n909,
    n239
  );


  not
  g459
  (
    n586,
    n321
  );


  not
  g460
  (
    n1046,
    n356
  );


  buf
  g461
  (
    n838,
    n282
  );


  buf
  g462
  (
    n622,
    n275
  );


  not
  g463
  (
    n971,
    n366
  );


  not
  g464
  (
    n1010,
    n251
  );


  not
  g465
  (
    n740,
    n240
  );


  buf
  g466
  (
    n415,
    n185
  );


  not
  g467
  (
    n861,
    n363
  );


  buf
  g468
  (
    n720,
    n274
  );


  buf
  g469
  (
    n912,
    n314
  );


  buf
  g470
  (
    n547,
    n333
  );


  buf
  g471
  (
    n651,
    n376
  );


  buf
  g472
  (
    n836,
    n324
  );


  not
  g473
  (
    n922,
    n301
  );


  not
  g474
  (
    n781,
    n275
  );


  buf
  g475
  (
    n852,
    n189
  );


  not
  g476
  (
    n1056,
    n237
  );


  buf
  g477
  (
    n565,
    n226
  );


  not
  g478
  (
    n481,
    n386
  );


  buf
  g479
  (
    n489,
    n181
  );


  buf
  g480
  (
    n983,
    n320
  );


  buf
  g481
  (
    n919,
    n397
  );


  buf
  g482
  (
    n722,
    n199
  );


  buf
  g483
  (
    n1020,
    n253
  );


  not
  g484
  (
    n550,
    n379
  );


  not
  g485
  (
    n731,
    n222
  );


  not
  g486
  (
    n539,
    n199
  );


  not
  g487
  (
    n528,
    n214
  );


  not
  g488
  (
    n710,
    n388
  );


  not
  g489
  (
    n906,
    n205
  );


  buf
  g490
  (
    n662,
    n376
  );


  not
  g491
  (
    n1007,
    n209
  );


  not
  g492
  (
    n1053,
    n250
  );


  not
  g493
  (
    n533,
    n323
  );


  buf
  g494
  (
    n799,
    n325
  );


  not
  g495
  (
    n583,
    n288
  );


  buf
  g496
  (
    n432,
    n191
  );


  not
  g497
  (
    n611,
    n393
  );


  not
  g498
  (
    n792,
    n372
  );


  buf
  g499
  (
    n608,
    n278
  );


  buf
  g500
  (
    n981,
    n233
  );


  not
  g501
  (
    n1019,
    n340
  );


  buf
  g502
  (
    n409,
    n178
  );


  not
  g503
  (
    n1052,
    n295
  );


  buf
  g504
  (
    n855,
    n360
  );


  buf
  g505
  (
    n1045,
    n286
  );


  not
  g506
  (
    n567,
    n230
  );


  buf
  g507
  (
    n926,
    n244
  );


  buf
  g508
  (
    n921,
    n270
  );


  buf
  g509
  (
    n478,
    n342
  );


  not
  g510
  (
    n523,
    n283
  );


  not
  g511
  (
    n494,
    n394
  );


  not
  g512
  (
    n614,
    n188
  );


  not
  g513
  (
    n411,
    n230
  );


  not
  g514
  (
    n837,
    n219
  );


  buf
  g515
  (
    n516,
    n259
  );


  buf
  g516
  (
    n561,
    n369
  );


  not
  g517
  (
    n576,
    n292
  );


  buf
  g518
  (
    n862,
    n180
  );


  buf
  g519
  (
    n421,
    n320
  );


  buf
  g520
  (
    n700,
    n331
  );


  not
  g521
  (
    n635,
    n322
  );


  buf
  g522
  (
    n461,
    n372
  );


  buf
  g523
  (
    n521,
    n224
  );


  not
  g524
  (
    n964,
    n300
  );


  buf
  g525
  (
    n470,
    n284
  );


  not
  g526
  (
    n616,
    n395
  );


  not
  g527
  (
    n745,
    n178
  );


  buf
  g528
  (
    n509,
    n191
  );


  not
  g529
  (
    n440,
    n357
  );


  not
  g530
  (
    n446,
    n222
  );


  not
  g531
  (
    n448,
    n275
  );


  buf
  g532
  (
    n1044,
    n320
  );


  not
  g533
  (
    n554,
    n217
  );


  not
  g534
  (
    n619,
    n257
  );


  buf
  g535
  (
    n659,
    n302
  );


  buf
  g536
  (
    n398,
    n199
  );


  buf
  g537
  (
    n988,
    n365
  );


  buf
  g538
  (
    n970,
    n319
  );


  not
  g539
  (
    n692,
    n321
  );


  buf
  g540
  (
    n897,
    n341
  );


  buf
  g541
  (
    n853,
    n208
  );


  not
  g542
  (
    n755,
    n396
  );


  not
  g543
  (
    n699,
    n337
  );


  not
  g544
  (
    n677,
    n304
  );


  buf
  g545
  (
    n1000,
    n285
  );


  not
  g546
  (
    n454,
    n356
  );


  buf
  g547
  (
    n707,
    n305
  );


  not
  g548
  (
    n491,
    n289
  );


  buf
  g549
  (
    n675,
    n355
  );


  not
  g550
  (
    n977,
    n193
  );


  not
  g551
  (
    n534,
    n243
  );


  buf
  g552
  (
    n1058,
    n366
  );


  not
  g553
  (
    n526,
    n186
  );


  buf
  g554
  (
    n883,
    n395
  );


  not
  g555
  (
    n472,
    n372
  );


  buf
  g556
  (
    n473,
    n233
  );


  not
  g557
  (
    n428,
    n241
  );


  buf
  g558
  (
    n546,
    n384
  );


  buf
  g559
  (
    n1036,
    n377
  );


  buf
  g560
  (
    n538,
    n255
  );


  buf
  g561
  (
    n1009,
    n265
  );


  buf
  g562
  (
    n517,
    n311
  );


  not
  g563
  (
    n789,
    n377
  );


  not
  g564
  (
    n673,
    n223
  );


  not
  g565
  (
    n525,
    n209
  );


  buf
  g566
  (
    n617,
    n302
  );


  not
  g567
  (
    n400,
    n358
  );


  not
  g568
  (
    n633,
    n342
  );


  not
  g569
  (
    n917,
    n246
  );


  not
  g570
  (
    n939,
    n289
  );


  not
  g571
  (
    n920,
    n347
  );


  not
  g572
  (
    n656,
    n252
  );


  buf
  g573
  (
    n911,
    n299
  );


  buf
  g574
  (
    n626,
    n280
  );


  buf
  g575
  (
    n930,
    n295
  );


  not
  g576
  (
    n637,
    n260
  );


  buf
  g577
  (
    n856,
    n194
  );


  buf
  g578
  (
    n902,
    n332
  );


  buf
  g579
  (
    n828,
    n282
  );


  not
  g580
  (
    n843,
    n380
  );


  not
  g581
  (
    n782,
    n389
  );


  not
  g582
  (
    n1011,
    n212
  );


  not
  g583
  (
    n725,
    n220
  );


  not
  g584
  (
    n864,
    n338
  );


  not
  g585
  (
    n992,
    n379
  );


  buf
  g586
  (
    n890,
    n328
  );


  not
  g587
  (
    n702,
    n228
  );


  buf
  g588
  (
    n447,
    n286
  );


  buf
  g589
  (
    n767,
    n179
  );


  buf
  g590
  (
    n773,
    n339
  );


  buf
  g591
  (
    n969,
    n219
  );


  not
  g592
  (
    n598,
    n371
  );


  not
  g593
  (
    n882,
    n273
  );


  buf
  g594
  (
    n660,
    n340
  );


  not
  g595
  (
    n935,
    n222
  );


  not
  g596
  (
    n972,
    n314
  );


  buf
  g597
  (
    n805,
    n312
  );


  not
  g598
  (
    n504,
    n218
  );


  not
  g599
  (
    n697,
    n240
  );


  buf
  g600
  (
    n798,
    n349
  );


  buf
  g601
  (
    n433,
    n285
  );


  buf
  g602
  (
    n910,
    n378
  );


  buf
  g603
  (
    n962,
    n307
  );


  not
  g604
  (
    n500,
    n235
  );


  buf
  g605
  (
    n928,
    n273
  );


  not
  g606
  (
    n787,
    n204
  );


  buf
  g607
  (
    n994,
    n221
  );


  not
  g608
  (
    n750,
    n290
  );


  buf
  g609
  (
    n519,
    n224
  );


  not
  g610
  (
    n795,
    n182
  );


  buf
  g611
  (
    n819,
    n352
  );


  not
  g612
  (
    n445,
    n204
  );


  buf
  g613
  (
    n587,
    n232
  );


  buf
  g614
  (
    KeyWire_0_15,
    n334
  );


  not
  g615
  (
    n427,
    n393
  );


  not
  g616
  (
    n634,
    n264
  );


  not
  g617
  (
    n718,
    n267
  );


  buf
  g618
  (
    n416,
    n388
  );


  buf
  g619
  (
    n495,
    n311
  );


  not
  g620
  (
    n987,
    n180
  );


  buf
  g621
  (
    n595,
    n370
  );


  not
  g622
  (
    n542,
    n245
  );


  buf
  g623
  (
    n899,
    n213
  );


  not
  g624
  (
    n548,
    n346
  );


  not
  g625
  (
    n701,
    n336
  );


  not
  g626
  (
    n758,
    n208
  );


  not
  g627
  (
    n893,
    n332
  );


  not
  g628
  (
    n744,
    n243
  );


  buf
  g629
  (
    n557,
    n272
  );


  not
  g630
  (
    n681,
    n270
  );


  buf
  g631
  (
    n483,
    n303
  );


  buf
  g632
  (
    KeyWire_0_6,
    n211
  );


  buf
  g633
  (
    n632,
    n228
  );


  buf
  g634
  (
    n698,
    n203
  );


  buf
  g635
  (
    n612,
    n246
  );


  buf
  g636
  (
    n621,
    n354
  );


  not
  g637
  (
    n628,
    n337
  );


  not
  g638
  (
    n484,
    n252
  );


  not
  g639
  (
    n674,
    n350
  );


  buf
  g640
  (
    n721,
    n263
  );


  buf
  g641
  (
    n426,
    n353
  );


  not
  g642
  (
    n954,
    n264
  );


  buf
  g643
  (
    n846,
    n303
  );


  not
  g644
  (
    n873,
    n206
  );


  not
  g645
  (
    n676,
    n215
  );


  buf
  g646
  (
    n610,
    n278
  );


  buf
  g647
  (
    n584,
    n242
  );


  buf
  g648
  (
    KeyWire_0_21,
    n310
  );


  not
  g649
  (
    n1034,
    n223
  );


  buf
  g650
  (
    n640,
    n287
  );


  buf
  g651
  (
    n459,
    n273
  );


  not
  g652
  (
    n502,
    n269
  );


  buf
  g653
  (
    n563,
    n371
  );


  buf
  g654
  (
    n984,
    n195
  );


  not
  g655
  (
    n742,
    n220
  );


  buf
  g656
  (
    KeyWire_0_16,
    n357
  );


  buf
  g657
  (
    n1012,
    n198
  );


  not
  g658
  (
    n671,
    n323
  );


  buf
  g659
  (
    n624,
    n258
  );


  not
  g660
  (
    n940,
    n208
  );


  buf
  g661
  (
    n747,
    n382
  );


  buf
  g662
  (
    KeyWire_0_31,
    n277
  );


  buf
  g663
  (
    n993,
    n362
  );


  not
  g664
  (
    n916,
    n278
  );


  buf
  g665
  (
    n809,
    n231
  );


  not
  g666
  (
    n961,
    n235
  );


  buf
  g667
  (
    n947,
    n328
  );


  not
  g668
  (
    n847,
    n271
  );


  not
  g669
  (
    n804,
    n264
  );


  buf
  g670
  (
    n915,
    n224
  );


  not
  g671
  (
    n402,
    n193
  );


  buf
  g672
  (
    n594,
    n358
  );


  not
  g673
  (
    n1002,
    n335
  );


  buf
  g674
  (
    n949,
    n358
  );


  buf
  g675
  (
    n403,
    n186
  );


  not
  g676
  (
    n946,
    n271
  );


  not
  g677
  (
    n726,
    n368
  );


  buf
  g678
  (
    n457,
    n306
  );


  not
  g679
  (
    n914,
    n293
  );


  not
  g680
  (
    n1028,
    n229
  );


  buf
  g681
  (
    n800,
    n332
  );


  not
  g682
  (
    n765,
    n306
  );


  buf
  g683
  (
    n412,
    n307
  );


  buf
  g684
  (
    n859,
    n342
  );


  not
  g685
  (
    n965,
    n310
  );


  buf
  g686
  (
    n844,
    n386
  );


  not
  g687
  (
    n686,
    n221
  );


  not
  g688
  (
    n401,
    n203
  );


  not
  g689
  (
    n762,
    n336
  );


  buf
  g690
  (
    n752,
    n348
  );


  not
  g691
  (
    n514,
    n336
  );


  not
  g692
  (
    n945,
    n345
  );


  buf
  g693
  (
    n575,
    n388
  );


  not
  g694
  (
    n1035,
    n262
  );


  not
  g695
  (
    n596,
    n274
  );


  not
  g696
  (
    n605,
    n233
  );


  buf
  g697
  (
    n406,
    n359
  );


  buf
  g698
  (
    n405,
    n378
  );


  not
  g699
  (
    n708,
    n211
  );


  not
  g700
  (
    n501,
    n326
  );


  buf
  g701
  (
    n486,
    n385
  );


  not
  g702
  (
    n803,
    n255
  );


  not
  g703
  (
    n763,
    n298
  );


  buf
  g704
  (
    n786,
    n195
  );


  buf
  g705
  (
    KeyWire_0_5,
    n234
  );


  not
  g706
  (
    n927,
    n225
  );


  buf
  g707
  (
    n887,
    n247
  );


  buf
  g708
  (
    n513,
    n384
  );


  not
  g709
  (
    n704,
    n314
  );


  not
  g710
  (
    n810,
    n387
  );


  not
  g711
  (
    n785,
    n232
  );


  not
  g712
  (
    n738,
    n308
  );


  buf
  g713
  (
    n858,
    n371
  );


  not
  g714
  (
    n817,
    n343
  );


  not
  g715
  (
    n1043,
    n217
  );


  not
  g716
  (
    n733,
    n383
  );


  not
  g717
  (
    n1026,
    n326
  );


  not
  g718
  (
    n452,
    n301
  );


  buf
  g719
  (
    n467,
    n346
  );


  not
  g720
  (
    n688,
    n234
  );


  not
  g721
  (
    KeyWire_0_7,
    n260
  );


  buf
  g722
  (
    n991,
    n325
  );


  not
  g723
  (
    n854,
    n355
  );


  not
  g724
  (
    n531,
    n322
  );


  buf
  g725
  (
    n772,
    n205
  );


  not
  g726
  (
    n820,
    n369
  );


  not
  g727
  (
    n463,
    n309
  );


  not
  g728
  (
    n978,
    n336
  );


  not
  g729
  (
    n1047,
    n257
  );


  not
  g730
  (
    n474,
    n269
  );


  buf
  g731
  (
    n724,
    n341
  );


  not
  g732
  (
    KeyWire_0_24,
    n378
  );


  not
  g733
  (
    n712,
    n374
  );


  buf
  g734
  (
    n1008,
    n331
  );


  not
  g735
  (
    n1055,
    n316
  );


  not
  g736
  (
    n597,
    n345
  );


  not
  g737
  (
    n668,
    n183
  );


  not
  g738
  (
    n591,
    n261
  );


  not
  g739
  (
    n572,
    n300
  );


  not
  g740
  (
    n1017,
    n338
  );


  buf
  g741
  (
    n540,
    n215
  );


  buf
  g742
  (
    n822,
    n229
  );


  buf
  g743
  (
    n477,
    n250
  );


  buf
  g744
  (
    n979,
    n183
  );


  not
  g745
  (
    n791,
    n196
  );


  buf
  g746
  (
    n573,
    n393
  );


  buf
  g747
  (
    n552,
    n383
  );


  not
  g748
  (
    n653,
    n325
  );


  not
  g749
  (
    n719,
    n291
  );


  not
  g750
  (
    n682,
    n292
  );


  buf
  g751
  (
    n754,
    n364
  );


  buf
  g752
  (
    n904,
    n237
  );


  not
  g753
  (
    n937,
    n194
  );


  buf
  g754
  (
    n757,
    n370
  );


  buf
  g755
  (
    n793,
    n198
  );


  not
  g756
  (
    n1033,
    n246
  );


  buf
  g757
  (
    n751,
    n208
  );


  not
  g758
  (
    n644,
    n214
  );


  not
  g759
  (
    n884,
    n270
  );


  buf
  g760
  (
    n963,
    n291
  );


  not
  g761
  (
    n530,
    n354
  );


  not
  g762
  (
    n960,
    n187
  );


  buf
  g763
  (
    n980,
    n296
  );


  buf
  g764
  (
    n1048,
    n324
  );


  not
  g765
  (
    KeyWire_0_2,
    n317
  );


  not
  g766
  (
    n689,
    n206
  );


  buf
  g767
  (
    n571,
    n196
  );


  buf
  g768
  (
    n766,
    n366
  );


  buf
  g769
  (
    n623,
    n361
  );


  not
  g770
  (
    n739,
    n392
  );


  not
  g771
  (
    n771,
    n256
  );


  buf
  g772
  (
    n680,
    n299
  );


  not
  g773
  (
    n652,
    n304
  );


  buf
  g774
  (
    n600,
    n241
  );


  buf
  g775
  (
    n1050,
    n321
  );


  not
  g776
  (
    n430,
    n396
  );


  buf
  g777
  (
    n549,
    n203
  );


  buf
  g778
  (
    n986,
    n190
  );


  buf
  g779
  (
    n580,
    n370
  );


  buf
  g780
  (
    n880,
    n329
  );


  not
  g781
  (
    n574,
    n353
  );


  buf
  g782
  (
    n606,
    n337
  );


  not
  g783
  (
    n641,
    n365
  );


  not
  g784
  (
    n434,
    n233
  );


  buf
  g785
  (
    n455,
    n376
  );


  not
  g786
  (
    n1025,
    n202
  );


  not
  g787
  (
    n734,
    n182
  );


  buf
  g788
  (
    n737,
    n280
  );


  buf
  g789
  (
    n441,
    n283
  );


  not
  g790
  (
    n685,
    n239
  );


  not
  g791
  (
    n556,
    n337
  );


  buf
  g792
  (
    n691,
    n363
  );


  not
  g793
  (
    n933,
    n268
  );


  buf
  g794
  (
    n955,
    n385
  );


  not
  g795
  (
    n818,
    n236
  );


  not
  g796
  (
    n438,
    n293
  );


  not
  g797
  (
    n876,
    n346
  );


  not
  g798
  (
    n578,
    n188
  );


  not
  g799
  (
    n604,
    n184
  );


  not
  g800
  (
    n631,
    n394
  );


  not
  g801
  (
    n1040,
    n209
  );


  buf
  g802
  (
    n907,
    n333
  );


  not
  g803
  (
    n825,
    n290
  );


  not
  g804
  (
    n664,
    n202
  );


  not
  g805
  (
    n996,
    n339
  );


  not
  g806
  (
    n823,
    n276
  );


  buf
  g807
  (
    n753,
    n238
  );


  not
  g808
  (
    n872,
    n245
  );


  not
  g809
  (
    n510,
    n365
  );


  buf
  g810
  (
    n518,
    n245
  );


  not
  g811
  (
    n683,
    n216
  );


  not
  g812
  (
    n953,
    n362
  );


  not
  g813
  (
    n1049,
    n358
  );


  buf
  g814
  (
    n666,
    n198
  );


  buf
  g815
  (
    n1032,
    n381
  );


  buf
  g816
  (
    n404,
    n204
  );


  buf
  g817
  (
    n588,
    n352
  );


  not
  g818
  (
    n670,
    n210
  );


  buf
  g819
  (
    n894,
    n222
  );


  buf
  g820
  (
    n776,
    n213
  );


  not
  g821
  (
    n493,
    n375
  );


  not
  g822
  (
    n694,
    n254
  );


  buf
  g823
  (
    n875,
    n363
  );


  not
  g824
  (
    n905,
    n362
  );


  buf
  g825
  (
    n931,
    n309
  );


  not
  g826
  (
    KeyWire_0_11,
    n348
  );


  buf
  g827
  (
    n422,
    n298
  );


  buf
  g828
  (
    n713,
    n312
  );


  not
  g829
  (
    n469,
    n382
  );


  buf
  g830
  (
    n827,
    n260
  );


  not
  g831
  (
    n1018,
    n191
  );


  not
  g832
  (
    n973,
    n196
  );


  buf
  g833
  (
    n638,
    n258
  );


  not
  g834
  (
    n399,
    n197
  );


  buf
  g835
  (
    n437,
    n186
  );


  buf
  g836
  (
    n761,
    n269
  );


  not
  g837
  (
    n480,
    n322
  );


  buf
  g838
  (
    n778,
    n184
  );


  buf
  g839
  (
    n942,
    n265
  );


  not
  g840
  (
    n952,
    n344
  );


  buf
  g841
  (
    n1038,
    n226
  );


  not
  g842
  (
    n989,
    n205
  );


  buf
  g843
  (
    n487,
    n185
  );


  not
  g844
  (
    n439,
    n278
  );


  buf
  g845
  (
    n735,
    n216
  );


  not
  g846
  (
    n545,
    n335
  );


  buf
  g847
  (
    n866,
    n214
  );


  not
  g848
  (
    n1039,
    n202
  );


  buf
  g849
  (
    n741,
    n200
  );


  not
  g850
  (
    n464,
    n375
  );


  buf
  g851
  (
    n496,
    n200
  );


  not
  g852
  (
    n1003,
    n242
  );


  not
  g853
  (
    n537,
    n244
  );


  buf
  g854
  (
    n515,
    n360
  );


  buf
  g855
  (
    n492,
    n218
  );


  buf
  g856
  (
    n886,
    n307
  );


  not
  g857
  (
    n642,
    n287
  );


  buf
  g858
  (
    n885,
    n321
  );


  buf
  g859
  (
    n1024,
    n225
  );


  buf
  g860
  (
    n497,
    n351
  );


  not
  g861
  (
    n589,
    n227
  );


  buf
  g862
  (
    n541,
    n391
  );


  buf
  g863
  (
    n669,
    n284
  );


  not
  g864
  (
    n488,
    n381
  );


  buf
  g865
  (
    n985,
    n285
  );


  buf
  g866
  (
    n975,
    n262
  );


  not
  g867
  (
    n609,
    n242
  );


  not
  g868
  (
    n654,
    n237
  );


  buf
  g869
  (
    n871,
    n226
  );


  not
  g870
  (
    n982,
    n258
  );


  not
  g871
  (
    n788,
    n384
  );


  not
  g872
  (
    n976,
    n254
  );


  not
  g873
  (
    n1022,
    n381
  );


  not
  g874
  (
    n410,
    n193
  );


  buf
  g875
  (
    n684,
    n330
  );


  not
  g876
  (
    n579,
    n296
  );


  not
  g877
  (
    n607,
    n369
  );


  not
  g878
  (
    n568,
    n274
  );


  not
  g879
  (
    n471,
    n357
  );


  not
  g880
  (
    n450,
    n188
  );


  not
  g881
  (
    n672,
    n236
  );


  not
  g882
  (
    n774,
    n360
  );


  buf
  g883
  (
    n913,
    n385
  );


  buf
  g884
  (
    n900,
    n397
  );


  not
  g885
  (
    n522,
    n351
  );


  not
  g886
  (
    n558,
    n211
  );


  buf
  g887
  (
    n941,
    n286
  );


  buf
  g888
  (
    n639,
    n190
  );


  buf
  g889
  (
    n889,
    n187
  );


  not
  g890
  (
    n466,
    n310
  );


  buf
  g891
  (
    n999,
    n353
  );


  not
  g892
  (
    n749,
    n297
  );


  not
  g893
  (
    n821,
    n218
  );


  not
  g894
  (
    n442,
    n374
  );


  not
  g895
  (
    n957,
    n216
  );


  not
  g896
  (
    KeyWire_0_10,
    n236
  );


  not
  g897
  (
    n695,
    n277
  );


  buf
  g898
  (
    n645,
    n384
  );


  not
  g899
  (
    n629,
    n201
  );


  buf
  g900
  (
    n566,
    n207
  );


  not
  g901
  (
    n829,
    n261
  );


  not
  g902
  (
    n990,
    n287
  );


  buf
  g903
  (
    n1030,
    n196
  );


  buf
  g904
  (
    n1013,
    n223
  );


  not
  g905
  (
    n601,
    n389
  );


  buf
  g906
  (
    n1054,
    n268
  );


  buf
  g907
  (
    n968,
    n180
  );


  not
  g908
  (
    n456,
    n346
  );


  buf
  g909
  (
    n998,
    n341
  );


  not
  g910
  (
    n663,
    n333
  );


  buf
  g911
  (
    n592,
    n325
  );


  buf
  g912
  (
    n729,
    n218
  );


  buf
  g913
  (
    n687,
    n214
  );


  buf
  g914
  (
    n1031,
    n228
  );


  not
  g915
  (
    n944,
    n377
  );


  not
  g916
  (
    n732,
    n281
  );


  buf
  g917
  (
    n764,
    n212
  );


  buf
  g918
  (
    n503,
    n181
  );


  not
  g919
  (
    n615,
    n374
  );


  buf
  g920
  (
    n903,
    n187
  );


  not
  g921
  (
    n775,
    n298
  );


  buf
  g922
  (
    n655,
    n294
  );


  not
  g923
  (
    n524,
    n327
  );


  not
  g924
  (
    n1023,
    n272
  );


  not
  g925
  (
    n535,
    n313
  );


  not
  g926
  (
    n559,
    n344
  );


  not
  g927
  (
    n850,
    n357
  );


  not
  g928
  (
    n728,
    n324
  );


  not
  g929
  (
    n618,
    n304
  );


  not
  g930
  (
    n790,
    n281
  );


  buf
  g931
  (
    n967,
    n351
  );


  buf
  g932
  (
    n693,
    n261
  );


  buf
  g933
  (
    n714,
    n207
  );


  not
  g934
  (
    n419,
    n352
  );


  buf
  g935
  (
    n485,
    n179
  );


  not
  g936
  (
    n874,
    n242
  );


  buf
  g937
  (
    n408,
    n354
  );


  buf
  g938
  (
    n436,
    n380
  );


  not
  g939
  (
    n1001,
    n387
  );


  not
  g940
  (
    n815,
    n338
  );


  buf
  g941
  (
    n1037,
    n257
  );


  not
  g942
  (
    n650,
    n355
  );


  buf
  g943
  (
    n924,
    n232
  );


  not
  g944
  (
    n679,
    n297
  );


  not
  g945
  (
    n831,
    n335
  );


  xnor
  g946
  (
    n860,
    n368,
    n397,
    n351,
    n339
  );


  xor
  g947
  (
    n736,
    n290,
    n295,
    n373,
    n230
  );


  nor
  g948
  (
    n560,
    n266,
    n305,
    n380,
    n289
  );


  or
  g949
  (
    n665,
    n290,
    n226,
    n255,
    n302
  );


  nor
  g950
  (
    n834,
    n318,
    n387,
    n207,
    n316
  );


  and
  g951
  (
    n462,
    n198,
    n181,
    n209,
    n253
  );


  nor
  g952
  (
    n458,
    n220,
    n291,
    n203,
    n363
  );


  or
  g953
  (
    n690,
    n230,
    n244,
    n315,
    n251
  );


  or
  g954
  (
    n716,
    n359,
    n345,
    n340,
    n194
  );


  nor
  g955
  (
    n938,
    n241,
    n354,
    n210,
    n280
  );


  xor
  g956
  (
    n505,
    n261,
    n368,
    n227,
    n293
  );


  and
  g957
  (
    n811,
    n389,
    n285,
    n376,
    n314
  );


  xnor
  g958
  (
    n784,
    n326,
    n372,
    n192,
    n267
  );


  or
  g959
  (
    n816,
    n220,
    n251,
    n350,
    n317
  );


  nand
  g960
  (
    n923,
    n225,
    n272,
    n183,
    n255
  );


  xnor
  g961
  (
    n630,
    n309,
    n381,
    n250,
    n268
  );


  or
  g962
  (
    n1006,
    n229,
    n245,
    n348,
    n394
  );


  or
  g963
  (
    n830,
    n394,
    n239,
    n344,
    n395
  );


  or
  g964
  (
    KeyWire_0_19,
    n333,
    n288,
    n247,
    n259
  );


  nor
  g965
  (
    n1016,
    n283,
    n199,
    n281,
    n201
  );


  xnor
  g966
  (
    n479,
    n320,
    n221,
    n343,
    n380
  );


  and
  g967
  (
    n468,
    n331,
    n340,
    n396,
    n364
  );


  nor
  g968
  (
    n925,
    n235,
    n280,
    n329,
    n215
  );


  or
  g969
  (
    n582,
    n181,
    n369,
    n313,
    n185
  );


  or
  g970
  (
    n603,
    n279,
    n390,
    n327,
    n322
  );


  nor
  g971
  (
    n892,
    n263,
    n194,
    n317,
    n299
  );


  and
  g972
  (
    n806,
    n217,
    n329,
    n324,
    n267
  );


  or
  g973
  (
    n867,
    n334,
    n188,
    n215,
    n201
  );


  xnor
  g974
  (
    n512,
    n232,
    n319,
    n249,
    n361
  );


  xor
  g975
  (
    n974,
    n288,
    n359,
    n382,
    n297
  );


  nor
  g976
  (
    n951,
    n266,
    n315,
    n300,
    n391
  );


  xor
  g977
  (
    n760,
    n248,
    n270,
    n249,
    n318
  );


  xor
  g978
  (
    n948,
    n276,
    n216,
    n294,
    n356
  );


  nand
  g979
  (
    n703,
    n265,
    n356,
    n392,
    n362
  );


  nand
  g980
  (
    n1057,
    n360,
    n311,
    n179,
    n332
  );


  or
  g981
  (
    n532,
    n182,
    n291,
    n307,
    n231
  );


  or
  g982
  (
    n759,
    n349,
    n189,
    n326,
    n289
  );


  xor
  g983
  (
    n646,
    n288,
    n374,
    n274,
    n293
  );


  nor
  g984
  (
    n490,
    n390,
    n344,
    n375,
    n189
  );


  xor
  g985
  (
    n413,
    n276,
    n292,
    n190,
    n224
  );


  nand
  g986
  (
    n966,
    n312,
    n191,
    n355,
    n309
  );


  nor
  g987
  (
    n756,
    n195,
    n223,
    n281,
    n316
  );


  xor
  g988
  (
    n1051,
    n338,
    n186,
    n313,
    n249
  );


  nand
  g989
  (
    n851,
    n365,
    n252,
    n238,
    n277
  );


  or
  g990
  (
    n425,
    n359,
    n253,
    n296,
    n367
  );


  nor
  g991
  (
    n555,
    n219,
    n349,
    n386,
    n301
  );


  xnor
  g992
  (
    n451,
    n328,
    n189,
    n347,
    n248
  );


  nor
  g993
  (
    n780,
    n387,
    n266,
    n271,
    n361
  );


  nand
  g994
  (
    n620,
    n258,
    n204,
    n368,
    n262
  );


  xor
  g995
  (
    n814,
    n347,
    n240,
    n279,
    n236
  );


  xor
  g996
  (
    n943,
    n373,
    n190,
    n377,
    n303
  );


  and
  g997
  (
    n870,
    n299,
    n330,
    n347,
    n317
  );


  xnor
  g998
  (
    n499,
    n334,
    n350,
    n328,
    n305
  );


  xnor
  g999
  (
    n869,
    n284,
    n247,
    n327,
    n275
  );


  or
  g1000
  (
    n730,
    n244,
    n375,
    n379,
    n249
  );


  xor
  g1001
  (
    n507,
    n262,
    n379,
    n212,
    n308
  );


  and
  g1002
  (
    n562,
    n323,
    n221,
    n201,
    n180
  );


  or
  g1003
  (
    n845,
    n318,
    n287,
    n342,
    n266
  );


  xor
  g1004
  (
    n661,
    n279,
    n395,
    n256,
    n330
  );


  xor
  g1005
  (
    n453,
    n294,
    n234,
    n390,
    n282
  );


  nand
  g1006
  (
    n877,
    n339,
    n200,
    n231,
    n276
  );


  xor
  g1007
  (
    n1029,
    n388,
    n343,
    n366,
    n385
  );


  xnor
  g1008
  (
    n443,
    n184,
    n294,
    n348,
    n345
  );


  xnor
  g1009
  (
    n423,
    n313,
    n334,
    n311,
    n382
  );


  nor
  g1010
  (
    n705,
    n185,
    n308,
    n323,
    n210
  );


  xnor
  g1011
  (
    KeyWire_0_29,
    n213,
    n225,
    n206,
    n303
  );


  nand
  g1012
  (
    n783,
    n331,
    n182,
    n210,
    n197
  );


  and
  g1013
  (
    n536,
    n282,
    n373,
    n300,
    n371
  );


  xor
  g1014
  (
    n465,
    n253,
    n227,
    n195,
    n272
  );


  nand
  g1015
  (
    n842,
    n213,
    n364,
    n286,
    n248
  );


  xor
  g1016
  (
    n417,
    n329,
    n304,
    n343,
    n259
  );


  xnor
  g1017
  (
    n932,
    n318,
    n241,
    n192,
    n235
  );


  xor
  g1018
  (
    n657,
    n361,
    n200,
    n187,
    n370
  );


  or
  g1019
  (
    n1074,
    n551,
    n457,
    n789,
    n429
  );


  xor
  g1020
  (
    n1085,
    n539,
    n683,
    n840,
    n553
  );


  nand
  g1021
  (
    n1121,
    n529,
    n795,
    n565,
    n451
  );


  xnor
  g1022
  (
    n1172,
    n721,
    n688,
    n643,
    n412
  );


  xnor
  g1023
  (
    n1160,
    n636,
    n908,
    n434,
    n816
  );


  xor
  g1024
  (
    n1153,
    n727,
    n562,
    n824,
    n420
  );


  nand
  g1025
  (
    n1127,
    n768,
    n668,
    n557,
    n530
  );


  nand
  g1026
  (
    n1155,
    n836,
    n411,
    n606,
    n613
  );


  or
  g1027
  (
    n1147,
    n733,
    n750,
    n794,
    n574
  );


  xnor
  g1028
  (
    KeyWire_0_4,
    n588,
    n525,
    n728,
    n575
  );


  xor
  g1029
  (
    n1063,
    n459,
    n738,
    n492,
    n855
  );


  xor
  g1030
  (
    n1099,
    n642,
    n475,
    n659,
    n616
  );


  xnor
  g1031
  (
    n1087,
    n674,
    n497,
    n503,
    n607
  );


  xnor
  g1032
  (
    n1165,
    n630,
    n481,
    n569,
    n909
  );


  nor
  g1033
  (
    n1122,
    n517,
    n414,
    n788,
    n784
  );


  xor
  g1034
  (
    n1175,
    n637,
    n640,
    n549,
    n535
  );


  nor
  g1035
  (
    n1174,
    n604,
    n558,
    n469,
    n678
  );


  and
  g1036
  (
    n1119,
    n744,
    n447,
    n591,
    n596
  );


  nor
  g1037
  (
    n1113,
    n899,
    n473,
    n739,
    n778
  );


  xnor
  g1038
  (
    n1167,
    n566,
    n590,
    n536,
    n452
  );


  xnor
  g1039
  (
    n1126,
    n781,
    n725,
    n737,
    n699
  );


  and
  g1040
  (
    n1186,
    n670,
    n743,
    n443,
    n520
  );


  nor
  g1041
  (
    n1089,
    n560,
    n757,
    n495,
    n809
  );


  or
  g1042
  (
    n1060,
    n792,
    n458,
    n564,
    n639
  );


  xnor
  g1043
  (
    n1073,
    n599,
    n779,
    n409,
    n417
  );


  xor
  g1044
  (
    n1177,
    n680,
    n446,
    n839,
    n532
  );


  or
  g1045
  (
    n1066,
    n405,
    n504,
    n499,
    n759
  );


  xnor
  g1046
  (
    n1136,
    n843,
    n402,
    n505,
    n802
  );


  xnor
  g1047
  (
    n1114,
    n877,
    n518,
    n437,
    n398
  );


  xnor
  g1048
  (
    n1168,
    n449,
    n807,
    n478,
    n825
  );


  nor
  g1049
  (
    n1183,
    n863,
    n658,
    n489,
    n468
  );


  nand
  g1050
  (
    n1094,
    n881,
    n701,
    n498,
    n656
  );


  nor
  g1051
  (
    n1143,
    n718,
    n764,
    n787,
    n598
  );


  nand
  g1052
  (
    n1170,
    n577,
    n521,
    n480,
    n772
  );


  or
  g1053
  (
    n1117,
    n651,
    n780,
    n608,
    n901
  );


  xnor
  g1054
  (
    n1163,
    n769,
    n586,
    n887,
    n399
  );


  xor
  g1055
  (
    n1148,
    n682,
    n485,
    n556,
    n488
  );


  xor
  g1056
  (
    n1071,
    n482,
    n403,
    n477,
    n888
  );


  xnor
  g1057
  (
    n1091,
    n673,
    n775,
    n548,
    n799
  );


  and
  g1058
  (
    n1161,
    n552,
    n430,
    n646,
    n878
  );


  xnor
  g1059
  (
    n1059,
    n634,
    n767,
    n490,
    n770
  );


  nand
  g1060
  (
    n1100,
    n442,
    n421,
    n664,
    n587
  );


  and
  g1061
  (
    n1134,
    n626,
    n568,
    n828,
    n419
  );


  and
  g1062
  (
    n1115,
    n487,
    n423,
    n837,
    n435
  );


  nand
  g1063
  (
    n1065,
    n691,
    n791,
    n461,
    n804
  );


  or
  g1064
  (
    n1109,
    n713,
    n415,
    n818,
    n748
  );


  nor
  g1065
  (
    n1144,
    n486,
    n508,
    n675,
    n669
  );


  xnor
  g1066
  (
    n1101,
    n885,
    n777,
    n582,
    n762
  );


  nor
  g1067
  (
    KeyWire_0_14,
    n677,
    n693,
    n635,
    n666
  );


  xor
  g1068
  (
    n1118,
    n621,
    n709,
    n690,
    n559
  );


  or
  g1069
  (
    n1107,
    n844,
    n722,
    n614,
    n679
  );


  nand
  g1070
  (
    n1124,
    n870,
    n823,
    n662,
    n858
  );


  nand
  g1071
  (
    n1080,
    n796,
    n879,
    n522,
    n790
  );


  xnor
  g1072
  (
    n1083,
    n861,
    n523,
    n502,
    n612
  );


  nor
  g1073
  (
    n1095,
    n627,
    n644,
    n515,
    n864
  );


  xor
  g1074
  (
    n1072,
    n715,
    n745,
    n689,
    n652
  );


  nand
  g1075
  (
    n1108,
    n866,
    n584,
    n544,
    n433
  );


  nor
  g1076
  (
    n1125,
    n625,
    n650,
    n705,
    n852
  );


  xor
  g1077
  (
    n1096,
    n793,
    n413,
    n467,
    n841
  );


  xnor
  g1078
  (
    n1164,
    n883,
    n734,
    n810,
    n550
  );


  xor
  g1079
  (
    n1162,
    n755,
    n814,
    n526,
    n519
  );


  xnor
  g1080
  (
    n1102,
    n661,
    n826,
    n890,
    n835
  );


  and
  g1081
  (
    n1176,
    n660,
    n753,
    n605,
    n867
  );


  or
  g1082
  (
    n1088,
    n479,
    n638,
    n424,
    n506
  );


  xor
  g1083
  (
    n1110,
    n484,
    n404,
    n408,
    n501
  );


  nand
  g1084
  (
    n1152,
    n869,
    n692,
    n578,
    n554
  );


  xnor
  g1085
  (
    n1068,
    n425,
    n533,
    n774,
    n902
  );


  nand
  g1086
  (
    n1184,
    n717,
    n573,
    n712,
    n834
  );


  or
  g1087
  (
    n1082,
    n815,
    n538,
    n724,
    n742
  );


  xnor
  g1088
  (
    n1070,
    n628,
    n454,
    n812,
    n471
  );


  xor
  g1089
  (
    n1141,
    n831,
    n561,
    n821,
    n893
  );


  or
  g1090
  (
    n1185,
    n440,
    n813,
    n543,
    n541
  );


  and
  g1091
  (
    n1106,
    n580,
    n747,
    n401,
    n703
  );


  nor
  g1092
  (
    n1157,
    n882,
    n589,
    n545,
    n464
  );


  nor
  g1093
  (
    n1146,
    n798,
    n624,
    n555,
    n672
  );


  nand
  g1094
  (
    n1064,
    n513,
    n845,
    n862,
    n752
  );


  nor
  g1095
  (
    n1061,
    n681,
    n671,
    n832,
    n460
  );


  nor
  g1096
  (
    n1138,
    n874,
    n428,
    n441,
    n426
  );


  nor
  g1097
  (
    n1062,
    n450,
    n884,
    n524,
    n579
  );


  nand
  g1098
  (
    n1097,
    n763,
    n886,
    n771,
    n811
  );


  xor
  g1099
  (
    n1151,
    n455,
    n773,
    n494,
    n629
  );


  and
  g1100
  (
    n1075,
    n406,
    n463,
    n873,
    n546
  );


  xnor
  g1101
  (
    n1137,
    n619,
    n740,
    n422,
    n849
  );


  xnor
  g1102
  (
    n1103,
    n857,
    n594,
    n694,
    n611
  );


  or
  g1103
  (
    n1086,
    n853,
    n697,
    n581,
    n714
  );


  nor
  g1104
  (
    n1181,
    n906,
    n766,
    n758,
    n645
  );


  xor
  g1105
  (
    n1178,
    n685,
    n500,
    n765,
    n407
  );


  or
  g1106
  (
    n1079,
    n601,
    n547,
    n410,
    n622
  );


  xnor
  g1107
  (
    n1179,
    n905,
    n817,
    n749,
    n875
  );


  xnor
  g1108
  (
    n1084,
    n527,
    n592,
    n702,
    n856
  );


  and
  g1109
  (
    n1081,
    n648,
    n760,
    n491,
    n465
  );


  and
  g1110
  (
    n1145,
    n438,
    n631,
    n496,
    n453
  );


  or
  g1111
  (
    n1123,
    n400,
    n667,
    n512,
    n756
  );


  and
  g1112
  (
    KeyWire_0_1,
    n829,
    n432,
    n830,
    n786
  );


  xnor
  g1113
  (
    n1182,
    n585,
    n716,
    n900,
    n860
  );


  and
  g1114
  (
    n1166,
    n448,
    n700,
    n708,
    n754
  );


  xnor
  g1115
  (
    n1171,
    n761,
    n903,
    n620,
    n618
  );


  xnor
  g1116
  (
    n1158,
    n597,
    n805,
    n583,
    n880
  );


  xnor
  g1117
  (
    n1140,
    n706,
    n483,
    n842,
    n665
  );


  nand
  g1118
  (
    n1116,
    n704,
    n735,
    n595,
    n808
  );


  nand
  g1119
  (
    n1169,
    n603,
    n470,
    n695,
    n531
  );


  and
  g1120
  (
    n1092,
    n570,
    n686,
    n609,
    n847
  );


  and
  g1121
  (
    n1090,
    n801,
    n472,
    n820,
    n846
  );


  or
  g1122
  (
    n1150,
    n466,
    n427,
    n436,
    n707
  );


  nor
  g1123
  (
    n1111,
    n797,
    n871,
    n782,
    n510
  );


  nor
  g1124
  (
    n1105,
    n563,
    n850,
    n439,
    n610
  );


  xor
  g1125
  (
    n1098,
    n676,
    n741,
    n444,
    n723
  );


  nor
  g1126
  (
    n1093,
    n615,
    n736,
    n868,
    n663
  );


  nor
  g1127
  (
    n1069,
    n567,
    n537,
    n746,
    n833
  );


  xnor
  g1128
  (
    n1076,
    n730,
    n800,
    n896,
    n571
  );


  or
  g1129
  (
    n1078,
    n848,
    n540,
    n516,
    n687
  );


  nand
  g1130
  (
    n1156,
    n593,
    n726,
    n456,
    n418
  );


  xor
  g1131
  (
    n1135,
    n576,
    n633,
    n649,
    n783
  );


  xor
  g1132
  (
    n1112,
    n719,
    n785,
    n416,
    n528
  );


  xnor
  g1133
  (
    n1159,
    n751,
    n872,
    n827,
    n865
  );


  or
  g1134
  (
    n1077,
    n534,
    n819,
    n710,
    n892
  );


  or
  g1135
  (
    n1142,
    n509,
    n895,
    n851,
    n776
  );


  xor
  g1136
  (
    n1131,
    n854,
    n696,
    n632,
    n889
  );


  or
  g1137
  (
    n1104,
    n898,
    n514,
    n654,
    n657
  );


  or
  g1138
  (
    n1180,
    n476,
    n907,
    n729,
    n838
  );


  or
  g1139
  (
    n1154,
    n623,
    n894,
    n431,
    n822
  );


  nor
  g1140
  (
    n1133,
    n655,
    n507,
    n462,
    n684
  );


  and
  g1141
  (
    n1129,
    n859,
    n653,
    n542,
    n641
  );


  nor
  g1142
  (
    n1067,
    n897,
    n803,
    n731,
    n904
  );


  or
  g1143
  (
    n1128,
    n602,
    n732,
    n600,
    n572
  );


  nor
  g1144
  (
    n1139,
    n493,
    n891,
    n711,
    n698
  );


  xnor
  g1145
  (
    n1149,
    n876,
    n806,
    n617,
    n720
  );


  and
  g1146
  (
    n1120,
    n511,
    n445,
    n474,
    n647
  );


  buf
  g1147
  (
    n1197,
    n1080
  );


  not
  g1148
  (
    n1205,
    n1081
  );


  not
  g1149
  (
    n1213,
    n1090
  );


  buf
  g1150
  (
    n1196,
    n1084
  );


  buf
  g1151
  (
    n1190,
    n1089
  );


  not
  g1152
  (
    n1218,
    n1066
  );


  buf
  g1153
  (
    n1195,
    n1060
  );


  buf
  g1154
  (
    n1212,
    n1078
  );


  not
  g1155
  (
    n1191,
    n1088
  );


  not
  g1156
  (
    n1192,
    n1075
  );


  not
  g1157
  (
    n1204,
    n1087
  );


  buf
  g1158
  (
    n1200,
    n1072
  );


  not
  g1159
  (
    n1187,
    n1070
  );


  buf
  g1160
  (
    n1211,
    n1077
  );


  not
  g1161
  (
    n1215,
    n1067
  );


  buf
  g1162
  (
    n1208,
    n1068
  );


  not
  g1163
  (
    n1210,
    n1074
  );


  buf
  g1164
  (
    n1203,
    n1061
  );


  buf
  g1165
  (
    n1199,
    n1079
  );


  buf
  g1166
  (
    n1189,
    n1083
  );


  not
  g1167
  (
    n1198,
    n1062
  );


  not
  g1168
  (
    n1206,
    n1064
  );


  not
  g1169
  (
    n1217,
    n1085
  );


  buf
  g1170
  (
    n1201,
    n1073
  );


  buf
  g1171
  (
    n1207,
    n1069
  );


  buf
  g1172
  (
    n1214,
    n1071
  );


  buf
  g1173
  (
    n1216,
    n1082
  );


  buf
  g1174
  (
    n1194,
    n1063
  );


  not
  g1175
  (
    n1188,
    n1065
  );


  buf
  g1176
  (
    n1193,
    n1076
  );


  buf
  g1177
  (
    n1202,
    n1086
  );


  buf
  g1178
  (
    n1209,
    n1059
  );


  xor
  g1179
  (
    n1226,
    n1193,
    n1189
  );


  nand
  g1180
  (
    n1220,
    n1190,
    n1091
  );


  nor
  g1181
  (
    n1222,
    n1199,
    n1198
  );


  xnor
  g1182
  (
    n1221,
    n1196,
    n1187
  );


  xor
  g1183
  (
    n1219,
    n1197,
    n1194
  );


  nand
  g1184
  (
    n1225,
    n1195,
    n1188
  );


  xnor
  g1185
  (
    n1224,
    n1192,
    n1200
  );


  and
  g1186
  (
    n1223,
    n1199,
    n1191
  );


  xnor
  g1187
  (
    n1235,
    n1221,
    n1225,
    n1226
  );


  nand
  g1188
  (
    n1234,
    n1204,
    n1206,
    n1226
  );


  or
  g1189
  (
    n1227,
    n1201,
    n1202,
    n1220
  );


  or
  g1190
  (
    n1231,
    n1204,
    n1225,
    n1203
  );


  and
  g1191
  (
    n1230,
    n1205,
    n1203,
    n1222
  );


  nor
  g1192
  (
    n1228,
    n1203,
    n1205,
    n1204
  );


  xor
  g1193
  (
    n1233,
    n1204,
    n1202
  );


  xnor
  g1194
  (
    n1232,
    n1202,
    n1203,
    n1201
  );


  or
  g1195
  (
    n1236,
    n1219,
    n1205,
    n1223
  );


  xnor
  g1196
  (
    n1229,
    n1200,
    n1201,
    n1224
  );


  xnor
  g1197
  (
    n1237,
    n943,
    n920,
    n1236,
    n933
  );


  xnor
  g1198
  (
    n1266,
    n991,
    n910,
    n1207
  );


  xnor
  g1199
  (
    n1272,
    n912,
    n1207,
    n930,
    n1229
  );


  and
  g1200
  (
    n1276,
    n1209,
    n1228,
    n1006,
    n934
  );


  xor
  g1201
  (
    n1273,
    n941,
    n927,
    n996,
    n1001
  );


  or
  g1202
  (
    n1253,
    n1228,
    n940,
    n924,
    n1231
  );


  xor
  g1203
  (
    n1249,
    n1231,
    n953,
    n952,
    n945
  );


  xor
  g1204
  (
    n1267,
    n981,
    n1230,
    n979,
    n1231
  );


  or
  g1205
  (
    n1268,
    n936,
    n970,
    n1003,
    n1227
  );


  xor
  g1206
  (
    n1247,
    n959,
    n928,
    n1209,
    n938
  );


  nand
  g1207
  (
    n1254,
    n1100,
    n1000,
    n966,
    n913
  );


  nor
  g1208
  (
    n1262,
    n963,
    n1207,
    n1098,
    n957
  );


  nand
  g1209
  (
    KeyWire_0_22,
    n990,
    n1229,
    n972,
    n977
  );


  or
  g1210
  (
    n1263,
    n998,
    n914,
    n931,
    n1206
  );


  or
  g1211
  (
    n1256,
    n1231,
    n932,
    n915,
    n971
  );


  and
  g1212
  (
    n1274,
    n988,
    n976,
    n1232,
    n1235
  );


  xnor
  g1213
  (
    n1240,
    n1234,
    n1233,
    n965,
    n978
  );


  or
  g1214
  (
    n1242,
    n1232,
    n1233,
    n958,
    n985
  );


  nand
  g1215
  (
    n1257,
    n946,
    n926,
    n1235,
    n984
  );


  xnor
  g1216
  (
    n1248,
    n1233,
    n989,
    n1235,
    n917
  );


  or
  g1217
  (
    n1271,
    n937,
    n935,
    n1096,
    n1004
  );


  or
  g1218
  (
    n1255,
    n918,
    n1206,
    n964
  );


  or
  g1219
  (
    n1261,
    n1208,
    n942,
    n925,
    n992
  );


  nor
  g1220
  (
    n1265,
    n929,
    n1228,
    n1002,
    n916
  );


  xor
  g1221
  (
    KeyWire_0_8,
    n1228,
    n1232,
    n987,
    n919
  );


  or
  g1222
  (
    n1260,
    n1233,
    n973,
    n962,
    n1230
  );


  or
  g1223
  (
    n1239,
    n999,
    n983,
    n967,
    n961
  );


  xnor
  g1224
  (
    n1259,
    n1094,
    n1229,
    n993
  );


  xnor
  g1225
  (
    n1270,
    n950,
    n1234,
    n982
  );


  or
  g1226
  (
    n1246,
    n923,
    n1230,
    n1093,
    n921
  );


  and
  g1227
  (
    n1245,
    n1236,
    n948,
    n974,
    n949
  );


  nor
  g1228
  (
    n1241,
    n1227,
    n975,
    n956,
    n944
  );


  or
  g1229
  (
    n1258,
    n980,
    n1007,
    n951,
    n939
  );


  nand
  g1230
  (
    n1244,
    n969,
    n1232,
    n994,
    n1230
  );


  or
  g1231
  (
    n1251,
    n1227,
    n955,
    n947,
    n1095
  );


  nor
  g1232
  (
    KeyWire_0_20,
    n1208,
    n1235,
    n968,
    n1099
  );


  or
  g1233
  (
    n1250,
    n1234,
    n1092,
    n1236,
    n1227
  );


  or
  g1234
  (
    n1252,
    n986,
    n954,
    n1005,
    n1097
  );


  xnor
  g1235
  (
    n1275,
    n960,
    n1208,
    n911
  );


  or
  g1236
  (
    n1238,
    n922,
    n995,
    n997,
    n1236
  );


  or
  g1237
  (
    n1280,
    n1115,
    n1111,
    n1106,
    n1237
  );


  nor
  g1238
  (
    n1282,
    n1104,
    n1114,
    n1112,
    n1238
  );


  xor
  g1239
  (
    n1277,
    n1238,
    n1117,
    n1237,
    n1110
  );


  xor
  g1240
  (
    n1279,
    n1237,
    n1101,
    n1113,
    n1109
  );


  and
  g1241
  (
    n1278,
    n1102,
    n1103,
    n1237,
    n1108
  );


  and
  g1242
  (
    n1281,
    n1116,
    n1105,
    n1118,
    n1107
  );


  buf
  g1243
  (
    n1295,
    n1280
  );


  not
  g1244
  (
    n1298,
    n1281
  );


  not
  g1245
  (
    n1283,
    n1282
  );


  not
  g1246
  (
    n1292,
    n1209
  );


  buf
  g1247
  (
    n1296,
    n1282
  );


  buf
  g1248
  (
    n1286,
    n1277
  );


  buf
  g1249
  (
    n1284,
    n1282
  );


  buf
  g1250
  (
    n1293,
    n1279
  );


  not
  g1251
  (
    n1285,
    n1281
  );


  not
  g1252
  (
    n1297,
    n1280
  );


  not
  g1253
  (
    n1290,
    n1281
  );


  buf
  g1254
  (
    n1289,
    n1280
  );


  not
  g1255
  (
    n1287,
    n1211
  );


  xor
  g1256
  (
    n1299,
    n1278,
    n1210
  );


  xnor
  g1257
  (
    n1291,
    n1279,
    n1210
  );


  xor
  g1258
  (
    n1294,
    n1282,
    n1281,
    n1210
  );


  xor
  g1259
  (
    n1288,
    n1209,
    n1278,
    n1280
  );


  buf
  g1260
  (
    n1310,
    n1298
  );


  buf
  g1261
  (
    n1343,
    n1294
  );


  buf
  g1262
  (
    n1355,
    n1284
  );


  not
  g1263
  (
    n1346,
    n1293
  );


  buf
  g1264
  (
    n1302,
    n1286
  );


  not
  g1265
  (
    n1321,
    n1213
  );


  buf
  g1266
  (
    n1304,
    n1296
  );


  buf
  g1267
  (
    n1354,
    n1297
  );


  buf
  g1268
  (
    n1352,
    n1299
  );


  not
  g1269
  (
    n1347,
    n1298
  );


  not
  g1270
  (
    n1309,
    n1287
  );


  buf
  g1271
  (
    n1327,
    n1286
  );


  not
  g1272
  (
    n1357,
    n1292
  );


  not
  g1273
  (
    n1341,
    n1286
  );


  not
  g1274
  (
    n1315,
    n1214
  );


  not
  g1275
  (
    n1349,
    n1285
  );


  buf
  g1276
  (
    n1319,
    n1213
  );


  not
  g1277
  (
    n1340,
    n1299
  );


  not
  g1278
  (
    n1313,
    n1211
  );


  buf
  g1279
  (
    n1350,
    n1295
  );


  not
  g1280
  (
    n1331,
    n1285
  );


  not
  g1281
  (
    n1308,
    n1287
  );


  not
  g1282
  (
    n1336,
    n1285
  );


  buf
  g1283
  (
    n1329,
    n1290
  );


  buf
  g1284
  (
    n1328,
    n1288
  );


  not
  g1285
  (
    n1306,
    n1212
  );


  buf
  g1286
  (
    KeyWire_0_28,
    n1295
  );


  not
  g1287
  (
    n1301,
    n1121
  );


  not
  g1288
  (
    n1317,
    n1284
  );


  not
  g1289
  (
    n1332,
    n1294
  );


  not
  g1290
  (
    n1324,
    n1293
  );


  not
  g1291
  (
    n1339,
    n1211
  );


  buf
  g1292
  (
    n1345,
    n1290
  );


  buf
  g1293
  (
    n1337,
    n1297
  );


  not
  g1294
  (
    n1359,
    n1287
  );


  not
  g1295
  (
    n1344,
    n1294
  );


  not
  g1296
  (
    n1322,
    n1295
  );


  not
  g1297
  (
    n1305,
    n1283
  );


  buf
  g1298
  (
    n1351,
    n1283
  );


  buf
  g1299
  (
    n1342,
    n1296
  );


  not
  g1300
  (
    n1353,
    n1287
  );


  buf
  g1301
  (
    n1318,
    n1296
  );


  not
  g1302
  (
    n1356,
    n1288
  );


  not
  g1303
  (
    n1333,
    n1285
  );


  buf
  g1304
  (
    n1316,
    n1212
  );


  not
  g1305
  (
    n1330,
    n1296
  );


  not
  g1306
  (
    n1323,
    n1299
  );


  buf
  g1307
  (
    n1307,
    n1214
  );


  buf
  g1308
  (
    n1334,
    n1289
  );


  buf
  g1309
  (
    n1325,
    n1293
  );


  and
  g1310
  (
    n1326,
    n1299,
    n1298,
    n1288
  );


  nor
  g1311
  (
    n1311,
    n1297,
    n1289,
    n1284
  );


  nor
  g1312
  (
    n1320,
    n1215,
    n1120,
    n1293,
    n1291
  );


  and
  g1313
  (
    n1338,
    n1286,
    n1291,
    n1290
  );


  or
  g1314
  (
    n1335,
    n1212,
    n1283,
    n1122,
    n1294
  );


  nor
  g1315
  (
    n1358,
    n1283,
    n1284,
    n1213,
    n1289
  );


  and
  g1316
  (
    n1312,
    n1295,
    n1298,
    n1292,
    n1212
  );


  or
  g1317
  (
    n1300,
    n1297,
    n1119,
    n1292
  );


  xor
  g1318
  (
    n1303,
    n1213,
    n1291,
    n1289,
    n1288
  );


  or
  g1319
  (
    n1348,
    n1211,
    n1290,
    n1214
  );


  buf
  g1320
  (
    n1366,
    n1305
  );


  buf
  g1321
  (
    n1379,
    n1308
  );


  not
  g1322
  (
    n1370,
    n1307
  );


  not
  g1323
  (
    n1369,
    n1309
  );


  buf
  g1324
  (
    n1363,
    n1300
  );


  buf
  g1325
  (
    n1372,
    n1304
  );


  not
  g1326
  (
    n1362,
    n1313
  );


  not
  g1327
  (
    n1377,
    n1302
  );


  not
  g1328
  (
    n1375,
    n1314
  );


  not
  g1329
  (
    n1368,
    n1319
  );


  not
  g1330
  (
    n1371,
    n1318
  );


  not
  g1331
  (
    n1365,
    n1303
  );


  buf
  g1332
  (
    n1361,
    n1310
  );


  buf
  g1333
  (
    n1376,
    n1317
  );


  buf
  g1334
  (
    n1367,
    n1315
  );


  not
  g1335
  (
    n1378,
    n1306
  );


  not
  g1336
  (
    n1360,
    n1312
  );


  buf
  g1337
  (
    n1364,
    n1301
  );


  not
  g1338
  (
    n1373,
    n1316
  );


  buf
  g1339
  (
    n1374,
    n1311
  );


  buf
  g1340
  (
    n1408,
    n1243
  );


  not
  g1341
  (
    n1418,
    n1257
  );


  buf
  g1342
  (
    n1428,
    n1248
  );


  buf
  g1343
  (
    n1425,
    n1215
  );


  buf
  g1344
  (
    n1387,
    n1255
  );


  not
  g1345
  (
    n1415,
    n1368
  );


  not
  g1346
  (
    n1419,
    n1369
  );


  not
  g1347
  (
    n1442,
    n1379
  );


  not
  g1348
  (
    n1396,
    n1372
  );


  not
  g1349
  (
    n1403,
    n1253
  );


  buf
  g1350
  (
    n1447,
    n1371
  );


  buf
  g1351
  (
    n1390,
    n1377
  );


  not
  g1352
  (
    n1431,
    n1374
  );


  not
  g1353
  (
    n1413,
    n1238
  );


  buf
  g1354
  (
    n1407,
    n1368
  );


  buf
  g1355
  (
    n1438,
    n1258
  );


  buf
  g1356
  (
    n1411,
    n1260
  );


  not
  g1357
  (
    n1454,
    n1365
  );


  not
  g1358
  (
    n1426,
    n1261
  );


  not
  g1359
  (
    n1414,
    n1271
  );


  buf
  g1360
  (
    n1436,
    n1372
  );


  not
  g1361
  (
    n1451,
    n1371
  );


  buf
  g1362
  (
    n1433,
    n1240
  );


  not
  g1363
  (
    n1424,
    n1366
  );


  buf
  g1364
  (
    n1391,
    n1266
  );


  buf
  g1365
  (
    n1420,
    n1369
  );


  buf
  g1366
  (
    n1402,
    n1249
  );


  buf
  g1367
  (
    n1455,
    n1262
  );


  not
  g1368
  (
    n1439,
    n1270
  );


  not
  g1369
  (
    n1380,
    n1264
  );


  not
  g1370
  (
    n1430,
    n1262
  );


  or
  g1371
  (
    n1384,
    n1364,
    n1251
  );


  nand
  g1372
  (
    n1457,
    n1260,
    n1245,
    n1370,
    n1374
  );


  xnor
  g1373
  (
    n1392,
    n1367,
    n1241,
    n1378,
    n1216
  );


  xnor
  g1374
  (
    n1445,
    n1374,
    n1245,
    n38,
    n1263
  );


  xnor
  g1375
  (
    n1459,
    n1253,
    n1242,
    n1240,
    n1269
  );


  nor
  g1376
  (
    n1409,
    n1269,
    n1255,
    n1365
  );


  or
  g1377
  (
    n1427,
    n1376,
    n1362,
    n1244,
    n1268
  );


  and
  g1378
  (
    n1429,
    n1258,
    n1361,
    n1371,
    n1379
  );


  and
  g1379
  (
    KeyWire_0_12,
    n37,
    n1266,
    n1257,
    n1375
  );


  xor
  g1380
  (
    n1386,
    n1362,
    n1363,
    n1250,
    n1373
  );


  xor
  g1381
  (
    KeyWire_0_26,
    n1372,
    n1268,
    n1244,
    n1260
  );


  nor
  g1382
  (
    n1404,
    n1369,
    n1361,
    n1241,
    n1370
  );


  nand
  g1383
  (
    n1458,
    n1248,
    n1251,
    n1216,
    n1364
  );


  and
  g1384
  (
    n1432,
    n1379,
    n1378,
    n1269,
    n1367
  );


  xor
  g1385
  (
    n1388,
    n1361,
    n1238,
    n1263,
    n1265
  );


  and
  g1386
  (
    n1441,
    n1370,
    n1270,
    n1264,
    n1261
  );


  nand
  g1387
  (
    n1406,
    n1360,
    n1366,
    n1255,
    n1249
  );


  xnor
  g1388
  (
    n1440,
    n1271,
    n1245,
    n1243,
    n1362
  );


  and
  g1389
  (
    n1383,
    n1375,
    n1364,
    n1374,
    n1271
  );


  nand
  g1390
  (
    n1456,
    n1270,
    n1267,
    n1363,
    n1245
  );


  nor
  g1391
  (
    n1382,
    n1253,
    n1259,
    n1250,
    n1264
  );


  nand
  g1392
  (
    n1412,
    n1241,
    n1363,
    n1378,
    n1377
  );


  nand
  g1393
  (
    n1422,
    n1259,
    n1247,
    n1377,
    n1373
  );


  nand
  g1394
  (
    n1434,
    n1251,
    n38,
    n1267,
    n1262
  );


  nand
  g1395
  (
    n1389,
    n1246,
    n1248,
    n1269,
    n1368
  );


  nand
  g1396
  (
    n1400,
    n1253,
    n1248,
    n1379,
    n1361
  );


  nor
  g1397
  (
    n1405,
    n1262,
    n1246,
    n1265,
    n1368
  );


  or
  g1398
  (
    n1453,
    n1267,
    n1244,
    n1360,
    n1367
  );


  and
  g1399
  (
    n1401,
    n1216,
    n1256,
    n1251,
    n1254
  );


  nor
  g1400
  (
    n1437,
    n1252,
    n1366,
    n1265,
    n1257
  );


  and
  g1401
  (
    n1416,
    n38,
    n1249,
    n1242,
    n1252
  );


  nor
  g1402
  (
    n1443,
    n1243,
    n1241,
    n1250,
    n1215
  );


  nor
  g1403
  (
    n1450,
    n1258,
    n1242,
    n1246,
    n1362
  );


  nand
  g1404
  (
    n1423,
    n1216,
    n1247,
    n1242,
    n1377
  );


  or
  g1405
  (
    n1410,
    n1260,
    n1256,
    n1378
  );


  and
  g1406
  (
    n1381,
    n1259,
    n1239,
    n1365,
    n1375
  );


  nor
  g1407
  (
    n1397,
    n1270,
    n1244,
    n1261,
    n1243
  );


  xor
  g1408
  (
    n1394,
    n38,
    n1268,
    n1370,
    n1376
  );


  or
  g1409
  (
    n1448,
    n1215,
    n1258,
    n1240,
    n1267
  );


  or
  g1410
  (
    n1399,
    n1239,
    n1252,
    n1246
  );


  or
  g1411
  (
    n1417,
    n1254,
    n1373,
    n1257,
    n1250
  );


  or
  g1412
  (
    n1385,
    n1366,
    n1254,
    n1264
  );


  xnor
  g1413
  (
    n1449,
    n1255,
    n1239,
    n1360
  );


  xnor
  g1414
  (
    n1395,
    n1263,
    n1364,
    n1265,
    n1363
  );


  nor
  g1415
  (
    n1398,
    n1240,
    n1268,
    n1261,
    n1263
  );


  and
  g1416
  (
    n1446,
    n1376,
    n1376,
    n1369,
    n1247
  );


  and
  g1417
  (
    KeyWire_0_25,
    n1249,
    n1367,
    n1266,
    n1373
  );


  xnor
  g1418
  (
    n1435,
    n1360,
    n1256,
    n1372,
    n1259
  );


  nor
  g1419
  (
    n1393,
    n1371,
    n1247,
    n1266,
    n1375
  );


  or
  g1420
  (
    n1462,
    n1387,
    n1413,
    n1447,
    n1431
  );


  nand
  g1421
  (
    n1463,
    n174,
    n1125,
    n1422,
    n1402
  );


  xnor
  g1422
  (
    n1471,
    n1400,
    n1380,
    n1396,
    n1453
  );


  and
  g1423
  (
    n1481,
    n1448,
    n175,
    n1434,
    n1384
  );


  xor
  g1424
  (
    n1467,
    n1451,
    n1127,
    n1425,
    n1391
  );


  xnor
  g1425
  (
    n1460,
    n1389,
    n174,
    n1420,
    n1430
  );


  or
  g1426
  (
    n1466,
    n1459,
    n1429,
    n1406,
    n1446
  );


  nor
  g1427
  (
    n1464,
    n1416,
    n1437,
    n1404,
    n1126
  );


  or
  g1428
  (
    n1473,
    n1458,
    n1428,
    n1418,
    n1442
  );


  nand
  g1429
  (
    n1483,
    n1455,
    n1439,
    n176,
    n1454
  );


  or
  g1430
  (
    n1475,
    n1441,
    n1426,
    n1397,
    n1394
  );


  nor
  g1431
  (
    n1482,
    n175,
    n1452,
    n1124,
    n1385
  );


  and
  g1432
  (
    n1469,
    n1438,
    n1412,
    n1427,
    n1392
  );


  xor
  g1433
  (
    n1470,
    n1423,
    n1386,
    n1382,
    n1398
  );


  xor
  g1434
  (
    n1465,
    n1433,
    n1410,
    n1393,
    n1432
  );


  nor
  g1435
  (
    n1479,
    n1415,
    n1405,
    n1436,
    n1390
  );


  and
  g1436
  (
    KeyWire_0_27,
    n1445,
    n1395,
    n1409,
    n1401
  );


  or
  g1437
  (
    n1478,
    n1435,
    n175,
    n1388,
    n1450
  );


  xor
  g1438
  (
    n1477,
    n1414,
    n1403,
    n1440,
    n1130
  );


  nor
  g1439
  (
    n1480,
    n175,
    n1381,
    n1123,
    n174
  );


  nor
  g1440
  (
    n1474,
    n1443,
    n1417,
    n1407,
    n1399
  );


  and
  g1441
  (
    n1476,
    n1457,
    n1128,
    n1411,
    n1456
  );


  xor
  g1442
  (
    n1461,
    n1444,
    n1129,
    n1408,
    n1383
  );


  nor
  g1443
  (
    n1468,
    n1424,
    n1419,
    n1421,
    n1449
  );


  not
  g1444
  (
    n1489,
    n1460
  );


  not
  g1445
  (
    n1488,
    n1462
  );


  buf
  g1446
  (
    n1485,
    n1463
  );


  not
  g1447
  (
    n1487,
    n1467
  );


  not
  g1448
  (
    n1491,
    n1465
  );


  buf
  g1449
  (
    n1484,
    n1464
  );


  buf
  g1450
  (
    n1486,
    n1461
  );


  buf
  g1451
  (
    n1490,
    n1466
  );


  and
  g1452
  (
    n1499,
    n1022,
    n1137,
    n1351,
    n1487
  );


  xor
  g1453
  (
    n1520,
    n1343,
    n1032,
    n1323,
    n1042
  );


  nand
  g1454
  (
    n1497,
    n1016,
    n1320,
    n1348,
    n1009
  );


  nand
  g1455
  (
    n1517,
    n1485,
    n1031,
    n1324,
    n1133
  );


  and
  g1456
  (
    n1495,
    n1035,
    n1048,
    n1484,
    n1029
  );


  xor
  g1457
  (
    n1500,
    n1008,
    n1134,
    n1488,
    n1346
  );


  xor
  g1458
  (
    n1513,
    n1484,
    n1036,
    n1488,
    n1034
  );


  nand
  g1459
  (
    n1507,
    n1025,
    n1038,
    n1027,
    n1056
  );


  nand
  g1460
  (
    n1501,
    n1039,
    n1030,
    n1028,
    n1023
  );


  nor
  g1461
  (
    n1522,
    n1331,
    n1329,
    n1024,
    n1486
  );


  xor
  g1462
  (
    n1511,
    n1490,
    n1043,
    n1349,
    n1013
  );


  nand
  g1463
  (
    n1508,
    n1340,
    n1347,
    n1350,
    n1490
  );


  xor
  g1464
  (
    n1503,
    n1046,
    n1138,
    n1332,
    n1049
  );


  xnor
  g1465
  (
    n1521,
    n1469,
    n1484,
    n1033,
    n1132
  );


  or
  g1466
  (
    n1510,
    n1487,
    n1055,
    n1490,
    n1135
  );


  xor
  g1467
  (
    n1523,
    n1470,
    n1136,
    n1342,
    n1486
  );


  xnor
  g1468
  (
    n1519,
    n1019,
    n1328,
    n1485,
    n1344
  );


  xor
  g1469
  (
    n1498,
    n1139,
    n1327,
    n1052,
    n1054
  );


  xnor
  g1470
  (
    n1516,
    n1336,
    n1491,
    n1489,
    n1050
  );


  or
  g1471
  (
    n1504,
    n1040,
    n1321,
    n1322,
    n1217
  );


  nor
  g1472
  (
    n1506,
    n1053,
    n1491,
    n1485
  );


  xor
  g1473
  (
    n1493,
    n1045,
    n1487,
    n1140,
    n1334
  );


  nor
  g1474
  (
    n1496,
    n1041,
    n1333,
    n1489,
    n1018
  );


  xnor
  g1475
  (
    n1518,
    n1012,
    n1486,
    n1491,
    n1341
  );


  xnor
  g1476
  (
    n1502,
    n1217,
    n1011,
    n1014,
    n1131
  );


  nand
  g1477
  (
    n1512,
    n1047,
    n1044,
    n1020,
    n1488
  );


  or
  g1478
  (
    n1509,
    n1490,
    n1017,
    n1488,
    n1489
  );


  xor
  g1479
  (
    n1505,
    n1345,
    n1026,
    n1335,
    n1010
  );


  or
  g1480
  (
    n1515,
    n1491,
    n1484,
    n1021,
    n1337
  );


  xnor
  g1481
  (
    n1514,
    n1015,
    n1339,
    n1051,
    n1487
  );


  xnor
  g1482
  (
    n1494,
    n1325,
    n1037,
    n1468,
    n1338
  );


  xor
  g1483
  (
    n1492,
    n1486,
    n1330,
    n1489,
    n1326
  );


  buf
  g1484
  (
    n1524,
    n1492
  );


  buf
  g1485
  (
    n1525,
    n1493
  );


  xor
  g1486
  (
    n1526,
    n1142,
    n1525,
    n1143,
    n1141
  );


  buf
  g1487
  (
    n1527,
    n1217
  );


  xnor
  g1488
  (
    n1528,
    n1217,
    n1526
  );


  buf
  g1489
  (
    n1535,
    n1528
  );


  buf
  g1490
  (
    n1529,
    n1527
  );


  buf
  g1491
  (
    n1536,
    n1058
  );


  buf
  g1492
  (
    n1534,
    n1528
  );


  not
  g1493
  (
    n1530,
    n1527
  );


  buf
  g1494
  (
    n1533,
    n1527
  );


  xor
  g1495
  (
    n1532,
    n1057,
    n1527
  );


  buf
  g1496
  (
    n1531,
    n1528
  );


  buf
  g1497
  (
    n1537,
    n1146
  );


  buf
  g1498
  (
    n1539,
    n1529
  );


  or
  g1499
  (
    n1540,
    n1147,
    n1145
  );


  or
  g1500
  (
    n1538,
    n1530,
    n1530,
    n1144,
    n1529
  );


  nor
  g1501
  (
    n1541,
    n1540,
    n1148
  );


  not
  g1502
  (
    KeyWire_0_23,
    n1541
  );


  nor
  g1503
  (
    n1542,
    n1541,
    n1218
  );


  not
  g1504
  (
    n1544,
    n1542
  );


  buf
  g1505
  (
    n1545,
    n1150
  );


  buf
  g1506
  (
    n1549,
    n1153
  );


  buf
  g1507
  (
    n1547,
    n1152
  );


  xnor
  g1508
  (
    n1546,
    n1542,
    n1149,
    n1543,
    n1151
  );


  nor
  g1509
  (
    n1548,
    n1154,
    n1543
  );


  not
  g1510
  (
    n1557,
    n1354
  );


  not
  g1511
  (
    n1559,
    n1536
  );


  not
  g1512
  (
    n1568,
    n1531
  );


  not
  g1513
  (
    n1567,
    n1549
  );


  not
  g1514
  (
    KeyWire_0_17,
    n1352
  );


  not
  g1515
  (
    n1556,
    n1534
  );


  xnor
  g1516
  (
    n1571,
    n1275,
    n1532
  );


  xnor
  g1517
  (
    n1566,
    n1534,
    n1536,
    n1545
  );


  xnor
  g1518
  (
    n1560,
    n1532,
    n1276,
    n1544
  );


  and
  g1519
  (
    n1555,
    n1273,
    n1276,
    n1535,
    n1546
  );


  nand
  g1520
  (
    n1554,
    n1535,
    n1548,
    n1533
  );


  nor
  g1521
  (
    n1551,
    n1533,
    n1534,
    n1272,
    n1549
  );


  and
  g1522
  (
    n1563,
    n1534,
    n1530,
    n1531
  );


  xor
  g1523
  (
    n1558,
    n1532,
    n1273,
    n1548,
    n1535
  );


  xnor
  g1524
  (
    n1553,
    n1533,
    n1273,
    n1531,
    n1218
  );


  xor
  g1525
  (
    n1565,
    n1547,
    n1273,
    n1274,
    n1272
  );


  or
  g1526
  (
    n1562,
    n1272,
    n1275,
    n1549,
    n1530
  );


  xor
  g1527
  (
    n1564,
    n1353,
    n1547,
    n1546,
    n1545
  );


  and
  g1528
  (
    n1570,
    n1544,
    n1274,
    n1545,
    n1549
  );


  and
  g1529
  (
    n1572,
    n1272,
    n1276,
    n1274,
    n1548
  );


  and
  g1530
  (
    n1550,
    n1546,
    n1536,
    n1545,
    n1275
  );


  or
  g1531
  (
    n1552,
    n1275,
    n1547,
    n1544,
    n1274
  );


  nand
  g1532
  (
    n1573,
    n1218,
    n1533,
    n1544,
    n1546
  );


  xnor
  g1533
  (
    n1569,
    n1271,
    n1547,
    n1535,
    n1532
  );


  not
  g1534
  (
    n1588,
    n1571
  );


  buf
  g1535
  (
    n1592,
    n1564
  );


  not
  g1536
  (
    n1593,
    n1562
  );


  buf
  g1537
  (
    n1597,
    n1553
  );


  not
  g1538
  (
    n1596,
    n1559
  );


  buf
  g1539
  (
    n1582,
    n1554
  );


  buf
  g1540
  (
    n1598,
    n1557
  );


  buf
  g1541
  (
    n1594,
    n1550
  );


  not
  g1542
  (
    n1605,
    n1561
  );


  not
  g1543
  (
    n1583,
    n1568
  );


  not
  g1544
  (
    n1578,
    n1558
  );


  buf
  g1545
  (
    n1595,
    n1572
  );


  not
  g1546
  (
    n1584,
    n1570
  );


  buf
  g1547
  (
    n1587,
    n1565
  );


  not
  g1548
  (
    n1579,
    n1571
  );


  buf
  g1549
  (
    n1586,
    n1563
  );


  not
  g1550
  (
    n1603,
    n1552
  );


  not
  g1551
  (
    n1602,
    n1569
  );


  not
  g1552
  (
    n1608,
    n1555
  );


  buf
  g1553
  (
    n1607,
    n1566
  );


  not
  g1554
  (
    n1604,
    n1551
  );


  not
  g1555
  (
    n1590,
    n1571
  );


  not
  g1556
  (
    n1577,
    n1560
  );


  buf
  g1557
  (
    n1600,
    n1556
  );


  buf
  g1558
  (
    n1609,
    n1570
  );


  buf
  g1559
  (
    n1576,
    n1572
  );


  buf
  g1560
  (
    n1581,
    n1570
  );


  not
  g1561
  (
    n1585,
    n1573
  );


  buf
  g1562
  (
    n1575,
    n1569
  );


  not
  g1563
  (
    n1599,
    n1570
  );


  buf
  g1564
  (
    n1591,
    n1567
  );


  not
  g1565
  (
    n1606,
    n1572
  );


  buf
  g1566
  (
    n1574,
    n1571
  );


  buf
  g1567
  (
    n1601,
    n1572
  );


  buf
  g1568
  (
    n1589,
    n1568
  );


  buf
  g1569
  (
    n1580,
    n1573
  );


  and
  g1570
  (
    n1613,
    n1594,
    n1574,
    n1605,
    n1606
  );


  xor
  g1571
  (
    n1615,
    n1595,
    n1591,
    n1597,
    n1606
  );


  nand
  g1572
  (
    n1619,
    n1600,
    n1586,
    n1596,
    n1478
  );


  nor
  g1573
  (
    n1621,
    n1593,
    n1583,
    n1576,
    n1473
  );


  nand
  g1574
  (
    n1620,
    n1580,
    n1604,
    n1480,
    n1592
  );


  xor
  g1575
  (
    n1614,
    n1585,
    n1471,
    n1606,
    n1588
  );


  nand
  g1576
  (
    n1616,
    n1602,
    n1578,
    n1155,
    n1156
  );


  nand
  g1577
  (
    n1618,
    n1606,
    n1475,
    n1477,
    n1598
  );


  and
  g1578
  (
    n1617,
    n1601,
    n1579,
    n1603,
    n1472
  );


  xor
  g1579
  (
    n1612,
    n1575,
    n1587,
    n1599,
    n1476
  );


  xnor
  g1580
  (
    n1611,
    n1577,
    n1479,
    n1590,
    n1584
  );


  xor
  g1581
  (
    n1610,
    n1582,
    n1474,
    n1589,
    n1581
  );


  not
  g1582
  (
    n1622,
    n1617
  );


  buf
  g1583
  (
    n1627,
    n1619
  );


  buf
  g1584
  (
    n1626,
    n1620
  );


  buf
  g1585
  (
    n1623,
    n1618
  );


  not
  g1586
  (
    n1624,
    n1483
  );


  xnor
  g1587
  (
    n1625,
    n1616,
    n1482,
    n1481,
    n1621
  );


  or
  g1588
  (
    n1633,
    n1498,
    n1357,
    n1497,
    n1521
  );


  nand
  g1589
  (
    n1641,
    n1496,
    n1625,
    n1626,
    n1506
  );


  nor
  g1590
  (
    n1637,
    n1626,
    n1522,
    n1627,
    n39
  );


  xor
  g1591
  (
    n1631,
    n1508,
    n1624,
    n39,
    n1503
  );


  xor
  g1592
  (
    n1632,
    n1515,
    n1509,
    n1514,
    n1495
  );


  xor
  g1593
  (
    n1638,
    n1520,
    n1523,
    n1519,
    n1627
  );


  or
  g1594
  (
    n1628,
    n1358,
    n1505,
    n176,
    n1624
  );


  xor
  g1595
  (
    n1640,
    n1626,
    n1623,
    n1511,
    n1507
  );


  nor
  g1596
  (
    n1635,
    n1356,
    n1500,
    n1523,
    n177
  );


  and
  g1597
  (
    n1643,
    n1513,
    n1359,
    n1517,
    n1494
  );


  xor
  g1598
  (
    n1636,
    n176,
    n1627,
    n177
  );


  or
  g1599
  (
    n1629,
    n1355,
    n1625,
    n1518,
    n39
  );


  nor
  g1600
  (
    n1642,
    n1512,
    n176,
    n39,
    n1499
  );


  nor
  g1601
  (
    n1634,
    n1622,
    n1501,
    n1523,
    n1625
  );


  xnor
  g1602
  (
    n1630,
    n1625,
    n1502,
    n1516,
    n1510
  );


  nand
  g1603
  (
    n1639,
    n177,
    n1504,
    n1626,
    n1523
  );


  nor
  g1604
  (
    n1644,
    n177,
    n1573,
    n1643
  );


  or
  g1605
  (
    n1645,
    n1644,
    n1609,
    n1607
  );


  xnor
  g1606
  (
    n1647,
    n1644,
    n1607,
    n1608
  );


  or
  g1607
  (
    n1646,
    n1609,
    n1608,
    n1607
  );


  and
  g1608
  (
    n1648,
    n1607,
    n1609,
    n1644
  );


  nor
  g1609
  (
    n1657,
    n1157,
    n1184,
    n1648,
    n1159
  );


  nand
  g1610
  (
    n1656,
    n1158,
    n1174,
    n1163,
    n1173
  );


  nor
  g1611
  (
    n1658,
    n1171,
    n1168,
    n1176,
    n1648
  );


  and
  g1612
  (
    n1649,
    n1175,
    n1167,
    n1180,
    n1169
  );


  or
  g1613
  (
    n1652,
    n1165,
    n1160,
    n1646,
    n1185
  );


  nand
  g1614
  (
    n1655,
    n1164,
    n1183,
    n1647,
    n1170
  );


  xor
  g1615
  (
    n1653,
    n1181,
    n1166,
    n1647,
    n1161
  );


  xor
  g1616
  (
    n1651,
    n1179,
    n1178,
    n1648,
    n1177
  );


  or
  g1617
  (
    n1650,
    n1172,
    n1162,
    n1186,
    n1645
  );


  nand
  g1618
  (
    n1654,
    n1648,
    n1182,
    n1647
  );


  xor
  KeyGate_0_0
  (
    n90,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1130,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1004,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n349,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1132,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n711,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n570,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n896,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1264,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n174,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n768,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n801,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1452,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n328,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1173,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n807,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n551,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1561,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n141,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n868,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1243,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n956,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1269,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1543,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n420,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1421,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1444,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1472,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1314,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n770,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n958,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n901,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


