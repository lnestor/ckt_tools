

module Stat_1728_18_5
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n725,
  n729,
  n734,
  n728,
  n723,
  n788,
  n780,
  n799,
  n1739,
  n1725,
  n1738,
  n1746,
  n1742,
  n1744,
  n1733,
  n1741,
  n1728,
  n1727,
  n1735,
  n1726,
  n1737,
  n1724,
  n1723,
  n1745,
  n1732,
  n1729,
  n1734,
  n1743,
  n1736,
  n1731,
  n1740,
  n1730,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n725;
  output n729;
  output n734;
  output n728;
  output n723;
  output n788;
  output n780;
  output n799;
  output n1739;
  output n1725;
  output n1738;
  output n1746;
  output n1742;
  output n1744;
  output n1733;
  output n1741;
  output n1728;
  output n1727;
  output n1735;
  output n1726;
  output n1737;
  output n1724;
  output n1723;
  output n1745;
  output n1732;
  output n1729;
  output n1734;
  output n1743;
  output n1736;
  output n1731;
  output n1740;
  output n1730;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n724;
  wire n726;
  wire n727;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    n75,
    n17
  );


  not
  g1
  (
    n49,
    n11
  );


  not
  g2
  (
    n64,
    n15
  );


  not
  g3
  (
    n50,
    n10
  );


  not
  g4
  (
    n76,
    n12
  );


  not
  g5
  (
    n39,
    n9
  );


  not
  g6
  (
    n66,
    n10
  );


  not
  g7
  (
    n70,
    n7
  );


  not
  g8
  (
    n90,
    n2
  );


  buf
  g9
  (
    n40,
    n4
  );


  buf
  g10
  (
    n22,
    n4
  );


  not
  g11
  (
    n58,
    n3
  );


  not
  g12
  (
    n79,
    n16
  );


  not
  g13
  (
    n62,
    n8
  );


  not
  g14
  (
    n21,
    n16
  );


  not
  g15
  (
    n82,
    n16
  );


  not
  g16
  (
    n63,
    n8
  );


  not
  g17
  (
    n71,
    n1
  );


  not
  g18
  (
    n69,
    n4
  );


  buf
  g19
  (
    n37,
    n13
  );


  buf
  g20
  (
    n88,
    n8
  );


  not
  g21
  (
    n42,
    n5
  );


  not
  g22
  (
    n26,
    n16
  );


  not
  g23
  (
    n87,
    n18
  );


  not
  g24
  (
    n72,
    n10
  );


  not
  g25
  (
    n28,
    n17
  );


  not
  g26
  (
    n77,
    n11
  );


  not
  g27
  (
    n20,
    n6
  );


  not
  g28
  (
    n51,
    n17
  );


  not
  g29
  (
    n33,
    n10
  );


  buf
  g30
  (
    n48,
    n6
  );


  buf
  g31
  (
    n85,
    n14
  );


  not
  g32
  (
    n84,
    n2
  );


  not
  g33
  (
    n34,
    n9
  );


  buf
  g34
  (
    n36,
    n5
  );


  not
  g35
  (
    n32,
    n6
  );


  not
  g36
  (
    n61,
    n13
  );


  buf
  g37
  (
    n25,
    n5
  );


  buf
  g38
  (
    n27,
    n1
  );


  not
  g39
  (
    n89,
    n8
  );


  buf
  g40
  (
    KeyWire_0_35,
    n15
  );


  not
  g41
  (
    KeyWire_0_15,
    n18
  );


  buf
  g42
  (
    n41,
    n4
  );


  not
  g43
  (
    n44,
    n3
  );


  not
  g44
  (
    n19,
    n14
  );


  not
  g45
  (
    n23,
    n13
  );


  not
  g46
  (
    n57,
    n3
  );


  buf
  g47
  (
    n60,
    n1
  );


  not
  g48
  (
    n30,
    n5
  );


  buf
  g49
  (
    n31,
    n11
  );


  not
  g50
  (
    n74,
    n9
  );


  not
  g51
  (
    n54,
    n1
  );


  buf
  g52
  (
    n52,
    n2
  );


  not
  g53
  (
    n73,
    n12
  );


  not
  g54
  (
    n67,
    n12
  );


  not
  g55
  (
    n45,
    n17
  );


  not
  g56
  (
    n56,
    n11
  );


  buf
  g57
  (
    n47,
    n7
  );


  not
  g58
  (
    n81,
    n18
  );


  buf
  g59
  (
    n65,
    n18
  );


  not
  g60
  (
    n24,
    n3
  );


  buf
  g61
  (
    n86,
    n13
  );


  buf
  g62
  (
    n35,
    n7
  );


  buf
  g63
  (
    n59,
    n14
  );


  not
  g64
  (
    n55,
    n9
  );


  buf
  g65
  (
    n46,
    n7
  );


  not
  g66
  (
    n68,
    n2
  );


  buf
  g67
  (
    n38,
    n14
  );


  not
  g68
  (
    n43,
    n12
  );


  not
  g69
  (
    n53,
    n6
  );


  buf
  g70
  (
    n80,
    n15
  );


  not
  g71
  (
    n29,
    n15
  );


  buf
  g72
  (
    n369,
    n40
  );


  not
  g73
  (
    n130,
    n32
  );


  buf
  g74
  (
    n265,
    n84
  );


  not
  g75
  (
    KeyWire_0_33,
    n23
  );


  not
  g76
  (
    n298,
    n35
  );


  not
  g77
  (
    n112,
    n65
  );


  buf
  g78
  (
    n118,
    n70
  );


  not
  g79
  (
    n260,
    n31
  );


  buf
  g80
  (
    n122,
    n74
  );


  buf
  g81
  (
    n251,
    n79
  );


  not
  g82
  (
    n315,
    n69
  );


  buf
  g83
  (
    n128,
    n66
  );


  buf
  g84
  (
    n196,
    n30
  );


  buf
  g85
  (
    KeyWire_0_11,
    n87
  );


  not
  g86
  (
    n328,
    n37
  );


  not
  g87
  (
    n349,
    n24
  );


  not
  g88
  (
    n204,
    n60
  );


  not
  g89
  (
    n212,
    n61
  );


  not
  g90
  (
    n318,
    n64
  );


  buf
  g91
  (
    n285,
    n75
  );


  not
  g92
  (
    n162,
    n36
  );


  not
  g93
  (
    n254,
    n61
  );


  buf
  g94
  (
    n160,
    n62
  );


  not
  g95
  (
    n290,
    n35
  );


  not
  g96
  (
    n355,
    n70
  );


  buf
  g97
  (
    n263,
    n69
  );


  not
  g98
  (
    n345,
    n32
  );


  buf
  g99
  (
    n173,
    n50
  );


  not
  g100
  (
    n375,
    n51
  );


  buf
  g101
  (
    n362,
    n45
  );


  not
  g102
  (
    n320,
    n82
  );


  buf
  g103
  (
    n361,
    n75
  );


  not
  g104
  (
    n257,
    n73
  );


  buf
  g105
  (
    n255,
    n73
  );


  not
  g106
  (
    n367,
    n63
  );


  buf
  g107
  (
    KeyWire_0_7,
    n46
  );


  buf
  g108
  (
    n153,
    n62
  );


  not
  g109
  (
    n226,
    n54
  );


  buf
  g110
  (
    n211,
    n73
  );


  not
  g111
  (
    n157,
    n38
  );


  not
  g112
  (
    n302,
    n82
  );


  not
  g113
  (
    n303,
    n45
  );


  buf
  g114
  (
    n334,
    n24
  );


  buf
  g115
  (
    n305,
    n84
  );


  buf
  g116
  (
    n216,
    n25
  );


  not
  g117
  (
    n124,
    n52
  );


  not
  g118
  (
    n267,
    n79
  );


  not
  g119
  (
    n322,
    n85
  );


  not
  g120
  (
    n219,
    n31
  );


  buf
  g121
  (
    n281,
    n35
  );


  not
  g122
  (
    n312,
    n64
  );


  not
  g123
  (
    n323,
    n83
  );


  buf
  g124
  (
    n228,
    n66
  );


  buf
  g125
  (
    KeyWire_0_16,
    n77
  );


  buf
  g126
  (
    n107,
    n58
  );


  buf
  g127
  (
    n270,
    n30
  );


  buf
  g128
  (
    n346,
    n19
  );


  not
  g129
  (
    n106,
    n81
  );


  not
  g130
  (
    n220,
    n72
  );


  not
  g131
  (
    n353,
    n83
  );


  buf
  g132
  (
    n374,
    n48
  );


  buf
  g133
  (
    n340,
    n41
  );


  buf
  g134
  (
    n368,
    n25
  );


  buf
  g135
  (
    n371,
    n54
  );


  buf
  g136
  (
    n174,
    n82
  );


  not
  g137
  (
    n206,
    n81
  );


  not
  g138
  (
    n332,
    n78
  );


  buf
  g139
  (
    n376,
    n84
  );


  not
  g140
  (
    n197,
    n43
  );


  buf
  g141
  (
    n360,
    n80
  );


  buf
  g142
  (
    n282,
    n49
  );


  not
  g143
  (
    n184,
    n74
  );


  not
  g144
  (
    n135,
    n55
  );


  buf
  g145
  (
    n287,
    n90
  );


  not
  g146
  (
    n199,
    n65
  );


  buf
  g147
  (
    n168,
    n85
  );


  not
  g148
  (
    n278,
    n22
  );


  buf
  g149
  (
    n109,
    n66
  );


  buf
  g150
  (
    n145,
    n87
  );


  buf
  g151
  (
    n294,
    n78
  );


  not
  g152
  (
    n231,
    n49
  );


  not
  g153
  (
    n170,
    n28
  );


  buf
  g154
  (
    n178,
    n83
  );


  buf
  g155
  (
    n137,
    n89
  );


  buf
  g156
  (
    n232,
    n89
  );


  buf
  g157
  (
    n261,
    n32
  );


  not
  g158
  (
    n177,
    n60
  );


  not
  g159
  (
    n306,
    n28
  );


  not
  g160
  (
    n291,
    n57
  );


  buf
  g161
  (
    n275,
    n47
  );


  not
  g162
  (
    KeyWire_0_60,
    n76
  );


  buf
  g163
  (
    n222,
    n22
  );


  buf
  g164
  (
    n165,
    n29
  );


  not
  g165
  (
    n325,
    n66
  );


  not
  g166
  (
    n300,
    n58
  );


  not
  g167
  (
    n195,
    n79
  );


  not
  g168
  (
    n279,
    n71
  );


  buf
  g169
  (
    n139,
    n21
  );


  not
  g170
  (
    n319,
    n76
  );


  buf
  g171
  (
    n317,
    n49
  );


  buf
  g172
  (
    n131,
    n69
  );


  not
  g173
  (
    n268,
    n80
  );


  buf
  g174
  (
    n351,
    n64
  );


  not
  g175
  (
    n344,
    n87
  );


  buf
  g176
  (
    n264,
    n55
  );


  buf
  g177
  (
    n108,
    n84
  );


  not
  g178
  (
    n227,
    n88
  );


  not
  g179
  (
    n166,
    n36
  );


  not
  g180
  (
    n101,
    n78
  );


  buf
  g181
  (
    n175,
    n42
  );


  not
  g182
  (
    n366,
    n44
  );


  not
  g183
  (
    n123,
    n86
  );


  buf
  g184
  (
    n329,
    n27
  );


  not
  g185
  (
    n239,
    n73
  );


  not
  g186
  (
    n299,
    n76
  );


  buf
  g187
  (
    n364,
    n52
  );


  not
  g188
  (
    n152,
    n25
  );


  not
  g189
  (
    n342,
    n27
  );


  not
  g190
  (
    n203,
    n38
  );


  buf
  g191
  (
    n167,
    n53
  );


  not
  g192
  (
    n377,
    n83
  );


  buf
  g193
  (
    n304,
    n22
  );


  buf
  g194
  (
    n314,
    n41
  );


  not
  g195
  (
    n243,
    n39
  );


  not
  g196
  (
    n125,
    n72
  );


  buf
  g197
  (
    n273,
    n47
  );


  not
  g198
  (
    n150,
    n52
  );


  not
  g199
  (
    n120,
    n80
  );


  not
  g200
  (
    n213,
    n52
  );


  not
  g201
  (
    n245,
    n49
  );


  not
  g202
  (
    n148,
    n56
  );


  not
  g203
  (
    n252,
    n56
  );


  buf
  g204
  (
    n223,
    n36
  );


  not
  g205
  (
    n350,
    n34
  );


  buf
  g206
  (
    n225,
    n45
  );


  not
  g207
  (
    n330,
    n41
  );


  not
  g208
  (
    n126,
    n48
  );


  buf
  g209
  (
    n230,
    n30
  );


  buf
  g210
  (
    n142,
    n25
  );


  not
  g211
  (
    n103,
    n51
  );


  not
  g212
  (
    n310,
    n67
  );


  buf
  g213
  (
    KeyWire_0_8,
    n46
  );


  not
  g214
  (
    n301,
    n53
  );


  buf
  g215
  (
    n187,
    n67
  );


  buf
  g216
  (
    n324,
    n41
  );


  not
  g217
  (
    n316,
    n63
  );


  not
  g218
  (
    n96,
    n39
  );


  not
  g219
  (
    n113,
    n88
  );


  not
  g220
  (
    n115,
    n48
  );


  buf
  g221
  (
    n338,
    n33
  );


  not
  g222
  (
    n233,
    n53
  );


  not
  g223
  (
    n180,
    n71
  );


  buf
  g224
  (
    n256,
    n23
  );


  buf
  g225
  (
    n246,
    n40
  );


  buf
  g226
  (
    n140,
    n58
  );


  buf
  g227
  (
    n333,
    n70
  );


  buf
  g228
  (
    n144,
    n21
  );


  not
  g229
  (
    n181,
    n26
  );


  buf
  g230
  (
    n248,
    n70
  );


  not
  g231
  (
    n365,
    n20
  );


  not
  g232
  (
    n104,
    n29
  );


  not
  g233
  (
    n276,
    n85
  );


  buf
  g234
  (
    n102,
    n51
  );


  buf
  g235
  (
    n262,
    n60
  );


  buf
  g236
  (
    n343,
    n57
  );


  buf
  g237
  (
    n117,
    n50
  );


  not
  g238
  (
    n176,
    n45
  );


  not
  g239
  (
    n215,
    n37
  );


  not
  g240
  (
    n163,
    n20
  );


  buf
  g241
  (
    n309,
    n80
  );


  not
  g242
  (
    n326,
    n44
  );


  not
  g243
  (
    n249,
    n55
  );


  not
  g244
  (
    n321,
    n71
  );


  buf
  g245
  (
    n158,
    n43
  );


  buf
  g246
  (
    n134,
    n47
  );


  not
  g247
  (
    n241,
    n74
  );


  buf
  g248
  (
    n224,
    n48
  );


  buf
  g249
  (
    n92,
    n50
  );


  buf
  g250
  (
    n132,
    n87
  );


  buf
  g251
  (
    n159,
    n74
  );


  buf
  g252
  (
    n202,
    n24
  );


  buf
  g253
  (
    n359,
    n86
  );


  buf
  g254
  (
    n286,
    n69
  );


  buf
  g255
  (
    n308,
    n26
  );


  not
  g256
  (
    n236,
    n46
  );


  not
  g257
  (
    n201,
    n27
  );


  buf
  g258
  (
    n114,
    n88
  );


  not
  g259
  (
    n151,
    n59
  );


  buf
  g260
  (
    n186,
    n67
  );


  buf
  g261
  (
    n266,
    n42
  );


  not
  g262
  (
    n147,
    n89
  );


  buf
  g263
  (
    n307,
    n68
  );


  buf
  g264
  (
    n280,
    n55
  );


  not
  g265
  (
    n182,
    n64
  );


  buf
  g266
  (
    n161,
    n37
  );


  not
  g267
  (
    n238,
    n21
  );


  buf
  g268
  (
    n214,
    n68
  );


  buf
  g269
  (
    n337,
    n90
  );


  buf
  g270
  (
    n179,
    n57
  );


  not
  g271
  (
    n149,
    n20
  );


  buf
  g272
  (
    n258,
    n22
  );


  not
  g273
  (
    n105,
    n67
  );


  not
  g274
  (
    n143,
    n40
  );


  not
  g275
  (
    n235,
    n31
  );


  buf
  g276
  (
    n98,
    n62
  );


  buf
  g277
  (
    n191,
    n72
  );


  not
  g278
  (
    n154,
    n77
  );


  not
  g279
  (
    n111,
    n39
  );


  buf
  g280
  (
    KeyWire_0_26,
    n56
  );


  not
  g281
  (
    n244,
    n72
  );


  buf
  g282
  (
    n356,
    n65
  );


  buf
  g283
  (
    KeyWire_0_14,
    n60
  );


  not
  g284
  (
    n110,
    n37
  );


  buf
  g285
  (
    n297,
    n28
  );


  buf
  g286
  (
    n221,
    n53
  );


  buf
  g287
  (
    n331,
    n19
  );


  not
  g288
  (
    n229,
    n61
  );


  not
  g289
  (
    n136,
    n63
  );


  not
  g290
  (
    KeyWire_0_27,
    n26
  );


  buf
  g291
  (
    n284,
    n57
  );


  buf
  g292
  (
    n363,
    n81
  );


  buf
  g293
  (
    n97,
    n20
  );


  not
  g294
  (
    n218,
    n86
  );


  not
  g295
  (
    n116,
    n82
  );


  not
  g296
  (
    n190,
    n78
  );


  buf
  g297
  (
    n240,
    n42
  );


  buf
  g298
  (
    n205,
    n23
  );


  not
  g299
  (
    n271,
    n59
  );


  not
  g300
  (
    n372,
    n21
  );


  not
  g301
  (
    n155,
    n28
  );


  not
  g302
  (
    n259,
    n24
  );


  buf
  g303
  (
    KeyWire_0_38,
    n30
  );


  not
  g304
  (
    n234,
    n31
  );


  not
  g305
  (
    n274,
    n43
  );


  buf
  g306
  (
    n129,
    n33
  );


  buf
  g307
  (
    KeyWire_0_34,
    n34
  );


  not
  g308
  (
    n295,
    n46
  );


  buf
  g309
  (
    n293,
    n65
  );


  buf
  g310
  (
    n313,
    n40
  );


  buf
  g311
  (
    n192,
    n39
  );


  buf
  g312
  (
    n146,
    n32
  );


  not
  g313
  (
    n95,
    n71
  );


  buf
  g314
  (
    n183,
    n50
  );


  buf
  g315
  (
    n193,
    n89
  );


  not
  g316
  (
    n341,
    n34
  );


  buf
  g317
  (
    n133,
    n68
  );


  buf
  g318
  (
    n292,
    n75
  );


  not
  g319
  (
    n207,
    n75
  );


  not
  g320
  (
    n141,
    n88
  );


  buf
  g321
  (
    n119,
    n23
  );


  not
  g322
  (
    n172,
    n51
  );


  buf
  g323
  (
    n209,
    n29
  );


  not
  g324
  (
    n247,
    n90
  );


  buf
  g325
  (
    n336,
    n54
  );


  buf
  g326
  (
    n277,
    n33
  );


  not
  g327
  (
    n358,
    n27
  );


  buf
  g328
  (
    n269,
    n59
  );


  buf
  g329
  (
    n94,
    n54
  );


  not
  g330
  (
    n91,
    n19
  );


  buf
  g331
  (
    n370,
    n68
  );


  not
  g332
  (
    n156,
    n38
  );


  not
  g333
  (
    n242,
    n33
  );


  not
  g334
  (
    n208,
    n42
  );


  not
  g335
  (
    n250,
    n26
  );


  buf
  g336
  (
    n171,
    n62
  );


  not
  g337
  (
    n217,
    n63
  );


  not
  g338
  (
    n335,
    n35
  );


  not
  g339
  (
    n327,
    n36
  );


  not
  g340
  (
    n288,
    n44
  );


  not
  g341
  (
    n354,
    n47
  );


  not
  g342
  (
    n194,
    n81
  );


  buf
  g343
  (
    n188,
    n29
  );


  buf
  g344
  (
    n348,
    n79
  );


  not
  g345
  (
    n237,
    n56
  );


  buf
  g346
  (
    n347,
    n86
  );


  buf
  g347
  (
    n189,
    n76
  );


  not
  g348
  (
    n185,
    n43
  );


  buf
  g349
  (
    n272,
    n34
  );


  not
  g350
  (
    n138,
    n77
  );


  buf
  g351
  (
    n253,
    n58
  );


  buf
  g352
  (
    n339,
    n59
  );


  buf
  g353
  (
    n373,
    n44
  );


  not
  g354
  (
    n99,
    n77
  );


  buf
  g355
  (
    n164,
    n38
  );


  buf
  g356
  (
    n283,
    n19
  );


  not
  g357
  (
    n311,
    n85
  );


  not
  g358
  (
    n100,
    n61
  );


  not
  g359
  (
    n449,
    n127
  );


  not
  g360
  (
    n424,
    n115
  );


  buf
  g361
  (
    n687,
    n105
  );


  buf
  g362
  (
    n499,
    n194
  );


  buf
  g363
  (
    n465,
    n224
  );


  not
  g364
  (
    n498,
    n228
  );


  not
  g365
  (
    n693,
    n264
  );


  buf
  g366
  (
    n488,
    n126
  );


  not
  g367
  (
    n559,
    n213
  );


  buf
  g368
  (
    n584,
    n134
  );


  buf
  g369
  (
    n598,
    n178
  );


  buf
  g370
  (
    n500,
    n342
  );


  buf
  g371
  (
    n599,
    n91
  );


  buf
  g372
  (
    n442,
    n183
  );


  buf
  g373
  (
    n624,
    n303
  );


  not
  g374
  (
    n415,
    n330
  );


  buf
  g375
  (
    n496,
    n288
  );


  not
  g376
  (
    n493,
    n214
  );


  buf
  g377
  (
    n565,
    n211
  );


  buf
  g378
  (
    n507,
    n167
  );


  buf
  g379
  (
    n515,
    n223
  );


  not
  g380
  (
    n631,
    n337
  );


  buf
  g381
  (
    n670,
    n303
  );


  not
  g382
  (
    n657,
    n187
  );


  buf
  g383
  (
    n528,
    n321
  );


  buf
  g384
  (
    n384,
    n353
  );


  not
  g385
  (
    n689,
    n181
  );


  not
  g386
  (
    n413,
    n307
  );


  not
  g387
  (
    n677,
    n311
  );


  not
  g388
  (
    n686,
    n339
  );


  buf
  g389
  (
    n616,
    n127
  );


  buf
  g390
  (
    n569,
    n256
  );


  buf
  g391
  (
    n523,
    n205
  );


  not
  g392
  (
    n640,
    n212
  );


  not
  g393
  (
    n471,
    n233
  );


  buf
  g394
  (
    n635,
    n188
  );


  not
  g395
  (
    n430,
    n251
  );


  not
  g396
  (
    n644,
    n330
  );


  not
  g397
  (
    n558,
    n255
  );


  buf
  g398
  (
    n634,
    n260
  );


  not
  g399
  (
    n426,
    n345
  );


  not
  g400
  (
    n382,
    n228
  );


  not
  g401
  (
    n590,
    n344
  );


  buf
  g402
  (
    n668,
    n327
  );


  buf
  g403
  (
    n683,
    n193
  );


  not
  g404
  (
    n655,
    n299
  );


  buf
  g405
  (
    n432,
    n345
  );


  not
  g406
  (
    n600,
    n251
  );


  not
  g407
  (
    n695,
    n322
  );


  buf
  g408
  (
    n630,
    n325
  );


  buf
  g409
  (
    n593,
    n232
  );


  not
  g410
  (
    n615,
    n207
  );


  buf
  g411
  (
    n535,
    n115
  );


  not
  g412
  (
    n632,
    n354
  );


  not
  g413
  (
    n556,
    n154
  );


  buf
  g414
  (
    n645,
    n349
  );


  not
  g415
  (
    n428,
    n332
  );


  not
  g416
  (
    n522,
    n323
  );


  not
  g417
  (
    n482,
    n249
  );


  buf
  g418
  (
    n472,
    n225
  );


  not
  g419
  (
    n563,
    n169
  );


  buf
  g420
  (
    n678,
    n195
  );


  buf
  g421
  (
    n444,
    n315
  );


  buf
  g422
  (
    n462,
    n202
  );


  not
  g423
  (
    n456,
    n315
  );


  buf
  g424
  (
    n652,
    n211
  );


  buf
  g425
  (
    n603,
    n236
  );


  buf
  g426
  (
    n682,
    n218
  );


  buf
  g427
  (
    n573,
    n152
  );


  not
  g428
  (
    n684,
    n273
  );


  not
  g429
  (
    n394,
    n330
  );


  buf
  g430
  (
    n418,
    n211
  );


  buf
  g431
  (
    n544,
    n202
  );


  not
  g432
  (
    n607,
    n185
  );


  buf
  g433
  (
    n551,
    n191
  );


  not
  g434
  (
    n529,
    n295
  );


  buf
  g435
  (
    n666,
    n133
  );


  not
  g436
  (
    n595,
    n281
  );


  buf
  g437
  (
    n495,
    n124
  );


  buf
  g438
  (
    n455,
    n208
  );


  buf
  g439
  (
    n427,
    n153
  );


  not
  g440
  (
    n450,
    n307
  );


  buf
  g441
  (
    n526,
    n344
  );


  buf
  g442
  (
    n660,
    n265
  );


  nand
  g443
  (
    n673,
    n165,
    n106,
    n335,
    n246
  );


  xor
  g444
  (
    n534,
    n161,
    n140,
    n175,
    n227
  );


  and
  g445
  (
    n393,
    n109,
    n312,
    n318,
    n280
  );


  nor
  g446
  (
    KeyWire_0_28,
    n334,
    n145,
    n184,
    n277
  );


  or
  g447
  (
    n699,
    n295,
    n141,
    n171,
    n241
  );


  nor
  g448
  (
    n613,
    n327,
    n247,
    n345,
    n323
  );


  xnor
  g449
  (
    n691,
    n272,
    n162,
    n274,
    n94
  );


  xor
  g450
  (
    n437,
    n175,
    n136,
    n121,
    n145
  );


  and
  g451
  (
    n397,
    n122,
    n178,
    n333,
    n360
  );


  or
  g452
  (
    n611,
    n237,
    n230,
    n125,
    n141
  );


  nand
  g453
  (
    n587,
    n214,
    n314,
    n322,
    n185
  );


  xor
  g454
  (
    n420,
    n267,
    n323,
    n213,
    n295
  );


  xor
  g455
  (
    n572,
    n304,
    n180,
    n266,
    n300
  );


  nor
  g456
  (
    n581,
    n155,
    n108,
    n292,
    n121
  );


  xnor
  g457
  (
    n548,
    n209,
    n128,
    n297,
    n319
  );


  nor
  g458
  (
    n486,
    n121,
    n164,
    n207,
    n142
  );


  nand
  g459
  (
    n416,
    n256,
    n301,
    n311,
    n103
  );


  xnor
  g460
  (
    n651,
    n282,
    n320,
    n297,
    n270
  );


  xor
  g461
  (
    n674,
    n324,
    n329,
    n220,
    n240
  );


  nand
  g462
  (
    KeyWire_0_56,
    n268,
    n318,
    n348,
    n144
  );


  xor
  g463
  (
    n386,
    n250,
    n274,
    n327,
    n114
  );


  and
  g464
  (
    n480,
    n269,
    n328,
    n287,
    n191
  );


  xnor
  g465
  (
    n509,
    n183,
    n139,
    n228,
    n203
  );


  xor
  g466
  (
    n469,
    n333,
    n166,
    n338,
    n289
  );


  and
  g467
  (
    n464,
    n357,
    n237,
    n204,
    n297
  );


  xnor
  g468
  (
    n560,
    n341,
    n299,
    n307,
    n316
  );


  xnor
  g469
  (
    n614,
    n342,
    n113,
    n145,
    n324
  );


  or
  g470
  (
    n606,
    n189,
    n96,
    n237,
    n196
  );


  nor
  g471
  (
    n467,
    n250,
    n151,
    n122,
    n169
  );


  nand
  g472
  (
    n574,
    n155,
    n167,
    n318,
    n334
  );


  or
  g473
  (
    n625,
    n270,
    n275,
    n340,
    n326
  );


  nand
  g474
  (
    n458,
    n265,
    n170,
    n358,
    n184
  );


  xor
  g475
  (
    n527,
    n204,
    n296,
    n259
  );


  xor
  g476
  (
    n445,
    n278,
    n277,
    n152,
    n220
  );


  nor
  g477
  (
    KeyWire_0_3,
    n122,
    n337,
    n138,
    n130
  );


  or
  g478
  (
    n566,
    n343,
    n231,
    n148,
    n216
  );


  and
  g479
  (
    n463,
    n179,
    n261,
    n176,
    n351
  );


  xor
  g480
  (
    n403,
    n97,
    n272,
    n128,
    n155
  );


  xnor
  g481
  (
    n435,
    n189,
    n126,
    n292,
    n291
  );


  xnor
  g482
  (
    n537,
    n132,
    n321,
    n351,
    n246
  );


  xor
  g483
  (
    n536,
    n313,
    n294,
    n253,
    n149
  );


  or
  g484
  (
    n505,
    n278,
    n160,
    n259,
    n118
  );


  nand
  g485
  (
    n654,
    n239,
    n137,
    n115,
    n278
  );


  xor
  g486
  (
    n454,
    n156,
    n275,
    n223,
    n274
  );


  nand
  g487
  (
    n609,
    n157,
    n164,
    n280,
    n289
  );


  nor
  g488
  (
    n398,
    n283,
    n147,
    n343,
    n357
  );


  nor
  g489
  (
    KeyWire_0_45,
    n219,
    n168,
    n156,
    n135
  );


  or
  g490
  (
    n494,
    n142,
    n110,
    n235,
    n201
  );


  or
  g491
  (
    n580,
    n181,
    n191,
    n132,
    n235
  );


  xnor
  g492
  (
    n491,
    n229,
    n221,
    n200,
    n95
  );


  and
  g493
  (
    KeyWire_0_37,
    n325,
    n338,
    n249,
    n196
  );


  nand
  g494
  (
    n696,
    n192,
    n340,
    n357,
    n329
  );


  nand
  g495
  (
    n410,
    n173,
    n99,
    n212,
    n248
  );


  or
  g496
  (
    n554,
    n336,
    n210,
    n279,
    n144
  );


  xor
  g497
  (
    n575,
    n298,
    n276,
    n236,
    n172
  );


  and
  g498
  (
    n502,
    n218,
    n230,
    n217,
    n264
  );


  and
  g499
  (
    n381,
    n245,
    n287,
    n347,
    n140
  );


  nor
  g500
  (
    n589,
    n291,
    n124,
    n336,
    n270
  );


  or
  g501
  (
    n530,
    n199,
    n114,
    n214,
    n112
  );


  nor
  g502
  (
    n648,
    n124,
    n203,
    n244,
    n186
  );


  xor
  g503
  (
    n588,
    n350,
    n257,
    n112,
    n217
  );


  nor
  g504
  (
    n661,
    n269,
    n210,
    n271,
    n182
  );


  or
  g505
  (
    n478,
    n248,
    n110,
    n288,
    n119
  );


  and
  g506
  (
    n436,
    n289,
    n162,
    n352,
    n250
  );


  and
  g507
  (
    n446,
    n104,
    n111,
    n243,
    n258
  );


  nand
  g508
  (
    n594,
    n184,
    n264,
    n229,
    n151
  );


  and
  g509
  (
    n545,
    n230,
    n242,
    n225,
    n304
  );


  xnor
  g510
  (
    n517,
    n190,
    n166,
    n232,
    n97
  );


  and
  g511
  (
    n601,
    n302,
    n301,
    n150,
    n232
  );


  and
  g512
  (
    n621,
    n309,
    n185,
    n195,
    n244
  );


  or
  g513
  (
    n380,
    n347,
    n210,
    n291,
    n174
  );


  xnor
  g514
  (
    n637,
    n206,
    n237,
    n159,
    n100
  );


  and
  g515
  (
    KeyWire_0_44,
    n346,
    n236,
    n234
  );


  nor
  g516
  (
    n567,
    n322,
    n180,
    n151,
    n92
  );


  nand
  g517
  (
    n385,
    n271,
    n341,
    n167,
    n351
  );


  or
  g518
  (
    n543,
    n162,
    n283,
    n216,
    n332
  );


  xnor
  g519
  (
    n667,
    n284,
    n98,
    n359,
    n331
  );


  xor
  g520
  (
    n685,
    n197,
    n273,
    n243,
    n198
  );


  nor
  g521
  (
    n383,
    n134,
    n313,
    n354,
    n130
  );


  nand
  g522
  (
    n562,
    n358,
    n119,
    n150,
    n164
  );


  nor
  g523
  (
    n447,
    n206,
    n267,
    n241,
    n240
  );


  xnor
  g524
  (
    n597,
    n332,
    n277,
    n335,
    n201
  );


  nor
  g525
  (
    n692,
    n172,
    n241,
    n293,
    n281
  );


  xnor
  g526
  (
    n697,
    n299,
    n349,
    n326,
    n344
  );


  and
  g527
  (
    n492,
    n285,
    n168,
    n281,
    n359
  );


  and
  g528
  (
    n516,
    n108,
    n210,
    n238,
    n311
  );


  xor
  g529
  (
    n407,
    n154,
    n221,
    n192,
    n144
  );


  nor
  g530
  (
    n514,
    n107,
    n113,
    n287,
    n219
  );


  and
  g531
  (
    n596,
    n341,
    n291,
    n166,
    n207
  );


  nor
  g532
  (
    n459,
    n219,
    n346,
    n178,
    n270
  );


  xor
  g533
  (
    n605,
    n178,
    n272,
    n243,
    n344
  );


  xnor
  g534
  (
    n421,
    n135,
    n123,
    n156,
    n208
  );


  or
  g535
  (
    n400,
    n159,
    n117,
    n113,
    n120
  );


  or
  g536
  (
    n391,
    n199,
    n165,
    n246,
    n273
  );


  xor
  g537
  (
    n675,
    n222,
    n127,
    n202,
    n264
  );


  xnor
  g538
  (
    n643,
    n253,
    n324,
    n153,
    n194
  );


  xor
  g539
  (
    n622,
    n177,
    n122,
    n307,
    n300
  );


  nand
  g540
  (
    n694,
    n314,
    n172,
    n134,
    n107
  );


  or
  g541
  (
    n577,
    n197,
    n101,
    n338,
    n255
  );


  nor
  g542
  (
    n379,
    n138,
    n261,
    n211,
    n158
  );


  nor
  g543
  (
    n629,
    n148,
    n276,
    n150,
    n258
  );


  nor
  g544
  (
    n490,
    n154,
    n287,
    n141,
    n143
  );


  or
  g545
  (
    n582,
    n151,
    n339,
    n204,
    n169
  );


  xnor
  g546
  (
    n489,
    n347,
    n206,
    n240,
    n360
  );


  or
  g547
  (
    n570,
    n298,
    n193,
    n202,
    n338
  );


  xnor
  g548
  (
    n402,
    n265,
    n233,
    n285,
    n356
  );


  nand
  g549
  (
    n612,
    n278,
    n227,
    n170,
    n326
  );


  xor
  g550
  (
    n404,
    n334,
    n230,
    n143,
    n163
  );


  xor
  g551
  (
    n513,
    n191,
    n279,
    n102,
    n179
  );


  and
  g552
  (
    n619,
    n279,
    n243,
    n284,
    n152
  );


  or
  g553
  (
    n389,
    n125,
    n284,
    n157,
    n241
  );


  nand
  g554
  (
    n409,
    n133,
    n215,
    n235,
    n142
  );


  xnor
  g555
  (
    n638,
    n262,
    n263,
    n91,
    n140
  );


  or
  g556
  (
    n628,
    n111,
    n106,
    n312,
    n262
  );


  xnor
  g557
  (
    n392,
    n186,
    n129,
    n195,
    n234
  );


  and
  g558
  (
    n451,
    n341,
    n193,
    n166,
    n315
  );


  xor
  g559
  (
    n477,
    n207,
    n102,
    n282,
    n114
  );


  xor
  g560
  (
    n608,
    n257,
    n251,
    n306,
    n170
  );


  and
  g561
  (
    n487,
    n201,
    n313,
    n184,
    n182
  );


  nand
  g562
  (
    n448,
    n119,
    n294,
    n246,
    n131
  );


  nand
  g563
  (
    n452,
    n336,
    n336,
    n161,
    n176
  );


  nor
  g564
  (
    n508,
    n139,
    n189,
    n304,
    n337
  );


  and
  g565
  (
    n610,
    n136,
    n123,
    n360,
    n321
  );


  nand
  g566
  (
    n656,
    n250,
    n267,
    n352,
    n312
  );


  xor
  g567
  (
    n519,
    n200,
    n348,
    n279,
    n129
  );


  nor
  g568
  (
    n460,
    n226,
    n128,
    n229,
    n231
  );


  nand
  g569
  (
    n497,
    n310,
    n139,
    n265,
    n248
  );


  nor
  g570
  (
    n592,
    n187,
    n294,
    n238,
    n357
  );


  xor
  g571
  (
    n623,
    n289,
    n254,
    n101,
    n99
  );


  nand
  g572
  (
    n602,
    n350,
    n257,
    n225
  );


  xnor
  g573
  (
    n378,
    n329,
    n208,
    n223,
    n245
  );


  xnor
  g574
  (
    n549,
    n160,
    n197,
    n93,
    n228
  );


  xnor
  g575
  (
    n422,
    n329,
    n159,
    n153,
    n266
  );


  and
  g576
  (
    KeyWire_0_41,
    n355,
    n306,
    n116,
    n220
  );


  xor
  g577
  (
    n676,
    n161,
    n212,
    n215,
    n352
  );


  nor
  g578
  (
    n503,
    n205,
    n299,
    n317,
    n325
  );


  xnor
  g579
  (
    n425,
    n354,
    n238,
    n247,
    n196
  );


  xnor
  g580
  (
    n440,
    n349,
    n258,
    n259,
    n109
  );


  and
  g581
  (
    n542,
    n309,
    n138,
    n227,
    n127
  );


  and
  g582
  (
    n501,
    n319,
    n267,
    n342,
    n286
  );


  nor
  g583
  (
    n443,
    n137,
    n216,
    n309,
    n295
  );


  nand
  g584
  (
    n531,
    n268,
    n117,
    n158,
    n162
  );


  nor
  g585
  (
    n476,
    n170,
    n304,
    n350,
    n260
  );


  or
  g586
  (
    n423,
    n239,
    n292,
    n224,
    n179
  );


  nor
  g587
  (
    n649,
    n248,
    n226,
    n253,
    n197
  );


  nand
  g588
  (
    n474,
    n266,
    n222,
    n339,
    n252
  );


  nor
  g589
  (
    n688,
    n310,
    n213,
    n105,
    n205
  );


  and
  g590
  (
    n561,
    n129,
    n231,
    n173,
    n315
  );


  xnor
  g591
  (
    n576,
    n314,
    n302,
    n293,
    n157
  );


  nor
  g592
  (
    n512,
    n114,
    n180,
    n158,
    n160
  );


  and
  g593
  (
    n564,
    n153,
    n117,
    n317,
    n200
  );


  and
  g594
  (
    n586,
    n206,
    n359,
    n355,
    n251
  );


  xor
  g595
  (
    n520,
    n298,
    n303,
    n343,
    n226
  );


  nand
  g596
  (
    n583,
    n138,
    n168,
    n189,
    n177
  );


  xnor
  g597
  (
    n396,
    n290,
    n176,
    n271,
    n346
  );


  or
  g598
  (
    n555,
    n174,
    n192,
    n346,
    n340
  );


  and
  g599
  (
    n641,
    n149,
    n252,
    n260,
    n305
  );


  and
  g600
  (
    n468,
    n118,
    n350,
    n332,
    n347
  );


  nand
  g601
  (
    n511,
    n133,
    n308,
    n275,
    n177
  );


  nor
  g602
  (
    KeyWire_0_12,
    n275,
    n253,
    n301,
    n302
  );


  xnor
  g603
  (
    n671,
    n190,
    n181,
    n224,
    n294
  );


  and
  g604
  (
    n639,
    n120,
    n182,
    n285,
    n339
  );


  nand
  g605
  (
    n479,
    n353,
    n215,
    n327,
    n290
  );


  xnor
  g606
  (
    n604,
    n196,
    n268,
    n193,
    n274
  );


  nand
  g607
  (
    n411,
    n116,
    n331,
    n254,
    n273
  );


  and
  g608
  (
    n647,
    n342,
    n147,
    n309,
    n190
  );


  xor
  g609
  (
    n510,
    n213,
    n348,
    n132,
    n171
  );


  and
  g610
  (
    n473,
    n301,
    n244,
    n100
  );


  nor
  g611
  (
    n550,
    n120,
    n348,
    n310,
    n245
  );


  or
  g612
  (
    KeyWire_0_32,
    n280,
    n186,
    n335,
    n145
  );


  nor
  g613
  (
    n431,
    n358,
    n222,
    n126,
    n263
  );


  and
  g614
  (
    n636,
    n152,
    n234,
    n165,
    n209
  );


  xor
  g615
  (
    n387,
    n224,
    n203,
    n254,
    n119
  );


  nor
  g616
  (
    n553,
    n143,
    n201,
    n272,
    n300
  );


  xor
  g617
  (
    n441,
    n104,
    n132,
    n276,
    n249
  );


  xor
  g618
  (
    n568,
    n174,
    n171,
    n280,
    n212
  );


  nor
  g619
  (
    n406,
    n181,
    n136,
    n356
  );


  xor
  g620
  (
    KeyWire_0_62,
    n198,
    n192,
    n195,
    n156
  );


  nor
  g621
  (
    n680,
    n354,
    n263,
    n320,
    n231
  );


  nor
  g622
  (
    n664,
    n163,
    n308,
    n194,
    n204
  );


  xnor
  g623
  (
    n571,
    n261,
    n328,
    n255,
    n245
  );


  nor
  g624
  (
    n483,
    n320,
    n136,
    n225,
    n305
  );


  and
  g625
  (
    n433,
    n159,
    n120,
    n345,
    n227
  );


  xnor
  g626
  (
    n524,
    n177,
    n306,
    n317,
    n175
  );


  xor
  g627
  (
    n405,
    n269,
    n263,
    n158,
    n239
  );


  xor
  g628
  (
    n525,
    n186,
    n296,
    n343,
    n266
  );


  xnor
  g629
  (
    n618,
    n259,
    n130,
    n129,
    n188
  );


  nand
  g630
  (
    n672,
    n305,
    n217,
    n288,
    n226
  );


  and
  g631
  (
    n466,
    n308,
    n168,
    n232,
    n113
  );


  and
  g632
  (
    n399,
    n217,
    n262,
    n200,
    n260
  );


  xor
  g633
  (
    n470,
    n98,
    n288,
    n123,
    n300
  );


  nand
  g634
  (
    n412,
    n355,
    n194,
    n233,
    n183
  );


  nor
  g635
  (
    n439,
    n351,
    n233,
    n125,
    n242
  );


  or
  g636
  (
    n627,
    n130,
    n276,
    n203,
    n310
  );


  nand
  g637
  (
    n665,
    n167,
    n216,
    n328,
    n185
  );


  nor
  g638
  (
    n690,
    n283,
    n116,
    n131,
    n282
  );


  xnor
  g639
  (
    n438,
    n256,
    n358,
    n296,
    n333
  );


  xor
  g640
  (
    n620,
    n290,
    n198,
    n199,
    n298
  );


  nand
  g641
  (
    n417,
    n187,
    n165,
    n116,
    n333
  );


  nand
  g642
  (
    KeyWire_0_22,
    n337,
    n146,
    n292,
    n256
  );


  nor
  g643
  (
    n698,
    n149,
    n218,
    n255,
    n219
  );


  xor
  g644
  (
    n485,
    n163,
    n252,
    n297,
    n220
  );


  or
  g645
  (
    n475,
    n209,
    n209,
    n334,
    n335
  );


  nand
  g646
  (
    n395,
    n316,
    n254,
    n360,
    n221
  );


  xor
  g647
  (
    n663,
    n115,
    n148,
    n199,
    n252
  );


  and
  g648
  (
    n681,
    n286,
    n271,
    n326,
    n268
  );


  xor
  g649
  (
    n579,
    n93,
    n281,
    n262,
    n308
  );


  nor
  g650
  (
    n617,
    n215,
    n121,
    n311,
    n117
  );


  xnor
  g651
  (
    n679,
    n277,
    n118,
    n331,
    n323
  );


  and
  g652
  (
    n401,
    n137,
    n161,
    n325,
    n284
  );


  or
  g653
  (
    n506,
    n355,
    n135,
    n155,
    n146
  );


  and
  g654
  (
    n539,
    n182,
    n269,
    n183,
    n313
  );


  and
  g655
  (
    n662,
    n128,
    n258,
    n188,
    n322
  );


  and
  g656
  (
    n429,
    n242,
    n124,
    n282,
    n144
  );


  xnor
  g657
  (
    n533,
    n148,
    n356,
    n143,
    n173
  );


  nand
  g658
  (
    n408,
    n94,
    n163,
    n92,
    n140
  );


  nor
  g659
  (
    n541,
    n221,
    n316,
    n150,
    n125
  );


  nand
  g660
  (
    n552,
    n103,
    n142,
    n190,
    n198
  );


  or
  g661
  (
    n414,
    n214,
    n293,
    n223,
    n187
  );


  nor
  g662
  (
    n484,
    n305,
    n247,
    n286,
    n172
  );


  nand
  g663
  (
    n591,
    n317,
    n146,
    n222,
    n286
  );


  xnor
  g664
  (
    n521,
    n290,
    n293,
    n218,
    n330
  );


  and
  g665
  (
    n659,
    n137,
    n242,
    n164,
    n126
  );


  xor
  g666
  (
    n538,
    n169,
    n96,
    n179,
    n352
  );


  and
  g667
  (
    n669,
    n131,
    n331,
    n302,
    n157
  );


  xnor
  g668
  (
    n419,
    n229,
    n312,
    n249,
    n149
  );


  xnor
  g669
  (
    n626,
    n123,
    n205,
    n235,
    n319
  );


  xor
  g670
  (
    n388,
    n359,
    n176,
    n285,
    n303
  );


  xnor
  g671
  (
    n642,
    n240,
    n318,
    n353,
    n171
  );


  or
  g672
  (
    KeyWire_0_6,
    n160,
    n324,
    n316,
    n349
  );


  nand
  g673
  (
    n390,
    n135,
    n319,
    n146,
    n139
  );


  nand
  g674
  (
    n546,
    n95,
    n131,
    n314,
    n188
  );


  nor
  g675
  (
    n658,
    n134,
    n328,
    n236,
    n133
  );


  nand
  g676
  (
    n540,
    n239,
    n175,
    n247,
    n283
  );


  nand
  g677
  (
    n653,
    n261,
    n321,
    n238,
    n353
  );


  nand
  g678
  (
    n457,
    n208,
    n320,
    n141,
    n147
  );


  xnor
  g679
  (
    n585,
    n118,
    n147,
    n306,
    n180
  );


  or
  g680
  (
    n646,
    n154,
    n340,
    n173,
    n174
  );


  not
  g681
  (
    KeyWire_0_59,
    n378
  );


  buf
  g682
  (
    n705,
    n402
  );


  not
  g683
  (
    n704,
    n389
  );


  not
  g684
  (
    n719,
    n382
  );


  buf
  g685
  (
    n700,
    n401
  );


  buf
  g686
  (
    n718,
    n385
  );


  buf
  g687
  (
    n711,
    n379
  );


  buf
  g688
  (
    n703,
    n398
  );


  buf
  g689
  (
    n701,
    n396
  );


  not
  g690
  (
    n710,
    n399
  );


  not
  g691
  (
    n721,
    n381
  );


  buf
  g692
  (
    n720,
    n405
  );


  not
  g693
  (
    n712,
    n392
  );


  not
  g694
  (
    n707,
    n403
  );


  not
  g695
  (
    n716,
    n383
  );


  buf
  g696
  (
    n702,
    n384
  );


  not
  g697
  (
    n709,
    n390
  );


  buf
  g698
  (
    n715,
    n400
  );


  buf
  g699
  (
    n713,
    n386
  );


  xnor
  g700
  (
    n708,
    n387,
    n395,
    n397
  );


  xor
  g701
  (
    n706,
    n391,
    n394,
    n393
  );


  xnor
  g702
  (
    n714,
    n404,
    n388,
    n380
  );


  not
  g703
  (
    n733,
    n703
  );


  buf
  g704
  (
    n735,
    n706
  );


  buf
  g705
  (
    n723,
    n410
  );


  buf
  g706
  (
    n734,
    n701
  );


  buf
  g707
  (
    n724,
    n707
  );


  buf
  g708
  (
    n726,
    n416
  );


  not
  g709
  (
    n736,
    n417
  );


  buf
  g710
  (
    n725,
    n415
  );


  not
  g711
  (
    n727,
    n418
  );


  buf
  g712
  (
    n732,
    n414
  );


  nor
  g713
  (
    n728,
    n708,
    n702,
    n705,
    n704
  );


  or
  g714
  (
    n730,
    n713,
    n420,
    n419,
    n411
  );


  nand
  g715
  (
    n729,
    n408,
    n714,
    n412,
    n711
  );


  or
  g716
  (
    n722,
    n413,
    n710,
    n712,
    n406
  );


  xor
  g717
  (
    n731,
    n700,
    n709,
    n409,
    n407
  );


  buf
  g718
  (
    n744,
    n728
  );


  not
  g719
  (
    n742,
    n730
  );


  buf
  g720
  (
    n740,
    n732
  );


  not
  g721
  (
    n745,
    n736
  );


  not
  g722
  (
    n739,
    n733
  );


  not
  g723
  (
    n737,
    n731
  );


  not
  g724
  (
    n741,
    n729
  );


  buf
  g725
  (
    n743,
    n735
  );


  not
  g726
  (
    n738,
    n734
  );


  not
  g727
  (
    n746,
    n727
  );


  buf
  g728
  (
    n752,
    n424
  );


  buf
  g729
  (
    n753,
    n740
  );


  buf
  g730
  (
    n747,
    n744
  );


  buf
  g731
  (
    n754,
    n743
  );


  not
  g732
  (
    n748,
    n739
  );


  not
  g733
  (
    n749,
    n738
  );


  xnor
  g734
  (
    n757,
    n427,
    n742,
    n737
  );


  xor
  g735
  (
    n759,
    n741,
    n741,
    n744,
    n423
  );


  nor
  g736
  (
    n762,
    n744,
    n429,
    n742,
    n422
  );


  nor
  g737
  (
    n761,
    n741,
    n739,
    n738
  );


  xor
  g738
  (
    n756,
    n739,
    n425,
    n745
  );


  and
  g739
  (
    n751,
    n741,
    n421,
    n426,
    n745
  );


  nand
  g740
  (
    n758,
    n744,
    n742,
    n739,
    n737
  );


  xor
  g741
  (
    n755,
    n428,
    n738,
    n740,
    n737
  );


  nor
  g742
  (
    KeyWire_0_42,
    n746,
    n743,
    n740
  );


  xor
  g743
  (
    n750,
    n740,
    n737,
    n743,
    n745
  );


  not
  g744
  (
    n763,
    n748
  );


  buf
  g745
  (
    n765,
    n749
  );


  not
  g746
  (
    n764,
    n751
  );


  buf
  g747
  (
    n767,
    n750
  );


  buf
  g748
  (
    n766,
    n747
  );


  buf
  g749
  (
    n778,
    n439
  );


  buf
  g750
  (
    n775,
    n436
  );


  buf
  g751
  (
    n777,
    n430
  );


  not
  g752
  (
    n774,
    n766
  );


  buf
  g753
  (
    n773,
    n764
  );


  buf
  g754
  (
    n772,
    n765
  );


  not
  g755
  (
    n771,
    n763
  );


  buf
  g756
  (
    n769,
    n763
  );


  or
  g757
  (
    n779,
    n438,
    n431,
    n765,
    n433
  );


  nand
  g758
  (
    n776,
    n765,
    n440,
    n764
  );


  nand
  g759
  (
    n768,
    n434,
    n765,
    n437,
    n435
  );


  and
  g760
  (
    n770,
    n432,
    n766,
    n441,
    n764
  );


  nor
  g761
  (
    n793,
    n777,
    n778,
    n717,
    n774
  );


  xor
  g762
  (
    n787,
    n363,
    n772,
    n771
  );


  nor
  g763
  (
    n786,
    n443,
    n361,
    n767,
    n774
  );


  nor
  g764
  (
    n799,
    n446,
    n448,
    n768,
    n361
  );


  and
  g765
  (
    n780,
    n779,
    n775,
    n719,
    n778
  );


  xor
  g766
  (
    n782,
    n770,
    n768,
    n716,
    n754
  );


  xnor
  g767
  (
    n791,
    n769,
    n769,
    n773,
    n776
  );


  and
  g768
  (
    n790,
    n445,
    n362,
    n777,
    n768
  );


  nor
  g769
  (
    n798,
    n758,
    n776,
    n775,
    n773
  );


  and
  g770
  (
    n800,
    n771,
    n773,
    n777,
    n774
  );


  xnor
  g771
  (
    n795,
    n769,
    n776,
    n779
  );


  nand
  g772
  (
    n797,
    n770,
    n362,
    n779
  );


  or
  g773
  (
    n792,
    n772,
    n362,
    n761,
    n363
  );


  or
  g774
  (
    n789,
    n449,
    n718,
    n767,
    n760
  );


  nor
  g775
  (
    n803,
    n778,
    n769,
    n454,
    n770
  );


  nor
  g776
  (
    n794,
    n772,
    n759,
    n450,
    n756
  );


  or
  g777
  (
    n785,
    n361,
    n771,
    n447,
    n720
  );


  xor
  g778
  (
    KeyWire_0_10,
    n768,
    n451,
    n770,
    n766
  );


  or
  g779
  (
    n783,
    n453,
    n455,
    n773,
    n442
  );


  and
  g780
  (
    n802,
    n774,
    n766,
    n721,
    n775
  );


  nand
  g781
  (
    n784,
    n755,
    n777,
    n753,
    n778
  );


  or
  g782
  (
    n788,
    n757,
    n767,
    n779,
    n762
  );


  xnor
  g783
  (
    n796,
    n444,
    n361,
    n775,
    n752
  );


  or
  g784
  (
    n801,
    n715,
    n767,
    n772,
    n452
  );


  buf
  g785
  (
    KeyWire_0_61,
    n456
  );


  not
  g786
  (
    n804,
    n364
  );


  not
  g787
  (
    n807,
    n783
  );


  not
  g788
  (
    n811,
    n787
  );


  not
  g789
  (
    n810,
    n791
  );


  not
  g790
  (
    n812,
    n786
  );


  not
  g791
  (
    n813,
    n364
  );


  not
  g792
  (
    n805,
    n794
  );


  nand
  g793
  (
    n815,
    n789,
    n364
  );


  and
  g794
  (
    n806,
    n365,
    n363,
    n793,
    n785
  );


  xnor
  g795
  (
    n808,
    n788,
    n363,
    n457,
    n364
  );


  xor
  g796
  (
    n814,
    n365,
    n784,
    n792,
    n790
  );


  buf
  g797
  (
    n818,
    n805
  );


  not
  g798
  (
    KeyWire_0_25,
    n804
  );


  not
  g799
  (
    n823,
    n458
  );


  not
  g800
  (
    n819,
    n806
  );


  not
  g801
  (
    n816,
    n807
  );


  buf
  g802
  (
    n817,
    n806
  );


  buf
  g803
  (
    n820,
    n804
  );


  not
  g804
  (
    n821,
    n808
  );


  buf
  g805
  (
    n822,
    n805
  );


  and
  g806
  (
    KeyWire_0_50,
    n459,
    n807,
    n808
  );


  and
  g807
  (
    n826,
    n368,
    n823,
    n376,
    n821
  );


  nand
  g808
  (
    KeyWire_0_39,
    n373,
    n811,
    n366,
    n371
  );


  nand
  g809
  (
    n845,
    n811,
    n369,
    n809,
    n824
  );


  nor
  g810
  (
    n831,
    n822,
    n373,
    n369,
    n365
  );


  or
  g811
  (
    n827,
    n377,
    n375,
    n366,
    n811
  );


  xor
  g812
  (
    n828,
    n375,
    n822,
    n371,
    n377
  );


  nand
  g813
  (
    n836,
    n372,
    n370,
    n368,
    n374
  );


  nor
  g814
  (
    n835,
    n365,
    n370,
    n816,
    n819
  );


  nand
  g815
  (
    n834,
    n820,
    n369,
    n372,
    n376
  );


  or
  g816
  (
    n833,
    n820,
    n825,
    n377,
    n824
  );


  nand
  g817
  (
    n840,
    n374,
    n809,
    n817,
    n810
  );


  and
  g818
  (
    n844,
    n810,
    n825,
    n823,
    n368
  );


  nand
  g819
  (
    n838,
    n374,
    n367,
    n373,
    n366
  );


  and
  g820
  (
    n841,
    n372,
    n810,
    n368,
    n817
  );


  xor
  g821
  (
    n830,
    n372,
    n810,
    n375,
    n374
  );


  xnor
  g822
  (
    n837,
    n371,
    n377,
    n376,
    n816
  );


  or
  g823
  (
    KeyWire_0_5,
    n818,
    n367,
    n371,
    n370
  );


  nor
  g824
  (
    n843,
    n819,
    n375,
    n373,
    n367
  );


  xor
  g825
  (
    n832,
    n376,
    n818,
    n811,
    n367
  );


  xor
  g826
  (
    n842,
    n821,
    n369,
    n366,
    n370
  );


  xor
  g827
  (
    n895,
    n603,
    n549,
    n591,
    n826
  );


  and
  g828
  (
    n864,
    n504,
    n568,
    n558,
    n837
  );


  nor
  g829
  (
    n909,
    n689,
    n697,
    n523,
    n594
  );


  xnor
  g830
  (
    n869,
    n670,
    n467,
    n536,
    n830
  );


  nand
  g831
  (
    n877,
    n526,
    n836,
    n831,
    n609
  );


  xnor
  g832
  (
    n919,
    n584,
    n469,
    n490,
    n593
  );


  xnor
  g833
  (
    n898,
    n648,
    n463,
    n472,
    n498
  );


  nor
  g834
  (
    n856,
    n838,
    n835,
    n840,
    n639
  );


  nor
  g835
  (
    n874,
    n843,
    n574,
    n642,
    n831
  );


  nand
  g836
  (
    n871,
    n841,
    n588,
    n559,
    n835
  );


  xnor
  g837
  (
    n882,
    n842,
    n634,
    n508,
    n845
  );


  or
  g838
  (
    n910,
    n630,
    n674,
    n649,
    n686
  );


  xnor
  g839
  (
    n904,
    n482,
    n519,
    n669,
    n628
  );


  nor
  g840
  (
    n851,
    n487,
    n570,
    n478,
    n622
  );


  xor
  g841
  (
    n860,
    n832,
    n605,
    n510,
    n585
  );


  nand
  g842
  (
    n907,
    n551,
    n481,
    n681,
    n842
  );


  xor
  g843
  (
    n892,
    n830,
    n600,
    n599,
    n460
  );


  or
  g844
  (
    n885,
    n627,
    n626,
    n483,
    n829
  );


  or
  g845
  (
    n918,
    n494,
    n631,
    n484,
    n563
  );


  and
  g846
  (
    n863,
    n667,
    n561,
    n839,
    n844
  );


  nor
  g847
  (
    n890,
    n629,
    n845,
    n534
  );


  or
  g848
  (
    n857,
    n842,
    n619,
    n830,
    n562
  );


  xnor
  g849
  (
    n881,
    n837,
    n655,
    n690,
    n607
  );


  xor
  g850
  (
    n862,
    n522,
    n625,
    n840,
    n533
  );


  and
  g851
  (
    n866,
    n836,
    n496,
    n583,
    n465
  );


  nor
  g852
  (
    n920,
    n592,
    n606,
    n473,
    n840
  );


  xor
  g853
  (
    n865,
    n844,
    n471,
    n571,
    n476
  );


  nand
  g854
  (
    n883,
    n596,
    n618,
    n462,
    n643
  );


  or
  g855
  (
    KeyWire_0_54,
    n497,
    n833,
    n615,
    n524
  );


  nor
  g856
  (
    n893,
    n545,
    n677,
    n513,
    n491
  );


  or
  g857
  (
    n913,
    n577,
    n663,
    n657,
    n698
  );


  xnor
  g858
  (
    n846,
    n586,
    n826,
    n833,
    n521
  );


  xnor
  g859
  (
    n897,
    n623,
    n612,
    n837,
    n687
  );


  or
  g860
  (
    n921,
    n838,
    n829,
    n500,
    n661
  );


  nand
  g861
  (
    n858,
    n516,
    n693,
    n515,
    n840
  );


  xor
  g862
  (
    n878,
    n832,
    n676,
    n839,
    n550
  );


  xnor
  g863
  (
    n894,
    n617,
    n553,
    n831,
    n844
  );


  xor
  g864
  (
    n879,
    n831,
    n837,
    n548,
    n828
  );


  xor
  g865
  (
    n888,
    n843,
    n517,
    n692,
    n488
  );


  or
  g866
  (
    n902,
    n827,
    n552,
    n554,
    n833
  );


  nor
  g867
  (
    n853,
    n645,
    n489,
    n486,
    n650
  );


  xnor
  g868
  (
    n906,
    n835,
    n503,
    n611,
    n509
  );


  xnor
  g869
  (
    n899,
    n827,
    n475,
    n841,
    n595
  );


  xor
  g870
  (
    n925,
    n679,
    n598,
    n646,
    n637
  );


  or
  g871
  (
    n861,
    n601,
    n699,
    n632,
    n839
  );


  xnor
  g872
  (
    n900,
    n544,
    n525,
    n613,
    n560
  );


  xor
  g873
  (
    n903,
    n836,
    n542,
    n529,
    n685
  );


  xor
  g874
  (
    n923,
    n535,
    n843,
    n573
  );


  nand
  g875
  (
    n854,
    n691,
    n507,
    n688,
    n479
  );


  or
  g876
  (
    n872,
    n835,
    n466,
    n581,
    n696
  );


  nor
  g877
  (
    n852,
    n575,
    n827,
    n682,
    n659
  );


  nor
  g878
  (
    n887,
    n566,
    n841,
    n511,
    n567
  );


  xor
  g879
  (
    n901,
    n638,
    n644,
    n633,
    n620
  );


  nor
  g880
  (
    n886,
    n501,
    n610,
    n537,
    n492
  );


  nand
  g881
  (
    n911,
    n464,
    n589,
    n624,
    n845
  );


  nand
  g882
  (
    n876,
    n532,
    n660,
    n541,
    n636
  );


  xnor
  g883
  (
    KeyWire_0_58,
    n652,
    n834,
    n461,
    n838
  );


  or
  g884
  (
    n915,
    n572,
    n662,
    n495,
    n485
  );


  nor
  g885
  (
    n848,
    n531,
    n505,
    n520,
    n833
  );


  or
  g886
  (
    n896,
    n654,
    n582,
    n512,
    n499
  );


  and
  g887
  (
    n875,
    n621,
    n836,
    n826,
    n828
  );


  xor
  g888
  (
    n889,
    n834,
    n514,
    n695,
    n608
  );


  xor
  g889
  (
    n867,
    n470,
    n543,
    n668,
    n834
  );


  xor
  g890
  (
    KeyWire_0_24,
    n656,
    n675,
    n826,
    n673
  );


  and
  g891
  (
    n912,
    n665,
    n556,
    n547,
    n842
  );


  xor
  g892
  (
    n868,
    n569,
    n832,
    n604,
    n678
  );


  and
  g893
  (
    n891,
    n590,
    n834,
    n579,
    n474
  );


  xnor
  g894
  (
    n849,
    n683,
    n578,
    n832,
    n538
  );


  nand
  g895
  (
    n916,
    n480,
    n651,
    n841,
    n602
  );


  and
  g896
  (
    n922,
    n565,
    n829,
    n664,
    n564
  );


  xor
  g897
  (
    n924,
    n502,
    n828,
    n587,
    n468
  );


  or
  g898
  (
    n917,
    n597,
    n830,
    n527,
    n658
  );


  nand
  g899
  (
    n855,
    n506,
    n838,
    n827,
    n555
  );


  xnor
  g900
  (
    n870,
    n557,
    n493,
    n653,
    n647
  );


  nand
  g901
  (
    n908,
    n839,
    n640,
    n684,
    n477
  );


  xnor
  g902
  (
    n847,
    n672,
    n530,
    n680,
    n641
  );


  or
  g903
  (
    n880,
    n539,
    n666,
    n580,
    n518
  );


  or
  g904
  (
    n905,
    n614,
    n844,
    n540,
    n616
  );


  nand
  g905
  (
    n884,
    n528,
    n635,
    n694,
    n546
  );


  nor
  g906
  (
    n850,
    n576,
    n828,
    n829,
    n671
  );


  not
  g907
  (
    n1072,
    n914
  );


  buf
  g908
  (
    n1220,
    n877
  );


  buf
  g909
  (
    n1213,
    n856
  );


  not
  g910
  (
    KeyWire_0_63,
    n925
  );


  buf
  g911
  (
    n944,
    n883
  );


  not
  g912
  (
    n1188,
    n860
  );


  not
  g913
  (
    n1132,
    n867
  );


  buf
  g914
  (
    n1051,
    n907
  );


  buf
  g915
  (
    n1119,
    n895
  );


  not
  g916
  (
    n1061,
    n853
  );


  not
  g917
  (
    n976,
    n846
  );


  not
  g918
  (
    KeyWire_0_4,
    n863
  );


  buf
  g919
  (
    n1084,
    n906
  );


  not
  g920
  (
    n1224,
    n910
  );


  not
  g921
  (
    n1242,
    n912
  );


  buf
  g922
  (
    n1212,
    n872
  );


  buf
  g923
  (
    n981,
    n874
  );


  not
  g924
  (
    n1234,
    n869
  );


  buf
  g925
  (
    n1029,
    n918
  );


  buf
  g926
  (
    n966,
    n901
  );


  not
  g927
  (
    n1148,
    n893
  );


  not
  g928
  (
    n1039,
    n916
  );


  buf
  g929
  (
    n984,
    n872
  );


  buf
  g930
  (
    n1187,
    n847
  );


  not
  g931
  (
    n1049,
    n920
  );


  buf
  g932
  (
    n1184,
    n871
  );


  buf
  g933
  (
    n1070,
    n900
  );


  not
  g934
  (
    n1133,
    n914
  );


  buf
  g935
  (
    n1062,
    n882
  );


  not
  g936
  (
    n1136,
    n863
  );


  buf
  g937
  (
    n1065,
    n859
  );


  buf
  g938
  (
    n1021,
    n908
  );


  not
  g939
  (
    n989,
    n855
  );


  buf
  g940
  (
    n1186,
    n858
  );


  not
  g941
  (
    n952,
    n902
  );


  not
  g942
  (
    n934,
    n862
  );


  not
  g943
  (
    n1205,
    n892
  );


  not
  g944
  (
    n930,
    n893
  );


  buf
  g945
  (
    n1128,
    n904
  );


  buf
  g946
  (
    n1019,
    n846
  );


  buf
  g947
  (
    n1001,
    n890
  );


  not
  g948
  (
    n975,
    n874
  );


  not
  g949
  (
    n932,
    n893
  );


  not
  g950
  (
    n1022,
    n883
  );


  buf
  g951
  (
    n946,
    n901
  );


  buf
  g952
  (
    n1056,
    n847
  );


  not
  g953
  (
    n1150,
    n904
  );


  not
  g954
  (
    n953,
    n897
  );


  not
  g955
  (
    n1174,
    n885
  );


  buf
  g956
  (
    n947,
    n912
  );


  not
  g957
  (
    n1141,
    n923
  );


  not
  g958
  (
    n1191,
    n870
  );


  buf
  g959
  (
    n1194,
    n922
  );


  not
  g960
  (
    n1211,
    n890
  );


  not
  g961
  (
    n977,
    n746
  );


  buf
  g962
  (
    n1083,
    n868
  );


  not
  g963
  (
    n948,
    n880
  );


  buf
  g964
  (
    n1091,
    n853
  );


  not
  g965
  (
    n1040,
    n898
  );


  not
  g966
  (
    n1153,
    n847
  );


  buf
  g967
  (
    n1202,
    n896
  );


  buf
  g968
  (
    n1203,
    n899
  );


  not
  g969
  (
    n1118,
    n914
  );


  not
  g970
  (
    n1121,
    n889
  );


  not
  g971
  (
    n1110,
    n886
  );


  not
  g972
  (
    n1164,
    n896
  );


  not
  g973
  (
    n1035,
    n901
  );


  buf
  g974
  (
    n1013,
    n876
  );


  buf
  g975
  (
    n1067,
    n857
  );


  not
  g976
  (
    n1077,
    n903
  );


  not
  g977
  (
    n1200,
    n913
  );


  not
  g978
  (
    n1126,
    n859
  );


  buf
  g979
  (
    n970,
    n904
  );


  not
  g980
  (
    n1243,
    n910
  );


  buf
  g981
  (
    n1076,
    n875
  );


  not
  g982
  (
    n1214,
    n865
  );


  not
  g983
  (
    n1099,
    n868
  );


  not
  g984
  (
    n962,
    n909
  );


  buf
  g985
  (
    n1221,
    n887
  );


  buf
  g986
  (
    n994,
    n920
  );


  buf
  g987
  (
    n1131,
    n862
  );


  not
  g988
  (
    n1219,
    n925
  );


  buf
  g989
  (
    n1055,
    n908
  );


  not
  g990
  (
    n1038,
    n860
  );


  buf
  g991
  (
    n1085,
    n859
  );


  not
  g992
  (
    n1011,
    n904
  );


  buf
  g993
  (
    n1017,
    n886
  );


  not
  g994
  (
    n1069,
    n852
  );


  buf
  g995
  (
    n1209,
    n918
  );


  not
  g996
  (
    n957,
    n876
  );


  not
  g997
  (
    n1223,
    n923
  );


  buf
  g998
  (
    n1037,
    n918
  );


  buf
  g999
  (
    n1168,
    n887
  );


  not
  g1000
  (
    n964,
    n746
  );


  buf
  g1001
  (
    n991,
    n868
  );


  buf
  g1002
  (
    n1016,
    n867
  );


  buf
  g1003
  (
    n1033,
    n889
  );


  buf
  g1004
  (
    n1095,
    n873
  );


  not
  g1005
  (
    n1192,
    n899
  );


  buf
  g1006
  (
    n945,
    n861
  );


  buf
  g1007
  (
    n1172,
    n856
  );


  not
  g1008
  (
    n1185,
    n884
  );


  not
  g1009
  (
    n980,
    n894
  );


  buf
  g1010
  (
    n1173,
    n881
  );


  buf
  g1011
  (
    n979,
    n850
  );


  buf
  g1012
  (
    n1103,
    n905
  );


  not
  g1013
  (
    n1031,
    n877
  );


  buf
  g1014
  (
    n963,
    n925
  );


  buf
  g1015
  (
    n1181,
    n923
  );


  not
  g1016
  (
    n1159,
    n851
  );


  buf
  g1017
  (
    n937,
    n849
  );


  buf
  g1018
  (
    n1167,
    n900
  );


  buf
  g1019
  (
    n1155,
    n883
  );


  not
  g1020
  (
    n1222,
    n875
  );


  not
  g1021
  (
    n998,
    n885
  );


  buf
  g1022
  (
    n1197,
    n850
  );


  not
  g1023
  (
    n1047,
    n919
  );


  buf
  g1024
  (
    n1127,
    n865
  );


  not
  g1025
  (
    n1079,
    n909
  );


  buf
  g1026
  (
    n1006,
    n886
  );


  not
  g1027
  (
    n972,
    n915
  );


  buf
  g1028
  (
    n993,
    n857
  );


  buf
  g1029
  (
    n1225,
    n876
  );


  buf
  g1030
  (
    n1052,
    n899
  );


  buf
  g1031
  (
    n1057,
    n922
  );


  buf
  g1032
  (
    n1180,
    n917
  );


  buf
  g1033
  (
    n992,
    n879
  );


  not
  g1034
  (
    n1044,
    n854
  );


  buf
  g1035
  (
    KeyWire_0_36,
    n882
  );


  not
  g1036
  (
    n1129,
    n858
  );


  not
  g1037
  (
    n1074,
    n867
  );


  buf
  g1038
  (
    n997,
    n864
  );


  not
  g1039
  (
    n1092,
    n848
  );


  buf
  g1040
  (
    n1160,
    n922
  );


  not
  g1041
  (
    n1170,
    n746
  );


  buf
  g1042
  (
    n1113,
    n881
  );


  not
  g1043
  (
    n1116,
    n878
  );


  not
  g1044
  (
    n1112,
    n917
  );


  buf
  g1045
  (
    n1000,
    n857
  );


  not
  g1046
  (
    n1165,
    n851
  );


  buf
  g1047
  (
    n974,
    n863
  );


  not
  g1048
  (
    n1097,
    n854
  );


  not
  g1049
  (
    n1054,
    n853
  );


  buf
  g1050
  (
    n1046,
    n912
  );


  not
  g1051
  (
    n985,
    n913
  );


  not
  g1052
  (
    n931,
    n870
  );


  buf
  g1053
  (
    n936,
    n855
  );


  not
  g1054
  (
    n1010,
    n882
  );


  buf
  g1055
  (
    n929,
    n855
  );


  buf
  g1056
  (
    n1124,
    n902
  );


  not
  g1057
  (
    n1012,
    n884
  );


  buf
  g1058
  (
    n1198,
    n864
  );


  not
  g1059
  (
    n967,
    n873
  );


  buf
  g1060
  (
    n1030,
    n867
  );


  not
  g1061
  (
    n1059,
    n902
  );


  not
  g1062
  (
    n1036,
    n888
  );


  buf
  g1063
  (
    n1082,
    n887
  );


  buf
  g1064
  (
    n1096,
    n878
  );


  buf
  g1065
  (
    n1080,
    n913
  );


  buf
  g1066
  (
    n1226,
    n847
  );


  buf
  g1067
  (
    n1195,
    n895
  );


  buf
  g1068
  (
    n1137,
    n921
  );


  not
  g1069
  (
    n961,
    n846
  );


  not
  g1070
  (
    n1125,
    n884
  );


  buf
  g1071
  (
    n1190,
    n894
  );


  buf
  g1072
  (
    n1115,
    n869
  );


  buf
  g1073
  (
    n1075,
    n915
  );


  buf
  g1074
  (
    n938,
    n916
  );


  buf
  g1075
  (
    n941,
    n920
  );


  buf
  g1076
  (
    n1064,
    n878
  );


  buf
  g1077
  (
    n1104,
    n861
  );


  not
  g1078
  (
    n1088,
    n871
  );


  not
  g1079
  (
    n1134,
    n874
  );


  buf
  g1080
  (
    n971,
    n922
  );


  not
  g1081
  (
    n1244,
    n911
  );


  not
  g1082
  (
    n1041,
    n899
  );


  not
  g1083
  (
    n1162,
    n921
  );


  buf
  g1084
  (
    n1149,
    n895
  );


  buf
  g1085
  (
    n1117,
    n898
  );


  buf
  g1086
  (
    n1239,
    n897
  );


  buf
  g1087
  (
    n940,
    n891
  );


  not
  g1088
  (
    n955,
    n857
  );


  buf
  g1089
  (
    n996,
    n849
  );


  buf
  g1090
  (
    n1229,
    n873
  );


  not
  g1091
  (
    n1098,
    n911
  );


  not
  g1092
  (
    n1063,
    n918
  );


  not
  g1093
  (
    n1023,
    n866
  );


  not
  g1094
  (
    n1108,
    n888
  );


  not
  g1095
  (
    n1086,
    n885
  );


  not
  g1096
  (
    n1178,
    n851
  );


  not
  g1097
  (
    n1025,
    n902
  );


  buf
  g1098
  (
    n1043,
    n891
  );


  not
  g1099
  (
    n1145,
    n860
  );


  buf
  g1100
  (
    n1105,
    n848
  );


  buf
  g1101
  (
    n960,
    n875
  );


  not
  g1102
  (
    n1120,
    n856
  );


  buf
  g1103
  (
    n1002,
    n905
  );


  buf
  g1104
  (
    n1045,
    n853
  );


  buf
  g1105
  (
    n999,
    n880
  );


  not
  g1106
  (
    n958,
    n916
  );


  not
  g1107
  (
    n1003,
    n903
  );


  not
  g1108
  (
    n1024,
    n848
  );


  buf
  g1109
  (
    n1210,
    n913
  );


  not
  g1110
  (
    n1179,
    n858
  );


  buf
  g1111
  (
    n1058,
    n895
  );


  buf
  g1112
  (
    n1007,
    n865
  );


  not
  g1113
  (
    n1216,
    n909
  );


  buf
  g1114
  (
    n1028,
    n916
  );


  not
  g1115
  (
    n1042,
    n881
  );


  not
  g1116
  (
    n965,
    n885
  );


  not
  g1117
  (
    n1094,
    n903
  );


  not
  g1118
  (
    n1235,
    n908
  );


  buf
  g1119
  (
    n943,
    n923
  );


  buf
  g1120
  (
    n1109,
    n909
  );


  buf
  g1121
  (
    n1166,
    n889
  );


  buf
  g1122
  (
    n1008,
    n878
  );


  buf
  g1123
  (
    n1230,
    n906
  );


  buf
  g1124
  (
    n1101,
    n888
  );


  not
  g1125
  (
    n1100,
    n848
  );


  not
  g1126
  (
    n951,
    n880
  );


  not
  g1127
  (
    n1199,
    n855
  );


  buf
  g1128
  (
    n982,
    n905
  );


  not
  g1129
  (
    n1154,
    n859
  );


  buf
  g1130
  (
    n990,
    n897
  );


  not
  g1131
  (
    n1169,
    n886
  );


  buf
  g1132
  (
    n1232,
    n919
  );


  not
  g1133
  (
    n1196,
    n870
  );


  not
  g1134
  (
    n1060,
    n892
  );


  not
  g1135
  (
    n935,
    n898
  );


  buf
  g1136
  (
    n1206,
    n868
  );


  buf
  g1137
  (
    n1143,
    n911
  );


  not
  g1138
  (
    n983,
    n891
  );


  not
  g1139
  (
    n978,
    n849
  );


  not
  g1140
  (
    n1176,
    n921
  );


  buf
  g1141
  (
    n1048,
    n917
  );


  buf
  g1142
  (
    n1147,
    n882
  );


  buf
  g1143
  (
    n1114,
    n852
  );


  buf
  g1144
  (
    n1102,
    n919
  );


  buf
  g1145
  (
    n1151,
    n864
  );


  not
  g1146
  (
    KeyWire_0_29,
    n854
  );


  not
  g1147
  (
    n1228,
    n863
  );


  not
  g1148
  (
    n1201,
    n890
  );


  buf
  g1149
  (
    n1161,
    n854
  );


  buf
  g1150
  (
    n1034,
    n915
  );


  not
  g1151
  (
    n1142,
    n849
  );


  buf
  g1152
  (
    n1171,
    n856
  );


  not
  g1153
  (
    n1053,
    n880
  );


  not
  g1154
  (
    n1090,
    n912
  );


  not
  g1155
  (
    n1111,
    n900
  );


  buf
  g1156
  (
    n988,
    n896
  );


  not
  g1157
  (
    n1018,
    n914
  );


  not
  g1158
  (
    n1093,
    n879
  );


  not
  g1159
  (
    n1004,
    n850
  );


  buf
  g1160
  (
    n949,
    n900
  );


  buf
  g1161
  (
    n1050,
    n850
  );


  buf
  g1162
  (
    n926,
    n920
  );


  buf
  g1163
  (
    n1233,
    n861
  );


  not
  g1164
  (
    n1130,
    n924
  );


  not
  g1165
  (
    n1218,
    n892
  );


  buf
  g1166
  (
    n1204,
    n869
  );


  buf
  g1167
  (
    n1005,
    n903
  );


  buf
  g1168
  (
    n1140,
    n894
  );


  buf
  g1169
  (
    n1014,
    n873
  );


  buf
  g1170
  (
    n939,
    n883
  );


  buf
  g1171
  (
    KeyWire_0_51,
    n852
  );


  buf
  g1172
  (
    n1177,
    n897
  );


  not
  g1173
  (
    n1020,
    n925
  );


  buf
  g1174
  (
    n927,
    n898
  );


  buf
  g1175
  (
    n1027,
    n864
  );


  buf
  g1176
  (
    n1107,
    n872
  );


  buf
  g1177
  (
    n950,
    n871
  );


  not
  g1178
  (
    n1026,
    n910
  );


  buf
  g1179
  (
    n1135,
    n851
  );


  not
  g1180
  (
    n956,
    n869
  );


  not
  g1181
  (
    n1241,
    n877
  );


  not
  g1182
  (
    n959,
    n865
  );


  buf
  g1183
  (
    n1208,
    n896
  );


  not
  g1184
  (
    n1071,
    n872
  );


  buf
  g1185
  (
    n928,
    n866
  );


  buf
  g1186
  (
    n987,
    n924
  );


  buf
  g1187
  (
    n1068,
    n862
  );


  not
  g1188
  (
    n1158,
    n877
  );


  not
  g1189
  (
    n1138,
    n894
  );


  buf
  g1190
  (
    n1078,
    n908
  );


  buf
  g1191
  (
    n1227,
    n911
  );


  buf
  g1192
  (
    n1175,
    n881
  );


  buf
  g1193
  (
    n1245,
    n866
  );


  not
  g1194
  (
    n1183,
    n919
  );


  not
  g1195
  (
    n968,
    n879
  );


  not
  g1196
  (
    n1032,
    n901
  );


  buf
  g1197
  (
    KeyWire_0_53,
    n874
  );


  buf
  g1198
  (
    n995,
    n892
  );


  not
  g1199
  (
    n942,
    n907
  );


  buf
  g1200
  (
    n973,
    n905
  );


  not
  g1201
  (
    n1106,
    n866
  );


  buf
  g1202
  (
    n1122,
    n870
  );


  not
  g1203
  (
    n1081,
    n924
  );


  buf
  g1204
  (
    n1182,
    n871
  );


  buf
  g1205
  (
    n986,
    n910
  );


  not
  g1206
  (
    n1146,
    n860
  );


  not
  g1207
  (
    n1066,
    n917
  );


  buf
  g1208
  (
    n1237,
    n862
  );


  buf
  g1209
  (
    n1240,
    n846
  );


  not
  g1210
  (
    n1087,
    n915
  );


  buf
  g1211
  (
    n1073,
    n884
  );


  not
  g1212
  (
    n1089,
    n891
  );


  not
  g1213
  (
    n1193,
    n924
  );


  not
  g1214
  (
    n933,
    n906
  );


  buf
  g1215
  (
    n1189,
    n888
  );


  not
  g1216
  (
    n1123,
    n879
  );


  not
  g1217
  (
    n1156,
    n893
  );


  buf
  g1218
  (
    n954,
    n875
  );


  not
  g1219
  (
    n1009,
    n861
  );


  not
  g1220
  (
    n1152,
    n907
  );


  not
  g1221
  (
    n1236,
    n887
  );


  not
  g1222
  (
    n1207,
    n889
  );


  not
  g1223
  (
    n969,
    n907
  );


  not
  g1224
  (
    KeyWire_0_17,
    n858
  );


  not
  g1225
  (
    n1238,
    n906
  );


  nor
  g1226
  (
    n1163,
    n921,
    n876,
    n852,
    n890
  );


  not
  g1227
  (
    n1543,
    n1218
  );


  not
  g1228
  (
    n1288,
    n1214
  );


  buf
  g1229
  (
    n1589,
    n1085
  );


  not
  g1230
  (
    n1553,
    n1070
  );


  buf
  g1231
  (
    n1426,
    n1129
  );


  not
  g1232
  (
    n1382,
    n1010
  );


  buf
  g1233
  (
    n1557,
    n1211
  );


  not
  g1234
  (
    n1263,
    n1116
  );


  buf
  g1235
  (
    n1345,
    n1105
  );


  not
  g1236
  (
    n1544,
    n1066
  );


  not
  g1237
  (
    n1403,
    n1100
  );


  buf
  g1238
  (
    n1281,
    n959
  );


  not
  g1239
  (
    n1620,
    n1036
  );


  not
  g1240
  (
    n1331,
    n1240
  );


  buf
  g1241
  (
    n1418,
    n1112
  );


  buf
  g1242
  (
    n1383,
    n1192
  );


  buf
  g1243
  (
    n1279,
    n1154
  );


  not
  g1244
  (
    n1249,
    n1159
  );


  buf
  g1245
  (
    n1457,
    n1141
  );


  buf
  g1246
  (
    n1365,
    n958
  );


  buf
  g1247
  (
    KeyWire_0_46,
    n977
  );


  buf
  g1248
  (
    n1539,
    n1218
  );


  not
  g1249
  (
    n1516,
    n1120
  );


  buf
  g1250
  (
    n1431,
    n1195
  );


  not
  g1251
  (
    n1491,
    n1156
  );


  not
  g1252
  (
    n1299,
    n1165
  );


  not
  g1253
  (
    n1573,
    n1041
  );


  not
  g1254
  (
    n1582,
    n1097
  );


  buf
  g1255
  (
    n1621,
    n1101
  );


  not
  g1256
  (
    KeyWire_0_52,
    n990
  );


  not
  g1257
  (
    n1294,
    n813
  );


  buf
  g1258
  (
    n1601,
    n1194
  );


  buf
  g1259
  (
    n1528,
    n931
  );


  buf
  g1260
  (
    n1465,
    n1155
  );


  not
  g1261
  (
    n1399,
    n935
  );


  not
  g1262
  (
    n1432,
    n963
  );


  buf
  g1263
  (
    n1260,
    n1075
  );


  not
  g1264
  (
    KeyWire_0_57,
    n962
  );


  not
  g1265
  (
    n1502,
    n977
  );


  buf
  g1266
  (
    KeyWire_0_23,
    n1065
  );


  not
  g1267
  (
    n1395,
    n1019
  );


  buf
  g1268
  (
    n1483,
    n1185
  );


  not
  g1269
  (
    n1257,
    n1143
  );


  not
  g1270
  (
    n1453,
    n992
  );


  not
  g1271
  (
    n1476,
    n952
  );


  not
  g1272
  (
    KeyWire_0_0,
    n1245
  );


  not
  g1273
  (
    n1380,
    n987
  );


  buf
  g1274
  (
    n1356,
    n989
  );


  not
  g1275
  (
    n1499,
    n965
  );


  buf
  g1276
  (
    n1473,
    n1080
  );


  not
  g1277
  (
    n1468,
    n1150
  );


  buf
  g1278
  (
    n1524,
    n1004
  );


  not
  g1279
  (
    n1459,
    n1095
  );


  buf
  g1280
  (
    n1298,
    n1045
  );


  not
  g1281
  (
    KeyWire_0_2,
    n1201
  );


  buf
  g1282
  (
    n1578,
    n1156
  );


  buf
  g1283
  (
    n1396,
    n1178
  );


  not
  g1284
  (
    n1277,
    n1051
  );


  buf
  g1285
  (
    n1333,
    n948
  );


  buf
  g1286
  (
    n1292,
    n1144
  );


  not
  g1287
  (
    n1291,
    n987
  );


  buf
  g1288
  (
    n1407,
    n956
  );


  buf
  g1289
  (
    n1314,
    n971
  );


  buf
  g1290
  (
    n1503,
    n1125
  );


  not
  g1291
  (
    n1306,
    n1080
  );


  buf
  g1292
  (
    n1551,
    n1072
  );


  not
  g1293
  (
    n1414,
    n1238
  );


  not
  g1294
  (
    n1246,
    n1074
  );


  not
  g1295
  (
    n1519,
    n1031
  );


  not
  g1296
  (
    n1265,
    n1229
  );


  buf
  g1297
  (
    n1247,
    n1059
  );


  buf
  g1298
  (
    n1509,
    n1135
  );


  not
  g1299
  (
    n1261,
    n1120
  );


  xor
  g1300
  (
    n1450,
    n1193,
    n991,
    n1121,
    n1056
  );


  nor
  g1301
  (
    n1445,
    n1169,
    n941,
    n1186,
    n1231
  );


  xnor
  g1302
  (
    n1375,
    n1212,
    n957,
    n1235,
    n984
  );


  nor
  g1303
  (
    n1506,
    n1234,
    n944,
    n1094,
    n1220
  );


  xnor
  g1304
  (
    n1487,
    n1015,
    n1099,
    n1067,
    n939
  );


  and
  g1305
  (
    n1255,
    n1031,
    n967,
    n1061,
    n1159
  );


  xnor
  g1306
  (
    n1355,
    n1053,
    n1173,
    n1029,
    n1146
  );


  nand
  g1307
  (
    n1612,
    n1122,
    n1030,
    n1100,
    n948
  );


  and
  g1308
  (
    n1317,
    n1216,
    n934,
    n1052,
    n1116
  );


  nand
  g1309
  (
    n1425,
    n1179,
    n1184,
    n1161,
    n1231
  );


  or
  g1310
  (
    n1325,
    n1166,
    n938,
    n1169,
    n1005
  );


  nand
  g1311
  (
    n1469,
    n1238,
    n1196,
    n1074,
    n1115
  );


  xnor
  g1312
  (
    n1262,
    n997,
    n978,
    n981,
    n1241
  );


  and
  g1313
  (
    KeyWire_0_18,
    n1168,
    n1001,
    n1171,
    n1209
  );


  nand
  g1314
  (
    n1283,
    n1038,
    n937,
    n1202,
    n1011
  );


  xor
  g1315
  (
    n1464,
    n1130,
    n1031,
    n936,
    n1139
  );


  nor
  g1316
  (
    n1477,
    n1141,
    n936,
    n948,
    n953
  );


  nand
  g1317
  (
    n1410,
    n1227,
    n1199,
    n1073,
    n1015
  );


  nor
  g1318
  (
    n1329,
    n1188,
    n1232,
    n1005,
    n1194
  );


  xnor
  g1319
  (
    n1254,
    n815,
    n1007,
    n983,
    n1188
  );


  xor
  g1320
  (
    n1598,
    n1133,
    n1132,
    n1076,
    n993
  );


  nand
  g1321
  (
    n1507,
    n1066,
    n992,
    n936,
    n1072
  );


  or
  g1322
  (
    n1388,
    n1208,
    n982,
    n1200,
    n1089
  );


  and
  g1323
  (
    n1344,
    n800,
    n931,
    n1030,
    n1092
  );


  or
  g1324
  (
    n1567,
    n1117,
    n803,
    n1108,
    n1163
  );


  nor
  g1325
  (
    n1374,
    n934,
    n1101,
    n1142,
    n1215
  );


  xor
  g1326
  (
    n1533,
    n1105,
    n1021,
    n1025,
    n986
  );


  nand
  g1327
  (
    n1293,
    n944,
    n999,
    n1010,
    n1043
  );


  or
  g1328
  (
    n1540,
    n1071,
    n1188,
    n1086,
    n1230
  );


  nor
  g1329
  (
    n1562,
    n955,
    n1214,
    n1211,
    n1131
  );


  or
  g1330
  (
    KeyWire_0_9,
    n1201,
    n977,
    n1238,
    n1151
  );


  and
  g1331
  (
    n1520,
    n1086,
    n990,
    n1207,
    n1145
  );


  and
  g1332
  (
    n1563,
    n1005,
    n1034,
    n1171,
    n1042
  );


  xnor
  g1333
  (
    n1327,
    n1150,
    n1111,
    n1028,
    n1241
  );


  and
  g1334
  (
    n1492,
    n814,
    n971,
    n1125,
    n1147
  );


  and
  g1335
  (
    n1347,
    n1026,
    n1064,
    n1186,
    n1200
  );


  or
  g1336
  (
    n1515,
    n983,
    n1042,
    n1222,
    n1031
  );


  nand
  g1337
  (
    n1367,
    n987,
    n1042,
    n1089,
    n927
  );


  xnor
  g1338
  (
    n1349,
    n944,
    n1162,
    n1195,
    n969
  );


  nor
  g1339
  (
    n1266,
    n1059,
    n993,
    n796,
    n957
  );


  and
  g1340
  (
    n1274,
    n933,
    n955,
    n1017,
    n1041
  );


  and
  g1341
  (
    n1276,
    n1225,
    n1085,
    n1119,
    n1223
  );


  xnor
  g1342
  (
    n1614,
    n934,
    n1240,
    n981,
    n1187
  );


  nand
  g1343
  (
    n1586,
    n1182,
    n1000,
    n1075,
    n949
  );


  xnor
  g1344
  (
    n1547,
    n1244,
    n953,
    n1173,
    n1050
  );


  xnor
  g1345
  (
    n1610,
    n1219,
    n1179,
    n1126,
    n1024
  );


  xor
  g1346
  (
    n1548,
    n1154,
    n1242,
    n930,
    n1244
  );


  nor
  g1347
  (
    n1555,
    n945,
    n1074,
    n1175,
    n999
  );


  and
  g1348
  (
    n1591,
    n1119,
    n946,
    n955,
    n1077
  );


  xnor
  g1349
  (
    n1311,
    n926,
    n982,
    n1069,
    n1191
  );


  nand
  g1350
  (
    n1273,
    n1204,
    n1189,
    n943,
    n1176
  );


  xnor
  g1351
  (
    n1359,
    n1171,
    n813,
    n948,
    n1057
  );


  nor
  g1352
  (
    n1438,
    n980,
    n1026,
    n1206,
    n985
  );


  xor
  g1353
  (
    n1310,
    n1128,
    n1157,
    n1163,
    n1167
  );


  nor
  g1354
  (
    n1518,
    n1105,
    n989,
    n1034,
    n1023
  );


  or
  g1355
  (
    n1575,
    n954,
    n1229,
    n1109,
    n1136
  );


  and
  g1356
  (
    n1510,
    n964,
    n984,
    n1047,
    n1152
  );


  nor
  g1357
  (
    n1566,
    n1197,
    n1129,
    n1182,
    n1071
  );


  nand
  g1358
  (
    n1618,
    n951,
    n1140,
    n1115,
    n1090
  );


  or
  g1359
  (
    n1448,
    n1034,
    n1209,
    n1054,
    n1173
  );


  xor
  g1360
  (
    n1489,
    n999,
    n1101,
    n960,
    n1114
  );


  or
  g1361
  (
    KeyWire_0_48,
    n1047,
    n1225,
    n983,
    n1048
  );


  xnor
  g1362
  (
    n1564,
    n1033,
    n1178,
    n1192,
    n1114
  );


  or
  g1363
  (
    n1400,
    n1036,
    n1169,
    n1128,
    n1087
  );


  or
  g1364
  (
    n1308,
    n1159,
    n1167,
    n1242,
    n1140
  );


  and
  g1365
  (
    n1424,
    n985,
    n1046,
    n1157,
    n1011
  );


  xnor
  g1366
  (
    n1581,
    n940,
    n1079,
    n927,
    n1172
  );


  nor
  g1367
  (
    n1606,
    n1052,
    n1210,
    n1107,
    n972
  );


  nand
  g1368
  (
    n1330,
    n976,
    n1032,
    n1122,
    n943
  );


  xnor
  g1369
  (
    n1398,
    n812,
    n1016,
    n1176,
    n1049
  );


  xor
  g1370
  (
    n1576,
    n1170,
    n1002,
    n947,
    n1139
  );


  xor
  g1371
  (
    n1337,
    n1098,
    n801,
    n975,
    n966
  );


  nand
  g1372
  (
    n1602,
    n1151,
    n1070,
    n1108,
    n1123
  );


  nand
  g1373
  (
    n1268,
    n1094,
    n1018,
    n1148,
    n982
  );


  or
  g1374
  (
    n1405,
    n1022,
    n1108,
    n1193,
    n1064
  );


  xnor
  g1375
  (
    n1286,
    n1190,
    n1027,
    n1045,
    n929
  );


  and
  g1376
  (
    n1622,
    n1120,
    n1020,
    n1067,
    n988
  );


  xnor
  g1377
  (
    n1433,
    n1158,
    n1118,
    n1007,
    n1046
  );


  xnor
  g1378
  (
    n1603,
    n1021,
    n1137,
    n1032,
    n1106
  );


  and
  g1379
  (
    n1530,
    n998,
    n1139,
    n1066,
    n1046
  );


  or
  g1380
  (
    n1542,
    n1220,
    n1108,
    n995,
    n952
  );


  nor
  g1381
  (
    n1363,
    n1014,
    n1069,
    n1161,
    n988
  );


  xor
  g1382
  (
    n1258,
    n954,
    n1106,
    n1177,
    n1112
  );


  xor
  g1383
  (
    n1318,
    n1085,
    n1037,
    n1143,
    n1211
  );


  or
  g1384
  (
    n1478,
    n1007,
    n1063,
    n1112,
    n1212
  );


  or
  g1385
  (
    n1437,
    n1004,
    n1165,
    n1208,
    n1140
  );


  nand
  g1386
  (
    n1590,
    n1017,
    n1187,
    n1016,
    n1204
  );


  xnor
  g1387
  (
    KeyWire_0_19,
    n1234,
    n1148,
    n1013,
    n1029
  );


  nand
  g1388
  (
    n1259,
    n1097,
    n1189,
    n1012,
    n1244
  );


  nand
  g1389
  (
    n1368,
    n1194,
    n1227,
    n1008,
    n978
  );


  and
  g1390
  (
    n1289,
    n957,
    n1018,
    n1020,
    n1023
  );


  nand
  g1391
  (
    n1313,
    n1096,
    n994,
    n966,
    n958
  );


  nand
  g1392
  (
    n1360,
    n1053,
    n1162,
    n1100,
    n1051
  );


  or
  g1393
  (
    n1419,
    n1226,
    n930,
    n962,
    n1013
  );


  and
  g1394
  (
    n1427,
    n984,
    n941,
    n1063,
    n1196
  );


  xor
  g1395
  (
    n1269,
    n965,
    n1232,
    n1134,
    n1236
  );


  xnor
  g1396
  (
    KeyWire_0_40,
    n1079,
    n1211,
    n933,
    n1143
  );


  nand
  g1397
  (
    n1511,
    n1105,
    n1224,
    n1094,
    n1231
  );


  nor
  g1398
  (
    n1532,
    n1165,
    n1065,
    n1050,
    n1000
  );


  or
  g1399
  (
    n1583,
    n1215,
    n1241,
    n1088,
    n1130
  );


  or
  g1400
  (
    n1334,
    n996,
    n1155,
    n1233,
    n1009
  );


  and
  g1401
  (
    n1357,
    n1180,
    n814,
    n1024,
    n966
  );


  xnor
  g1402
  (
    n1596,
    n939,
    n1118,
    n1098,
    n1171
  );


  or
  g1403
  (
    n1434,
    n1168,
    n1069,
    n1058,
    n1084
  );


  xnor
  g1404
  (
    n1324,
    n1185,
    n976,
    n1018,
    n928
  );


  and
  g1405
  (
    n1541,
    n1227,
    n1152,
    n1079,
    n1216
  );


  xor
  g1406
  (
    n1381,
    n1162,
    n1175,
    n1136,
    n1047
  );


  xnor
  g1407
  (
    n1546,
    n967,
    n798,
    n1149,
    n1155
  );


  xor
  g1408
  (
    n1336,
    n958,
    n1010,
    n1154,
    n1060
  );


  nor
  g1409
  (
    n1561,
    n1158,
    n1061,
    n978,
    n1060
  );


  and
  g1410
  (
    n1471,
    n1210,
    n1025,
    n971,
    n1158
  );


  xor
  g1411
  (
    n1462,
    n1080,
    n1197,
    n1009,
    n1148
  );


  xor
  g1412
  (
    n1393,
    n930,
    n963,
    n1156,
    n945
  );


  or
  g1413
  (
    n1369,
    n965,
    n1043,
    n1141,
    n975
  );


  nand
  g1414
  (
    n1538,
    n1180,
    n1060,
    n1206,
    n1088
  );


  xnor
  g1415
  (
    n1415,
    n1198,
    n1010,
    n963,
    n1025
  );


  xor
  g1416
  (
    n1529,
    n1049,
    n945,
    n1023,
    n955
  );


  xnor
  g1417
  (
    n1625,
    n813,
    n1030,
    n1135,
    n1158
  );


  or
  g1418
  (
    n1332,
    n1039,
    n1116,
    n993,
    n931
  );


  xnor
  g1419
  (
    n1303,
    n1127,
    n1000,
    n1024,
    n1100
  );


  nor
  g1420
  (
    n1456,
    n1029,
    n1083,
    n1153,
    n1133
  );


  xor
  g1421
  (
    n1467,
    n1066,
    n1187,
    n1138,
    n999
  );


  or
  g1422
  (
    n1421,
    n1222,
    n1230,
    n1086,
    n970
  );


  or
  g1423
  (
    n1508,
    n1215,
    n1081,
    n941,
    n1137
  );


  xor
  g1424
  (
    n1420,
    n938,
    n1151,
    n1206,
    n1065
  );


  xnor
  g1425
  (
    n1585,
    n1186,
    n1243,
    n1198,
    n991
  );


  or
  g1426
  (
    n1423,
    n1164,
    n1038,
    n1094,
    n1087
  );


  nor
  g1427
  (
    n1446,
    n1228,
    n1077,
    n1225,
    n1137
  );


  nand
  g1428
  (
    n1376,
    n1182,
    n1001,
    n928,
    n1073
  );


  and
  g1429
  (
    n1615,
    n1204,
    n1027,
    n1172,
    n1020
  );


  or
  g1430
  (
    KeyWire_0_1,
    n1036,
    n1220,
    n1129,
    n956
  );


  xor
  g1431
  (
    n1411,
    n996,
    n1199,
    n932,
    n1221
  );


  nor
  g1432
  (
    n1304,
    n1087,
    n1087,
    n1210,
    n1033
  );


  and
  g1433
  (
    n1402,
    n950,
    n1191,
    n1190,
    n1168
  );


  xor
  g1434
  (
    n1290,
    n986,
    n1206,
    n1067,
    n949
  );


  or
  g1435
  (
    n1505,
    n1179,
    n1210,
    n1245,
    n1199
  );


  xor
  g1436
  (
    n1430,
    n1141,
    n1208,
    n802,
    n1059
  );


  and
  g1437
  (
    n1394,
    n1091,
    n815,
    n1040,
    n1226
  );


  nor
  g1438
  (
    n1364,
    n1051,
    n1232,
    n1160,
    n1043
  );


  xnor
  g1439
  (
    n1439,
    n998,
    n1028,
    n1109,
    n1122
  );


  nand
  g1440
  (
    n1624,
    n974,
    n976,
    n956,
    n1006
  );


  nand
  g1441
  (
    n1305,
    n1023,
    n1102,
    n1068,
    n1197
  );


  or
  g1442
  (
    n1417,
    n1076,
    n1183,
    n1044,
    n1113
  );


  xor
  g1443
  (
    n1301,
    n1002,
    n991,
    n969,
    n1104
  );


  or
  g1444
  (
    n1514,
    n1103,
    n1151,
    n1051,
    n1008
  );


  xnor
  g1445
  (
    n1341,
    n1003,
    n1233,
    n1102,
    n1142
  );


  xor
  g1446
  (
    n1250,
    n1134,
    n1128,
    n960,
    n968
  );


  or
  g1447
  (
    n1593,
    n1190,
    n1040,
    n1062,
    n1113
  );


  or
  g1448
  (
    n1626,
    n1128,
    n1053,
    n1236,
    n1003
  );


  or
  g1449
  (
    n1587,
    n1070,
    n1172,
    n957,
    n962
  );


  xor
  g1450
  (
    n1335,
    n1004,
    n1117,
    n1097,
    n1091
  );


  nand
  g1451
  (
    n1323,
    n1032,
    n973,
    n951,
    n1121
  );


  xor
  g1452
  (
    n1338,
    n1213,
    n1040,
    n1146,
    n1006
  );


  xnor
  g1453
  (
    n1390,
    n1237,
    n950,
    n1002,
    n1043
  );


  and
  g1454
  (
    n1389,
    n1140,
    n938,
    n972,
    n1208
  );


  nand
  g1455
  (
    n1379,
    n1135,
    n1195,
    n979,
    n932
  );


  xor
  g1456
  (
    n1574,
    n983,
    n1132,
    n1138,
    n940
  );


  nand
  g1457
  (
    n1353,
    n1005,
    n1219,
    n1121,
    n1242
  );


  or
  g1458
  (
    n1623,
    n942,
    n814,
    n1181,
    n1035
  );


  xnor
  g1459
  (
    n1535,
    n1103,
    n1037,
    n1233,
    n985
  );


  or
  g1460
  (
    n1588,
    n1149,
    n1149,
    n1056,
    n1223
  );


  and
  g1461
  (
    n1251,
    n815,
    n1239,
    n1166,
    n937
  );


  xnor
  g1462
  (
    n1495,
    n1088,
    n1132,
    n1004,
    n1184
  );


  nor
  g1463
  (
    n1316,
    n1053,
    n931,
    n961,
    n1132
  );


  nor
  g1464
  (
    n1497,
    n1075,
    n1217,
    n926,
    n1102
  );


  nand
  g1465
  (
    n1454,
    n975,
    n941,
    n952,
    n997
  );


  nor
  g1466
  (
    n1531,
    n932,
    n1096,
    n1146,
    n970
  );


  xnor
  g1467
  (
    n1609,
    n1033,
    n1070,
    n1224,
    n812
  );


  nor
  g1468
  (
    n1354,
    n1081,
    n946,
    n1083,
    n1109
  );


  nor
  g1469
  (
    n1493,
    n1078,
    n1143,
    n1213,
    n949
  );


  nand
  g1470
  (
    n1406,
    n1124,
    n1037,
    n1209,
    n1014
  );


  nand
  g1471
  (
    n1608,
    n1239,
    n1202,
    n1190,
    n1147
  );


  xnor
  g1472
  (
    n1577,
    n1177,
    n1212,
    n995,
    n994
  );


  xnor
  g1473
  (
    n1348,
    n1205,
    n1194,
    n967,
    n1209
  );


  xnor
  g1474
  (
    n1455,
    n1045,
    n1207,
    n934,
    n1133
  );


  or
  g1475
  (
    n1267,
    n1201,
    n1178,
    n1081,
    n1073
  );


  xor
  g1476
  (
    n1319,
    n795,
    n1176,
    n1002,
    n1006
  );


  or
  g1477
  (
    n1440,
    n1136,
    n1134,
    n1191,
    n973
  );


  xor
  g1478
  (
    n1253,
    n1181,
    n1019,
    n953,
    n1065
  );


  xor
  g1479
  (
    n1297,
    n1229,
    n1057,
    n1137,
    n1230
  );


  xor
  g1480
  (
    n1580,
    n1032,
    n942,
    n1076,
    n1089
  );


  xnor
  g1481
  (
    n1568,
    n986,
    n1219,
    n1174,
    n1014
  );


  and
  g1482
  (
    n1328,
    n1228,
    n953,
    n1124,
    n1062
  );


  xor
  g1483
  (
    n1412,
    n975,
    n1041,
    n1034,
    n1121
  );


  and
  g1484
  (
    KeyWire_0_13,
    n1039,
    n1058,
    n980,
    n1111
  );


  xnor
  g1485
  (
    n1560,
    n982,
    n1117,
    n926,
    n1144
  );


  xor
  g1486
  (
    n1436,
    n1022,
    n990,
    n1238,
    n1024
  );


  nor
  g1487
  (
    n1550,
    n1123,
    n1075,
    n1035,
    n1203
  );


  nor
  g1488
  (
    n1604,
    n1198,
    n946,
    n1020,
    n1203
  );


  xor
  g1489
  (
    n1616,
    n1203,
    n961,
    n1104,
    n1074
  );


  and
  g1490
  (
    n1256,
    n1188,
    n962,
    n1027,
    n1178
  );


  or
  g1491
  (
    n1248,
    n1203,
    n1003,
    n1009,
    n996
  );


  nand
  g1492
  (
    n1472,
    n1042,
    n959,
    n1035,
    n998
  );


  nor
  g1493
  (
    n1504,
    n1205,
    n1060,
    n973,
    n1035
  );


  nand
  g1494
  (
    n1361,
    n1022,
    n1222,
    n1110,
    n947
  );


  xnor
  g1495
  (
    n1285,
    n1218,
    n1170,
    n974,
    n1038
  );


  xnor
  g1496
  (
    n1458,
    n1124,
    n1199,
    n1163,
    n968
  );


  nor
  g1497
  (
    n1534,
    n972,
    n981,
    n1236,
    n1226
  );


  xnor
  g1498
  (
    n1312,
    n935,
    n1142,
    n1056,
    n1243
  );


  nand
  g1499
  (
    n1416,
    n1007,
    n954,
    n950,
    n1184
  );


  or
  g1500
  (
    n1558,
    n1078,
    n1059,
    n986,
    n1011
  );


  or
  g1501
  (
    n1377,
    n1014,
    n1142,
    n1125,
    n1221
  );


  xor
  g1502
  (
    n1385,
    n980,
    n1122,
    n1085,
    n1223
  );


  and
  g1503
  (
    n1490,
    n1090,
    n1077,
    n1113,
    n970
  );


  nor
  g1504
  (
    n1397,
    n1177,
    n977,
    n1148,
    n1119
  );


  nor
  g1505
  (
    n1463,
    n1044,
    n1078,
    n1167,
    n939
  );


  xnor
  g1506
  (
    n1461,
    n1082,
    n937,
    n964,
    n1225
  );


  xnor
  g1507
  (
    n1321,
    n1050,
    n1117,
    n1073,
    n958
  );


  and
  g1508
  (
    n1552,
    n952,
    n1200,
    n1243,
    n997
  );


  or
  g1509
  (
    n1442,
    n1086,
    n979,
    n1013,
    n1044
  );


  nor
  g1510
  (
    n1282,
    n1160,
    n1000,
    n1164,
    n929
  );


  or
  g1511
  (
    n1549,
    n1088,
    n1072,
    n1135,
    n1196
  );


  xnor
  g1512
  (
    n1449,
    n1106,
    n1048,
    n970,
    n943
  );


  nor
  g1513
  (
    KeyWire_0_20,
    n1093,
    n1114,
    n933,
    n981
  );


  xor
  g1514
  (
    n1466,
    n1131,
    n960,
    n1150,
    n1154
  );


  nand
  g1515
  (
    n1300,
    n959,
    n935,
    n1124,
    n1092
  );


  or
  g1516
  (
    n1351,
    n1039,
    n928,
    n971,
    n1217
  );


  nor
  g1517
  (
    n1527,
    n1054,
    n1054,
    n1182,
    n813
  );


  xor
  g1518
  (
    n1302,
    n1116,
    n1177,
    n976,
    n1183
  );


  or
  g1519
  (
    KeyWire_0_21,
    n1037,
    n1099,
    n1127,
    n947
  );


  nand
  g1520
  (
    KeyWire_0_43,
    n1138,
    n933,
    n1164,
    n1092
  );


  nor
  g1521
  (
    n1545,
    n1025,
    n1239,
    n1084,
    n993
  );


  nor
  g1522
  (
    n1392,
    n1245,
    n959,
    n935,
    n994
  );


  xor
  g1523
  (
    n1480,
    n968,
    n1012,
    n1168,
    n974
  );


  xor
  g1524
  (
    KeyWire_0_49,
    n1235,
    n1241,
    n1054,
    n1017
  );


  xnor
  g1525
  (
    n1287,
    n1039,
    n1111,
    n1013,
    n1058
  );


  xnor
  g1526
  (
    n1441,
    n1175,
    n1017,
    n1163,
    n1016
  );


  nand
  g1527
  (
    n1343,
    n1026,
    n1089,
    n943,
    n1166
  );


  and
  g1528
  (
    n1486,
    n1069,
    n1131,
    n815,
    n1198
  );


  xnor
  g1529
  (
    n1309,
    n1106,
    n1189,
    n1201,
    n1062
  );


  xor
  g1530
  (
    n1460,
    n1145,
    n1110,
    n1123,
    n954
  );


  and
  g1531
  (
    n1401,
    n1077,
    n1055,
    n1244,
    n973
  );


  nor
  g1532
  (
    n1371,
    n928,
    n1159,
    n1152,
    n1207
  );


  nand
  g1533
  (
    n1370,
    n1126,
    n988,
    n1224,
    n1233
  );


  and
  g1534
  (
    n1350,
    n1172,
    n1221,
    n1021,
    n1019
  );


  and
  g1535
  (
    n1435,
    n1003,
    n1107,
    n1237,
    n1055
  );


  nor
  g1536
  (
    n1597,
    n950,
    n1152,
    n1186,
    n1115
  );


  xor
  g1537
  (
    n1362,
    n1204,
    n1084,
    n1230,
    n1217
  );


  and
  g1538
  (
    n1565,
    n1214,
    n1101,
    n945,
    n1162
  );


  xnor
  g1539
  (
    n1512,
    n1245,
    n1080,
    n1192,
    n1015
  );


  or
  g1540
  (
    KeyWire_0_47,
    n1107,
    n1240,
    n929,
    n1083
  );


  nor
  g1541
  (
    n1513,
    n1029,
    n1161,
    n963,
    n979
  );


  and
  g1542
  (
    n1366,
    n1011,
    n1028,
    n998,
    n1110
  );


  nor
  g1543
  (
    n1373,
    n1118,
    n1019,
    n812,
    n1071
  );


  xnor
  g1544
  (
    n1409,
    n969,
    n964,
    n990,
    n949
  );


  xnor
  g1545
  (
    n1594,
    n1068,
    n940,
    n1111,
    n946
  );


  or
  g1546
  (
    n1500,
    n1057,
    n1160,
    n995,
    n964
  );


  nor
  g1547
  (
    n1443,
    n1056,
    n1183,
    n1119,
    n1191
  );


  nor
  g1548
  (
    n1592,
    n1103,
    n1064,
    n1202,
    n1219
  );


  and
  g1549
  (
    n1485,
    n1092,
    n1015,
    n1063,
    n1130
  );


  xor
  g1550
  (
    n1340,
    n947,
    n1144,
    n1181,
    n967
  );


  xnor
  g1551
  (
    n1451,
    n1091,
    n1062,
    n1167,
    n1228
  );


  xnor
  g1552
  (
    n1619,
    n1237,
    n1096,
    n1200,
    n1175
  );


  and
  g1553
  (
    n1613,
    n1129,
    n1130,
    n1099,
    n1098
  );


  or
  g1554
  (
    n1559,
    n1095,
    n985,
    n1220,
    n1041
  );


  or
  g1555
  (
    n1498,
    n1104,
    n1216,
    n1048,
    n936
  );


  nand
  g1556
  (
    n1494,
    n1138,
    n1242,
    n1016,
    n1153
  );


  nand
  g1557
  (
    n1372,
    n1179,
    n932,
    n1227,
    n1174
  );


  and
  g1558
  (
    n1295,
    n1049,
    n1012,
    n979,
    n997
  );


  xnor
  g1559
  (
    n1326,
    n1145,
    n1082,
    n1110,
    n1235
  );


  xnor
  g1560
  (
    n1413,
    n1114,
    n1076,
    n989,
    n1153
  );


  nor
  g1561
  (
    n1342,
    n937,
    n1103,
    n1192,
    n1064
  );


  xor
  g1562
  (
    n1278,
    n1125,
    n1149,
    n1237,
    n1170
  );


  xor
  g1563
  (
    n1599,
    n1126,
    n1202,
    n1022,
    n1102
  );


  xor
  g1564
  (
    n1272,
    n1118,
    n965,
    n1008,
    n1112
  );


  or
  g1565
  (
    n1320,
    n1196,
    n1187,
    n1050,
    n944
  );


  xnor
  g1566
  (
    n1386,
    n1126,
    n1055,
    n939,
    n1213
  );


  xnor
  g1567
  (
    n1475,
    n1049,
    n1038,
    n1232,
    n1174
  );


  nand
  g1568
  (
    n1556,
    n1215,
    n1217,
    n1185,
    n966
  );


  xor
  g1569
  (
    n1554,
    n1107,
    n994,
    n1040,
    n951
  );


  xor
  g1570
  (
    n1526,
    n1109,
    n938,
    n814,
    n1221
  );


  and
  g1571
  (
    n1346,
    n1240,
    n1183,
    n1058,
    n1184
  );


  xor
  g1572
  (
    n1275,
    n1157,
    n1095,
    n1127,
    n1048
  );


  or
  g1573
  (
    n1339,
    n992,
    n1052,
    n1006,
    n1093
  );


  xor
  g1574
  (
    n1572,
    n1176,
    n1091,
    n1018,
    n1071
  );


  xnor
  g1575
  (
    n1484,
    n1180,
    n1197,
    n1078,
    n1047
  );


  xnor
  g1576
  (
    n1570,
    n1222,
    n956,
    n1147,
    n1063
  );


  xnor
  g1577
  (
    n1387,
    n1213,
    n1084,
    n1055,
    n1226
  );


  xnor
  g1578
  (
    n1252,
    n961,
    n1133,
    n1235,
    n927
  );


  xor
  g1579
  (
    n1607,
    n1021,
    n1026,
    n1083,
    n1243
  );


  and
  g1580
  (
    n1501,
    n988,
    n1229,
    n1081,
    n1115
  );


  or
  g1581
  (
    n1315,
    n1212,
    n1123,
    n927,
    n1001
  );


  xnor
  g1582
  (
    n1595,
    n1193,
    n1216,
    n1214,
    n1134
  );


  xnor
  g1583
  (
    n1522,
    n1150,
    n968,
    n989,
    n978
  );


  nor
  g1584
  (
    n1605,
    n987,
    n1228,
    n1205,
    n1234
  );


  nand
  g1585
  (
    n1280,
    n1223,
    n1146,
    n1099,
    n1155
  );


  nand
  g1586
  (
    n1271,
    n1169,
    n1090,
    n1173,
    n1145
  );


  xor
  g1587
  (
    n1404,
    n1095,
    n797,
    n1189,
    n991
  );


  xor
  g1588
  (
    n1579,
    n1044,
    n1170,
    n1057,
    n1131
  );


  nand
  g1589
  (
    n1264,
    n1161,
    n1205,
    n929,
    n1234
  );


  nand
  g1590
  (
    n1378,
    n972,
    n1061,
    n1068,
    n1096
  );


  or
  g1591
  (
    n1611,
    n1052,
    n1036,
    n969,
    n942
  );


  nand
  g1592
  (
    n1571,
    n1113,
    n974,
    n1166,
    n1156
  );


  nand
  g1593
  (
    n1517,
    n1093,
    n1068,
    n1033,
    n942
  );


  nand
  g1594
  (
    n1322,
    n930,
    n1008,
    n1165,
    n1139
  );


  or
  g1595
  (
    n1536,
    n1136,
    n1153,
    n799,
    n1174
  );


  xnor
  g1596
  (
    n1521,
    n1072,
    n1144,
    n1097,
    n995
  );


  xnor
  g1597
  (
    n1284,
    n1001,
    n940,
    n1045,
    n984
  );


  or
  g1598
  (
    n1479,
    n1090,
    n1218,
    n996,
    n1160
  );


  nand
  g1599
  (
    n1447,
    n951,
    n1082,
    n1157,
    n1030
  );


  nor
  g1600
  (
    n1488,
    n1207,
    n1181,
    n1185,
    n1195
  );


  and
  g1601
  (
    n1296,
    n1147,
    n1224,
    n1046,
    n1082
  );


  xor
  g1602
  (
    n1384,
    n926,
    n1061,
    n1012,
    n1239
  );


  xnor
  g1603
  (
    n1358,
    n1236,
    n1104,
    n1127,
    n1067
  );


  xor
  g1604
  (
    n1481,
    n1180,
    n1120,
    n1027,
    n961
  );


  and
  g1605
  (
    n1569,
    n1093,
    n1028,
    n1098,
    n1231
  );


  xor
  g1606
  (
    n1391,
    n980,
    n1009,
    n812,
    n960
  );


  nor
  g1607
  (
    n1600,
    n992,
    n1079,
    n1193,
    n1164
  );


  and
  g1608
  (
    n1697,
    n1618,
    n1256,
    n1444,
    n1246
  );


  nand
  g1609
  (
    n1641,
    n1250,
    n1291,
    n1577,
    n1488
  );


  nor
  g1610
  (
    n1706,
    n1484,
    n1481,
    n1616,
    n1525
  );


  nor
  g1611
  (
    n1717,
    n1528,
    n1380,
    n1561,
    n1409
  );


  or
  g1612
  (
    n1655,
    n1415,
    n1248,
    n1324,
    n1391
  );


  nor
  g1613
  (
    KeyWire_0_31,
    n1563,
    n1257,
    n1464,
    n1449
  );


  nand
  g1614
  (
    n1700,
    n1424,
    n1573,
    n1412,
    n1593
  );


  xor
  g1615
  (
    n1710,
    n1318,
    n1556,
    n1378,
    n1604
  );


  xnor
  g1616
  (
    n1720,
    n1457,
    n1429,
    n1471,
    n1352
  );


  and
  g1617
  (
    n1685,
    n1569,
    n1520,
    n1564,
    n1443
  );


  nand
  g1618
  (
    n1681,
    n1326,
    n1451,
    n1452,
    n1552
  );


  nand
  g1619
  (
    n1644,
    n1411,
    n1548,
    n1508,
    n1494
  );


  or
  g1620
  (
    n1696,
    n1358,
    n1251,
    n1592,
    n1435
  );


  xor
  g1621
  (
    KeyWire_0_30,
    n1428,
    n1566,
    n1472,
    n1296
  );


  and
  g1622
  (
    n1659,
    n1364,
    n1538,
    n1606,
    n1350
  );


  or
  g1623
  (
    n1633,
    n1375,
    n1276,
    n1254,
    n1419
  );


  and
  g1624
  (
    n1638,
    n1377,
    n1547,
    n1260,
    n1614
  );


  nor
  g1625
  (
    n1677,
    n1440,
    n1626,
    n1591,
    n1293
  );


  xnor
  g1626
  (
    n1647,
    n1524,
    n1615,
    n1413,
    n1550
  );


  and
  g1627
  (
    n1675,
    n1423,
    n1517,
    n1587,
    n1497
  );


  nand
  g1628
  (
    n1645,
    n1322,
    n1342,
    n1455,
    n1258
  );


  xnor
  g1629
  (
    KeyWire_0_55,
    n1295,
    n1536,
    n1405,
    n1625
  );


  xnor
  g1630
  (
    n1684,
    n1321,
    n1347,
    n1427,
    n1337
  );


  nand
  g1631
  (
    n1669,
    n1344,
    n1479,
    n1594,
    n1283
  );


  xor
  g1632
  (
    n1713,
    n1530,
    n1568,
    n1394,
    n1316
  );


  xor
  g1633
  (
    n1672,
    n1459,
    n1314,
    n1466,
    n1359
  );


  or
  g1634
  (
    n1693,
    n1274,
    n1447,
    n1626,
    n1448
  );


  or
  g1635
  (
    n1686,
    n1289,
    n1417,
    n1619,
    n1330
  );


  nor
  g1636
  (
    n1646,
    n1507,
    n1581,
    n1487,
    n1589
  );


  xnor
  g1637
  (
    n1694,
    n1303,
    n1298,
    n1384,
    n1288
  );


  and
  g1638
  (
    n1702,
    n1306,
    n1601,
    n1625,
    n1403
  );


  xor
  g1639
  (
    n1719,
    n1374,
    n1308,
    n1387,
    n1467
  );


  xnor
  g1640
  (
    n1716,
    n1402,
    n1502,
    n1586,
    n1348
  );


  and
  g1641
  (
    n1636,
    n1571,
    n1431,
    n1259,
    n1621
  );


  and
  g1642
  (
    n1656,
    n1372,
    n1310,
    n1263,
    n1247
  );


  nor
  g1643
  (
    n1652,
    n1277,
    n1559,
    n1255,
    n1468
  );


  or
  g1644
  (
    n1648,
    n1500,
    n1408,
    n1425,
    n1505
  );


  nand
  g1645
  (
    n1709,
    n1271,
    n1332,
    n1560,
    n1323
  );


  xor
  g1646
  (
    n1704,
    n1265,
    n1478,
    n1301,
    n1551
  );


  xnor
  g1647
  (
    n1721,
    n1325,
    n1532,
    n1341,
    n1462
  );


  and
  g1648
  (
    n1707,
    n1445,
    n1386,
    n1404,
    n1623
  );


  or
  g1649
  (
    n1663,
    n1420,
    n1537,
    n1516,
    n1362
  );


  nand
  g1650
  (
    n1695,
    n1454,
    n1521,
    n1609,
    n1590
  );


  and
  g1651
  (
    n1722,
    n1543,
    n1588,
    n1510,
    n1300
  );


  and
  g1652
  (
    n1654,
    n1328,
    n1514,
    n1284,
    n1311
  );


  nor
  g1653
  (
    n1631,
    n1434,
    n1458,
    n1275,
    n1607
  );


  nor
  g1654
  (
    n1689,
    n1582,
    n1489,
    n1441,
    n1357
  );


  xor
  g1655
  (
    n1691,
    n1622,
    n1385,
    n1473,
    n1290
  );


  nand
  g1656
  (
    n1634,
    n1426,
    n1361,
    n1414,
    n1585
  );


  or
  g1657
  (
    n1674,
    n1562,
    n1309,
    n1605,
    n1483
  );


  or
  g1658
  (
    n1653,
    n1546,
    n1558,
    n1612,
    n1529
  );


  xor
  g1659
  (
    n1643,
    n1365,
    n1437,
    n1453,
    n1280
  );


  nand
  g1660
  (
    n1651,
    n1430,
    n1482,
    n1476,
    n1511
  );


  nand
  g1661
  (
    n1701,
    n1596,
    n1268,
    n1613,
    n1401
  );


  and
  g1662
  (
    n1637,
    n1307,
    n1381,
    n1282,
    n1266
  );


  nor
  g1663
  (
    n1688,
    n1576,
    n1533,
    n1349,
    n1599
  );


  and
  g1664
  (
    n1649,
    n1299,
    n1304,
    n1345,
    n1356
  );


  and
  g1665
  (
    n1666,
    n1475,
    n1392,
    n1565,
    n1287
  );


  or
  g1666
  (
    n1714,
    n1580,
    n1395,
    n1253,
    n1540
  );


  nand
  g1667
  (
    n1635,
    n1315,
    n1351,
    n1495,
    n1353
  );


  xor
  g1668
  (
    n1630,
    n1509,
    n1432,
    n1264,
    n1603
  );


  xor
  g1669
  (
    n1665,
    n1579,
    n1598,
    n1393,
    n1512
  );


  or
  g1670
  (
    n1715,
    n1442,
    n1397,
    n1269,
    n1570
  );


  or
  g1671
  (
    n1682,
    n1519,
    n1279,
    n1285,
    n1327
  );


  xor
  g1672
  (
    n1660,
    n1480,
    n1331,
    n1486,
    n1410
  );


  xnor
  g1673
  (
    n1673,
    n1595,
    n1366,
    n1273,
    n1583
  );


  xnor
  g1674
  (
    n1692,
    n1608,
    n1346,
    n1336,
    n1544
  );


  xnor
  g1675
  (
    n1632,
    n1504,
    n1343,
    n1574,
    n1281
  );


  xor
  g1676
  (
    n1703,
    n1624,
    n1422,
    n1382,
    n1553
  );


  nor
  g1677
  (
    n1627,
    n1438,
    n1389,
    n1557,
    n1278
  );


  or
  g1678
  (
    n1679,
    n1535,
    n1355,
    n1534,
    n90
  );


  xnor
  g1679
  (
    n1657,
    n1496,
    n1567,
    n1400,
    n1398
  );


  xnor
  g1680
  (
    n1671,
    n1294,
    n1379,
    n1485,
    n1305
  );


  xor
  g1681
  (
    n1680,
    n1433,
    n1249,
    n1418,
    n1491
  );


  xor
  g1682
  (
    n1699,
    n1446,
    n1542,
    n1383,
    n1545
  );


  nand
  g1683
  (
    n1662,
    n1262,
    n1272,
    n1503,
    n1526
  );


  or
  g1684
  (
    n1642,
    n1261,
    n1320,
    n1317,
    n1368
  );


  nand
  g1685
  (
    n1629,
    n1554,
    n1388,
    n1539,
    n1312
  );


  and
  g1686
  (
    n1664,
    n1555,
    n1340,
    n1523,
    n1597
  );


  nand
  g1687
  (
    n1640,
    n1406,
    n1572,
    n1286,
    n1363
  );


  xnor
  g1688
  (
    n1690,
    n1371,
    n1329,
    n1333,
    n1370
  );


  xor
  g1689
  (
    n1678,
    n1541,
    n1334,
    n1292,
    n1501
  );


  xnor
  g1690
  (
    n1687,
    n1584,
    n1513,
    n1270,
    n1367
  );


  or
  g1691
  (
    n1670,
    n1469,
    n1617,
    n1515,
    n1470
  );


  and
  g1692
  (
    n1705,
    n1575,
    n1602,
    n1267,
    n1461
  );


  nor
  g1693
  (
    n1711,
    n1436,
    n1506,
    n1252,
    n1578
  );


  nand
  g1694
  (
    n1683,
    n1610,
    n1474,
    n1450,
    n1302
  );


  and
  g1695
  (
    n1708,
    n1460,
    n1439,
    n1354,
    n1549
  );


  xor
  g1696
  (
    n1676,
    n1399,
    n1369,
    n1490,
    n1600
  );


  nor
  g1697
  (
    n1712,
    n1492,
    n1376,
    n1527,
    n1360
  );


  nor
  g1698
  (
    n1698,
    n1531,
    n1465,
    n1421,
    n1416
  );


  nor
  g1699
  (
    n1667,
    n1498,
    n1396,
    n1297,
    n1499
  );


  nand
  g1700
  (
    n1661,
    n1313,
    n1319,
    n1477,
    n1407
  );


  and
  g1701
  (
    n1668,
    n1620,
    n1463,
    n1373,
    n1518
  );


  and
  g1702
  (
    n1639,
    n1456,
    n1522,
    n1493,
    n1338
  );


  nand
  g1703
  (
    n1650,
    n1339,
    n1611,
    n1335,
    n1390
  );


  and
  g1704
  (
    n1742,
    n1640,
    n1702,
    n1685,
    n1720
  );


  and
  g1705
  (
    n1733,
    n1633,
    n1690,
    n1695,
    n1694
  );


  xnor
  g1706
  (
    n1737,
    n1644,
    n1708,
    n1660,
    n1657
  );


  or
  g1707
  (
    n1731,
    n1629,
    n1712,
    n1673,
    n1700
  );


  or
  g1708
  (
    n1739,
    n1682,
    n1704,
    n1698,
    n1709
  );


  nor
  g1709
  (
    n1725,
    n1666,
    n1675,
    n1665,
    n1689
  );


  and
  g1710
  (
    n1734,
    n1677,
    n1638,
    n1688,
    n1715
  );


  nand
  g1711
  (
    n1738,
    n1662,
    n1703,
    n1710,
    n1641
  );


  nand
  g1712
  (
    n1732,
    n1628,
    n1699,
    n1631,
    n1687
  );


  xnor
  g1713
  (
    n1729,
    n1645,
    n1655,
    n1692,
    n1671
  );


  nand
  g1714
  (
    n1726,
    n1707,
    n1691,
    n1701,
    n1643
  );


  nor
  g1715
  (
    n1723,
    n1718,
    n1683,
    n1668,
    n1648
  );


  xnor
  g1716
  (
    n1735,
    n1674,
    n1667,
    n1649,
    n1678
  );


  nand
  g1717
  (
    n1744,
    n1693,
    n1696,
    n1656,
    n1653
  );


  or
  g1718
  (
    n1736,
    n1679,
    n1652,
    n1713,
    n1705
  );


  and
  g1719
  (
    n1730,
    n1659,
    n1635,
    n1706,
    n1636
  );


  xor
  g1720
  (
    n1746,
    n1719,
    n1721,
    n1664,
    n1634
  );


  and
  g1721
  (
    n1745,
    n1663,
    n1646,
    n1716,
    n1632
  );


  nand
  g1722
  (
    n1740,
    n1654,
    n1637,
    n1630,
    n1651
  );


  xor
  g1723
  (
    n1741,
    n1680,
    n1714,
    n1684,
    n1642
  );


  xor
  g1724
  (
    n1743,
    n1669,
    n1681,
    n1650,
    n1647
  );


  and
  g1725
  (
    n1728,
    n1627,
    n1672,
    n1658,
    n1676
  );


  xnor
  g1726
  (
    n1727,
    n1639,
    n1711,
    n1722,
    n1717
  );


  and
  g1727
  (
    n1724,
    n1670,
    n1661,
    n1686,
    n1697
  );


  xor
  KeyGate_0_0
  (
    n1470,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1444,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1537,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n578,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1139,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n839,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n557,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n169,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n352,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1307,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n781,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n296,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n518,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1523,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n121,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n78,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n210,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1015,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n1408,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1525,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1482,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1270,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n547,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n1584,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n873,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n824,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n357,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n289,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n453,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1144,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1718,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1628,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n532,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n198,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n127,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n83,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1157,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n633,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n200,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n829,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n1429,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n481,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n760,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n1452,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n504,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n461,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n1428,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n1496,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n1474,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n1422,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n825,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n1215,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n1617,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1217,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n914,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n1658,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n650,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n1352,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n859,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n717,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n93,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n809,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n434,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n1231,
    KeyNOTWire_0_63
  );


endmodule

