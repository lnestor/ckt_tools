// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_923_296 written by SynthGen on 2021/05/24 19:48:31
module Stat_923_296( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19,
 n75, n35, n54, n22, n67, n21, n45, n87,
 n56, n52, n23, n29, n84, n92, n33, n487,
 n637, n635, n640, n634, n802, n799, n914, n940,
 n936, n939, n938, n942, n941, n937);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19;

output n75, n35, n54, n22, n67, n21, n45, n87,
 n56, n52, n23, n29, n84, n92, n33, n487,
 n637, n635, n640, n634, n802, n799, n914, n940,
 n936, n939, n938, n942, n941, n937;

wire n20, n24, n25, n26, n27, n28, n30, n31,
 n32, n34, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n46, n47, n48, n49, n50,
 n51, n53, n55, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n68, n69, n70,
 n71, n72, n73, n74, n76, n77, n78, n79,
 n80, n81, n82, n83, n85, n86, n88, n89,
 n90, n91, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n636, n638,
 n639, n641, n642, n643, n644, n645, n646, n647,
 n648, n649, n650, n651, n652, n653, n654, n655,
 n656, n657, n658, n659, n660, n661, n662, n663,
 n664, n665, n666, n667, n668, n669, n670, n671,
 n672, n673, n674, n675, n676, n677, n678, n679,
 n680, n681, n682, n683, n684, n685, n686, n687,
 n688, n689, n690, n691, n692, n693, n694, n695,
 n696, n697, n698, n699, n700, n701, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735,
 n736, n737, n738, n739, n740, n741, n742, n743,
 n744, n745, n746, n747, n748, n749, n750, n751,
 n752, n753, n754, n755, n756, n757, n758, n759,
 n760, n761, n762, n763, n764, n765, n766, n767,
 n768, n769, n770, n771, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n794, n795, n796, n797, n798, n800,
 n801, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935;

buf  g0 (n37, n6);
not  g1 (n57, n2);
not  g2 (n79, n18);
not  g3 (n26, n15);
not  g4 (n88, n16);
not  g5 (n49, n12);
buf  g6 (n74, n13);
not  g7 (n80, n6);
buf  g8 (n82, n10);
not  g9 (n70, n7);
not  g10 (n63, n1);
not  g11 (n62, n11);
not  g12 (n39, n19);
not  g13 (n87, n7);
buf  g14 (n34, n3);
not  g15 (n89, n19);
buf  g16 (n25, n14);
not  g17 (n23, n4);
buf  g18 (n29, n8);
buf  g19 (n85, n10);
not  g20 (n51, n15);
buf  g21 (n61, n13);
not  g22 (n94, n9);
not  g23 (n44, n19);
buf  g24 (n90, n10);
buf  g25 (n67, n15);
buf  g26 (n35, n13);
buf  g27 (n28, n17);
not  g28 (n45, n5);
not  g29 (n38, n9);
not  g30 (n43, n16);
not  g31 (n33, n7);
buf  g32 (n55, n4);
buf  g33 (n47, n18);
buf  g34 (n32, n4);
not  g35 (n66, n17);
buf  g36 (n22, n11);
buf  g37 (n54, n18);
not  g38 (n72, n17);
not  g39 (n50, n7);
buf  g40 (n59, n1);
buf  g41 (n24, n3);
not  g42 (n42, n1);
not  g43 (n91, n6);
not  g44 (n36, n3);
buf  g45 (n69, n12);
not  g46 (n68, n14);
not  g47 (n20, n10);
not  g48 (n71, n14);
not  g49 (n40, n8);
not  g50 (n46, n3);
not  g51 (n77, n16);
buf  g52 (n75, n14);
not  g53 (n53, n13);
not  g54 (n81, n9);
buf  g55 (n58, n16);
not  g56 (n30, n18);
not  g57 (n78, n1);
not  g58 (n27, n11);
buf  g59 (n56, n9);
buf  g60 (n48, n17);
buf  g61 (n60, n8);
not  g62 (n76, n6);
buf  g63 (n41, n12);
not  g64 (n95, n5);
not  g65 (n65, n2);
buf  g66 (n84, n2);
buf  g67 (n52, n11);
not  g68 (n86, n5);
buf  g69 (n92, n8);
not  g70 (n31, n2);
buf  g71 (n83, n4);
not  g72 (n64, n12);
buf  g73 (n21, n5);
not  g74 (n93, n15);
not  g75 (n73, n19);
buf  g76 (n161, n39);
buf  g77 (n280, n65);
not  g78 (n267, n36);
buf  g79 (n151, n26);
not  g80 (n154, n36);
buf  g81 (n218, n50);
not  g82 (n129, n69);
buf  g83 (n201, n39);
not  g84 (n254, n29);
not  g85 (n176, n63);
buf  g86 (n114, n35);
not  g87 (n204, n73);
not  g88 (n236, n27);
buf  g89 (n233, n36);
buf  g90 (n131, n43);
buf  g91 (n99, n71);
not  g92 (n196, n53);
buf  g93 (n211, n43);
not  g94 (n110, n71);
not  g95 (n147, n49);
not  g96 (n266, n53);
buf  g97 (n251, n46);
buf  g98 (n222, n57);
buf  g99 (n288, n41);
not  g100 (n127, n73);
not  g101 (n173, n46);
not  g102 (n213, n66);
not  g103 (n136, n53);
buf  g104 (n121, n42);
buf  g105 (n191, n32);
not  g106 (n225, n55);
buf  g107 (n111, n38);
not  g108 (n192, n29);
not  g109 (n115, n67);
not  g110 (n123, n44);
buf  g111 (n199, n27);
not  g112 (n168, n61);
not  g113 (n250, n56);
buf  g114 (n295, n39);
buf  g115 (n263, n52);
buf  g116 (n108, n49);
buf  g117 (n120, n30);
buf  g118 (n239, n56);
buf  g119 (n246, n52);
buf  g120 (n112, n33);
not  g121 (n142, n63);
not  g122 (n242, n52);
buf  g123 (n207, n31);
not  g124 (n149, n71);
not  g125 (n195, n23);
buf  g126 (n96, n26);
not  g127 (n128, n73);
not  g128 (n103, n58);
not  g129 (n274, n69);
buf  g130 (n157, n65);
not  g131 (n180, n30);
not  g132 (n182, n27);
not  g133 (n107, n35);
not  g134 (n156, n67);
buf  g135 (n163, n37);
not  g136 (n208, n68);
buf  g137 (n158, n29);
buf  g138 (n134, n28);
buf  g139 (n243, n41);
not  g140 (n257, n48);
not  g141 (n184, n23);
not  g142 (n241, n33);
buf  g143 (n290, n58);
buf  g144 (n109, n54);
buf  g145 (n200, n54);
buf  g146 (n279, n51);
buf  g147 (n193, n51);
buf  g148 (n183, n69);
buf  g149 (n268, n64);
buf  g150 (n130, n41);
not  g151 (n140, n53);
not  g152 (n169, n47);
buf  g153 (n231, n37);
buf  g154 (n247, n37);
buf  g155 (n138, n46);
buf  g156 (n178, n47);
not  g157 (n287, n27);
buf  g158 (n116, n50);
not  g159 (n126, n60);
buf  g160 (n118, n40);
not  g161 (n276, n60);
not  g162 (n152, n55);
not  g163 (n113, n44);
not  g164 (n235, n57);
buf  g165 (n162, n33);
not  g166 (n133, n48);
not  g167 (n296, n67);
buf  g168 (n175, n60);
not  g169 (n124, n37);
not  g170 (n212, n47);
not  g171 (n214, n65);
buf  g172 (n281, n66);
buf  g173 (n260, n68);
buf  g174 (n240, n72);
not  g175 (n277, n30);
buf  g176 (n269, n42);
buf  g177 (n203, n41);
buf  g178 (n285, n25);
not  g179 (n186, n55);
buf  g180 (n237, n48);
not  g181 (n283, n73);
buf  g182 (n153, n64);
buf  g183 (n232, n67);
not  g184 (n286, n46);
buf  g185 (n137, n68);
not  g186 (n119, n45);
buf  g187 (n171, n40);
buf  g188 (n261, n62);
buf  g189 (n229, n62);
buf  g190 (n262, n59);
buf  g191 (n284, n59);
not  g192 (n282, n64);
not  g193 (n275, n71);
buf  g194 (n234, n32);
not  g195 (n185, n44);
buf  g196 (n172, n25);
not  g197 (n294, n28);
buf  g198 (n139, n52);
buf  g199 (n228, n66);
not  g200 (n141, n48);
not  g201 (n219, n65);
buf  g202 (n259, n45);
buf  g203 (n217, n34);
not  g204 (n272, n58);
not  g205 (n170, n72);
buf  g206 (n244, n63);
not  g207 (n144, n20);
buf  g208 (n252, n57);
buf  g209 (n98, n69);
buf  g210 (n164, n24);
buf  g211 (n177, n51);
buf  g212 (n206, n38);
not  g213 (n155, n61);
buf  g214 (n205, n68);
not  g215 (n255, n47);
not  g216 (n224, n50);
buf  g217 (n181, n54);
buf  g218 (n264, n44);
buf  g219 (n245, n45);
buf  g220 (n291, n31);
not  g221 (n293, n72);
not  g222 (n197, n58);
not  g223 (n278, n32);
not  g224 (n146, n43);
buf  g225 (n117, n31);
buf  g226 (n189, n49);
buf  g227 (n179, n49);
buf  g228 (n227, n21);
buf  g229 (n194, n64);
buf  g230 (n249, n40);
buf  g231 (n150, n62);
not  g232 (n166, n61);
not  g233 (n265, n56);
not  g234 (n148, n60);
not  g235 (n105, n51);
not  g236 (n216, n42);
buf  g237 (n238, n24);
not  g238 (n188, n34);
buf  g239 (n165, n70);
not  g240 (n273, n32);
buf  g241 (n220, n70);
buf  g242 (n190, n21);
not  g243 (n292, n22);
buf  g244 (n256, n22);
buf  g245 (n270, n59);
buf  g246 (n160, n34);
buf  g247 (n106, n40);
not  g248 (n122, n56);
not  g249 (n215, n35);
buf  g250 (n253, n62);
not  g251 (n143, n31);
buf  g252 (n125, n63);
buf  g253 (n132, n38);
buf  g254 (n101, n28);
buf  g255 (n135, n29);
not  g256 (n187, n61);
not  g257 (n289, n66);
buf  g258 (n159, n70);
not  g259 (n221, n59);
not  g260 (n248, n43);
buf  g261 (n258, n30);
buf  g262 (n230, n34);
not  g263 (n104, n35);
not  g264 (n271, n28);
not  g265 (n97, n39);
not  g266 (n145, n36);
not  g267 (n209, n57);
not  g268 (n100, n50);
not  g269 (n223, n54);
not  g270 (n167, n42);
buf  g271 (n210, n33);
not  g272 (n202, n55);
not  g273 (n198, n45);
not  g274 (n226, n38);
buf  g275 (n174, n72);
not  g276 (n102, n70);
not  g277 (n361, n231);
buf  g278 (n511, n212);
not  g279 (n478, n138);
not  g280 (n335, n177);
not  g281 (n494, n182);
not  g282 (n540, n81);
not  g283 (n325, n75);
buf  g284 (n433, n83);
not  g285 (n422, n260);
buf  g286 (n405, n229);
not  g287 (n340, n195);
not  g288 (n376, n188);
not  g289 (n455, n240);
buf  g290 (n524, n263);
not  g291 (n472, n262);
buf  g292 (n582, n236);
not  g293 (n305, n112);
buf  g294 (n467, n223);
buf  g295 (n375, n190);
buf  g296 (n423, n187);
buf  g297 (n513, n143);
buf  g298 (n509, n88);
buf  g299 (n410, n279);
not  g300 (n548, n212);
buf  g301 (n407, n91);
not  g302 (n574, n224);
not  g303 (n382, n75);
buf  g304 (n420, n167);
buf  g305 (n475, n170);
buf  g306 (n299, n206);
not  g307 (n387, n255);
not  g308 (n326, n156);
not  g309 (n590, n273);
not  g310 (n490, n261);
buf  g311 (n435, n104);
not  g312 (n452, n152);
not  g313 (n303, n127);
buf  g314 (n512, n253);
not  g315 (n364, n91);
not  g316 (n487, n255);
buf  g317 (n576, n101);
buf  g318 (n496, n112);
buf  g319 (n370, n165);
not  g320 (n585, n141);
buf  g321 (n533, n93);
not  g322 (n308, n258);
buf  g323 (n543, n265);
buf  g324 (n411, n202);
buf  g325 (n324, n263);
not  g326 (n421, n85);
not  g327 (n371, n79);
buf  g328 (n347, n133);
buf  g329 (n507, n184);
not  g330 (n379, n203);
not  g331 (n330, n276);
not  g332 (n355, n254);
not  g333 (n301, n246);
buf  g334 (n541, n82);
buf  g335 (n357, n243);
buf  g336 (n395, n262);
buf  g337 (n484, n148);
not  g338 (n537, n80);
not  g339 (n454, n200);
buf  g340 (n529, n217);
not  g341 (n327, n276);
buf  g342 (n317, n187);
not  g343 (n456, n266);
buf  g344 (n432, n229);
not  g345 (n604, n74);
buf  g346 (n545, n140);
not  g347 (n337, n151);
not  g348 (n489, n117);
not  g349 (n481, n77);
not  g350 (n469, n124);
buf  g351 (n413, n204);
not  g352 (n431, n227);
buf  g353 (n560, n205);
buf  g354 (n448, n228);
not  g355 (n390, n269);
buf  g356 (n373, n253);
buf  g357 (n600, n251);
buf  g358 (n602, n114);
buf  g359 (n446, n209);
buf  g360 (n306, n160);
buf  g361 (n599, n84);
buf  g362 (n316, n193);
buf  g363 (n417, n81);
not  g364 (n346, n192);
not  g365 (n447, n189);
not  g366 (n596, n201);
not  g367 (n384, n275);
buf  g368 (n499, n145);
buf  g369 (n385, n224);
buf  g370 (n312, n267);
buf  g371 (n441, n218);
buf  g372 (n535, n204);
buf  g373 (n424, n162);
not  g374 (n597, n223);
not  g375 (n608, n138);
buf  g376 (n404, n266);
buf  g377 (n366, n85);
not  g378 (n434, n236);
buf  g379 (n505, n216);
not  g380 (n436, n213);
not  g381 (n307, n221);
buf  g382 (n315, n275);
not  g383 (n297, n105);
not  g384 (n348, n230);
not  g385 (n464, n269);
buf  g386 (n501, n226);
buf  g387 (n443, n82);
buf  g388 (n563, n240);
not  g389 (n402, n227);
not  g390 (n453, n189);
not  g391 (n523, n242);
not  g392 (n566, n111);
buf  g393 (n587, n221);
not  g394 (n372, n258);
buf  g395 (n525, n274);
not  g396 (n569, n78);
not  g397 (n396, n90);
buf  g398 (n442, n273);
buf  g399 (n439, n83);
not  g400 (n437, n75);
buf  g401 (n398, n204);
not  g402 (n592, n212);
not  g403 (n408, n252);
buf  g404 (n532, n109);
buf  g405 (n504, n131);
buf  g406 (n440, n78);
not  g407 (n580, n269);
buf  g408 (n471, n260);
buf  g409 (n333, n87);
buf  g410 (n581, n245);
not  g411 (n589, n209);
not  g412 (n332, n117);
buf  g413 (n329, n115);
buf  g414 (n611, n105);
buf  g415 (n538, n164);
not  g416 (n457, n231);
buf  g417 (n528, n246);
not  g418 (n601, n258);
not  g419 (n531, n177);
buf  g420 (n321, n172);
buf  g421 (n350, n136);
not  g422 (n362, n199);
buf  g423 (n320, n132);
not  g424 (n359, n153);
not  g425 (n502, n140);
buf  g426 (n377, n244);
not  g427 (n520, n241);
not  g428 (n342, n212);
not  g429 (n383, n211);
buf  g430 (n577, n268);
buf  g431 (n415, n88);
buf  g432 (n522, n205);
buf  g433 (n555, n198);
not  g434 (n483, n215);
not  g435 (n336, n270);
buf  g436 (n338, n86);
not  g437 (n527, n116);
not  g438 (n318, n209);
buf  g439 (n334, n77);
buf  g440 (n603, n153);
not  g441 (n341, n191);
buf  g442 (n412, n215);
buf  g443 (n607, n235);
buf  g444 (n488, n220);
not  g445 (n530, n179);
buf  g446 (n465, n123);
not  g447 (n418, n206);
buf  g448 (n473, n256);
not  g449 (n610, n224);
buf  g450 (n319, n147);
not  g451 (n508, n244);
not  g452 (n500, n249);
not  g453 (n598, n86);
not  g454 (n539, n206);
buf  g455 (n344, n195);
buf  g456 (n356, n108);
not  g457 (n367, n265);
buf  g458 (n427, n237);
not  g459 (n298, n166);
not  g460 (n451, n256);
not  g461 (n426, n275);
buf  g462 (n514, n259);
not  g463 (n479, n85);
not  g464 (n595, n130);
not  g465 (n491, n139);
not  g466 (n572, n169);
not  g467 (n605, n221);
buf  g468 (n503, n163);
buf  g469 (n445, n220);
buf  g470 (n510, n93);
not  g471 (n526, n133);
not  g472 (n459, n149);
buf  g473 (n518, n264);
not  g474 (n463, n277);
buf  g475 (n380, n277);
not  g476 (n461, n226);
not  g477 (n575, n251);
buf  g478 (n409, n136);
buf  g479 (n568, n264);
buf  g480 (n571, n239);
not  g481 (n609, n231);
buf  g482 (n552, n275);
not  g483 (n358, n222);
not  g484 (n517, n79);
nor  g485 (n567, n84, n134, n250, n223);
and  g486 (n542, n86, n164, n148, n183);
and  g487 (n558, n247, n90, n232, n122);
and  g488 (n345, n239, n80, n181, n193);
and  g489 (n393, n128, n202, n248, n246);
nor  g490 (n515, n255, n259, n192, n203);
and  g491 (n388, n257, n107, n269, n173);
nor  g492 (n492, n74, n197, n87, n178);
nand g493 (n425, n216, n194, n219, n218);
nor  g494 (n544, n205, n232, n235, n265);
xor  g495 (n462, n89, n274, n279, n187);
and  g496 (n328, n185, n225, n219, n227);
nand g497 (n343, n276, n178, n271, n198);
xnor g498 (n360, n220, n214, n215, n155);
xnor g499 (n365, n200, n225, n75, n238);
xor  g500 (n363, n268, n222, n99, n168);
xor  g501 (n394, n144, n217, n225, n243);
nor  g502 (n476, n227, n247, n226, n81);
xor  g503 (n564, n176, n274, n152, n100);
and  g504 (n458, n214, n77, n271, n121);
xor  g505 (n579, n278, n199, n229);
and  g506 (n416, n256, n234, n161, n150);
xor  g507 (n482, n194, n141, n244, n193);
nor  g508 (n583, n270, n266, n200, n163);
xnor g509 (n349, n254, n280, n113, n237);
nand g510 (n428, n250, n259, n268, n165);
xnor g511 (n309, n137, n93, n193, n249);
xor  g512 (n606, n208, n232, n268, n180);
and  g513 (n406, n252, n234, n98, n84);
xor  g514 (n438, n191, n276, n187, n109);
xnor g515 (n485, n86, n88, n127, n211);
nand g516 (n313, n126, n248, n233, n207);
nand g517 (n553, n201, n78, n216, n245);
nand g518 (n429, n201, n169, n188, n248);
xnor g519 (n497, n150, n90, n207, n215);
nor  g520 (n351, n198, n256, n210);
xor  g521 (n536, n239, n199, n196, n106);
and  g522 (n323, n262, n245, n257, n144);
or   g523 (n551, n97, n261, n175, n93);
and  g524 (n399, n242, n214, n240, n196);
nand g525 (n310, n273, n211, n79, n198);
xor  g526 (n403, n151, n263, n166, n106);
nand g527 (n554, n158, n242, n206, n222);
and  g528 (n466, n274, n244, n161, n210);
xor  g529 (n450, n88, n192, n80, n191);
xnor g530 (n419, n192, n254, n203, n189);
nand g531 (n392, n139, n252, n213, n271);
xor  g532 (n397, n247, n76, n214, n101);
xor  g533 (n588, n243, n156, n135, n186);
xor  g534 (n322, n181, n87, n107, n154);
xor  g535 (n547, n203, n119, n270, n84);
xor  g536 (n559, n226, n235, n257);
and  g537 (n546, n185, n111, n80, n222);
nand g538 (n352, n110, n128, n265, n79);
or   g539 (n369, n237, n242, n145, n238);
xnor g540 (n314, n182, n255, n186, n123);
or   g541 (n486, n134, n132, n247, n92);
nor  g542 (n444, n175, n102, n197, n146);
and  g543 (n381, n82, n218, n76, n202);
and  g544 (n353, n129, n125, n120, n238);
xor  g545 (n430, n202, n216, n232, n149);
or   g546 (n557, n208, n191, n159, n211);
or   g547 (n562, n267, n267, n179, n218);
xor  g548 (n449, n172, n262, n188, n104);
xnor g549 (n516, n121, n130, n190, n233);
xor  g550 (n460, n273, n233, n230, n83);
or   g551 (n561, n180, n157, n98, n260);
or   g552 (n391, n260, n219, n110, n251);
xnor g553 (n591, n190, n170, n85, n272);
xnor g554 (n506, n108, n115, n280, n174);
xor  g555 (n570, n238, n116, n125, n131);
nor  g556 (n386, n261, n249, n272, n99);
nand g557 (n556, n82, n261, n246, n213);
xnor g558 (n474, n173, n230, n228, n97);
xor  g559 (n401, n195, n168, n277, n91);
or   g560 (n498, n230, n76, n279, n201);
xor  g561 (n300, n167, n213, n81, n102);
nor  g562 (n477, n92, n89, n229, n278);
or   g563 (n468, n114, n135, n184, n272);
nor  g564 (n549, n236, n188, n267, n77);
and  g565 (n339, n118, n234, n159, n252);
xor  g566 (n374, n245, n217, n209, n143);
xor  g567 (n584, n155, n189, n118, n237);
nand g568 (n578, n196, n147, n280, n266);
xnor g569 (n519, n194, n278, n91, n190);
nor  g570 (n331, n90, n103, n83, n250);
and  g571 (n573, n142, n142, n76, n250);
xor  g572 (n304, n239, n241, n254, n89);
or   g573 (n470, n176, n122, n87, n270);
xnor g574 (n368, n183, n234, n220, n92);
nor  g575 (n400, n204, n74, n257, n263);
xnor g576 (n354, n233, n264, n208, n207);
nor  g577 (n414, n74, n171, n224, n196);
and  g578 (n593, n219, n113, n119, n280);
or   g579 (n534, n207, n146, n228, n120);
nor  g580 (n565, n137, n258, n249, n100);
and  g581 (n495, n228, n200, n174, n154);
or   g582 (n493, n194, n162, n89, n271);
and  g583 (n378, n92, n129, n243, n205);
nor  g584 (n302, n241, n231, n157, n197);
xor  g585 (n311, n278, n171, n277, n253);
xnor g586 (n550, n259, n210, n248, n225);
and  g587 (n594, n236, n158, n124, n160);
xor  g588 (n480, n217, n251, n195, n264);
nand g589 (n389, n253, n221, n223, n103);
or   g590 (n521, n272, n78, n208, n240);
nor  g591 (n586, n126, n279, n197, n241);
not  g592 (n619, n309);
not  g593 (n626, n301);
buf  g594 (n623, n304);
buf  g595 (n628, n323);
buf  g596 (n621, n310);
buf  g597 (n624, n319);
buf  g598 (n616, n316);
buf  g599 (n627, n298);
buf  g600 (n614, n321);
not  g601 (n625, n303);
buf  g602 (n613, n299);
buf  g603 (n633, n313);
not  g604 (n630, n314);
buf  g605 (n632, n308);
not  g606 (n618, n307);
buf  g607 (n615, n312);
buf  g608 (n617, n318);
not  g609 (n620, n311);
buf  g610 (n629, n300);
not  g611 (n612, n315);
nor  g612 (n631, n306, n325, n305, n324);
nand g613 (n622, n320, n317, n302, n322);
xnor g614 (n635, n625, n356, n331, n339);
xor  g615 (n647, n335, n336, n355, n328);
or   g616 (n636, n345, n326, n358, n334);
nor  g617 (n643, n338, n350, n341, n621);
nor  g618 (n641, n618, n615, n340, n333);
and  g619 (n646, n361, n366, n351, n332);
or   g620 (n638, n364, n349, n617, n363);
or   g621 (n644, n616, n352, n614, n330);
or   g622 (n642, n613, n622, n347, n362);
nand g623 (n637, n342, n348, n619, n343);
or   g624 (n634, n329, n357, n354, n359);
nand g625 (n640, n367, n353, n337, n365);
nand g626 (n645, n612, n346, n620, n344);
nor  g627 (n639, n624, n327, n360, n623);
and  g628 (n654, n284, n283, n377, n642);
nor  g629 (n651, n379, n370, n643, n281);
nand g630 (n657, n281, n641, n283, n376);
or   g631 (n649, n371, n284, n283, n378);
xnor g632 (n653, n646, n647, n282, n283);
xor  g633 (n656, n284, n281, n645, n373);
xor  g634 (n655, n285, n369, n640, n282);
and  g635 (n650, n282, n285, n281, n644);
xnor g636 (n648, n284, n638, n372, n282);
xnor g637 (n652, n368, n639, n374, n375);
not  g638 (n661, n388);
buf  g639 (n658, n387);
nand g640 (n659, n649, n384);
xnor g641 (n662, n392, n386, n648, n383);
nor  g642 (n664, n654, n385, n381, n653);
nand g643 (n660, n380, n391, n652, n651);
or   g644 (n663, n389, n390, n650, n382);
and  g645 (n665, n406, n660, n659, n428);
or   g646 (n669, n417, n410, n403, n421);
nand g647 (n679, n661, n409, n402, n659);
nor  g648 (n666, n423, n405, n401, n659);
or   g649 (n677, n437, n658, n418, n411);
xor  g650 (n672, n661, n424, n658, n434);
or   g651 (n671, n431, n432, n661, n659);
nor  g652 (n678, n397, n414, n420, n660);
or   g653 (n673, n419, n399, n661, n436);
xor  g654 (n667, n662, n430, n407, n433);
nor  g655 (n668, n413, n426, n394, n415);
or   g656 (n670, n412, n396, n398, n422);
xnor g657 (n676, n395, n660, n425, n393);
nand g658 (n674, n400, n660, n427, n435);
xor  g659 (n675, n404, n416, n429, n408);
xor  g660 (n689, n285, n664, n667);
nand g661 (n693, n679, n628, n655, n666);
and  g662 (n682, n678, n675, n676, n632);
xnor g663 (n681, n94, n288, n679, n626);
xor  g664 (n686, n286, n440, n663, n629);
nand g665 (n695, n673, n630, n672, n288);
nand g666 (n683, n657, n663, n627, n662);
or   g667 (n680, n289, n286, n438);
or   g668 (n684, n671, n287, n285, n442);
or   g669 (n694, n288, n289, n439);
nand g670 (n690, n286, n633, n631, n670);
xor  g671 (n688, n287, n663, n664, n443);
nand g672 (n685, n665, n674, n287, n662);
and  g673 (n691, n668, n287, n664, n669);
nand g674 (n687, n677, n656, n663, n94);
nand g675 (n692, n441, n289, n288, n662);
not  g676 (n698, n680);
buf  g677 (n718, n682);
not  g678 (n707, n682);
not  g679 (n699, n684);
not  g680 (n710, n685);
buf  g681 (n717, n685);
not  g682 (n716, n684);
not  g683 (n709, n684);
buf  g684 (n702, n686);
not  g685 (n711, n680);
not  g686 (n703, n682);
buf  g687 (n715, n686);
not  g688 (n700, n683);
buf  g689 (n704, n683);
buf  g690 (n712, n683);
not  g691 (n719, n684);
not  g692 (n706, n681);
buf  g693 (n701, n681);
buf  g694 (n705, n685);
buf  g695 (n708, n686);
buf  g696 (n713, n683);
not  g697 (n714, n682);
not  g698 (n697, n685);
buf  g699 (n696, n686);
buf  g700 (n725, n697);
buf  g701 (n727, n699);
not  g702 (n721, n698);
buf  g703 (n726, n696);
not  g704 (n728, n687);
not  g705 (n724, n700);
xor  g706 (n720, n699, n687);
nand g707 (n729, n449, n697, n687, n698);
nand g708 (n723, n447, n448, n696, n445);
xor  g709 (n722, n444, n446, n700, n687);
not  g710 (n730, n720);
xnor g711 (n732, n701, n451, n454);
and  g712 (n733, n721, n456, n450, n722);
xnor g713 (n731, n721, n453, n452, n455);
buf  g714 (n740, n731);
not  g715 (n736, n730);
not  g716 (n738, n688);
not  g717 (n735, n688);
not  g718 (n737, n732);
nand g719 (n739, n689, n730, n731);
and  g720 (n741, n732, n689, n731);
xor  g721 (n734, n731, n688, n689);
buf  g722 (n748, n741);
buf  g723 (n745, n739);
not  g724 (n743, n735);
buf  g725 (n747, n741);
buf  g726 (n750, n734);
buf  g727 (n746, n737);
buf  g728 (n749, n736);
buf  g729 (n744, n738);
nand g730 (n742, n732, n740);
nand g731 (n777, n745, n712, n727, n716);
or   g732 (n770, n742, n744, n458, n728);
or   g733 (n758, n706, n746, n724);
nand g734 (n785, n722, n723, n705, n725);
xor  g735 (n762, n729, n723, n702, n750);
nor  g736 (n764, n722, n710, n723, n749);
xnor g737 (n759, n750, n750, n717, n713);
xnor g738 (n778, n728, n747, n290, n702);
xnor g739 (n771, n291, n709, n743, n742);
or   g740 (n767, n711, n711, n746, n712);
xor  g741 (n765, n729, n716, n709, n727);
or   g742 (n780, n457, n462, n722, n290);
or   g743 (n784, n744, n715, n714, n725);
xnor g744 (n761, n742, n744, n711, n723);
xnor g745 (n753, n465, n466, n748, n706);
xor  g746 (n782, n713, n708, n710, n742);
or   g747 (n786, n709, n705, n715);
and  g748 (n773, n726, n708, n707, n728);
nand g749 (n752, n710, n464, n714, n745);
nor  g750 (n781, n704, n290, n712, n743);
xnor g751 (n760, n746, n749, n291, n463);
xnor g752 (n783, n726, n748, n706, n747);
nand g753 (n776, n717, n744, n749, n707);
xor  g754 (n755, n714, n710, n290, n717);
and  g755 (n754, n291, n724, n715, n705);
nand g756 (n768, n727, n459, n743, n712);
xor  g757 (n769, n749, n708, n745, n746);
nand g758 (n766, n715, n726, n748, n724);
or   g759 (n763, n460, n725, n461, n709);
xor  g760 (n775, n727, n703, n748, n729);
xor  g761 (n757, n726, n716, n728, n713);
nand g762 (n774, n713, n706, n745, n708);
xor  g763 (n779, n750, n704, n711, n729);
xnor g764 (n772, n716, n747, n714, n703);
and  g765 (n751, n704, n743, n707, n701);
and  g766 (n756, n747, n707, n704, n725);
not  g767 (n789, n754);
not  g768 (n793, n753);
buf  g769 (n788, n754);
buf  g770 (n792, n752);
not  g771 (n795, n755);
buf  g772 (n790, n751);
buf  g773 (n791, n752);
buf  g774 (n794, n755);
not  g775 (n787, n753);
not  g776 (n796, n751);
xnor g777 (n798, n474, n475, n477, n467);
nand g778 (n800, n468, n760, n476, n759);
xnor g779 (n799, n471, n760, n787, n473);
nand g780 (n801, n469, n472, n758, n757);
nand g781 (n802, n787, n787, n788, n756);
and  g782 (n797, n756, n759, n758, n788);
nand g783 (n803, n757, n787, n470, n788);
nor  g784 (n808, n690, n691, n692);
xnor g785 (n805, n802, n690, n692, n691);
nor  g786 (n807, n788, n690, n799);
xor  g787 (n804, n693, n691, n789, n803);
xor  g788 (n806, n800, n801, n692);
nor  g789 (n816, n762, n783, n775, n808);
xnor g790 (n822, n804, n782, n779, n766);
xor  g791 (n812, n779, n806, n781, n763);
xnor g792 (n814, n783, n805, n807);
xnor g793 (n821, n806, n808, n769);
nand g794 (n826, n776, n774, n808, n806);
or   g795 (n818, n808, n807, n766, n782);
or   g796 (n823, n780, n765, n805, n778);
nor  g797 (n810, n807, n768, n780, n763);
nor  g798 (n811, n761, n768, n804, n771);
nand g799 (n824, n783, n770, n807, n775);
xnor g800 (n820, n764, n780, n762, n805);
and  g801 (n815, n783, n776, n774, n771);
or   g802 (n817, n806, n780, n772, n782);
or   g803 (n819, n773, n777, n764, n767);
xnor g804 (n813, n765, n778, n773, n777);
xnor g805 (n825, n761, n772, n782, n767);
xnor g806 (n809, n770, n781);
xor  g807 (n846, n816, n786, n823, n792);
nand g808 (n845, n789, n824, n794, n785);
nor  g809 (n835, n789, n732, n785, n811);
xnor g810 (n828, n794, n791, n795);
xor  g811 (n844, n790, n796, n821, n791);
or   g812 (n827, n478, n95, n795, n792);
nand g813 (n847, n824, n820, n826, n789);
and  g814 (n833, n796, n784, n794);
xnor g815 (n829, n718, n815, n793, n693);
xnor g816 (n841, n786, n793, n95, n826);
nor  g817 (n830, n814, n785, n813, n733);
nor  g818 (n838, n796, n479, n693, n784);
nor  g819 (n849, n786, n94, n822);
nor  g820 (n840, n733, n95, n693, n786);
nor  g821 (n839, n809, n822, n718, n792);
and  g822 (n850, n823, n821, n795, n733);
nand g823 (n832, n733, n718, n819, n694);
xnor g824 (n843, n717, n481, n718, n95);
and  g825 (n831, n485, n791, n793, n790);
or   g826 (n837, n794, n790, n817);
and  g827 (n848, n484, n825, n818, n784);
xor  g828 (n836, n812, n483, n810, n482);
and  g829 (n842, n719, n480, n793, n791);
nor  g830 (n834, n796, n792, n825, n785);
or   g831 (n865, n845, n519, n573, n539);
xor  g832 (n863, n526, n506, n491, n493);
or   g833 (n874, n546, n848, n495, n521);
or   g834 (n881, n499, n515, n568, n848);
and  g835 (n852, n842, n831, n516, n553);
xor  g836 (n867, n517, n846, n534, n505);
nor  g837 (n878, n508, n549, n528, n850);
xnor g838 (n851, n843, n532, n494, n844);
and  g839 (n873, n522, n838, n525, n575);
nor  g840 (n879, n832, n489, n510, n828);
nand g841 (n861, n847, n541, n574, n502);
xor  g842 (n876, n488, n529, n840, n846);
and  g843 (n869, n511, n538, n847, n556);
xor  g844 (n857, n837, n567, n514, n554);
xor  g845 (n859, n542, n512, n555, n503);
nand g846 (n854, n500, n490, n518, n536);
and  g847 (n858, n835, n487, n513, n560);
and  g848 (n868, n527, n545, n558, n486);
nor  g849 (n880, n830, n829, n850, n572);
nor  g850 (n855, n849, n523, n566, n497);
or   g851 (n862, n827, n533, n509, n559);
nor  g852 (n871, n548, n552, n520, n849);
nand g853 (n866, n577, n565, n547, n496);
nor  g854 (n877, n564, n498, n845, n841);
nand g855 (n856, n844, n543, n833, n569);
xnor g856 (n864, n836, n551, n507, n557);
xor  g857 (n860, n578, n540, n537, n501);
or   g858 (n853, n530, n561, n504, n563);
xor  g859 (n872, n492, n570, n535, n524);
nor  g860 (n870, n562, n576, n531, n544);
nor  g861 (n875, n839, n571, n834, n550);
buf  g862 (n885, n857);
not  g863 (n883, n856);
buf  g864 (n882, n858);
buf  g865 (n884, n855);
not  g866 (n890, n866);
not  g867 (n895, n883);
buf  g868 (n888, n861);
not  g869 (n886, n882);
xor  g870 (n893, n864, n579, n585, n884);
xor  g871 (n894, n883, n581, n862, n882);
and  g872 (n887, n586, n884, n583, n582);
xnor g873 (n891, n867, n580, n882, n863);
xnor g874 (n889, n865, n860, n584, n882);
and  g875 (n892, n859, n883, n587);
xor  g876 (n908, n872, n888, n886, n876);
or   g877 (n911, n886, n889);
xor  g878 (n900, n890, n885, n879, n869);
xnor g879 (n898, n889, n878, n887, n293);
xor  g880 (n904, n295, n293, n888, n886);
and  g881 (n896, n292, n873, n876, n293);
nand g882 (n902, n873, n872, n291, n887);
xnor g883 (n897, n294, n296, n867, n884);
nor  g884 (n899, n889, n871, n294, n875);
nand g885 (n901, n294, n884, n878, n870);
and  g886 (n910, n875, n888, n871, n885);
nand g887 (n907, n295, n890, n885, n292);
or   g888 (n909, n885, n292, n296, n294);
nor  g889 (n912, n888, n295, n874, n877);
or   g890 (n905, n292, n887, n877);
nand g891 (n906, n293, n869, n296, n874);
nand g892 (n903, n868, n868, n870, n295);
not  g893 (n913, n896);
nor  g894 (n914, n880, n897, n879);
or   g895 (n915, n914, n881, n880);
nor  g896 (n917, n890, n915, n891);
xor  g897 (n916, n892, n893, n915);
or   g898 (n918, n892, n891);
nor  g899 (n919, n915, n892, n893, n890);
or   g900 (n925, n895, n903, n916, n917);
xnor g901 (n922, n591, n589, n919, n893);
xor  g902 (n930, n609, n917, n608, n916);
and  g903 (n928, n595, n895, n917, n893);
or   g904 (n923, n603, n909, n592, n602);
or   g905 (n927, n894, n901, n590, n604);
nand g906 (n934, n597, n904, n919, n900);
xnor g907 (n935, n912, n894, n593, n594);
xnor g908 (n924, n905, n898, n599, n600);
nand g909 (n932, n908, n899, n606, n919);
xnor g910 (n933, n918, n911, n588, n895);
nor  g911 (n931, n916, n902, n601, n919);
or   g912 (n929, n894, n907, n918, n906);
nand g913 (n920, n610, n598, n894, n916);
and  g914 (n926, n596, n605, n918, n895);
or   g915 (n921, n917, n910, n918, n607);
or   g916 (n938, n695, n924, n935, n931);
xnor g917 (n939, n920, n694, n927);
xor  g918 (n941, n611, n695, n921);
and  g919 (n936, n719, n932, n933, n695);
xor  g920 (n942, n928, n930, n926, n719);
and  g921 (n940, n925, n934, n923, n719);
nor  g922 (n937, n694, n929, n296, n922);
endmodule
