// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_679_1333 written by SynthGen on 2021/05/24 19:48:29
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_679_1333 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31,
 n558, n685, n682, n702, n695, n686, n692, n690,
 n701, n683, n699, n687, n696, n689, n688, n703,
 n680, n691, n697, n684, n700, n694, n698, n708,
 n710, n709, n707);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31;

output n558, n685, n682, n702, n695, n686, n692, n690,
 n701, n683, n699, n687, n696, n689, n688, n703,
 n680, n691, n697, n684, n700, n694, n698, n708,
 n710, n709, n707;

wire n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n402, n403, n404, n405, n406, n407,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n425, n426, n427, n428, n429, n430, n431,
 n432, n433, n434, n435, n436, n437, n438, n439,
 n440, n441, n442, n443, n444, n445, n446, n447,
 n448, n449, n450, n451, n452, n453, n454, n455,
 n456, n457, n458, n459, n460, n461, n462, n463,
 n464, n465, n466, n467, n468, n469, n470, n471,
 n472, n473, n474, n475, n476, n477, n478, n479,
 n480, n481, n482, n483, n484, n485, n486, n487,
 n488, n489, n490, n491, n492, n493, n494, n495,
 n496, n497, n498, n499, n500, n501, n502, n503,
 n504, n505, n506, n507, n508, n509, n510, n511,
 n512, n513, n514, n515, n516, n517, n518, n519,
 n520, n521, n522, n523, n524, n525, n526, n527,
 n528, n529, n530, n531, n532, n533, n534, n535,
 n536, n537, n538, n539, n540, n541, n542, n543,
 n544, n545, n546, n547, n548, n549, n550, n551,
 n552, n553, n554, n555, n556, n557, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n681,
 n693, n704, n705, n706;

not  g0 (n38, n4);
buf  g1 (n76, n15);
not  g2 (n65, n10);
not  g3 (n40, n7);
buf  g4 (n55, n11);
not  g5 (n32, n25);
buf  g6 (n48, n21);
not  g7 (n78, n13);
not  g8 (n46, n11);
not  g9 (n68, n19);
not  g10 (n62, n26);
not  g11 (n47, n26);
nor  g12 (n42, n8, n12, n5);
xor  g13 (n58, n26, n22, n2);
and  g14 (n67, n20, n19, n29);
nand g15 (n60, n4, n9, n18);
xnor g16 (n70, n28, n21, n16);
nand g17 (n33, n16, n6, n4);
or   g18 (n45, n2, n28, n29);
and  g19 (n41, n30, n5, n24);
xor  g20 (n35, n16, n26, n12);
nand g21 (n79, n27, n14, n24);
or   g22 (n72, n16, n6, n15);
nor  g23 (n57, n14, n17, n5);
xor  g24 (n73, n8, n1);
nand g25 (n75, n23, n17, n30);
nor  g26 (n74, n27, n13, n7);
nor  g27 (n56, n29, n2, n9);
nand g28 (n52, n21, n28, n2);
or   g29 (n36, n30, n22, n7);
and  g30 (n43, n25, n9, n6);
nor  g31 (n53, n3, n20, n23);
and  g32 (n77, n15, n20, n4);
or   g33 (n34, n7, n20, n25);
and  g34 (n50, n12, n1, n19);
or   g35 (n49, n23, n25, n18);
xnor g36 (n63, n10, n23, n8);
or   g37 (n39, n27, n10, n29);
nor  g38 (n59, n3, n27, n24);
xor  g39 (n51, n12, n11, n17);
or   g40 (n37, n10, n18, n22);
xnor g41 (n44, n28, n14);
xor  g42 (n69, n19, n21, n24);
xnor g43 (n66, n3, n9, n13);
and  g44 (n54, n22, n3, n1);
and  g45 (n71, n15, n8, n30);
xor  g46 (n61, n13, n18, n17);
nor  g47 (n64, n11, n5, n6);
not  g48 (n213, n72);
buf  g49 (n238, n46);
buf  g50 (n125, n39);
not  g51 (n138, n49);
not  g52 (n197, n56);
not  g53 (n90, n62);
buf  g54 (n177, n69);
buf  g55 (n102, n68);
not  g56 (n106, n61);
buf  g57 (n232, n64);
not  g58 (n104, n70);
not  g59 (n235, n60);
not  g60 (n131, n74);
not  g61 (n250, n64);
buf  g62 (n246, n45);
buf  g63 (n247, n71);
not  g64 (n216, n45);
not  g65 (n231, n47);
not  g66 (n249, n64);
not  g67 (n180, n69);
buf  g68 (n243, n58);
not  g69 (n118, n44);
not  g70 (n183, n68);
not  g71 (n127, n73);
buf  g72 (n209, n75);
not  g73 (n217, n67);
not  g74 (n142, n33);
not  g75 (n140, n75);
buf  g76 (n190, n33);
buf  g77 (n199, n51);
not  g78 (n129, n32);
buf  g79 (n103, n71);
not  g80 (n178, n38);
buf  g81 (n229, n40);
not  g82 (n83, n57);
not  g83 (n164, n63);
not  g84 (n248, n52);
buf  g85 (n113, n74);
not  g86 (n114, n42);
not  g87 (n214, n66);
buf  g88 (n207, n50);
not  g89 (n244, n54);
buf  g90 (n210, n39);
not  g91 (n84, n70);
not  g92 (n234, n53);
buf  g93 (n116, n60);
not  g94 (n161, n55);
not  g95 (n171, n44);
not  g96 (n175, n52);
not  g97 (n100, n53);
not  g98 (n219, n33);
buf  g99 (n148, n73);
buf  g100 (n174, n69);
not  g101 (n122, n37);
buf  g102 (n223, n70);
buf  g103 (n211, n72);
buf  g104 (n176, n59);
buf  g105 (n241, n45);
not  g106 (n156, n55);
not  g107 (n123, n44);
buf  g108 (n86, n56);
not  g109 (n158, n36);
not  g110 (n237, n35);
not  g111 (n124, n32);
buf  g112 (n81, n61);
buf  g113 (n94, n36);
not  g114 (n144, n65);
buf  g115 (n132, n34);
not  g116 (n182, n73);
buf  g117 (n133, n59);
not  g118 (n119, n74);
buf  g119 (n224, n73);
not  g120 (n80, n36);
not  g121 (n188, n56);
not  g122 (n126, n68);
not  g123 (n220, n46);
not  g124 (n87, n61);
buf  g125 (n189, n32);
not  g126 (n115, n53);
buf  g127 (n121, n42);
not  g128 (n193, n43);
not  g129 (n151, n45);
buf  g130 (n198, n37);
buf  g131 (n205, n39);
buf  g132 (n251, n72);
not  g133 (n149, n56);
not  g134 (n203, n66);
buf  g135 (n165, n58);
not  g136 (n169, n48);
not  g137 (n163, n54);
buf  g138 (n112, n67);
buf  g139 (n96, n52);
buf  g140 (n194, n33);
buf  g141 (n97, n52);
buf  g142 (n105, n42);
not  g143 (n173, n41);
not  g144 (n155, n50);
buf  g145 (n166, n46);
not  g146 (n110, n63);
buf  g147 (n141, n41);
buf  g148 (n82, n71);
buf  g149 (n245, n75);
buf  g150 (n191, n60);
buf  g151 (n212, n58);
not  g152 (n146, n39);
buf  g153 (n107, n68);
not  g154 (n252, n51);
not  g155 (n215, n54);
buf  g156 (n147, n35);
buf  g157 (n185, n70);
buf  g158 (n85, n54);
not  g159 (n88, n47);
buf  g160 (n150, n48);
not  g161 (n91, n44);
not  g162 (n172, n47);
buf  g163 (n240, n71);
not  g164 (n134, n61);
not  g165 (n93, n62);
buf  g166 (n204, n37);
buf  g167 (n227, n63);
buf  g168 (n195, n66);
not  g169 (n128, n69);
not  g170 (n208, n57);
buf  g171 (n228, n67);
buf  g172 (n130, n67);
not  g173 (n225, n49);
not  g174 (n157, n35);
not  g175 (n236, n49);
not  g176 (n184, n72);
not  g177 (n226, n42);
buf  g178 (n162, n34);
buf  g179 (n221, n50);
not  g180 (n201, n40);
buf  g181 (n145, n34);
buf  g182 (n239, n51);
not  g183 (n187, n34);
buf  g184 (n120, n49);
not  g185 (n222, n50);
not  g186 (n153, n55);
buf  g187 (n111, n37);
buf  g188 (n186, n38);
not  g189 (n95, n55);
buf  g190 (n143, n53);
not  g191 (n109, n43);
buf  g192 (n137, n74);
buf  g193 (n108, n32);
not  g194 (n192, n57);
buf  g195 (n99, n47);
buf  g196 (n101, n40);
not  g197 (n202, n65);
buf  g198 (n152, n59);
buf  g199 (n167, n58);
buf  g200 (n181, n48);
not  g201 (n230, n38);
buf  g202 (n200, n57);
buf  g203 (n159, n35);
buf  g204 (n168, n48);
not  g205 (n179, n41);
not  g206 (n233, n65);
not  g207 (n242, n60);
not  g208 (n92, n51);
buf  g209 (n89, n59);
buf  g210 (n218, n40);
buf  g211 (n160, n63);
not  g212 (n170, n66);
buf  g213 (n135, n62);
buf  g214 (n154, n64);
buf  g215 (n98, n41);
not  g216 (n139, n36);
buf  g217 (n196, n38);
not  g218 (n206, n46);
buf  g219 (n136, n43);
and  g220 (n117, n65, n62, n43);
xnor g221 (n351, n241, n176, n164, n123);
or   g222 (n415, n190, n249, n127, n138);
xor  g223 (n413, n228, n132, n121, n206);
xor  g224 (n389, n164, n133, n124, n215);
xor  g225 (n382, n174, n146, n138, n143);
nand g226 (n293, n119, n128, n195, n226);
and  g227 (n321, n179, n117, n83);
or   g228 (n358, n176, n131, n157, n216);
nand g229 (n277, n236, n104, n126, n230);
xor  g230 (n305, n226, n206, n159, n134);
and  g231 (n341, n207, n200, n85, n242);
and  g232 (n334, n167, n241, n80, n160);
or   g233 (n324, n247, n137, n88, n100);
and  g234 (n279, n171, n140, n167, n93);
nand g235 (n278, n162, n192, n232, n89);
nor  g236 (n295, n95, n240, n188, n123);
nor  g237 (n374, n184, n130, n170, n231);
xor  g238 (n397, n207, n150, n218, n232);
nand g239 (n355, n196, n117, n203, n207);
xnor g240 (n298, n108, n128, n102, n111);
nor  g241 (n276, n168, n205, n118, n210);
or   g242 (n263, n228, n210, n196, n89);
xnor g243 (n347, n103, n152, n241, n127);
xor  g244 (n253, n201, n213, n122, n217);
nand g245 (n272, n123, n198, n189, n208);
xnor g246 (n302, n160, n157, n194, n202);
or   g247 (n292, n225, n110, n195, n226);
and  g248 (n337, n178, n99, n81, n182);
nand g249 (n289, n156, n156, n113, n213);
or   g250 (n317, n98, n175, n112, n177);
nor  g251 (n310, n163, n187, n138, n133);
xnor g252 (n412, n99, n215, n237, n236);
nand g253 (n303, n225, n172, n210, n153);
xnor g254 (n268, n234, n186, n224, n110);
and  g255 (n286, n122, n113, n191, n141);
nor  g256 (n265, n110, n158, n85, n245);
or   g257 (n312, n218, n139, n220, n111);
or   g258 (n256, n129, n239, n188, n120);
and  g259 (n345, n246, n129, n110, n197);
xnor g260 (n364, n189, n101, n198, n197);
nand g261 (n308, n195, n130, n220, n112);
or   g262 (n274, n120, n149, n180, n109);
or   g263 (n313, n248, n212, n98, n115);
nand g264 (n326, n237, n94, n199, n80);
xor  g265 (n332, n165, n171, n151, n141);
nand g266 (n311, n230, n205, n185, n101);
and  g267 (n319, n150, n139, n243, n116);
and  g268 (n375, n162, n82, n191, n229);
and  g269 (n410, n143, n193, n106, n108);
nor  g270 (n281, n216, n164, n202, n244);
nand g271 (n376, n148, n214, n172, n160);
nor  g272 (n390, n140, n223, n203, n171);
xor  g273 (n336, n223, n137, n109, n173);
and  g274 (n359, n166, n98, n200, n94);
xor  g275 (n384, n166, n149, n108, n193);
and  g276 (n349, n152, n129, n204, n125);
xnor g277 (n366, n191, n243, n123, n234);
xor  g278 (n309, n214, n234, n182, n205);
xor  g279 (n370, n90, n232, n88, n142);
nand g280 (n378, n231, n179, n186, n152);
xnor g281 (n283, n151, n244, n178);
xnor g282 (n372, n105, n101, n194, n136);
xnor g283 (n264, n127, n202, n114, n136);
nand g284 (n421, n141, n183, n168, n178);
and  g285 (n342, n153, n91, n243, n204);
nor  g286 (n393, n209, n96, n188, n189);
nand g287 (n354, n134, n186, n175, n185);
or   g288 (n338, n199, n198, n219, n91);
xor  g289 (n325, n145, n246, n238, n222);
nand g290 (n282, n82, n242, n145, n184);
xor  g291 (n383, n144, n193, n149, n246);
xnor g292 (n315, n159, n107, n81, n239);
nor  g293 (n320, n161, n163, n135, n165);
nor  g294 (n363, n176, n164, n124, n144);
or   g295 (n368, n103, n119, n231, n221);
or   g296 (n299, n90, n182, n213, n94);
xnor g297 (n411, n99, n223, n209, n181);
xnor g298 (n409, n229, n124, n96, n122);
nor  g299 (n314, n157, n105, n120, n223);
xor  g300 (n357, n245, n102, n177, n109);
or   g301 (n333, n244, n102, n165, n181);
xor  g302 (n356, n211, n245, n187, n106);
xnor g303 (n304, n93, n249, n146, n237);
or   g304 (n377, n120, n86, n144, n84);
xnor g305 (n416, n118, n177, n95, n88);
xnor g306 (n371, n86, n170, n143, n216);
xor  g307 (n287, n224, n173, n227, n191);
and  g308 (n266, n200, n133, n196, n205);
xnor g309 (n296, n220, n127, n187, n224);
xnor g310 (n400, n105, n181, n211, n218);
nand g311 (n380, n96, n242, n121, n153);
xor  g312 (n300, n128, n154, n136, n217);
and  g313 (n254, n207, n101, n169, n183);
nor  g314 (n406, n239, n179, n85, n232);
xnor g315 (n395, n201, n142, n81, n104);
and  g316 (n362, n229, n199, n235, n186);
xnor g317 (n306, n175, n118, n103, n239);
xor  g318 (n353, n222, n224, n88, n162);
and  g319 (n316, n148, n235, n135, n189);
nor  g320 (n343, n242, n86, n166, n97);
nor  g321 (n290, n233, n230, n126, n94);
xnor g322 (n294, n154, n92, n201, n225);
or   g323 (n407, n150, n93, n161, n206);
or   g324 (n420, n165, n217, n184, n175);
nand g325 (n402, n99, n247, n111, n168);
nor  g326 (n346, n196, n184, n201, n107);
xor  g327 (n301, n135, n100, n220, n96);
and  g328 (n327, n193, n132, n157, n147);
nor  g329 (n331, n113, n154, n235, n203);
xor  g330 (n352, n248, n162, n187, n146);
nor  g331 (n271, n116, n236, n132, n90);
nand g332 (n369, n217, n109, n176, n200);
and  g333 (n350, n208, n158, n151, n190);
nand g334 (n261, n182, n142, n185, n174);
nor  g335 (n348, n219, n240, n163, n86);
xnor g336 (n405, n240, n134, n124, n212);
or   g337 (n259, n215, n235, n112, n161);
nor  g338 (n291, n82, n227, n84);
xor  g339 (n367, n169, n185, n156, n209);
nand g340 (n257, n208, n155, n154, n172);
xor  g341 (n269, n130, n117, n126, n161);
and  g342 (n323, n219, n195, n245, n214);
nor  g343 (n361, n233, n108, n181, n212);
xnor g344 (n392, n83, n247, n130, n90);
xor  g345 (n381, n198, n93, n118, n194);
nor  g346 (n340, n97, n80, n113, n199);
nand g347 (n388, n197, n114, n84, n210);
or   g348 (n270, n159, n148, n231, n153);
nor  g349 (n418, n179, n208, n160, n97);
xnor g350 (n297, n115, n228, n221, n173);
xor  g351 (n267, n131, n114, n222, n145);
nand g352 (n330, n140, n211, n237, n180);
xnor g353 (n260, n214, n219, n163, n202);
and  g354 (n262, n150, n194, n248, n206);
nand g355 (n335, n111, n117, n133, n143);
and  g356 (n404, n119, n89, n138, n249);
xor  g357 (n391, n114, n103, n87, n246);
xor  g358 (n344, n129, n166, n238, n213);
nor  g359 (n373, n243, n171, n183, n136);
xor  g360 (n280, n105, n159, n225, n215);
and  g361 (n275, n180, n142, n91, n141);
xor  g362 (n360, n107, n158, n152, n170);
nand g363 (n322, n89, n131, n132, n148);
nor  g364 (n403, n98, n221, n106, n147);
and  g365 (n284, n100, n149, n247, n236);
xnor g366 (n285, n172, n167, n174, n95);
nand g367 (n385, n158, n92, n234, n155);
or   g368 (n419, n229, n126, n183, n249);
or   g369 (n339, n155, n125, n222, n209);
and  g370 (n328, n107, n233, n240, n134);
xor  g371 (n394, n115, n146, n87, n137);
nor  g372 (n379, n156, n92, n167, n87);
nor  g373 (n288, n116, n115, n188, n233);
nor  g374 (n387, n100, n104, n112, n83);
nor  g375 (n365, n190, n122, n203, n211);
and  g376 (n399, n104, n151, n87, n244);
and  g377 (n255, n125, n197, n192, n147);
nor  g378 (n307, n106, n145, n228, n218);
xor  g379 (n258, n128, n230, n177, n204);
nand g380 (n318, n212, n80, n95, n135);
nor  g381 (n401, n155, n121, n125, n169);
nor  g382 (n273, n192, n85, n139, n131);
xnor g383 (n422, n241, n121, n248, n147);
xnor g384 (n398, n238, n204, n180, n174);
xnor g385 (n408, n226, n170, n81, n102);
and  g386 (n417, n238, n173, n139, n119);
nand g387 (n414, n137, n116, n92, n144);
or   g388 (n396, n82, n192, n97, n227);
xnor g389 (n386, n190, n84, n168, n216);
nand g390 (n329, n140, n91, n221, n169);
xnor g391 (n450, n372, n340, n403, n365);
xnor g392 (n469, n382, n398, n328, n368);
or   g393 (n433, n390, n354, n397, n336);
or   g394 (n451, n348, n388, n386, n383);
nand g395 (n431, n256, n280, n357, n306);
nand g396 (n472, n356, n379, n363, n375);
nand g397 (n525, n400, n366, n383, n392);
and  g398 (n442, n300, n371, n334, n384);
nor  g399 (n502, n391, n339, n368, n344);
xnor g400 (n437, n399, n290, n377, n403);
or   g401 (n486, n322, n278, n392, n377);
xor  g402 (n493, n341, n384, n382, n376);
or   g403 (n441, n310, n288, n343, n321);
xnor g404 (n464, n335, n289, n318, n344);
xor  g405 (n424, n382, n295, n394, n327);
xor  g406 (n489, n402, n350, n344, n286);
nand g407 (n466, n353, n330, n383, n357);
xnor g408 (n481, n323, n379, n341, n353);
xor  g409 (n468, n402, n374, n389, n322);
or   g410 (n427, n338, n391, n404);
xor  g411 (n523, n334, n397, n354, n339);
xor  g412 (n478, n347, n366, n291, n375);
or   g413 (n454, n335, n357, n340, n380);
and  g414 (n459, n370, n388, n390, n275);
or   g415 (n444, n379, n384, n325, n371);
nand g416 (n463, n284, n349, n260, n287);
and  g417 (n447, n346, n267, n338, n305);
nor  g418 (n471, n400, n276, n401, n398);
nand g419 (n518, n322, n407, n380, n346);
xnor g420 (n425, n327, n374, n352, n345);
nand g421 (n434, n331, n351, n268, n324);
and  g422 (n443, n353, n402, n320, n332);
nand g423 (n482, n271, n263, n316, n296);
xnor g424 (n500, n317, n342, n348, n253);
xnor g425 (n495, n405, n323, n369, n395);
and  g426 (n491, n330, n266, n361, n335);
xnor g427 (n497, n390, n324, n397, n358);
nor  g428 (n456, n361, n354, n321, n325);
and  g429 (n438, n337, n362, n405, n328);
and  g430 (n490, n356, n281, n338, n401);
nor  g431 (n423, n352, n395, n269, n313);
or   g432 (n499, n405, n394, n332, n307);
xor  g433 (n504, n370, n254, n406, n355);
nand g434 (n439, n374, n380, n343, n349);
xor  g435 (n496, n365, n385, n376, n262);
nor  g436 (n506, n344, n385, n326, n405);
xnor g437 (n453, n369, n282, n361, n332);
nor  g438 (n524, n283, n294, n377, n315);
nand g439 (n460, n329, n398, n400, n331);
xnor g440 (n465, n397, n360, n392, n375);
xnor g441 (n457, n390, n343, n342, n399);
xor  g442 (n484, n265, n351, n385, n373);
nor  g443 (n435, n309, n364, n371, n264);
xnor g444 (n473, n387, n387, n386, n355);
nand g445 (n516, n298, n347, n357, n273);
xnor g446 (n494, n393, n326, n272, n327);
xor  g447 (n477, n365, n391, n327, n406);
or   g448 (n507, n339, n362, n335, n261);
nor  g449 (n487, n329, n330, n370, n346);
xor  g450 (n461, n377, n347, n325, n359);
xor  g451 (n514, n338, n396, n333, n363);
and  g452 (n479, n369, n323, n328, n372);
and  g453 (n498, n367, n375, n311, n274);
nor  g454 (n470, n364, n381, n402, n337);
xnor g455 (n501, n404, n382, n349, n352);
or   g456 (n488, n391, n378, n342, n400);
xor  g457 (n474, n350, n355, n326, n376);
and  g458 (n476, n403, n347, n399, n333);
nand g459 (n426, n312, n388, n372, n356);
or   g460 (n448, n325, n350, n367, n393);
or   g461 (n458, n320, n308, n373, n359);
xnor g462 (n508, n345, n387, n336, n366);
and  g463 (n480, n323, n270, n329, n337);
nand g464 (n475, n367, n334, n340, n368);
or   g465 (n462, n398, n331, n401, n301);
xor  g466 (n429, n341, n304, n381, n374);
nor  g467 (n455, n399, n322, n376, n358);
and  g468 (n509, n319, n362, n359, n406);
xnor g469 (n520, n360, n363, n393, n326);
xnor g470 (n436, n277, n392, n360, n334);
nor  g471 (n519, n350, n383, n324, n320);
xnor g472 (n440, n314, n354, n346, n396);
nand g473 (n428, n388, n360, n303, n353);
or   g474 (n483, n330, n386, n385, n379);
xnor g475 (n446, n401, n339, n386, n395);
nand g476 (n526, n378, n369, n359, n329);
nor  g477 (n511, n258, n372, n321, n336);
or   g478 (n492, n404, n302, n358, n355);
xor  g479 (n452, n394, n371, n364, n341);
xor  g480 (n521, n363, n362, n259, n403);
nand g481 (n503, n387, n361, n293, n366);
nand g482 (n430, n396, n348, n255, n337);
and  g483 (n515, n320, n349, n340, n352);
or   g484 (n522, n384, n394, n333, n380);
nand g485 (n505, n285, n365, n378, n343);
nor  g486 (n517, n378, n292, n279, n389);
nor  g487 (n445, n351, n333, n336, n395);
or   g488 (n467, n328, n364, n356, n370);
xor  g489 (n512, n381, n348, n342, n324);
nor  g490 (n449, n368, n389, n332, n331);
or   g491 (n510, n406, n345, n358, n396);
nor  g492 (n432, n345, n381, n299, n321);
nand g493 (n513, n389, n373, n297);
xor  g494 (n485, n367, n351, n257, n393);
or   g495 (n543, n450, n480, n485, n448);
nand g496 (n591, n436, n505, n452, n473);
nand g497 (n571, n472, n456, n517, n501);
xnor g498 (n588, n489, n455, n519, n501);
nor  g499 (n595, n484, n491, n470, n429);
xor  g500 (n555, n512, n453, n509, n496);
or   g501 (n563, n468, n443, n508, n466);
xor  g502 (n557, n450, n448, n479, n452);
nand g503 (n602, n491, n458, n478, n474);
xor  g504 (n566, n493, n499, n455, n473);
nand g505 (n551, n445, n510, n447, n499);
or   g506 (n560, n501, n514, n513, n474);
xor  g507 (n553, n504, n433, n435, n424);
nor  g508 (n583, n519, n480, n454, n461);
nand g509 (n558, n491, n470, n502, n520);
nor  g510 (n584, n469, n456, n459, n443);
or   g511 (n586, n463, n516, n492, n460);
and  g512 (n592, n461, n465, n518, n504);
and  g513 (n550, n475, n484, n480);
or   g514 (n562, n432, n514, n520, n468);
or   g515 (n547, n449, n515, n479, n507);
nor  g516 (n594, n446, n466, n502, n496);
xnor g517 (n601, n450, n490, n445, n465);
or   g518 (n608, n494, n514, n475, n471);
or   g519 (n537, n513, n430, n499, n516);
xor  g520 (n536, n494, n466, n482, n472);
xnor g521 (n570, n485, n510, n471, n518);
and  g522 (n542, n489, n487, n479, n450);
nand g523 (n577, n518, n490, n482, n444);
or   g524 (n582, n507, n489, n447);
and  g525 (n548, n465, n467, n511, n472);
and  g526 (n531, n470, n483, n485, n454);
nor  g527 (n580, n462, n483, n497, n488);
nand g528 (n596, n506, n474, n477, n454);
nand g529 (n535, n427, n426, n481, n495);
or   g530 (n576, n506, n457, n464, n439);
or   g531 (n552, n503, n493, n457, n486);
xor  g532 (n567, n467, n453, n458);
and  g533 (n530, n520, n483, n470, n515);
and  g534 (n539, n519, n497, n458, n472);
or   g535 (n593, n479, n468, n464, n478);
or   g536 (n534, n499, n477, n512, n448);
xor  g537 (n574, n443, n511, n487, n505);
nor  g538 (n532, n494, n441, n498, n490);
or   g539 (n575, n497, n498, n452, n475);
and  g540 (n579, n437, n478, n503, n518);
nand g541 (n607, n463, n423, n442, n517);
or   g542 (n587, n477, n476, n434, n455);
xor  g543 (n581, n456, n496, n492, n469);
nor  g544 (n564, n500, n516, n515, n446);
and  g545 (n538, n463, n507, n447, n477);
nand g546 (n556, n494, n454, n481);
nor  g547 (n578, n497, n449, n460, n512);
xor  g548 (n559, n495, n511, n449);
nor  g549 (n554, n463, n495, n489, n488);
or   g550 (n569, n505, n443, n480, n428);
xnor g551 (n598, n506, n506, n516, n466);
and  g552 (n572, n487, n487, n453, n478);
and  g553 (n528, n459, n476, n491, n498);
and  g554 (n605, n493, n507, n440, n459);
and  g555 (n527, n519, n444, n474, n508);
nand g556 (n600, n455, n464, n510, n457);
nand g557 (n606, n509, n514, n445, n503);
xor  g558 (n540, n500, n473, n503, n460);
nor  g559 (n590, n446, n490, n486, n475);
nor  g560 (n565, n502, n451, n517, n473);
and  g561 (n568, n465, n471, n452, n485);
xor  g562 (n597, n492, n512, n484, n445);
xor  g563 (n585, n500, n467, n513, n493);
nor  g564 (n561, n476, n464, n471, n504);
nor  g565 (n589, n446, n482, n456);
and  g566 (n549, n520, n444, n462, n451);
and  g567 (n533, n517, n510, n448, n476);
xor  g568 (n604, n508, n461, n449, n498);
xor  g569 (n573, n469, n500, n457, n467);
xor  g570 (n603, n515, n488, n501, n459);
xor  g571 (n541, n508, n488, n481, n468);
or   g572 (n609, n453, n469, n513, n504);
nand g573 (n529, n509, n451, n431, n461);
xor  g574 (n544, n495, n462, n444, n492);
nor  g575 (n546, n483, n496, n425, n486);
and  g576 (n599, n509, n502, n462, n451);
xor  g577 (n545, n486, n460, n505, n438);
xor  g578 (n611, n556, n536, n558);
and  g579 (n618, n528, n544, n537);
xor  g580 (n628, n593, n549, n533);
nand g581 (n624, n548, n571, n562);
or   g582 (n621, n586, n567, n577);
xnor g583 (n631, n547, n589, n574);
or   g584 (n627, n590, n582, n568);
nand g585 (n623, n569, n539, n565);
and  g586 (n616, n572, n588, n575);
nand g587 (n617, n591, n579, n543);
or   g588 (n620, n554, n583, n532);
nor  g589 (n614, n535, n578, n534);
xnor g590 (n619, n538, n545, n550);
or   g591 (n626, n531, n540, n559);
and  g592 (n613, n553, n552, n561);
nor  g593 (n630, n587, n592, n564);
xor  g594 (n610, n576, n581, n563);
nor  g595 (n622, n542, n580, n585);
xnor g596 (n629, n529, n570, n555);
nand g597 (n625, n546, n595, n541);
xor  g598 (n612, n530, n584, n557, n560);
xnor g599 (n615, n551, n594, n566, n573);
xor  g600 (n644, n407, n411, n618, n614);
nand g601 (n638, n623, n614, n411, n410);
nand g602 (n639, n414, n627, n620, n616);
nand g603 (n641, n413, n616, n624, n611);
xnor g604 (n636, n616, n626, n618, n624);
nand g605 (n646, n413, n617, n408, n407);
nand g606 (n634, n623, n621, n612);
nand g607 (n648, n612, n626, n628, n620);
or   g608 (n657, n612, n407, n611, n410);
xnor g609 (n635, n412, n619, n613, n620);
nand g610 (n650, n623, n625, n619, n626);
nand g611 (n637, n408, n409, n610, n615);
and  g612 (n647, n622, n621, n615, n627);
nand g613 (n643, n627, n622, n409, n624);
nor  g614 (n633, n621, n410, n414);
and  g615 (n651, n412, n409, n611, n411);
xor  g616 (n640, n408, n617, n613, n411);
xnor g617 (n645, n610, n613, n623, n614);
nor  g618 (n649, n614, n413, n619, n613);
or   g619 (n652, n409, n625, n610, n627);
xnor g620 (n632, n408, n622, n626, n612);
and  g621 (n656, n620, n622, n618, n414);
nor  g622 (n653, n624, n617, n615);
and  g623 (n654, n619, n412, n618, n414);
and  g624 (n655, n611, n625, n615, n616);
nand g625 (n642, n625, n610, n412, n413);
and  g626 (n670, n416, n522, n415, n419);
and  g627 (n665, n647, n657, n633, n521);
xnor g628 (n662, n416, n31, n250, n635);
and  g629 (n668, n636, n522, n521);
nand g630 (n658, n416, n523, n522);
nand g631 (n669, n634, n417, n415, n524);
nand g632 (n667, n645, n597, n415, n642);
and  g633 (n673, n640, n641, n650, n31);
nor  g634 (n660, n654, n648, n632, n418);
xnor g635 (n661, n644, n418, n250, n653);
nand g636 (n659, n655, n418, n416, n417);
or   g637 (n666, n637, n417, n523, n596);
or   g638 (n672, n521, n656, n31);
nor  g639 (n663, n415, n521, n651, n638);
nor  g640 (n664, n523, n649, n417, n643);
or   g641 (n671, n639, n652, n418, n646);
not  g642 (n674, n662);
buf  g643 (n677, n660);
buf  g644 (n678, n658);
not  g645 (n675, n663);
buf  g646 (n676, n659);
not  g647 (n679, n661);
xor  g648 (n680, n629, n252, n75, n251);
nand g649 (n691, n629, n600, n664, n631);
xnor g650 (n685, n674, n78, n250);
or   g651 (n696, n631, n676, n251, n421);
nor  g652 (n701, n599, n678, n670, n250);
nand g653 (n700, n525, n677, n629, n524);
xor  g654 (n681, n251, n77, n674, n79);
nor  g655 (n702, n421, n677, n679, n79);
and  g656 (n694, n252, n76, n631, n630);
and  g657 (n697, n628, n628, n630, n601);
xnor g658 (n689, n675, n525, n677, n77);
nand g659 (n684, n679, n630, n419, n598);
xnor g660 (n698, n419, n674, n676, n631);
nor  g661 (n687, n76, n420, n669, n679);
nand g662 (n693, n251, n674, n678, n79);
nand g663 (n695, n252, n524, n679, n678);
xnor g664 (n683, n676, n78, n76);
nor  g665 (n699, n79, n675, n676, n420);
or   g666 (n703, n602, n252, n419, n675);
or   g667 (n692, n76, n667, n668, n420);
nand g668 (n688, n420, n628, n77, n629);
xor  g669 (n686, n666, n77, n526, n677);
nand g670 (n682, n603, n525, n630, n665);
xnor g671 (n690, n675, n524, n525, n678);
nand g672 (n705, n703, n422);
or   g673 (n704, n422, n421, n702);
or   g674 (n706, n704, n705);
xnor g675 (n708, n526, n607, n608, n672);
nand g676 (n707, n609, n706, n605, n604);
xor  g677 (n710, n673, n706, n526, n606);
xnor g678 (n709, n671, n706, n526);
endmodule
