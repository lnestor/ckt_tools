

module Stat_1000_101
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n754,
  n964,
  n941,
  n992,
  n972,
  n958,
  n981,
  n973,
  n977,
  n987,
  n978,
  n980,
  n996,
  n942,
  n983,
  n985,
  n962,
  n947,
  n967,
  n1027,
  n1030,
  n1024,
  n1021,
  n1023,
  n1029,
  n1031,
  n1028,
  n1032,
  n1025,
  n1020,
  n1026,
  n1022
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n754;output n964;output n941;output n992;output n972;output n958;output n981;output n973;output n977;output n987;output n978;output n980;output n996;output n942;output n983;output n985;output n962;output n947;output n967;output n1027;output n1030;output n1024;output n1021;output n1023;output n1029;output n1031;output n1028;output n1032;output n1025;output n1020;output n1026;output n1022;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n943;wire n944;wire n945;wire n946;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n959;wire n960;wire n961;wire n963;wire n965;wire n966;wire n968;wire n969;wire n970;wire n971;wire n974;wire n975;wire n976;wire n979;wire n982;wire n984;wire n986;wire n988;wire n989;wire n990;wire n991;wire n993;wire n994;wire n995;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n117,
    n26
  );


  buf
  g1
  (
    n93,
    n27
  );


  not
  g2
  (
    n138,
    n29
  );


  not
  g3
  (
    n153,
    n11
  );


  not
  g4
  (
    n131,
    n29
  );


  buf
  g5
  (
    n75,
    n28
  );


  buf
  g6
  (
    n88,
    n21
  );


  not
  g7
  (
    n154,
    n19
  );


  buf
  g8
  (
    n127,
    n5
  );


  buf
  g9
  (
    n54,
    n21
  );


  buf
  g10
  (
    n87,
    n8
  );


  buf
  g11
  (
    n37,
    n30
  );


  buf
  g12
  (
    KeyWire_0_22,
    n27
  );


  buf
  g13
  (
    n136,
    n7
  );


  not
  g14
  (
    n125,
    n32
  );


  buf
  g15
  (
    n147,
    n21
  );


  not
  g16
  (
    n106,
    n23
  );


  not
  g17
  (
    KeyWire_0_3,
    n7
  );


  not
  g18
  (
    n134,
    n12
  );


  buf
  g19
  (
    n142,
    n31
  );


  buf
  g20
  (
    n148,
    n14
  );


  buf
  g21
  (
    n109,
    n9
  );


  not
  g22
  (
    n120,
    n29
  );


  not
  g23
  (
    n144,
    n23
  );


  buf
  g24
  (
    n76,
    n25
  );


  not
  g25
  (
    n99,
    n30
  );


  buf
  g26
  (
    KeyWire_0_10,
    n6
  );


  buf
  g27
  (
    n50,
    n25
  );


  not
  g28
  (
    n51,
    n17
  );


  not
  g29
  (
    n52,
    n26
  );


  buf
  g30
  (
    n133,
    n23
  );


  buf
  g31
  (
    n55,
    n10
  );


  buf
  g32
  (
    n95,
    n31
  );


  not
  g33
  (
    n152,
    n12
  );


  buf
  g34
  (
    n139,
    n24
  );


  buf
  g35
  (
    n126,
    n11
  );


  not
  g36
  (
    n141,
    n2
  );


  buf
  g37
  (
    n112,
    n4
  );


  buf
  g38
  (
    n128,
    n12
  );


  not
  g39
  (
    n90,
    n17
  );


  not
  g40
  (
    n62,
    n14
  );


  buf
  g41
  (
    n123,
    n24
  );


  buf
  g42
  (
    n145,
    n1
  );


  not
  g43
  (
    n130,
    n24
  );


  not
  g44
  (
    n39,
    n15
  );


  not
  g45
  (
    n105,
    n28
  );


  buf
  g46
  (
    n104,
    n11
  );


  buf
  g47
  (
    n149,
    n20
  );


  buf
  g48
  (
    n44,
    n16
  );


  buf
  g49
  (
    n40,
    n18
  );


  not
  g50
  (
    n96,
    n4
  );


  buf
  g51
  (
    n66,
    n3
  );


  buf
  g52
  (
    n57,
    n18
  );


  buf
  g53
  (
    n92,
    n16
  );


  not
  g54
  (
    n111,
    n20
  );


  not
  g55
  (
    n59,
    n9
  );


  buf
  g56
  (
    n42,
    n18
  );


  not
  g57
  (
    n83,
    n22
  );


  buf
  g58
  (
    n122,
    n4
  );


  not
  g59
  (
    n78,
    n3
  );


  not
  g60
  (
    n118,
    n24
  );


  buf
  g61
  (
    n121,
    n4
  );


  buf
  g62
  (
    n101,
    n8
  );


  buf
  g63
  (
    n102,
    n13
  );


  buf
  g64
  (
    n103,
    n10
  );


  not
  g65
  (
    n69,
    n7
  );


  buf
  g66
  (
    n34,
    n20
  );


  buf
  g67
  (
    n65,
    n14
  );


  buf
  g68
  (
    n71,
    n10
  );


  not
  g69
  (
    n61,
    n5
  );


  buf
  g70
  (
    n143,
    n11
  );


  not
  g71
  (
    n58,
    n3
  );


  not
  g72
  (
    n132,
    n13
  );


  buf
  g73
  (
    n47,
    n8
  );


  not
  g74
  (
    n98,
    n14
  );


  buf
  g75
  (
    n115,
    n25
  );


  not
  g76
  (
    n100,
    n15
  );


  buf
  g77
  (
    n107,
    n32
  );


  buf
  g78
  (
    n129,
    n6
  );


  not
  g79
  (
    n86,
    n3
  );


  not
  g80
  (
    n33,
    n30
  );


  not
  g81
  (
    n68,
    n15
  );


  buf
  g82
  (
    n36,
    n9
  );


  not
  g83
  (
    n91,
    n32
  );


  buf
  g84
  (
    n79,
    n31
  );


  buf
  g85
  (
    n84,
    n17
  );


  not
  g86
  (
    n81,
    n26
  );


  buf
  g87
  (
    n85,
    n26
  );


  not
  g88
  (
    n46,
    n29
  );


  buf
  g89
  (
    n74,
    n25
  );


  buf
  g90
  (
    n151,
    n31
  );


  buf
  g91
  (
    n135,
    n22
  );


  not
  g92
  (
    n137,
    n8
  );


  buf
  g93
  (
    n80,
    n28
  );


  not
  g94
  (
    n45,
    n16
  );


  not
  g95
  (
    n63,
    n19
  );


  buf
  g96
  (
    n110,
    n6
  );


  buf
  g97
  (
    n94,
    n7
  );


  buf
  g98
  (
    n150,
    n9
  );


  not
  g99
  (
    n67,
    n28
  );


  buf
  g100
  (
    n119,
    n19
  );


  not
  g101
  (
    n146,
    n12
  );


  not
  g102
  (
    n43,
    n20
  );


  buf
  g103
  (
    n124,
    n22
  );


  buf
  g104
  (
    n41,
    n5
  );


  not
  g105
  (
    n113,
    n22
  );


  not
  g106
  (
    n116,
    n2
  );


  buf
  g107
  (
    n97,
    n6
  );


  buf
  g108
  (
    n72,
    n23
  );


  buf
  g109
  (
    n108,
    n5
  );


  not
  g110
  (
    n70,
    n13
  );


  not
  g111
  (
    KeyWire_0_26,
    n27
  );


  buf
  g112
  (
    n89,
    n17
  );


  not
  g113
  (
    n48,
    n10
  );


  not
  g114
  (
    n114,
    n27
  );


  buf
  g115
  (
    n53,
    n19
  );


  buf
  g116
  (
    n82,
    n16
  );


  buf
  g117
  (
    n60,
    n21
  );


  buf
  g118
  (
    n56,
    n32
  );


  buf
  g119
  (
    n155,
    n13
  );


  not
  g120
  (
    n38,
    n18
  );


  buf
  g121
  (
    n49,
    n15
  );


  buf
  g122
  (
    n140,
    n30
  );


  not
  g123
  (
    n317,
    n138
  );


  buf
  g124
  (
    n364,
    n73
  );


  not
  g125
  (
    n312,
    n120
  );


  not
  g126
  (
    n282,
    n127
  );


  not
  g127
  (
    n380,
    n108
  );


  buf
  g128
  (
    n384,
    n104
  );


  buf
  g129
  (
    n227,
    n129
  );


  not
  g130
  (
    n291,
    n51
  );


  buf
  g131
  (
    n389,
    n133
  );


  not
  g132
  (
    n329,
    n52
  );


  buf
  g133
  (
    n328,
    n97
  );


  buf
  g134
  (
    n321,
    n131
  );


  buf
  g135
  (
    n315,
    n79
  );


  not
  g136
  (
    n357,
    n115
  );


  not
  g137
  (
    KeyWire_0_15,
    n60
  );


  buf
  g138
  (
    n375,
    n74
  );


  buf
  g139
  (
    n269,
    n66
  );


  not
  g140
  (
    n297,
    n128
  );


  buf
  g141
  (
    n214,
    n112
  );


  buf
  g142
  (
    n287,
    n143
  );


  buf
  g143
  (
    n366,
    n90
  );


  buf
  g144
  (
    n230,
    n52
  );


  not
  g145
  (
    n318,
    n117
  );


  not
  g146
  (
    n196,
    n40
  );


  not
  g147
  (
    n293,
    n127
  );


  buf
  g148
  (
    n217,
    n70
  );


  buf
  g149
  (
    n212,
    n111
  );


  not
  g150
  (
    n285,
    n63
  );


  not
  g151
  (
    n268,
    n145
  );


  buf
  g152
  (
    n181,
    n92
  );


  not
  g153
  (
    n204,
    n62
  );


  not
  g154
  (
    n347,
    n136
  );


  not
  g155
  (
    n337,
    n65
  );


  buf
  g156
  (
    n359,
    n140
  );


  not
  g157
  (
    n231,
    n103
  );


  buf
  g158
  (
    KeyWire_0_9,
    n80
  );


  buf
  g159
  (
    n259,
    n128
  );


  not
  g160
  (
    n166,
    n114
  );


  buf
  g161
  (
    n260,
    n114
  );


  not
  g162
  (
    n201,
    n119
  );


  buf
  g163
  (
    KeyWire_0_29,
    n85
  );


  buf
  g164
  (
    n284,
    n40
  );


  not
  g165
  (
    n341,
    n36
  );


  buf
  g166
  (
    n197,
    n76
  );


  buf
  g167
  (
    n275,
    n39
  );


  buf
  g168
  (
    n250,
    n125
  );


  not
  g169
  (
    n186,
    n57
  );


  not
  g170
  (
    n294,
    n119
  );


  buf
  g171
  (
    n261,
    n61
  );


  buf
  g172
  (
    n283,
    n51
  );


  buf
  g173
  (
    n270,
    n104
  );


  buf
  g174
  (
    n264,
    n47
  );


  not
  g175
  (
    n199,
    n60
  );


  not
  g176
  (
    n180,
    n99
  );


  not
  g177
  (
    n332,
    n132
  );


  not
  g178
  (
    n185,
    n116
  );


  not
  g179
  (
    n156,
    n143
  );


  not
  g180
  (
    n158,
    n87
  );


  not
  g181
  (
    n326,
    n50
  );


  not
  g182
  (
    n225,
    n76
  );


  not
  g183
  (
    n295,
    n48
  );


  buf
  g184
  (
    n289,
    n61
  );


  buf
  g185
  (
    n376,
    n138
  );


  not
  g186
  (
    n184,
    n76
  );


  buf
  g187
  (
    n393,
    n41
  );


  not
  g188
  (
    n216,
    n120
  );


  not
  g189
  (
    n363,
    n42
  );


  not
  g190
  (
    n333,
    n60
  );


  buf
  g191
  (
    n383,
    n93
  );


  buf
  g192
  (
    n267,
    n62
  );


  not
  g193
  (
    n345,
    n118
  );


  not
  g194
  (
    n313,
    n117
  );


  not
  g195
  (
    n162,
    n147
  );


  buf
  g196
  (
    n195,
    n41
  );


  not
  g197
  (
    n336,
    n135
  );


  buf
  g198
  (
    n170,
    n133
  );


  not
  g199
  (
    n203,
    n92
  );


  buf
  g200
  (
    n266,
    n107
  );


  buf
  g201
  (
    n374,
    n73
  );


  not
  g202
  (
    n343,
    n81
  );


  buf
  g203
  (
    n373,
    n50
  );


  not
  g204
  (
    n258,
    n141
  );


  not
  g205
  (
    n278,
    n93
  );


  buf
  g206
  (
    n299,
    n46
  );


  buf
  g207
  (
    n247,
    n36
  );


  buf
  g208
  (
    n213,
    n144
  );


  buf
  g209
  (
    n371,
    n96
  );


  buf
  g210
  (
    n390,
    n106
  );


  not
  g211
  (
    n233,
    n100
  );


  not
  g212
  (
    n339,
    n140
  );


  not
  g213
  (
    n369,
    n79
  );


  buf
  g214
  (
    n396,
    n132
  );


  not
  g215
  (
    n226,
    n53
  );


  not
  g216
  (
    n273,
    n59
  );


  buf
  g217
  (
    n327,
    n144
  );


  not
  g218
  (
    n171,
    n95
  );


  buf
  g219
  (
    n169,
    n116
  );


  buf
  g220
  (
    n340,
    n93
  );


  not
  g221
  (
    n159,
    n77
  );


  buf
  g222
  (
    n338,
    n83
  );


  not
  g223
  (
    n193,
    n147
  );


  not
  g224
  (
    n367,
    n140
  );


  buf
  g225
  (
    n237,
    n131
  );


  not
  g226
  (
    n161,
    n99
  );


  not
  g227
  (
    n308,
    n51
  );


  not
  g228
  (
    KeyWire_0_14,
    n81
  );


  buf
  g229
  (
    n311,
    n90
  );


  not
  g230
  (
    n342,
    n125
  );


  buf
  g231
  (
    n382,
    n72
  );


  buf
  g232
  (
    n157,
    n57
  );


  not
  g233
  (
    n290,
    n142
  );


  buf
  g234
  (
    n190,
    n109
  );


  not
  g235
  (
    n254,
    n62
  );


  buf
  g236
  (
    n306,
    n69
  );


  not
  g237
  (
    n272,
    n106
  );


  buf
  g238
  (
    n256,
    n124
  );


  not
  g239
  (
    n277,
    n118
  );


  buf
  g240
  (
    n292,
    n124
  );


  buf
  g241
  (
    n319,
    n80
  );


  not
  g242
  (
    KeyWire_0_4,
    n69
  );


  buf
  g243
  (
    n219,
    n68
  );


  not
  g244
  (
    n245,
    n134
  );


  not
  g245
  (
    n351,
    n124
  );


  not
  g246
  (
    n222,
    n66
  );


  buf
  g247
  (
    n198,
    n76
  );


  not
  g248
  (
    n235,
    n125
  );


  buf
  g249
  (
    n324,
    n136
  );


  not
  g250
  (
    KeyWire_0_6,
    n53
  );


  buf
  g251
  (
    n206,
    n137
  );


  buf
  g252
  (
    n350,
    n55
  );


  buf
  g253
  (
    n301,
    n121
  );


  not
  g254
  (
    n236,
    n84
  );


  buf
  g255
  (
    n160,
    n33
  );


  not
  g256
  (
    n271,
    n100
  );


  not
  g257
  (
    n187,
    n61
  );


  buf
  g258
  (
    n176,
    n147
  );


  not
  g259
  (
    n330,
    n119
  );


  buf
  g260
  (
    n228,
    n33
  );


  buf
  g261
  (
    n234,
    n46
  );


  not
  g262
  (
    KeyWire_0_16,
    n71
  );


  buf
  g263
  (
    n362,
    n43
  );


  buf
  g264
  (
    n361,
    n143
  );


  buf
  g265
  (
    n207,
    n103
  );


  buf
  g266
  (
    n265,
    n58
  );


  not
  g267
  (
    n249,
    n53
  );


  not
  g268
  (
    n279,
    n94
  );


  not
  g269
  (
    n177,
    n108
  );


  buf
  g270
  (
    n302,
    n68
  );


  not
  g271
  (
    n334,
    n91
  );


  buf
  g272
  (
    n253,
    n112
  );


  not
  g273
  (
    n335,
    n122
  );


  not
  g274
  (
    n370,
    n94
  );


  buf
  g275
  (
    n163,
    n123
  );


  buf
  g276
  (
    n288,
    n119
  );


  buf
  g277
  (
    n360,
    n69
  );


  buf
  g278
  (
    n244,
    n98
  );


  buf
  g279
  (
    n178,
    n135
  );


  buf
  g280
  (
    n188,
    n82
  );


  buf
  g281
  (
    n358,
    n55
  );


  buf
  g282
  (
    n232,
    n64
  );


  not
  g283
  (
    n323,
    n67
  );


  not
  g284
  (
    n377,
    n45
  );


  buf
  g285
  (
    n257,
    n35
  );


  buf
  g286
  (
    n368,
    n65
  );


  buf
  g287
  (
    n286,
    n88
  );


  not
  g288
  (
    n242,
    n146
  );


  buf
  g289
  (
    n356,
    n143
  );


  buf
  g290
  (
    n173,
    n79
  );


  nor
  g291
  (
    n394,
    n89,
    n43
  );


  and
  g292
  (
    n174,
    n90,
    n54,
    n141,
    n48
  );


  or
  g293
  (
    n325,
    n55,
    n141,
    n145,
    n118
  );


  xnor
  g294
  (
    n309,
    n106,
    n77,
    n61,
    n139
  );


  and
  g295
  (
    n240,
    n33,
    n146,
    n111,
    n115
  );


  xor
  g296
  (
    n388,
    n39,
    n46,
    n142,
    n74
  );


  or
  g297
  (
    n305,
    n105,
    n84,
    n58,
    n44
  );


  and
  g298
  (
    n179,
    n55,
    n56,
    n86,
    n48
  );


  nor
  g299
  (
    n220,
    n80,
    n35,
    n147,
    n64
  );


  or
  g300
  (
    n182,
    n63,
    n84,
    n123,
    n126
  );


  or
  g301
  (
    n310,
    n130,
    n45,
    n114,
    n134
  );


  or
  g302
  (
    n239,
    n108,
    n63,
    n116,
    n128
  );


  xor
  g303
  (
    n243,
    n114,
    n102,
    n68,
    n64
  );


  xor
  g304
  (
    n385,
    n104,
    n110,
    n44,
    n113
  );


  or
  g305
  (
    n189,
    n52,
    n94,
    n105,
    n75
  );


  xnor
  g306
  (
    n221,
    n122,
    n111,
    n105,
    n87
  );


  nand
  g307
  (
    n164,
    n102,
    n53,
    n110,
    n105
  );


  and
  g308
  (
    n353,
    n121,
    n95,
    n92,
    n80
  );


  or
  g309
  (
    n200,
    n139,
    n90,
    n103,
    n62
  );


  xor
  g310
  (
    n211,
    n129,
    n96,
    n78,
    n59
  );


  xor
  g311
  (
    n229,
    n82,
    n85,
    n40,
    n120
  );


  and
  g312
  (
    n349,
    n71,
    n58,
    n135,
    n84
  );


  and
  g313
  (
    n348,
    n121,
    n49,
    n133,
    n75
  );


  nor
  g314
  (
    n175,
    n52,
    n43,
    n101
  );


  or
  g315
  (
    n246,
    n41,
    n136,
    n49
  );


  xor
  g316
  (
    n194,
    n54,
    n78,
    n97,
    n110
  );


  or
  g317
  (
    n192,
    n111,
    n56,
    n81,
    n89
  );


  or
  g318
  (
    n172,
    n92,
    n99,
    n57,
    n117
  );


  xnor
  g319
  (
    n223,
    n140,
    n130,
    n96,
    n145
  );


  xnor
  g320
  (
    n202,
    n83,
    n124,
    n49,
    n71
  );


  nand
  g321
  (
    n274,
    n38,
    n51,
    n118,
    n145
  );


  nand
  g322
  (
    n191,
    n79,
    n64,
    n95,
    n73
  );


  or
  g323
  (
    n241,
    n131,
    n38,
    n91,
    n41
  );


  and
  g324
  (
    n387,
    n50,
    n42,
    n115,
    n97
  );


  xnor
  g325
  (
    n263,
    n88,
    n107,
    n78,
    n106
  );


  or
  g326
  (
    n314,
    n113,
    n109,
    n57,
    n65
  );


  and
  g327
  (
    n183,
    n47,
    n126,
    n72,
    n95
  );


  and
  g328
  (
    n281,
    n89,
    n67,
    n138,
    n116
  );


  and
  g329
  (
    n303,
    n134,
    n37,
    n45,
    n130
  );


  nand
  g330
  (
    n165,
    n74,
    n59,
    n146,
    n68
  );


  nor
  g331
  (
    n296,
    n141,
    n117,
    n60,
    n91
  );


  or
  g332
  (
    n255,
    n83,
    n99,
    n70,
    n97
  );


  xnor
  g333
  (
    n378,
    n65,
    n127,
    n39,
    n75
  );


  xor
  g334
  (
    n215,
    n98,
    n44,
    n123,
    n109
  );


  xor
  g335
  (
    n344,
    n71,
    n148,
    n66,
    n139
  );


  xor
  g336
  (
    n168,
    n115,
    n88,
    n34,
    n130
  );


  nand
  g337
  (
    n251,
    n78,
    n142,
    n38,
    n112
  );


  and
  g338
  (
    n238,
    n35,
    n103,
    n82,
    n48
  );


  nor
  g339
  (
    n365,
    n122,
    n83,
    n37,
    n50
  );


  xor
  g340
  (
    n280,
    n120,
    n113,
    n137,
    n102
  );


  and
  g341
  (
    n210,
    n75,
    n45,
    n86,
    n101
  );


  nand
  g342
  (
    n320,
    n112,
    n132,
    n137,
    n56
  );


  or
  g343
  (
    n276,
    n122,
    n54,
    n129
  );


  nor
  g344
  (
    n224,
    n134,
    n35,
    n89,
    n93
  );


  or
  g345
  (
    n372,
    n36,
    n69,
    n139,
    n77
  );


  xnor
  g346
  (
    n208,
    n133,
    n49,
    n126,
    n59
  );


  xnor
  g347
  (
    n205,
    n67,
    n43,
    n108,
    n126
  );


  xor
  g348
  (
    n331,
    n100,
    n104,
    n38,
    n82
  );


  or
  g349
  (
    n167,
    n98,
    n129,
    n107,
    n123
  );


  nor
  g350
  (
    n379,
    n96,
    n100,
    n34,
    n40
  );


  xnor
  g351
  (
    n346,
    n144,
    n63,
    n94,
    n46
  );


  nor
  g352
  (
    n381,
    n87,
    n98,
    n128,
    n47
  );


  nand
  g353
  (
    n395,
    n121,
    n33,
    n86,
    n34
  );


  and
  g354
  (
    n304,
    n146,
    n72,
    n37,
    n81
  );


  xor
  g355
  (
    n391,
    n138,
    n56,
    n131,
    n148
  );


  and
  g356
  (
    n355,
    n91,
    n39,
    n77,
    n66
  );


  or
  g357
  (
    n392,
    n37,
    n73,
    n70,
    n72
  );


  nand
  g358
  (
    n262,
    n88,
    n74,
    n85
  );


  nor
  g359
  (
    n248,
    n132,
    n67,
    n101,
    n36
  );


  nor
  g360
  (
    n300,
    n125,
    n102,
    n107,
    n109
  );


  or
  g361
  (
    n307,
    n70,
    n58,
    n135,
    n47
  );


  nor
  g362
  (
    n397,
    n137,
    n113,
    n42,
    n44
  );


  xnor
  g363
  (
    n386,
    n110,
    n42,
    n87,
    n144
  );


  or
  g364
  (
    n252,
    n127,
    n142,
    n86,
    n34
  );


  buf
  g365
  (
    n551,
    n249
  );


  buf
  g366
  (
    n428,
    n198
  );


  buf
  g367
  (
    n456,
    n337
  );


  not
  g368
  (
    KeyWire_0_27,
    n221
  );


  not
  g369
  (
    n543,
    n343
  );


  not
  g370
  (
    n478,
    n254
  );


  buf
  g371
  (
    n501,
    n342
  );


  buf
  g372
  (
    n514,
    n187
  );


  buf
  g373
  (
    n559,
    n306
  );


  not
  g374
  (
    n483,
    n342
  );


  buf
  g375
  (
    n536,
    n288
  );


  buf
  g376
  (
    n479,
    n331
  );


  buf
  g377
  (
    n448,
    n292
  );


  not
  g378
  (
    n517,
    n226
  );


  not
  g379
  (
    n408,
    n174
  );


  buf
  g380
  (
    n557,
    n170
  );


  not
  g381
  (
    n529,
    n315
  );


  buf
  g382
  (
    n413,
    n300
  );


  buf
  g383
  (
    n490,
    n255
  );


  buf
  g384
  (
    n430,
    n196
  );


  buf
  g385
  (
    n444,
    n180
  );


  not
  g386
  (
    n398,
    n350
  );


  buf
  g387
  (
    n455,
    n193
  );


  buf
  g388
  (
    n465,
    n318
  );


  not
  g389
  (
    n470,
    n237
  );


  not
  g390
  (
    n486,
    n286
  );


  buf
  g391
  (
    n422,
    n231
  );


  not
  g392
  (
    n482,
    n164
  );


  not
  g393
  (
    n527,
    n194
  );


  buf
  g394
  (
    n499,
    n279
  );


  buf
  g395
  (
    n519,
    n317
  );


  not
  g396
  (
    n457,
    n234
  );


  not
  g397
  (
    n513,
    n174
  );


  buf
  g398
  (
    n516,
    n185
  );


  not
  g399
  (
    n468,
    n200
  );


  not
  g400
  (
    n426,
    n345
  );


  not
  g401
  (
    n412,
    n320
  );


  buf
  g402
  (
    n460,
    n282
  );


  not
  g403
  (
    n498,
    n355
  );


  buf
  g404
  (
    n542,
    n196
  );


  not
  g405
  (
    n452,
    n259
  );


  not
  g406
  (
    n553,
    n241
  );


  buf
  g407
  (
    n561,
    n182
  );


  buf
  g408
  (
    n562,
    n192
  );


  buf
  g409
  (
    n535,
    n202
  );


  buf
  g410
  (
    n548,
    n258
  );


  buf
  g411
  (
    n447,
    n265
  );


  not
  g412
  (
    n491,
    n260
  );


  buf
  g413
  (
    KeyWire_0_31,
    n236
  );


  buf
  g414
  (
    n420,
    n157
  );


  buf
  g415
  (
    n492,
    n159
  );


  not
  g416
  (
    n511,
    n346
  );


  buf
  g417
  (
    n442,
    n334
  );


  not
  g418
  (
    n541,
    n227
  );


  buf
  g419
  (
    n435,
    n214
  );


  not
  g420
  (
    n532,
    n172
  );


  not
  g421
  (
    n488,
    n279
  );


  not
  g422
  (
    n480,
    n299
  );


  buf
  g423
  (
    n495,
    n171
  );


  buf
  g424
  (
    n552,
    n168
  );


  not
  g425
  (
    n494,
    n333
  );


  not
  g426
  (
    n484,
    n307
  );


  not
  g427
  (
    n510,
    n206
  );


  buf
  g428
  (
    n407,
    n288
  );


  buf
  g429
  (
    n520,
    n328
  );


  not
  g430
  (
    n410,
    n284
  );


  buf
  g431
  (
    n477,
    n160
  );


  not
  g432
  (
    KeyWire_0_25,
    n222
  );


  not
  g433
  (
    n487,
    n277
  );


  buf
  g434
  (
    n506,
    n340
  );


  buf
  g435
  (
    n540,
    n269
  );


  not
  g436
  (
    n555,
    n192
  );


  buf
  g437
  (
    n463,
    n283
  );


  not
  g438
  (
    n421,
    n332
  );


  not
  g439
  (
    n450,
    n266
  );


  not
  g440
  (
    n545,
    n198
  );


  buf
  g441
  (
    n515,
    n186
  );


  buf
  g442
  (
    n414,
    n228
  );


  buf
  g443
  (
    n489,
    n254
  );


  buf
  g444
  (
    n474,
    n179
  );


  buf
  g445
  (
    n454,
    n237
  );


  not
  g446
  (
    n546,
    n322
  );


  buf
  g447
  (
    n423,
    n185
  );


  buf
  g448
  (
    n524,
    n188
  );


  not
  g449
  (
    n503,
    n319
  );


  not
  g450
  (
    n473,
    n308
  );


  buf
  g451
  (
    n526,
    n177
  );


  not
  g452
  (
    n432,
    n205
  );


  nor
  g453
  (
    n453,
    n327,
    n337,
    n246,
    n239
  );


  xnor
  g454
  (
    n443,
    n274,
    n258,
    n214,
    n240
  );


  xor
  g455
  (
    n475,
    n199,
    n281,
    n335,
    n290
  );


  nor
  g456
  (
    n400,
    n211,
    n312,
    n326,
    n341
  );


  xnor
  g457
  (
    n550,
    n332,
    n291,
    n167,
    n350
  );


  xor
  g458
  (
    n451,
    n256,
    n351,
    n303,
    n225
  );


  nor
  g459
  (
    n462,
    n308,
    n316,
    n191,
    n218
  );


  nand
  g460
  (
    n433,
    n348,
    n262,
    n289,
    n166
  );


  xnor
  g461
  (
    n538,
    n225,
    n215,
    n184,
    n194
  );


  xnor
  g462
  (
    n512,
    n321,
    n335,
    n298,
    n344
  );


  nand
  g463
  (
    n505,
    n327,
    n338,
    n272,
    n309
  );


  nor
  g464
  (
    n415,
    n277,
    n201,
    n259,
    n184
  );


  nand
  g465
  (
    n533,
    n201,
    n224,
    n162,
    n341
  );


  xor
  g466
  (
    n431,
    n268,
    n208,
    n244,
    n219
  );


  nor
  g467
  (
    n445,
    n253,
    n242,
    n222,
    n167
  );


  xnor
  g468
  (
    n560,
    n317,
    n352,
    n347,
    n294
  );


  or
  g469
  (
    n481,
    n313,
    n273,
    n285,
    n181
  );


  nand
  g470
  (
    n528,
    n311,
    n281,
    n301,
    n266
  );


  or
  g471
  (
    n525,
    n305,
    n289,
    n257,
    n160
  );


  or
  g472
  (
    n472,
    n349,
    n212,
    n352,
    n252
  );


  or
  g473
  (
    n449,
    n190,
    n293,
    n253,
    n176
  );


  nor
  g474
  (
    n471,
    n276,
    n300,
    n295,
    n264
  );


  nor
  g475
  (
    n416,
    n219,
    n193,
    n285,
    n190
  );


  xnor
  g476
  (
    n507,
    n205,
    n215,
    n297,
    n339
  );


  xnor
  g477
  (
    n436,
    n234,
    n243,
    n159,
    n284
  );


  or
  g478
  (
    n530,
    n311,
    n336,
    n183,
    n178
  );


  nor
  g479
  (
    n417,
    n188,
    n228,
    n346,
    n181
  );


  or
  g480
  (
    n554,
    n257,
    n345,
    n301,
    n310
  );


  xor
  g481
  (
    n404,
    n280,
    n197,
    n325,
    n239
  );


  and
  g482
  (
    n437,
    n170,
    n209,
    n238,
    n230
  );


  and
  g483
  (
    n440,
    n263,
    n316,
    n274,
    n353
  );


  nand
  g484
  (
    n493,
    n206,
    n325,
    n313,
    n236
  );


  or
  g485
  (
    n434,
    n256,
    n231,
    n246,
    n168
  );


  or
  g486
  (
    n469,
    n334,
    n200,
    n216,
    n324
  );


  xor
  g487
  (
    n508,
    n278,
    n213,
    n263,
    n280
  );


  nand
  g488
  (
    n537,
    n243,
    n208,
    n304,
    n233
  );


  and
  g489
  (
    n500,
    n333,
    n261,
    n169,
    n264
  );


  or
  g490
  (
    n419,
    n220,
    n340,
    n339,
    n329
  );


  nor
  g491
  (
    n402,
    n261,
    n163,
    n197,
    n171
  );


  or
  g492
  (
    n496,
    n207,
    n306,
    n158,
    n312
  );


  nor
  g493
  (
    n467,
    n195,
    n164,
    n156,
    n294
  );


  nand
  g494
  (
    n518,
    n158,
    n295,
    n283,
    n348
  );


  nor
  g495
  (
    n521,
    n218,
    n189,
    n271,
    n269
  );


  nor
  g496
  (
    n534,
    n297,
    n296,
    n252,
    n330
  );


  nor
  g497
  (
    n459,
    n249,
    n235,
    n355,
    n173
  );


  nand
  g498
  (
    n405,
    n287,
    n211,
    n302,
    n203
  );


  xnor
  g499
  (
    n409,
    n291,
    n275,
    n232,
    n270
  );


  xnor
  g500
  (
    n539,
    n318,
    n344,
    n241,
    n250
  );


  or
  g501
  (
    n399,
    n186,
    n189,
    n329,
    n267
  );


  nand
  g502
  (
    n466,
    n157,
    n354,
    n165,
    n278
  );


  xnor
  g503
  (
    KeyWire_0_2,
    n309,
    n240,
    n251,
    n250
  );


  xnor
  g504
  (
    n461,
    n302,
    n161,
    n305,
    n177
  );


  and
  g505
  (
    n563,
    n262,
    n331,
    n226,
    n247
  );


  xnor
  g506
  (
    n427,
    n319,
    n229,
    n199,
    n349
  );


  and
  g507
  (
    n401,
    n267,
    n230,
    n314,
    n173
  );


  and
  g508
  (
    n502,
    n320,
    n265,
    n165,
    n175
  );


  xor
  g509
  (
    n522,
    n245,
    n182,
    n353,
    n203
  );


  nor
  g510
  (
    n476,
    n169,
    n271,
    n163,
    n290
  );


  xor
  g511
  (
    n424,
    n275,
    n270,
    n220,
    n282
  );


  xor
  g512
  (
    n509,
    n161,
    n328,
    n248,
    n354
  );


  or
  g513
  (
    n438,
    n324,
    n191,
    n175,
    n223
  );


  xnor
  g514
  (
    n441,
    n268,
    n315,
    n223,
    n276
  );


  xnor
  g515
  (
    n549,
    n351,
    n292,
    n326,
    n247
  );


  xor
  g516
  (
    n544,
    n233,
    n238,
    n299,
    n204
  );


  xor
  g517
  (
    n558,
    n343,
    n293,
    n204,
    n183
  );


  nor
  g518
  (
    n497,
    n287,
    n273,
    n244,
    n229
  );


  and
  g519
  (
    n439,
    n323,
    n272,
    n213,
    n207
  );


  and
  g520
  (
    n429,
    n232,
    n255,
    n178,
    n227
  );


  nor
  g521
  (
    n406,
    n212,
    n162,
    n323,
    n322
  );


  xor
  g522
  (
    n446,
    n321,
    n224,
    n235,
    n166
  );


  and
  g523
  (
    n523,
    n209,
    n298,
    n245,
    n251
  );


  xor
  g524
  (
    n403,
    n217,
    n210,
    n221,
    n172
  );


  xor
  g525
  (
    n418,
    n314,
    n248,
    n304,
    n202
  );


  nand
  g526
  (
    n425,
    n180,
    n216,
    n296,
    n156
  );


  or
  g527
  (
    n464,
    n176,
    n217,
    n260,
    n195
  );


  and
  g528
  (
    n556,
    n210,
    n187,
    n310,
    n336
  );


  and
  g529
  (
    n547,
    n242,
    n303,
    n286,
    n330
  );


  nand
  g530
  (
    n504,
    n338,
    n307,
    n347,
    n179
  );


  or
  g531
  (
    n719,
    n501,
    n426,
    n428,
    n405
  );


  nor
  g532
  (
    n695,
    n453,
    n546,
    n513,
    n461
  );


  xnor
  g533
  (
    n705,
    n504,
    n520,
    n497,
    n508
  );


  nor
  g534
  (
    n619,
    n530,
    n519,
    n459,
    n534
  );


  nand
  g535
  (
    n648,
    n434,
    n503,
    n556,
    n428
  );


  and
  g536
  (
    n623,
    n410,
    n524,
    n416,
    n511
  );


  xnor
  g537
  (
    n689,
    n489,
    n423,
    n521,
    n455
  );


  and
  g538
  (
    n699,
    n454,
    n512,
    n449,
    n559
  );


  xor
  g539
  (
    n618,
    n414,
    n514,
    n542,
    n472
  );


  and
  g540
  (
    n692,
    n492,
    n430,
    n558,
    n468
  );


  xnor
  g541
  (
    n637,
    n423,
    n407,
    n452,
    n500
  );


  nand
  g542
  (
    n702,
    n509,
    n413,
    n531,
    n486
  );


  and
  g543
  (
    n602,
    n539,
    n537,
    n535,
    n534
  );


  nand
  g544
  (
    n590,
    n427,
    n401,
    n432,
    n470
  );


  nand
  g545
  (
    n672,
    n489,
    n403,
    n442,
    n482
  );


  nand
  g546
  (
    n633,
    n426,
    n462,
    n463,
    n496
  );


  or
  g547
  (
    n625,
    n534,
    n533,
    n434,
    n399
  );


  or
  g548
  (
    n632,
    n466,
    n483,
    n494,
    n527
  );


  nand
  g549
  (
    n600,
    n508,
    n516,
    n490,
    n450
  );


  or
  g550
  (
    n697,
    n444,
    n417,
    n496,
    n421
  );


  nor
  g551
  (
    n654,
    n467,
    n425,
    n497,
    n486
  );


  nand
  g552
  (
    n640,
    n536,
    n511,
    n523,
    n466
  );


  xor
  g553
  (
    n713,
    n468,
    n475,
    n498,
    n537
  );


  xor
  g554
  (
    n634,
    n562,
    n524,
    n544,
    n504
  );


  xor
  g555
  (
    n645,
    n525,
    n409,
    n526,
    n484
  );


  and
  g556
  (
    n596,
    n442,
    n458,
    n486,
    n551
  );


  nand
  g557
  (
    n574,
    n518,
    n509,
    n542,
    n531
  );


  and
  g558
  (
    n593,
    n435,
    n433,
    n455,
    n479
  );


  or
  g559
  (
    n598,
    n557,
    n443,
    n514,
    n478
  );


  nor
  g560
  (
    n662,
    n430,
    n415,
    n490,
    n530
  );


  xnor
  g561
  (
    n579,
    n465,
    n476,
    n437,
    n528
  );


  and
  g562
  (
    n639,
    n405,
    n417,
    n439,
    n401
  );


  or
  g563
  (
    n668,
    n546,
    n525,
    n501,
    n418
  );


  nand
  g564
  (
    n711,
    n556,
    n479,
    n418,
    n417
  );


  xor
  g565
  (
    n708,
    n464,
    n445,
    n401,
    n430
  );


  nor
  g566
  (
    n567,
    n535,
    n487,
    n478,
    n485
  );


  nor
  g567
  (
    n678,
    n552,
    n468,
    n436,
    n424
  );


  or
  g568
  (
    n686,
    n423,
    n403,
    n540,
    n467
  );


  nand
  g569
  (
    n690,
    n555,
    n547,
    n421,
    n406
  );


  nor
  g570
  (
    n671,
    n410,
    n441,
    n529,
    n509
  );


  nand
  g571
  (
    n608,
    n512,
    n435,
    n513,
    n424
  );


  nand
  g572
  (
    n725,
    n501,
    n411,
    n521,
    n515
  );


  nand
  g573
  (
    n566,
    n546,
    n553,
    n449,
    n443
  );


  xnor
  g574
  (
    n657,
    n550,
    n442,
    n519,
    n483
  );


  and
  g575
  (
    n594,
    n527,
    n520,
    n433,
    n409
  );


  and
  g576
  (
    n685,
    n416,
    n553,
    n556,
    n560
  );


  and
  g577
  (
    n643,
    n457,
    n415,
    n516,
    n479
  );


  xor
  g578
  (
    n724,
    n439,
    n492,
    n403,
    n559
  );


  or
  g579
  (
    n649,
    n482,
    n398,
    n559,
    n444
  );


  nand
  g580
  (
    n712,
    n558,
    n400,
    n541,
    n493
  );


  nor
  g581
  (
    n624,
    n557,
    n412,
    n436,
    n473
  );


  or
  g582
  (
    n586,
    n499,
    n497,
    n407,
    n507
  );


  xnor
  g583
  (
    n622,
    n526,
    n464,
    n528,
    n553
  );


  xor
  g584
  (
    n709,
    n539,
    n481,
    n411,
    n536
  );


  nor
  g585
  (
    n569,
    n529,
    n470,
    n560,
    n485
  );


  and
  g586
  (
    n614,
    n411,
    n447,
    n414,
    n500
  );


  xnor
  g587
  (
    n588,
    n518,
    n423,
    n480,
    n445
  );


  xor
  g588
  (
    n621,
    n437,
    n422,
    n549,
    n404
  );


  xor
  g589
  (
    n651,
    n436,
    n495,
    n492,
    n508
  );


  and
  g590
  (
    n714,
    n414,
    n462,
    n408,
    n426
  );


  and
  g591
  (
    KeyWire_0_1,
    n554,
    n477,
    n543,
    n544
  );


  nor
  g592
  (
    n684,
    n457,
    n420,
    n464,
    n456
  );


  nor
  g593
  (
    n706,
    n491,
    n438,
    n517,
    n503
  );


  nor
  g594
  (
    n568,
    n522,
    n441,
    n444,
    n487
  );


  xnor
  g595
  (
    n580,
    n454,
    n429,
    n474,
    n413
  );


  nor
  g596
  (
    n642,
    n402,
    n541,
    n547,
    n498
  );


  nand
  g597
  (
    n669,
    n477,
    n552,
    n474,
    n417
  );


  or
  g598
  (
    n635,
    n440,
    n443,
    n561,
    n444
  );


  or
  g599
  (
    KeyWire_0_19,
    n549,
    n402,
    n483,
    n494
  );


  nor
  g600
  (
    n707,
    n484,
    n544,
    n424,
    n533
  );


  or
  g601
  (
    n627,
    n523,
    n472,
    n510,
    n502
  );


  nand
  g602
  (
    n572,
    n454,
    n412,
    n517,
    n533
  );


  or
  g603
  (
    n630,
    n427,
    n508,
    n458,
    n524
  );


  nand
  g604
  (
    n595,
    n552,
    n473,
    n441,
    n538
  );


  xnor
  g605
  (
    n565,
    n510,
    n453,
    n461,
    n421
  );


  nand
  g606
  (
    n607,
    n522,
    n563,
    n404
  );


  xnor
  g607
  (
    n599,
    n555,
    n539,
    n528,
    n447
  );


  nor
  g608
  (
    n670,
    n408,
    n479,
    n517,
    n446
  );


  nand
  g609
  (
    n661,
    n517,
    n438,
    n500,
    n463
  );


  nand
  g610
  (
    n680,
    n499,
    n527,
    n428,
    n543
  );


  and
  g611
  (
    n652,
    n419,
    n419,
    n413,
    n435
  );


  or
  g612
  (
    n570,
    n563,
    n557,
    n495,
    n538
  );


  nand
  g613
  (
    n606,
    n472,
    n475,
    n420,
    n481
  );


  or
  g614
  (
    n679,
    n524,
    n557,
    n520,
    n455
  );


  nor
  g615
  (
    KeyWire_0_17,
    n445,
    n450,
    n551,
    n433
  );


  or
  g616
  (
    n592,
    n430,
    n412,
    n531,
    n446
  );


  xnor
  g617
  (
    n675,
    n475,
    n425,
    n495,
    n465
  );


  xnor
  g618
  (
    n710,
    n555,
    n445,
    n450,
    n534
  );


  xor
  g619
  (
    n658,
    n440,
    n522,
    n451,
    n426
  );


  or
  g620
  (
    n718,
    n460,
    n469,
    n505,
    n453
  );


  or
  g621
  (
    n585,
    n446,
    n505,
    n550,
    n477
  );


  or
  g622
  (
    n665,
    n477,
    n493,
    n543,
    n506
  );


  xnor
  g623
  (
    n603,
    n519,
    n441,
    n463,
    n556
  );


  and
  g624
  (
    n609,
    n452,
    n507,
    n439,
    n489
  );


  nand
  g625
  (
    n676,
    n504,
    n514,
    n516,
    n513
  );


  xor
  g626
  (
    n617,
    n523,
    n436,
    n419,
    n422
  );


  xor
  g627
  (
    n723,
    n478,
    n442,
    n465,
    n548
  );


  or
  g628
  (
    n610,
    n428,
    n432,
    n490,
    n476
  );


  xnor
  g629
  (
    n631,
    n506,
    n413,
    n434,
    n448
  );


  or
  g630
  (
    n583,
    n521,
    n512,
    n509,
    n434
  );


  nand
  g631
  (
    n700,
    n497,
    n537,
    n480,
    n528
  );


  nand
  g632
  (
    n666,
    n494,
    n415,
    n405,
    n531
  );


  and
  g633
  (
    n691,
    n537,
    n553,
    n549,
    n511
  );


  xor
  g634
  (
    n674,
    n406,
    n539,
    n535,
    n467
  );


  and
  g635
  (
    n693,
    n491,
    n421,
    n466,
    n465
  );


  xnor
  g636
  (
    n577,
    n527,
    n469,
    n487
  );


  nor
  g637
  (
    n571,
    n405,
    n476,
    n561,
    n456
  );


  xor
  g638
  (
    n722,
    n510,
    n452,
    n504,
    n410
  );


  nor
  g639
  (
    n591,
    n431,
    n411,
    n464,
    n499
  );


  xor
  g640
  (
    n660,
    n448,
    n407,
    n429,
    n457
  );


  and
  g641
  (
    n728,
    n470,
    n432,
    n476,
    n408
  );


  nand
  g642
  (
    KeyWire_0_23,
    n447,
    n402,
    n491,
    n473
  );


  nand
  g643
  (
    n601,
    n440,
    n538,
    n485,
    n429
  );


  xnor
  g644
  (
    n636,
    n462,
    n466,
    n469,
    n470
  );


  and
  g645
  (
    n694,
    n481,
    n404,
    n440,
    n545
  );


  nand
  g646
  (
    n573,
    n400,
    n489,
    n538,
    n480
  );


  xor
  g647
  (
    n673,
    n533,
    n548,
    n447,
    n482
  );


  nand
  g648
  (
    n703,
    n400,
    n409,
    n560,
    n437
  );


  and
  g649
  (
    n629,
    n562,
    n526,
    n529,
    n400
  );


  and
  g650
  (
    n704,
    n502,
    n555,
    n474,
    n532
  );


  xnor
  g651
  (
    n647,
    n496,
    n562,
    n431,
    n461
  );


  xnor
  g652
  (
    n721,
    n469,
    n558,
    n438,
    n523
  );


  xor
  g653
  (
    n612,
    n409,
    n554,
    n454,
    n451
  );


  xor
  g654
  (
    n646,
    n456,
    n512,
    n551,
    n503
  );


  nor
  g655
  (
    n582,
    n474,
    n425,
    n416,
    n561
  );


  nor
  g656
  (
    n664,
    n506,
    n438,
    n483,
    n502
  );


  nand
  g657
  (
    n696,
    n505,
    n467,
    n408,
    n516
  );


  nand
  g658
  (
    n613,
    n455,
    n505,
    n398,
    n427
  );


  and
  g659
  (
    n663,
    n540,
    n446,
    n532,
    n542
  );


  xnor
  g660
  (
    n687,
    n501,
    n425,
    n536,
    n418
  );


  xor
  g661
  (
    n650,
    n547,
    n521,
    n471,
    n532
  );


  nand
  g662
  (
    n587,
    n507,
    n485,
    n492,
    n541
  );


  or
  g663
  (
    n720,
    n541,
    n412,
    n443,
    n490
  );


  xnor
  g664
  (
    n701,
    n419,
    n458,
    n563,
    n493
  );


  xor
  g665
  (
    n620,
    n500,
    n540,
    n433,
    n460
  );


  xor
  g666
  (
    n564,
    n540,
    n420,
    n542,
    n513
  );


  xor
  g667
  (
    n626,
    n545,
    n431,
    n498,
    n486
  );


  xor
  g668
  (
    n638,
    n416,
    n526,
    n545,
    n482
  );


  xor
  g669
  (
    n717,
    n488,
    n530,
    n432,
    n472
  );


  nand
  g670
  (
    n655,
    n404,
    n559,
    n450,
    n448
  );


  or
  g671
  (
    n641,
    n536,
    n515,
    n520,
    n529
  );


  xnor
  g672
  (
    n715,
    n449,
    n422,
    n562,
    n552
  );


  or
  g673
  (
    n656,
    n437,
    n550,
    n460,
    n481
  );


  or
  g674
  (
    n698,
    n459,
    n402,
    n549,
    n493
  );


  xor
  g675
  (
    n653,
    n431,
    n420,
    n456,
    n459
  );


  or
  g676
  (
    n605,
    n488,
    n475,
    n515,
    n424
  );


  and
  g677
  (
    n616,
    n414,
    n554,
    n502,
    n452
  );


  xor
  g678
  (
    KeyWire_0_30,
    n530,
    n511,
    n543,
    n506
  );


  and
  g679
  (
    n726,
    n453,
    n525,
    n551,
    n495
  );


  nand
  g680
  (
    n667,
    n449,
    n418,
    n406
  );


  nand
  g681
  (
    n683,
    n525,
    n435,
    n471,
    n488
  );


  xnor
  g682
  (
    n604,
    n478,
    n507,
    n471,
    n499
  );


  nand
  g683
  (
    n727,
    n554,
    n510,
    n403,
    n401
  );


  xnor
  g684
  (
    n659,
    n451,
    n399,
    n522,
    n459
  );


  xor
  g685
  (
    n681,
    n415,
    n550,
    n427,
    n532
  );


  or
  g686
  (
    n682,
    n496,
    n462,
    n518,
    n451
  );


  xor
  g687
  (
    n575,
    n491,
    n558,
    n410,
    n518
  );


  or
  g688
  (
    n611,
    n448,
    n519,
    n494,
    n498
  );


  nand
  g689
  (
    n576,
    n460,
    n484,
    n514,
    n458
  );


  xor
  g690
  (
    n677,
    n548,
    n560,
    n484,
    n463
  );


  xnor
  g691
  (
    n716,
    n546,
    n457,
    n407,
    n561
  );


  or
  g692
  (
    n578,
    n547,
    n548,
    n422,
    n471
  );


  xnor
  g693
  (
    n688,
    n439,
    n515,
    n535,
    n461
  );


  xor
  g694
  (
    n584,
    n544,
    n468,
    n429,
    n488
  );


  nor
  g695
  (
    KeyWire_0_0,
    n473,
    n545,
    n503,
    n480
  );


  buf
  g696
  (
    n748,
    n567
  );


  not
  g697
  (
    n764,
    n565
  );


  buf
  g698
  (
    n765,
    n598
  );


  not
  g699
  (
    n729,
    n573
  );


  buf
  g700
  (
    n772,
    n590
  );


  not
  g701
  (
    n751,
    n576
  );


  not
  g702
  (
    n776,
    n602
  );


  buf
  g703
  (
    n747,
    n578
  );


  buf
  g704
  (
    n756,
    n575
  );


  not
  g705
  (
    n738,
    n605
  );


  not
  g706
  (
    n775,
    n608
  );


  buf
  g707
  (
    n750,
    n604
  );


  buf
  g708
  (
    n752,
    n592
  );


  not
  g709
  (
    n768,
    n583
  );


  not
  g710
  (
    n735,
    n593
  );


  buf
  g711
  (
    n766,
    n611
  );


  not
  g712
  (
    n746,
    n603
  );


  not
  g713
  (
    n733,
    n581
  );


  not
  g714
  (
    n744,
    n566
  );


  buf
  g715
  (
    n741,
    n588
  );


  buf
  g716
  (
    n754,
    n610
  );


  not
  g717
  (
    n742,
    n579
  );


  not
  g718
  (
    n771,
    n564
  );


  not
  g719
  (
    n773,
    n591
  );


  not
  g720
  (
    n734,
    n585
  );


  not
  g721
  (
    n753,
    n599
  );


  not
  g722
  (
    n760,
    n568
  );


  not
  g723
  (
    n757,
    n586
  );


  not
  g724
  (
    n761,
    n571
  );


  not
  g725
  (
    n769,
    n597
  );


  not
  g726
  (
    n759,
    n589
  );


  buf
  g727
  (
    n749,
    n577
  );


  not
  g728
  (
    n770,
    n587
  );


  buf
  g729
  (
    n763,
    n584
  );


  buf
  g730
  (
    n740,
    n601
  );


  buf
  g731
  (
    n737,
    n596
  );


  not
  g732
  (
    n762,
    n609
  );


  buf
  g733
  (
    n739,
    n595
  );


  buf
  g734
  (
    n774,
    n606
  );


  buf
  g735
  (
    n758,
    n580
  );


  buf
  g736
  (
    n731,
    n569
  );


  not
  g737
  (
    n755,
    n594
  );


  buf
  g738
  (
    n767,
    n600
  );


  buf
  g739
  (
    n736,
    n574
  );


  buf
  g740
  (
    n743,
    n570
  );


  not
  g741
  (
    KeyWire_0_11,
    n582
  );


  buf
  g742
  (
    n732,
    n607
  );


  not
  g743
  (
    n730,
    n572
  );


  xnor
  g744
  (
    n841,
    n365,
    n770,
    n774,
    n366
  );


  or
  g745
  (
    n791,
    n624,
    n377,
    n732,
    n645
  );


  and
  g746
  (
    n813,
    n744,
    n390,
    n380,
    n612
  );


  xor
  g747
  (
    n853,
    n372,
    n671,
    n684,
    n629
  );


  and
  g748
  (
    KeyWire_0_24,
    n360,
    n395,
    n737,
    n377
  );


  xor
  g749
  (
    n817,
    n377,
    n391,
    n739,
    n372
  );


  xor
  g750
  (
    n802,
    n362,
    n771,
    n766,
    n393
  );


  xnor
  g751
  (
    n884,
    n615,
    n382,
    n774,
    n394
  );


  or
  g752
  (
    n808,
    n700,
    n384,
    n381,
    n674
  );


  xor
  g753
  (
    n834,
    n746,
    n369,
    n383,
    n767
  );


  or
  g754
  (
    KeyWire_0_7,
    n381,
    n737,
    n357,
    n644
  );


  xor
  g755
  (
    n805,
    n390,
    n698,
    n731,
    n631
  );


  or
  g756
  (
    n777,
    n677,
    n396,
    n676,
    n759
  );


  nor
  g757
  (
    n879,
    n743,
    n632,
    n388,
    n649
  );


  nand
  g758
  (
    n866,
    n683,
    n752,
    n382,
    n383
  );


  and
  g759
  (
    n819,
    n634,
    n689,
    n362,
    n357
  );


  xnor
  g760
  (
    n872,
    n397,
    n368,
    n746,
    n741
  );


  nor
  g761
  (
    n787,
    n385,
    n772,
    n379,
    n374
  );


  xor
  g762
  (
    n781,
    n669,
    n729,
    n774,
    n754
  );


  xor
  g763
  (
    n789,
    n696,
    n395,
    n756,
    n382
  );


  nor
  g764
  (
    n830,
    n748,
    n745,
    n659,
    n376
  );


  or
  g765
  (
    n799,
    n397,
    n394,
    n364,
    n733
  );


  and
  g766
  (
    n850,
    n741,
    n371,
    n755,
    n746
  );


  nor
  g767
  (
    n793,
    n768,
    n384,
    n766,
    n699
  );


  nand
  g768
  (
    n867,
    n375,
    n769,
    n753,
    n752
  );


  nor
  g769
  (
    n859,
    n750,
    n765,
    n379,
    n738
  );


  nor
  g770
  (
    n803,
    n637,
    n383,
    n731,
    n384
  );


  nand
  g771
  (
    n810,
    n747,
    n370,
    n773,
    n655
  );


  nand
  g772
  (
    n875,
    n744,
    n759,
    n730,
    n692
  );


  and
  g773
  (
    n863,
    n685,
    n735,
    n758,
    n762
  );


  xnor
  g774
  (
    n874,
    n668,
    n763,
    n379,
    n749
  );


  nor
  g775
  (
    n855,
    n390,
    n366,
    n768,
    n386
  );


  nor
  g776
  (
    n807,
    n371,
    n750,
    n642,
    n365
  );


  xor
  g777
  (
    n838,
    n739,
    n733,
    n380,
    n769
  );


  nor
  g778
  (
    n857,
    n761,
    n766,
    n759,
    n378
  );


  nand
  g779
  (
    n881,
    n757,
    n690,
    n743,
    n733
  );


  nor
  g780
  (
    n852,
    n761,
    n392,
    n776,
    n374
  );


  nor
  g781
  (
    n824,
    n369,
    n613,
    n758,
    n393
  );


  and
  g782
  (
    n860,
    n653,
    n678,
    n378,
    n762
  );


  and
  g783
  (
    n883,
    n745,
    n758,
    n749
  );


  nand
  g784
  (
    n816,
    n737,
    n757,
    n731,
    n368
  );


  xor
  g785
  (
    n780,
    n370,
    n376,
    n765
  );


  xnor
  g786
  (
    n809,
    n734,
    n736,
    n614,
    n748
  );


  nand
  g787
  (
    n815,
    n744,
    n773,
    n776,
    n770
  );


  nand
  g788
  (
    n783,
    n747,
    n697,
    n364,
    n370
  );


  nand
  g789
  (
    n837,
    n369,
    n654,
    n664,
    n391
  );


  or
  g790
  (
    KeyWire_0_13,
    n386,
    n735,
    n772,
    n740
  );


  xor
  g791
  (
    n826,
    n749,
    n675,
    n640,
    n688
  );


  xor
  g792
  (
    n858,
    n356,
    n751,
    n361,
    n657
  );


  xnor
  g793
  (
    n794,
    n373,
    n756,
    n771,
    n738
  );


  nor
  g794
  (
    n862,
    n395,
    n356,
    n628,
    n371
  );


  xor
  g795
  (
    n845,
    n680,
    n376,
    n764,
    n756
  );


  xor
  g796
  (
    n868,
    n764,
    n769,
    n742,
    n691
  );


  xnor
  g797
  (
    n878,
    n373,
    n754,
    n770,
    n763
  );


  or
  g798
  (
    n842,
    n380,
    n391,
    n742,
    n367
  );


  nand
  g799
  (
    n812,
    n662,
    n391,
    n365,
    n378
  );


  and
  g800
  (
    n836,
    n383,
    n647,
    n766,
    n757
  );


  and
  g801
  (
    n847,
    n754,
    n368,
    n378,
    n392
  );


  nand
  g802
  (
    n811,
    n372,
    n735,
    n730,
    n732
  );


  xor
  g803
  (
    n825,
    n638,
    n387,
    n760,
    n392
  );


  or
  g804
  (
    n796,
    n364,
    n767,
    n739,
    n673
  );


  nand
  g805
  (
    n851,
    n630,
    n741,
    n761,
    n687
  );


  nor
  g806
  (
    n797,
    n367,
    n682,
    n751,
    n775
  );


  or
  g807
  (
    n880,
    n667,
    n742,
    n770,
    n648
  );


  nand
  g808
  (
    n829,
    n750,
    n775,
    n737,
    n773
  );


  xor
  g809
  (
    n792,
    n776,
    n375,
    n775,
    n394
  );


  nand
  g810
  (
    n865,
    n389,
    n752,
    n753,
    n744
  );


  nand
  g811
  (
    n844,
    n772,
    n381,
    n760,
    n658
  );


  xnor
  g812
  (
    n790,
    n732,
    n765,
    n672,
    n774
  );


  xor
  g813
  (
    n814,
    n767,
    n771,
    n775,
    n760
  );


  xor
  g814
  (
    n795,
    n359,
    n360,
    n623,
    n758
  );


  xor
  g815
  (
    n820,
    n363,
    n776,
    n373,
    n379
  );


  and
  g816
  (
    n786,
    n367,
    n740,
    n396,
    n377
  );


  xnor
  g817
  (
    n877,
    n670,
    n750,
    n733,
    n387
  );


  and
  g818
  (
    n800,
    n643,
    n625,
    n639,
    n368
  );


  nand
  g819
  (
    n832,
    n732,
    n617,
    n393,
    n385
  );


  xor
  g820
  (
    n839,
    n626,
    n755,
    n771
  );


  xnor
  g821
  (
    n818,
    n396,
    n394,
    n681,
    n397
  );


  xnor
  g822
  (
    n835,
    n734,
    n627,
    n679,
    n748
  );


  or
  g823
  (
    n806,
    n372,
    n772,
    n367,
    n763
  );


  nor
  g824
  (
    n778,
    n366,
    n382,
    n389,
    n384
  );


  nor
  g825
  (
    n864,
    n762,
    n753,
    n388,
    n663
  );


  and
  g826
  (
    n779,
    n748,
    n745,
    n358,
    n755
  );


  nor
  g827
  (
    n843,
    n741,
    n395,
    n371,
    n621
  );


  and
  g828
  (
    n821,
    n616,
    n736,
    n618,
    n388
  );


  nand
  g829
  (
    n827,
    n641,
    n747,
    n739,
    n753
  );


  or
  g830
  (
    n861,
    n633,
    n743,
    n764
  );


  nand
  g831
  (
    n801,
    n389,
    n763,
    n695,
    n635
  );


  xnor
  g832
  (
    n784,
    n366,
    n729,
    n636,
    n363
  );


  xor
  g833
  (
    n788,
    n373,
    n736,
    n380,
    n386
  );


  xor
  g834
  (
    n823,
    n767,
    n742,
    n359,
    n757
  );


  nor
  g835
  (
    n873,
    n773,
    n385,
    n387,
    n376
  );


  nand
  g836
  (
    n833,
    n760,
    n361,
    n740,
    n650
  );


  or
  g837
  (
    n856,
    n738,
    n651,
    n751,
    n385
  );


  nand
  g838
  (
    n882,
    n768,
    n693,
    n746,
    n388
  );


  nor
  g839
  (
    n785,
    n769,
    n374,
    n752,
    n738
  );


  nor
  g840
  (
    n822,
    n622,
    n764,
    n652,
    n734
  );


  nor
  g841
  (
    n876,
    n661,
    n386,
    n375,
    n694
  );


  nor
  g842
  (
    n804,
    n389,
    n358,
    n392,
    n666
  );


  nor
  g843
  (
    n840,
    n734,
    n375,
    n730,
    n701
  );


  or
  g844
  (
    n848,
    n761,
    n646,
    n730,
    n735
  );


  nand
  g845
  (
    n854,
    n364,
    n381,
    n387,
    n759
  );


  xor
  g846
  (
    n871,
    n619,
    n660,
    n751,
    n369
  );


  nand
  g847
  (
    n849,
    n365,
    n740,
    n686,
    n736
  );


  nor
  g848
  (
    n831,
    n397,
    n665,
    n768,
    n396
  );


  nand
  g849
  (
    n828,
    n393,
    n762,
    n745,
    n620
  );


  nand
  g850
  (
    n869,
    n390,
    n370,
    n656,
    n754
  );


  xnor
  g851
  (
    n798,
    n747,
    n374,
    n731,
    n756
  );


  or
  g852
  (
    KeyWire_0_28,
    n815,
    n868,
    n814,
    n793
  );


  or
  g853
  (
    n929,
    n883,
    n803,
    n791,
    n848
  );


  nor
  g854
  (
    n925,
    n808,
    n798,
    n828,
    n865
  );


  and
  g855
  (
    n912,
    n791,
    n800,
    n818,
    n847
  );


  and
  g856
  (
    n890,
    n880,
    n826,
    n852,
    n868
  );


  nor
  g857
  (
    n896,
    n879,
    n863,
    n805,
    n820
  );


  xor
  g858
  (
    n909,
    n810,
    n843,
    n881,
    n839
  );


  and
  g859
  (
    n918,
    n798,
    n866,
    n841,
    n838
  );


  nand
  g860
  (
    n891,
    n794,
    n840,
    n779,
    n843
  );


  and
  g861
  (
    n937,
    n855,
    n865,
    n880,
    n819
  );


  xor
  g862
  (
    KeyWire_0_8,
    n789,
    n851,
    n869,
    n803
  );


  xnor
  g863
  (
    KeyWire_0_20,
    n851,
    n802,
    n796,
    n792
  );


  nor
  g864
  (
    KeyWire_0_21,
    n797,
    n790,
    n824,
    n848
  );


  or
  g865
  (
    n913,
    n850,
    n785,
    n783,
    n837
  );


  and
  g866
  (
    n902,
    n784,
    n831,
    n882,
    n801
  );


  or
  g867
  (
    n924,
    n849,
    n826,
    n840,
    n873
  );


  nor
  g868
  (
    n922,
    n852,
    n844,
    n819,
    n867
  );


  nand
  g869
  (
    n915,
    n812,
    n825,
    n800,
    n778
  );


  and
  g870
  (
    n885,
    n834,
    n824,
    n881,
    n861
  );


  nand
  g871
  (
    n927,
    n847,
    n790,
    n817,
    n799
  );


  xor
  g872
  (
    n934,
    n795,
    n834,
    n858,
    n862
  );


  xor
  g873
  (
    n907,
    n777,
    n871,
    n835,
    n815
  );


  nor
  g874
  (
    n888,
    n849,
    n877,
    n870,
    n802
  );


  or
  g875
  (
    n893,
    n801,
    n878,
    n871,
    n828
  );


  xnor
  g876
  (
    n900,
    n782,
    n816,
    n827,
    n876
  );


  or
  g877
  (
    n936,
    n805,
    n837,
    n804,
    n782
  );


  nor
  g878
  (
    n904,
    n811,
    n846,
    n793,
    n862
  );


  nor
  g879
  (
    n919,
    n807,
    n838,
    n812,
    n817
  );


  nor
  g880
  (
    n901,
    n853,
    n807,
    n799,
    n783
  );


  nand
  g881
  (
    n928,
    n836,
    n858,
    n833,
    n857
  );


  or
  g882
  (
    n932,
    n842,
    n856,
    n822,
    n806
  );


  nor
  g883
  (
    n897,
    n780,
    n882,
    n788,
    n860
  );


  nor
  g884
  (
    n905,
    n778,
    n787,
    n809,
    n854
  );


  or
  g885
  (
    n935,
    n795,
    n861,
    n869,
    n810
  );


  or
  g886
  (
    n916,
    n873,
    n816,
    n874,
    n830
  );


  and
  g887
  (
    n931,
    n859,
    n845,
    n857,
    n813
  );


  xor
  g888
  (
    n898,
    n780,
    n794,
    n860,
    n832
  );


  or
  g889
  (
    n889,
    n844,
    n875,
    n839,
    n796
  );


  xnor
  g890
  (
    n921,
    n831,
    n822,
    n821,
    n867
  );


  nand
  g891
  (
    n917,
    n784,
    n797,
    n820,
    n781
  );


  nand
  g892
  (
    n903,
    n787,
    n835,
    n789,
    n874
  );


  nand
  g893
  (
    n886,
    n877,
    n813,
    n825,
    n853
  );


  nand
  g894
  (
    n911,
    n823,
    n841,
    n872,
    n811
  );


  xor
  g895
  (
    n887,
    n850,
    n870,
    n809,
    n830
  );


  and
  g896
  (
    n926,
    n866,
    n823,
    n878,
    n846
  );


  xor
  g897
  (
    n908,
    n829,
    n786,
    n856,
    n842
  );


  xnor
  g898
  (
    n923,
    n845,
    n792,
    n829,
    n827
  );


  nor
  g899
  (
    n914,
    n875,
    n818,
    n786,
    n781
  );


  and
  g900
  (
    n892,
    n814,
    n821,
    n833,
    n788
  );


  xor
  g901
  (
    n899,
    n836,
    n879,
    n779,
    n872
  );


  or
  g902
  (
    n930,
    n863,
    n832,
    n876,
    n785
  );


  nor
  g903
  (
    n920,
    n859,
    n808,
    n855,
    n806
  );


  xor
  g904
  (
    KeyWire_0_18,
    n804,
    n864,
    n854
  );


  buf
  g905
  (
    n981,
    n899
  );


  not
  g906
  (
    n971,
    n907
  );


  not
  g907
  (
    n982,
    n914
  );


  not
  g908
  (
    n995,
    n927
  );


  not
  g909
  (
    n954,
    n933
  );


  buf
  g910
  (
    n978,
    n915
  );


  not
  g911
  (
    n974,
    n898
  );


  not
  g912
  (
    n983,
    n921
  );


  not
  g913
  (
    n962,
    n922
  );


  not
  g914
  (
    n957,
    n902
  );


  not
  g915
  (
    KeyWire_0_12,
    n924
  );


  buf
  g916
  (
    n985,
    n915
  );


  buf
  g917
  (
    n958,
    n936
  );


  buf
  g918
  (
    n948,
    n902
  );


  not
  g919
  (
    n989,
    n928
  );


  not
  g920
  (
    n991,
    n896
  );


  not
  g921
  (
    n960,
    n907
  );


  buf
  g922
  (
    n944,
    n931
  );


  buf
  g923
  (
    n977,
    n891
  );


  not
  g924
  (
    n945,
    n928
  );


  not
  g925
  (
    n946,
    n910
  );


  buf
  g926
  (
    n990,
    n910
  );


  buf
  g927
  (
    n963,
    n893
  );


  not
  g928
  (
    n939,
    n899
  );


  buf
  g929
  (
    n947,
    n930
  );


  not
  g930
  (
    n965,
    n916
  );


  buf
  g931
  (
    n968,
    n916
  );


  buf
  g932
  (
    n997,
    n918
  );


  buf
  g933
  (
    n987,
    n906
  );


  not
  g934
  (
    n967,
    n936
  );


  not
  g935
  (
    n964,
    n895
  );


  buf
  g936
  (
    n952,
    n927
  );


  not
  g937
  (
    n959,
    n894
  );


  buf
  g938
  (
    KeyWire_0_5,
    n887
  );


  not
  g939
  (
    n943,
    n934
  );


  buf
  g940
  (
    n969,
    n896
  );


  buf
  g941
  (
    n972,
    n909
  );


  not
  g942
  (
    n993,
    n913
  );


  not
  g943
  (
    n941,
    n929
  );


  not
  g944
  (
    n940,
    n933
  );


  buf
  g945
  (
    n950,
    n909
  );


  not
  g946
  (
    n980,
    n922
  );


  not
  g947
  (
    n953,
    n934
  );


  buf
  g948
  (
    n979,
    n906
  );


  buf
  g949
  (
    n961,
    n919
  );


  not
  g950
  (
    n975,
    n917
  );


  buf
  g951
  (
    n938,
    n929
  );


  buf
  g952
  (
    n986,
    n932
  );


  and
  g953
  (
    n992,
    n923,
    n908,
    n914,
    n911
  );


  xnor
  g954
  (
    n951,
    n918,
    n892,
    n895,
    n917
  );


  nand
  g955
  (
    n996,
    n897,
    n908,
    n921,
    n889
  );


  and
  g956
  (
    n949,
    n926,
    n913,
    n900,
    n931
  );


  nand
  g957
  (
    n966,
    n935,
    n904,
    n901,
    n890
  );


  nor
  g958
  (
    n994,
    n894,
    n904,
    n897,
    n920
  );


  xor
  g959
  (
    n942,
    n901,
    n924,
    n912,
    n888
  );


  nand
  g960
  (
    n956,
    n925,
    n919,
    n920,
    n893
  );


  and
  g961
  (
    n988,
    n903,
    n905,
    n930,
    n886
  );


  xor
  g962
  (
    n984,
    n923,
    n900,
    n892,
    n932
  );


  nand
  g963
  (
    n970,
    n925,
    n898,
    n935,
    n903
  );


  xnor
  g964
  (
    n973,
    n912,
    n926,
    n905,
    n911
  );


  xnor
  g965
  (
    n1000,
    n988,
    n975,
    n153,
    n984
  );


  xor
  g966
  (
    n1009,
    n972,
    n986,
    n150,
    n970
  );


  nor
  g967
  (
    n1002,
    n976,
    n971,
    n155,
    n703
  );


  xnor
  g968
  (
    n1010,
    n713,
    n964,
    n987,
    n996
  );


  and
  g969
  (
    n1003,
    n149,
    n993,
    n982,
    n994
  );


  or
  g970
  (
    n1017,
    n956,
    n153,
    n150,
    n714
  );


  xnor
  g971
  (
    n1004,
    n997,
    n154,
    n989,
    n974
  );


  and
  g972
  (
    n1012,
    n152,
    n706,
    n708,
    n717
  );


  and
  g973
  (
    n1005,
    n148,
    n712,
    n705,
    n150
  );


  xnor
  g974
  (
    n1016,
    n965,
    n980,
    n152,
    n154
  );


  and
  g975
  (
    n1007,
    n153,
    n152,
    n702,
    n148
  );


  nand
  g976
  (
    n1008,
    n150,
    n958,
    n960,
    n151
  );


  nand
  g977
  (
    n1006,
    n992,
    n710,
    n973,
    n995
  );


  and
  g978
  (
    n999,
    n154,
    n154,
    n716,
    n962
  );


  and
  g979
  (
    n1011,
    n155,
    n155,
    n957,
    n707
  );


  nand
  g980
  (
    n1015,
    n149,
    n711,
    n961,
    n983
  );


  xor
  g981
  (
    n1001,
    n967,
    n978,
    n155,
    n151
  );


  xnor
  g982
  (
    n1018,
    n153,
    n959,
    n977,
    n709
  );


  nand
  g983
  (
    n998,
    n969,
    n979,
    n991,
    n966
  );


  nor
  g984
  (
    n1014,
    n963,
    n704,
    n151,
    n715
  );


  nand
  g985
  (
    n1013,
    n981,
    n990,
    n968,
    n149
  );


  nand
  g986
  (
    n1019,
    n149,
    n985,
    n152,
    n151
  );


  nor
  g987
  (
    n1028,
    n883,
    n728,
    n1012,
    n1011
  );


  nor
  g988
  (
    n1022,
    n1007,
    n1015,
    n999,
    n1000
  );


  or
  g989
  (
    n1029,
    n722,
    n1017,
    n1016,
    n1019
  );


  xor
  g990
  (
    n1026,
    n1014,
    n725,
    n1004,
    n723
  );


  or
  g991
  (
    n1025,
    n719,
    n1014,
    n884,
    n1018
  );


  nor
  g992
  (
    n1031,
    n1015,
    n884,
    n1011,
    n1018
  );


  nand
  g993
  (
    n1020,
    n724,
    n1006,
    n1003,
    n1008
  );


  or
  g994
  (
    n1027,
    n1016,
    n1013,
    n1005,
    n1017
  );


  or
  g995
  (
    n1030,
    n727,
    n1012,
    n1013,
    n1009
  );


  xor
  g996
  (
    n1023,
    n726,
    n998,
    n937,
    n1007
  );


  nand
  g997
  (
    n1032,
    n720,
    n1006,
    n937,
    n1002
  );


  nand
  g998
  (
    n1024,
    n718,
    n1010,
    n1009,
    n721
  );


  and
  g999
  (
    n1021,
    n1019,
    n1001,
    n1008,
    n1010
  );


  xnor
  KeyGate_0_0
  (
    n628,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n589,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n531,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n35,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n352,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n955,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n316,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n782,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n933,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n209,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n77,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n745,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n976,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n870,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n298,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n218,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n322,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n644,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n894,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n597,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n895,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n910,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n64,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n581,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n846,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n485,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n73,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n411,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n906,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n354,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n615,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n458,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


