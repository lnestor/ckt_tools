

module Stat_655_65
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n669,
  n665,
  n666,
  n664,
  n674,
  n676,
  n672,
  n663,
  n660,
  n658,
  n671,
  n680,
  n662,
  n678,
  n679,
  n667,
  n675,
  n659,
  n673,
  n668,
  n677,
  n661,
  n681,
  n670,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;
  output n669;output n665;output n666;output n664;output n674;output n676;output n672;output n663;output n660;output n658;output n671;output n680;output n662;output n678;output n679;output n667;output n675;output n659;output n673;output n668;output n677;output n661;output n681;output n670;
  wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n39,
    n6
  );


  not
  g1
  (
    n44,
    n1
  );


  not
  g2
  (
    n41,
    n3
  );


  not
  g3
  (
    n30,
    n4
  );


  not
  g4
  (
    n34,
    n6
  );


  buf
  g5
  (
    n36,
    n2
  );


  not
  g6
  (
    n37,
    n3
  );


  not
  g7
  (
    n33,
    n5
  );


  buf
  g8
  (
    n40,
    n4
  );


  buf
  g9
  (
    n45,
    n3
  );


  not
  g10
  (
    n38,
    n7
  );


  not
  g11
  (
    n42,
    n2
  );


  not
  g12
  (
    n31,
    n1
  );


  not
  g13
  (
    n28,
    n2
  );


  not
  g14
  (
    n32,
    n5
  );


  not
  g15
  (
    n27,
    n5
  );


  not
  g16
  (
    n43,
    n4
  );


  buf
  g17
  (
    n29,
    n6
  );


  not
  g18
  (
    n35,
    n1
  );


  not
  g19
  (
    n67,
    n41
  );


  not
  g20
  (
    n52,
    n34
  );


  not
  g21
  (
    n61,
    n38
  );


  not
  g22
  (
    n66,
    n45
  );


  not
  g23
  (
    n69,
    n30
  );


  not
  g24
  (
    n96,
    n42
  );


  buf
  g25
  (
    n51,
    n28
  );


  buf
  g26
  (
    n65,
    n29
  );


  not
  g27
  (
    n70,
    n35
  );


  not
  g28
  (
    n71,
    n42
  );


  buf
  g29
  (
    n68,
    n36
  );


  buf
  g30
  (
    n85,
    n37
  );


  buf
  g31
  (
    n84,
    n36
  );


  not
  g32
  (
    n95,
    n44
  );


  not
  g33
  (
    n58,
    n43
  );


  not
  g34
  (
    n74,
    n36
  );


  buf
  g35
  (
    n93,
    n31
  );


  buf
  g36
  (
    n59,
    n34
  );


  not
  g37
  (
    n55,
    n35
  );


  buf
  g38
  (
    n81,
    n29
  );


  not
  g39
  (
    n90,
    n40
  );


  not
  g40
  (
    n97,
    n38
  );


  buf
  g41
  (
    n62,
    n30
  );


  buf
  g42
  (
    n50,
    n45
  );


  buf
  g43
  (
    n82,
    n34
  );


  buf
  g44
  (
    n57,
    n43
  );


  buf
  g45
  (
    n99,
    n40
  );


  buf
  g46
  (
    n101,
    n39
  );


  buf
  g47
  (
    n86,
    n28
  );


  buf
  g48
  (
    n63,
    n43
  );


  not
  g49
  (
    n100,
    n29
  );


  not
  g50
  (
    n64,
    n44
  );


  buf
  g51
  (
    n89,
    n37
  );


  buf
  g52
  (
    n53,
    n45
  );


  buf
  g53
  (
    n92,
    n35
  );


  not
  g54
  (
    n79,
    n39
  );


  not
  g55
  (
    n46,
    n30
  );


  not
  g56
  (
    n83,
    n31
  );


  buf
  g57
  (
    n49,
    n33
  );


  not
  g58
  (
    n77,
    n41
  );


  not
  g59
  (
    n56,
    n44
  );


  buf
  g60
  (
    n73,
    n33
  );


  not
  g61
  (
    n78,
    n27
  );


  not
  g62
  (
    n94,
    n42
  );


  not
  g63
  (
    n87,
    n41
  );


  not
  g64
  (
    n98,
    n40
  );


  not
  g65
  (
    n60,
    n33
  );


  buf
  g66
  (
    n88,
    n32
  );


  buf
  g67
  (
    n54,
    n39
  );


  buf
  g68
  (
    n76,
    n32
  );


  buf
  g69
  (
    n47,
    n37
  );


  buf
  g70
  (
    n48,
    n38
  );


  buf
  g71
  (
    n80,
    n31
  );


  buf
  g72
  (
    n75,
    n28
  );


  not
  g73
  (
    n72,
    n32
  );


  not
  g74
  (
    n91,
    n27
  );


  not
  g75
  (
    n278,
    n95
  );


  buf
  g76
  (
    n323,
    n59
  );


  buf
  g77
  (
    n200,
    n63
  );


  not
  g78
  (
    n195,
    n61
  );


  not
  g79
  (
    n281,
    n46
  );


  not
  g80
  (
    n257,
    n85
  );


  buf
  g81
  (
    n293,
    n65
  );


  buf
  g82
  (
    n148,
    n84
  );


  buf
  g83
  (
    n309,
    n90
  );


  not
  g84
  (
    n306,
    n92
  );


  not
  g85
  (
    n274,
    n52
  );


  not
  g86
  (
    n238,
    n54
  );


  buf
  g87
  (
    n196,
    n80
  );


  buf
  g88
  (
    n128,
    n49
  );


  not
  g89
  (
    n299,
    n94
  );


  buf
  g90
  (
    n258,
    n99
  );


  not
  g91
  (
    n172,
    n97
  );


  buf
  g92
  (
    n152,
    n81
  );


  not
  g93
  (
    n129,
    n63
  );


  not
  g94
  (
    n302,
    n88
  );


  buf
  g95
  (
    n248,
    n51
  );


  buf
  g96
  (
    n255,
    n101
  );


  buf
  g97
  (
    n256,
    n77
  );


  not
  g98
  (
    n230,
    n86
  );


  not
  g99
  (
    n113,
    n60
  );


  buf
  g100
  (
    n177,
    n57
  );


  not
  g101
  (
    n202,
    n80
  );


  buf
  g102
  (
    n186,
    n91
  );


  buf
  g103
  (
    n160,
    n101
  );


  buf
  g104
  (
    n304,
    n82
  );


  not
  g105
  (
    n144,
    n73
  );


  not
  g106
  (
    n296,
    n85
  );


  buf
  g107
  (
    n307,
    n78
  );


  not
  g108
  (
    n125,
    n62
  );


  not
  g109
  (
    n167,
    n72
  );


  buf
  g110
  (
    n142,
    n95
  );


  buf
  g111
  (
    n140,
    n59
  );


  buf
  g112
  (
    n243,
    n82
  );


  buf
  g113
  (
    n156,
    n82
  );


  not
  g114
  (
    n265,
    n76
  );


  not
  g115
  (
    n103,
    n87
  );


  not
  g116
  (
    n280,
    n67
  );


  not
  g117
  (
    n316,
    n58
  );


  not
  g118
  (
    n189,
    n77
  );


  not
  g119
  (
    n127,
    n91
  );


  not
  g120
  (
    n203,
    n48
  );


  buf
  g121
  (
    n292,
    n48
  );


  buf
  g122
  (
    n241,
    n84
  );


  not
  g123
  (
    n181,
    n60
  );


  not
  g124
  (
    n108,
    n70
  );


  not
  g125
  (
    n194,
    n93
  );


  not
  g126
  (
    n282,
    n49
  );


  buf
  g127
  (
    n318,
    n49
  );


  not
  g128
  (
    n111,
    n94
  );


  not
  g129
  (
    n251,
    n86
  );


  buf
  g130
  (
    n310,
    n81
  );


  buf
  g131
  (
    n246,
    n64
  );


  buf
  g132
  (
    n224,
    n89
  );


  buf
  g133
  (
    n188,
    n58
  );


  buf
  g134
  (
    n253,
    n87
  );


  not
  g135
  (
    n229,
    n50
  );


  buf
  g136
  (
    n176,
    n76
  );


  not
  g137
  (
    n222,
    n87
  );


  buf
  g138
  (
    n155,
    n46
  );


  buf
  g139
  (
    n239,
    n54
  );


  buf
  g140
  (
    n204,
    n89
  );


  buf
  g141
  (
    n175,
    n55
  );


  not
  g142
  (
    n105,
    n100
  );


  buf
  g143
  (
    n150,
    n50
  );


  not
  g144
  (
    n117,
    n71
  );


  buf
  g145
  (
    n232,
    n83
  );


  buf
  g146
  (
    n171,
    n68
  );


  not
  g147
  (
    n219,
    n79
  );


  buf
  g148
  (
    n139,
    n83
  );


  not
  g149
  (
    n114,
    n94
  );


  buf
  g150
  (
    n269,
    n77
  );


  buf
  g151
  (
    n234,
    n99
  );


  not
  g152
  (
    n221,
    n47
  );


  not
  g153
  (
    n178,
    n95
  );


  buf
  g154
  (
    n291,
    n97
  );


  not
  g155
  (
    n104,
    n84
  );


  not
  g156
  (
    n240,
    n65
  );


  buf
  g157
  (
    n143,
    n69
  );


  not
  g158
  (
    n185,
    n66
  );


  not
  g159
  (
    n235,
    n74
  );


  not
  g160
  (
    n149,
    n56
  );


  buf
  g161
  (
    n187,
    n98
  );


  buf
  g162
  (
    n211,
    n64
  );


  not
  g163
  (
    n270,
    n52
  );


  not
  g164
  (
    n135,
    n60
  );


  not
  g165
  (
    n207,
    n90
  );


  buf
  g166
  (
    n163,
    n100
  );


  buf
  g167
  (
    n109,
    n65
  );


  buf
  g168
  (
    n294,
    n86
  );


  not
  g169
  (
    n169,
    n88
  );


  not
  g170
  (
    n107,
    n46
  );


  not
  g171
  (
    n166,
    n100
  );


  not
  g172
  (
    n218,
    n78
  );


  not
  g173
  (
    n151,
    n81
  );


  buf
  g174
  (
    n225,
    n68
  );


  not
  g175
  (
    n170,
    n61
  );


  buf
  g176
  (
    n223,
    n87
  );


  buf
  g177
  (
    n324,
    n57
  );


  not
  g178
  (
    n191,
    n72
  );


  not
  g179
  (
    n220,
    n62
  );


  buf
  g180
  (
    n317,
    n59
  );


  buf
  g181
  (
    n277,
    n86
  );


  not
  g182
  (
    n271,
    n53
  );


  buf
  g183
  (
    n173,
    n58
  );


  buf
  g184
  (
    n242,
    n48
  );


  buf
  g185
  (
    n209,
    n52
  );


  not
  g186
  (
    n227,
    n78
  );


  buf
  g187
  (
    n279,
    n90
  );


  not
  g188
  (
    n138,
    n67
  );


  not
  g189
  (
    n289,
    n97
  );


  buf
  g190
  (
    n260,
    n89
  );


  buf
  g191
  (
    n315,
    n75
  );


  buf
  g192
  (
    n244,
    n74
  );


  buf
  g193
  (
    n213,
    n77
  );


  buf
  g194
  (
    n120,
    n66
  );


  buf
  g195
  (
    n147,
    n69
  );


  not
  g196
  (
    n198,
    n80
  );


  buf
  g197
  (
    n158,
    n75
  );


  not
  g198
  (
    n300,
    n50
  );


  buf
  g199
  (
    n308,
    n99
  );


  not
  g200
  (
    n206,
    n66
  );


  buf
  g201
  (
    n133,
    n69
  );


  buf
  g202
  (
    n283,
    n47
  );


  buf
  g203
  (
    n285,
    n51
  );


  not
  g204
  (
    n199,
    n52
  );


  not
  g205
  (
    n216,
    n85
  );


  buf
  g206
  (
    n153,
    n69
  );


  not
  g207
  (
    n273,
    n76
  );


  buf
  g208
  (
    n141,
    n47
  );


  not
  g209
  (
    n303,
    n71
  );


  buf
  g210
  (
    n137,
    n55
  );


  buf
  g211
  (
    n183,
    n84
  );


  buf
  g212
  (
    n136,
    n79
  );


  buf
  g213
  (
    n272,
    n76
  );


  buf
  g214
  (
    n112,
    n91
  );


  buf
  g215
  (
    n157,
    n90
  );


  buf
  g216
  (
    n311,
    n71
  );


  not
  g217
  (
    n184,
    n63
  );


  not
  g218
  (
    n250,
    n49
  );


  not
  g219
  (
    n305,
    n53
  );


  buf
  g220
  (
    n275,
    n68
  );


  not
  g221
  (
    n102,
    n92
  );


  buf
  g222
  (
    n210,
    n53
  );


  not
  g223
  (
    n226,
    n68
  );


  buf
  g224
  (
    n268,
    n79
  );


  not
  g225
  (
    n287,
    n92
  );


  buf
  g226
  (
    n284,
    n73
  );


  buf
  g227
  (
    n201,
    n94
  );


  not
  g228
  (
    n233,
    n80
  );


  not
  g229
  (
    n118,
    n101
  );


  not
  g230
  (
    n197,
    n56
  );


  buf
  g231
  (
    n110,
    n89
  );


  buf
  g232
  (
    n252,
    n75
  );


  buf
  g233
  (
    n115,
    n73
  );


  buf
  g234
  (
    n212,
    n92
  );


  not
  g235
  (
    n237,
    n82
  );


  buf
  g236
  (
    n320,
    n66
  );


  buf
  g237
  (
    n261,
    n95
  );


  buf
  g238
  (
    n245,
    n56
  );


  buf
  g239
  (
    n276,
    n55
  );


  not
  g240
  (
    n123,
    n47
  );


  buf
  g241
  (
    n121,
    n54
  );


  not
  g242
  (
    n168,
    n96
  );


  not
  g243
  (
    n231,
    n57
  );


  not
  g244
  (
    n162,
    n72
  );


  not
  g245
  (
    n266,
    n61
  );


  not
  g246
  (
    n217,
    n85
  );


  buf
  g247
  (
    n236,
    n64
  );


  not
  g248
  (
    n301,
    n91
  );


  buf
  g249
  (
    n159,
    n93
  );


  not
  g250
  (
    n126,
    n78
  );


  not
  g251
  (
    n124,
    n70
  );


  not
  g252
  (
    n145,
    n88
  );


  not
  g253
  (
    n214,
    n98
  );


  not
  g254
  (
    n262,
    n96
  );


  not
  g255
  (
    n228,
    n65
  );


  not
  g256
  (
    n288,
    n99
  );


  not
  g257
  (
    n174,
    n62
  );


  buf
  g258
  (
    n254,
    n96
  );


  buf
  g259
  (
    n205,
    n57
  );


  not
  g260
  (
    n165,
    n79
  );


  not
  g261
  (
    n263,
    n48
  );


  buf
  g262
  (
    n131,
    n56
  );


  not
  g263
  (
    n182,
    n101
  );


  buf
  g264
  (
    n319,
    n97
  );


  not
  g265
  (
    n247,
    n51
  );


  not
  g266
  (
    n119,
    n46
  );


  buf
  g267
  (
    n290,
    n60
  );


  not
  g268
  (
    n193,
    n73
  );


  buf
  g269
  (
    n297,
    n93
  );


  buf
  g270
  (
    n190,
    n59
  );


  buf
  g271
  (
    n122,
    n74
  );


  buf
  g272
  (
    n314,
    n70
  );


  buf
  g273
  (
    n321,
    n67
  );


  not
  g274
  (
    n116,
    n83
  );


  not
  g275
  (
    n249,
    n58
  );


  buf
  g276
  (
    n295,
    n81
  );


  not
  g277
  (
    n106,
    n74
  );


  not
  g278
  (
    n264,
    n51
  );


  not
  g279
  (
    n146,
    n93
  );


  buf
  g280
  (
    n132,
    n53
  );


  buf
  g281
  (
    n325,
    n62
  );


  not
  g282
  (
    n313,
    n64
  );


  not
  g283
  (
    n164,
    n63
  );


  not
  g284
  (
    n130,
    n96
  );


  buf
  g285
  (
    n179,
    n98
  );


  not
  g286
  (
    n298,
    n67
  );


  not
  g287
  (
    n267,
    n98
  );


  not
  g288
  (
    n134,
    n50
  );


  not
  g289
  (
    n161,
    n83
  );


  buf
  g290
  (
    n215,
    n61
  );


  not
  g291
  (
    n259,
    n70
  );


  not
  g292
  (
    n312,
    n75
  );


  not
  g293
  (
    n322,
    n88
  );


  buf
  g294
  (
    n180,
    n100
  );


  buf
  g295
  (
    n154,
    n55
  );


  buf
  g296
  (
    n286,
    n54
  );


  buf
  g297
  (
    n192,
    n71
  );


  not
  g298
  (
    n208,
    n72
  );


  buf
  g299
  (
    n520,
    n144
  );


  buf
  g300
  (
    n490,
    n103
  );


  not
  g301
  (
    n553,
    n266
  );


  buf
  g302
  (
    n543,
    n186
  );


  buf
  g303
  (
    n405,
    n163
  );


  not
  g304
  (
    n452,
    n208
  );


  buf
  g305
  (
    n431,
    n235
  );


  buf
  g306
  (
    n498,
    n177
  );


  buf
  g307
  (
    n380,
    n244
  );


  not
  g308
  (
    n326,
    n134
  );


  xnor
  g309
  (
    n513,
    n102,
    n210,
    n143,
    n238
  );


  and
  g310
  (
    n400,
    n179,
    n299,
    n167,
    n310
  );


  nand
  g311
  (
    n499,
    n144,
    n260,
    n183,
    n222
  );


  xnor
  g312
  (
    n428,
    n169,
    n301,
    n256,
    n128
  );


  or
  g313
  (
    n554,
    n293,
    n11,
    n225,
    n147
  );


  and
  g314
  (
    n476,
    n240,
    n103,
    n145,
    n278
  );


  xnor
  g315
  (
    n447,
    n321,
    n25,
    n113,
    n291
  );


  nor
  g316
  (
    n371,
    n177,
    n249,
    n194,
    n304
  );


  nand
  g317
  (
    n509,
    n8,
    n233,
    n161,
    n323
  );


  xor
  g318
  (
    n484,
    n266,
    n224,
    n160,
    n20
  );


  nand
  g319
  (
    n423,
    n26,
    n280,
    n259,
    n179
  );


  xnor
  g320
  (
    n327,
    n314,
    n176,
    n243,
    n189
  );


  xor
  g321
  (
    n467,
    n152,
    n107,
    n236,
    n321
  );


  xnor
  g322
  (
    n464,
    n169,
    n244,
    n142,
    n14
  );


  or
  g323
  (
    n552,
    n159,
    n140,
    n118,
    n203
  );


  nor
  g324
  (
    n348,
    n19,
    n184,
    n150,
    n18
  );


  nand
  g325
  (
    n518,
    n131,
    n243,
    n249,
    n264
  );


  or
  g326
  (
    n459,
    n261,
    n251,
    n148,
    n315
  );


  or
  g327
  (
    n514,
    n246,
    n253,
    n195,
    n187
  );


  nand
  g328
  (
    n491,
    n228,
    n299,
    n325,
    n183
  );


  and
  g329
  (
    n451,
    n276,
    n217,
    n181,
    n260
  );


  xor
  g330
  (
    n503,
    n144,
    n232,
    n214,
    n174
  );


  or
  g331
  (
    n354,
    n192,
    n157,
    n156,
    n207
  );


  nand
  g332
  (
    n382,
    n165,
    n271,
    n170,
    n301
  );


  nand
  g333
  (
    n448,
    n14,
    n16,
    n167,
    n188
  );


  nor
  g334
  (
    n379,
    n171,
    n170,
    n235,
    n161
  );


  xnor
  g335
  (
    n512,
    n204,
    n300,
    n236,
    n241
  );


  nand
  g336
  (
    n536,
    n274,
    n15,
    n256,
    n314
  );


  and
  g337
  (
    n439,
    n108,
    n235,
    n252,
    n289
  );


  nor
  g338
  (
    n540,
    n309,
    n204,
    n155,
    n200
  );


  nand
  g339
  (
    n483,
    n297,
    n160,
    n132,
    n128
  );


  nand
  g340
  (
    n349,
    n254,
    n258,
    n267,
    n281
  );


  nand
  g341
  (
    n559,
    n169,
    n239,
    n230,
    n308
  );


  and
  g342
  (
    n424,
    n143,
    n239,
    n194,
    n117
  );


  nor
  g343
  (
    n436,
    n156,
    n322,
    n165,
    n116
  );


  or
  g344
  (
    n343,
    n237,
    n175,
    n111,
    n182
  );


  nand
  g345
  (
    n361,
    n270,
    n19,
    n272,
    n284
  );


  and
  g346
  (
    n369,
    n187,
    n292,
    n159,
    n171
  );


  xor
  g347
  (
    n481,
    n316,
    n236,
    n228,
    n106
  );


  or
  g348
  (
    n365,
    n303,
    n239,
    n140,
    n265
  );


  xnor
  g349
  (
    n383,
    n21,
    n180,
    n279,
    n24
  );


  nor
  g350
  (
    n386,
    n13,
    n211,
    n157,
    n220
  );


  nor
  g351
  (
    n442,
    n311,
    n174,
    n235,
    n212
  );


  xnor
  g352
  (
    n511,
    n214,
    n304,
    n209,
    n300
  );


  xor
  g353
  (
    n549,
    n291,
    n221,
    n120,
    n178
  );


  xor
  g354
  (
    n435,
    n297,
    n7,
    n115,
    n288
  );


  or
  g355
  (
    n555,
    n211,
    n218,
    n226,
    n310
  );


  nand
  g356
  (
    n544,
    n145,
    n220,
    n156,
    n202
  );


  xor
  g357
  (
    n482,
    n240,
    n275,
    n264,
    n305
  );


  and
  g358
  (
    n440,
    n244,
    n298,
    n323,
    n212
  );


  nand
  g359
  (
    n360,
    n168,
    n261,
    n271,
    n147
  );


  xor
  g360
  (
    n495,
    n316,
    n136,
    n257,
    n197
  );


  and
  g361
  (
    n561,
    n254,
    n113,
    n213,
    n231
  );


  and
  g362
  (
    n480,
    n117,
    n176,
    n164,
    n296
  );


  nand
  g363
  (
    n376,
    n121,
    n223,
    n170,
    n251
  );


  nor
  g364
  (
    n533,
    n301,
    n12,
    n18,
    n197
  );


  nor
  g365
  (
    n449,
    n12,
    n175,
    n294,
    n110
  );


  xor
  g366
  (
    n384,
    n185,
    n234,
    n247,
    n224
  );


  xor
  g367
  (
    n438,
    n118,
    n288,
    n196,
    n318
  );


  nand
  g368
  (
    n515,
    n260,
    n156,
    n302,
    n183
  );


  xnor
  g369
  (
    n505,
    n184,
    n317,
    n323,
    n201
  );


  xor
  g370
  (
    n517,
    n124,
    n230,
    n289,
    n208
  );


  or
  g371
  (
    n419,
    n132,
    n295,
    n233,
    n199
  );


  xor
  g372
  (
    n357,
    n253,
    n322,
    n280,
    n8
  );


  xnor
  g373
  (
    n410,
    n290,
    n224,
    n248,
    n168
  );


  or
  g374
  (
    n450,
    n243,
    n112,
    n153,
    n183
  );


  nand
  g375
  (
    n526,
    n250,
    n197,
    n294,
    n232
  );


  xor
  g376
  (
    n425,
    n190,
    n180,
    n260,
    n270
  );


  xnor
  g377
  (
    n395,
    n216,
    n11,
    n203,
    n269
  );


  xnor
  g378
  (
    n550,
    n237,
    n146,
    n135,
    n151
  );


  xor
  g379
  (
    n530,
    n212,
    n215,
    n134,
    n166
  );


  nand
  g380
  (
    n488,
    n168,
    n273,
    n155,
    n158
  );


  nor
  g381
  (
    n407,
    n306,
    n259,
    n146,
    n186
  );


  xnor
  g382
  (
    n471,
    n220,
    n309,
    n314,
    n23
  );


  nand
  g383
  (
    n453,
    n178,
    n21,
    n17,
    n202
  );


  nor
  g384
  (
    n364,
    n142,
    n238,
    n277,
    n140
  );


  or
  g385
  (
    n463,
    n286,
    n141,
    n193,
    n306
  );


  xor
  g386
  (
    n350,
    n205,
    n108,
    n225,
    n196
  );


  and
  g387
  (
    n389,
    n169,
    n321,
    n216,
    n257
  );


  and
  g388
  (
    n329,
    n199,
    n292,
    n22,
    n278
  );


  and
  g389
  (
    n539,
    n264,
    n185,
    n252,
    n139
  );


  nand
  g390
  (
    n433,
    n289,
    n273,
    n209,
    n317
  );


  xor
  g391
  (
    n532,
    n269,
    n155,
    n161,
    n240
  );


  xor
  g392
  (
    n502,
    n220,
    n219,
    n247,
    n209
  );


  nand
  g393
  (
    n342,
    n231,
    n319,
    n129,
    n163
  );


  xnor
  g394
  (
    n470,
    n10,
    n286,
    n150,
    n120
  );


  nand
  g395
  (
    n426,
    n300,
    n245,
    n11,
    n126
  );


  xor
  g396
  (
    n510,
    n208,
    n137,
    n142,
    n17
  );


  nand
  g397
  (
    n516,
    n190,
    n143,
    n324,
    n193
  );


  xor
  g398
  (
    n501,
    n258,
    n180,
    n250,
    n151
  );


  and
  g399
  (
    n475,
    n290,
    n205,
    n172,
    n150
  );


  xor
  g400
  (
    n506,
    n272,
    n155,
    n216,
    n313
  );


  nor
  g401
  (
    n385,
    n221,
    n305,
    n139,
    n131
  );


  or
  g402
  (
    n353,
    n320,
    n230,
    n250,
    n158
  );


  nor
  g403
  (
    n560,
    n112,
    n10,
    n237,
    n201
  );


  nor
  g404
  (
    n394,
    n131,
    n304,
    n312,
    n288
  );


  xnor
  g405
  (
    n397,
    n268,
    n249,
    n258,
    n271
  );


  nand
  g406
  (
    n489,
    n305,
    n9,
    n259,
    n222
  );


  and
  g407
  (
    n356,
    n242,
    n293,
    n106,
    n234
  );


  xor
  g408
  (
    n422,
    n276,
    n23,
    n255,
    n119
  );


  nand
  g409
  (
    n456,
    n225,
    n105,
    n158,
    n238
  );


  xor
  g410
  (
    n359,
    n269,
    n195,
    n151,
    n238
  );


  xor
  g411
  (
    n372,
    n164,
    n276,
    n223,
    n206
  );


  xor
  g412
  (
    n373,
    n214,
    n315,
    n104,
    n319
  );


  or
  g413
  (
    n341,
    n210,
    n198,
    n279,
    n218
  );


  xnor
  g414
  (
    n333,
    n166,
    n168,
    n184,
    n240
  );


  nand
  g415
  (
    n377,
    n270,
    n172,
    n227,
    n130
  );


  nor
  g416
  (
    n537,
    n242,
    n135,
    n124,
    n200
  );


  or
  g417
  (
    n331,
    n313,
    n152,
    n234,
    n232
  );


  or
  g418
  (
    n330,
    n213,
    n199,
    n325,
    n204
  );


  nor
  g419
  (
    n455,
    n322,
    n167,
    n290,
    n219
  );


  or
  g420
  (
    n412,
    n252,
    n300,
    n9
  );


  xnor
  g421
  (
    n528,
    n253,
    n284,
    n323,
    n248
  );


  or
  g422
  (
    n340,
    n190,
    n202,
    n251,
    n296
  );


  nor
  g423
  (
    n427,
    n267,
    n10,
    n234,
    n114
  );


  nand
  g424
  (
    n420,
    n274,
    n290,
    n208,
    n294
  );


  and
  g425
  (
    n415,
    n307,
    n172,
    n154,
    n254
  );


  nand
  g426
  (
    n558,
    n8,
    n144,
    n296,
    n320
  );


  and
  g427
  (
    n535,
    n196,
    n285,
    n263,
    n127
  );


  nor
  g428
  (
    n391,
    n257,
    n210,
    n215,
    n312
  );


  or
  g429
  (
    n351,
    n292,
    n205,
    n219,
    n309
  );


  and
  g430
  (
    n486,
    n296,
    n316,
    n222,
    n279
  );


  xnor
  g431
  (
    n403,
    n121,
    n299,
    n14,
    n321
  );


  or
  g432
  (
    n406,
    n268,
    n162,
    n130,
    n279
  );


  xor
  g433
  (
    n468,
    n248,
    n205,
    n117,
    n188
  );


  or
  g434
  (
    n396,
    n298,
    n130,
    n229,
    n227
  );


  and
  g435
  (
    n335,
    n174,
    n310,
    n241,
    n186
  );


  nand
  g436
  (
    n414,
    n258,
    n213,
    n241,
    n318
  );


  nand
  g437
  (
    n507,
    n181,
    n226,
    n112,
    n324
  );


  xnor
  g438
  (
    n465,
    n132,
    n125,
    n149,
    n223
  );


  xor
  g439
  (
    n339,
    n102,
    n147,
    n195,
    n161
  );


  nor
  g440
  (
    n344,
    n273,
    n277,
    n214,
    n113
  );


  nor
  g441
  (
    n352,
    n307,
    n191,
    n284,
    n271
  );


  xnor
  g442
  (
    n444,
    n20,
    n206,
    n237,
    n26
  );


  and
  g443
  (
    n527,
    n286,
    n211,
    n262,
    n189
  );


  or
  g444
  (
    n346,
    n311,
    n267,
    n133,
    n243
  );


  nand
  g445
  (
    n460,
    n256,
    n231,
    n283,
    n226
  );


  nor
  g446
  (
    n429,
    n263,
    n275,
    n105,
    n203
  );


  and
  g447
  (
    n393,
    n241,
    n153,
    n159,
    n7
  );


  and
  g448
  (
    n478,
    n107,
    n285,
    n129,
    n148
  );


  and
  g449
  (
    n336,
    n319,
    n272,
    n122,
    n233
  );


  nor
  g450
  (
    n443,
    n251,
    n174,
    n115,
    n213
  );


  xor
  g451
  (
    n500,
    n162,
    n267,
    n103,
    n301
  );


  xnor
  g452
  (
    n374,
    n215,
    n227,
    n320,
    n143
  );


  and
  g453
  (
    n529,
    n184,
    n255,
    n182,
    n173
  );


  xnor
  g454
  (
    n531,
    n297,
    n163,
    n282,
    n175
  );


  or
  g455
  (
    n434,
    n287,
    n318,
    n281,
    n120
  );


  nand
  g456
  (
    n522,
    n202,
    n16,
    n149,
    n148
  );


  nand
  g457
  (
    n367,
    n158,
    n189,
    n181,
    n311
  );


  nor
  g458
  (
    n474,
    n135,
    n316,
    n115,
    n137
  );


  xor
  g459
  (
    n493,
    n188,
    n312,
    n176,
    n139
  );


  nand
  g460
  (
    n545,
    n170,
    n200,
    n206,
    n22
  );


  and
  g461
  (
    n454,
    n303,
    n261,
    n293,
    n319
  );


  nand
  g462
  (
    n347,
    n163,
    n280,
    n275,
    n248
  );


  nor
  g463
  (
    n418,
    n191,
    n160,
    n185
  );


  xor
  g464
  (
    n366,
    n288,
    n246,
    n126,
    n125
  );


  xor
  g465
  (
    n411,
    n128,
    n284,
    n109,
    n134
  );


  xor
  g466
  (
    n404,
    n270,
    n282,
    n302,
    n141
  );


  xnor
  g467
  (
    n473,
    n109,
    n171,
    n295,
    n254
  );


  or
  g468
  (
    n355,
    n242,
    n221,
    n171,
    n266
  );


  and
  g469
  (
    n519,
    n308,
    n317,
    n245,
    n150
  );


  nand
  g470
  (
    n525,
    n230,
    n295,
    n229,
    n109
  );


  nand
  g471
  (
    n485,
    n149,
    n178,
    n137,
    n285
  );


  nor
  g472
  (
    n402,
    n310,
    n154,
    n263,
    n18
  );


  and
  g473
  (
    n534,
    n133,
    n23,
    n201,
    n165
  );


  nand
  g474
  (
    n328,
    n24,
    n268,
    n253,
    n187
  );


  and
  g475
  (
    n421,
    n315,
    n307,
    n262,
    n122
  );


  or
  g476
  (
    n387,
    n165,
    n265,
    n211,
    n164
  );


  and
  g477
  (
    n446,
    n166,
    n233,
    n127,
    n242
  );


  and
  g478
  (
    n399,
    n292,
    n278,
    n246,
    n179
  );


  xor
  g479
  (
    n381,
    n249,
    n148,
    n177,
    n193
  );


  and
  g480
  (
    n548,
    n304,
    n125,
    n122,
    n147
  );


  nor
  g481
  (
    n375,
    n108,
    n221,
    n247,
    n194
  );


  xor
  g482
  (
    n523,
    n287,
    n277,
    n157,
    n149
  );


  nor
  g483
  (
    n398,
    n261,
    n305,
    n15,
    n302
  );


  xor
  g484
  (
    n477,
    n255,
    n247,
    n207,
    n282
  );


  nand
  g485
  (
    n487,
    n116,
    n119,
    n277,
    n20
  );


  xor
  g486
  (
    n551,
    n167,
    n293,
    n111,
    n190
  );


  or
  g487
  (
    n358,
    n19,
    n186,
    n136,
    n152
  );


  nand
  g488
  (
    n494,
    n278,
    n15,
    n203,
    n179
  );


  xnor
  g489
  (
    n547,
    n227,
    n308,
    n256,
    n116
  );


  nand
  g490
  (
    n524,
    n138,
    n268,
    n245,
    n263
  );


  and
  g491
  (
    n472,
    n244,
    n201,
    n182,
    n286
  );


  nand
  g492
  (
    n388,
    n124,
    n276,
    n146,
    n104
  );


  xnor
  g493
  (
    n466,
    n308,
    n123,
    n225,
    n306
  );


  and
  g494
  (
    n362,
    n229,
    n285,
    n287,
    n162
  );


  or
  g495
  (
    n538,
    n198,
    n246,
    n110,
    n265
  );


  or
  g496
  (
    n437,
    n281,
    n317,
    n250,
    n25
  );


  nand
  g497
  (
    n408,
    n182,
    n217,
    n166,
    n262
  );


  xor
  g498
  (
    n338,
    n313,
    n218,
    n180,
    n255
  );


  or
  g499
  (
    n409,
    n226,
    n266,
    n105,
    n129
  );


  and
  g500
  (
    n542,
    n280,
    n126,
    n141,
    n164
  );


  nand
  g501
  (
    n417,
    n252,
    n218,
    n153,
    n106
  );


  nand
  g502
  (
    n416,
    n274,
    n154,
    n324,
    n151
  );


  or
  g503
  (
    n508,
    n207,
    n318,
    n312,
    n309
  );


  and
  g504
  (
    n370,
    n192,
    n191,
    n198,
    n210
  );


  xor
  g505
  (
    n504,
    n191,
    n307,
    n114,
    n281
  );


  nor
  g506
  (
    n462,
    n272,
    n294,
    n102,
    n13
  );


  nand
  g507
  (
    n445,
    n181,
    n111,
    n189,
    n162
  );


  or
  g508
  (
    n457,
    n206,
    n236,
    n303,
    n222
  );


  nand
  g509
  (
    n492,
    n262,
    n289,
    n175,
    n283
  );


  nand
  g510
  (
    n556,
    n298,
    n138,
    n153,
    n257
  );


  and
  g511
  (
    n378,
    n283,
    n133,
    n193,
    n303
  );


  nor
  g512
  (
    n337,
    n219,
    n177,
    n172,
    n136
  );


  nand
  g513
  (
    n541,
    n212,
    n325,
    n324,
    n17
  );


  or
  g514
  (
    n479,
    n195,
    n197,
    n297,
    n217
  );


  nand
  g515
  (
    n430,
    n24,
    n107,
    n264,
    n198
  );


  and
  g516
  (
    n334,
    n245,
    n188,
    n154,
    n119
  );


  xnor
  g517
  (
    n557,
    n13,
    n282,
    n123,
    n302
  );


  or
  g518
  (
    n441,
    n176,
    n25,
    n325,
    n104
  );


  or
  g519
  (
    n432,
    n12,
    n274,
    n187,
    n228
  );


  xnor
  g520
  (
    n496,
    n123,
    n207,
    n298,
    n306
  );


  or
  g521
  (
    n497,
    n152,
    n232,
    n224,
    n223
  );


  and
  g522
  (
    n413,
    n21,
    n311,
    n320,
    n185
  );


  nand
  g523
  (
    n461,
    n239,
    n295,
    n231,
    n192
  );


  or
  g524
  (
    n458,
    n209,
    n228,
    n322,
    n269
  );


  or
  g525
  (
    n392,
    n199,
    n157,
    n22,
    n173
  );


  xor
  g526
  (
    n521,
    n138,
    n291,
    n26,
    n283
  );


  nor
  g527
  (
    n390,
    n16,
    n192,
    n173,
    n273
  );


  and
  g528
  (
    n368,
    n127,
    n217,
    n299,
    n287
  );


  xor
  g529
  (
    n469,
    n314,
    n315,
    n114,
    n110
  );


  nor
  g530
  (
    n345,
    n229,
    n215,
    n275,
    n159
  );


  xor
  g531
  (
    n363,
    n118,
    n259,
    n313,
    n121
  );


  xor
  g532
  (
    n546,
    n200,
    n216,
    n145,
    n204
  );


  nand
  g533
  (
    n332,
    n291,
    n265,
    n178,
    n196
  );


  or
  g534
  (
    n401,
    n145,
    n146,
    n194,
    n173
  );


  nand
  g535
  (
    n579,
    n472,
    n531,
    n509,
    n384
  );


  or
  g536
  (
    n603,
    n502,
    n539,
    n420,
    n375
  );


  xnor
  g537
  (
    n636,
    n424,
    n413,
    n529,
    n549
  );


  or
  g538
  (
    n596,
    n338,
    n426,
    n471,
    n329
  );


  or
  g539
  (
    n631,
    n512,
    n527,
    n507,
    n558
  );


  xor
  g540
  (
    n627,
    n538,
    n414,
    n508,
    n493
  );


  xnor
  g541
  (
    n598,
    n487,
    n345,
    n343,
    n434
  );


  nand
  g542
  (
    n615,
    n418,
    n530,
    n524,
    n455
  );


  nand
  g543
  (
    n641,
    n494,
    n503,
    n463,
    n428
  );


  xnor
  g544
  (
    n614,
    n510,
    n543,
    n466,
    n534
  );


  xnor
  g545
  (
    n640,
    n515,
    n429,
    n482,
    n404
  );


  xnor
  g546
  (
    n570,
    n533,
    n450,
    n496,
    n556
  );


  and
  g547
  (
    n578,
    n532,
    n493,
    n469,
    n399
  );


  and
  g548
  (
    n650,
    n395,
    n555,
    n553,
    n519
  );


  and
  g549
  (
    n593,
    n503,
    n537,
    n550,
    n505
  );


  xor
  g550
  (
    n567,
    n389,
    n385,
    n355,
    n349
  );


  xnor
  g551
  (
    n583,
    n545,
    n487,
    n341,
    n353
  );


  nor
  g552
  (
    n604,
    n439,
    n543,
    n541,
    n528
  );


  nand
  g553
  (
    n656,
    n359,
    n407,
    n517,
    n508
  );


  xnor
  g554
  (
    n613,
    n509,
    n430,
    n523,
    n484
  );


  nor
  g555
  (
    n625,
    n363,
    n396,
    n342,
    n528
  );


  nand
  g556
  (
    n584,
    n511,
    n531,
    n410,
    n422
  );


  and
  g557
  (
    n587,
    n554,
    n480,
    n490,
    n541
  );


  and
  g558
  (
    n623,
    n401,
    n516,
    n548,
    n361
  );


  or
  g559
  (
    n621,
    n348,
    n415,
    n505,
    n529
  );


  and
  g560
  (
    n564,
    n556,
    n552,
    n505,
    n512
  );


  and
  g561
  (
    n626,
    n339,
    n398,
    n440,
    n506
  );


  or
  g562
  (
    n600,
    n539,
    n477,
    n392,
    n465
  );


  xnor
  g563
  (
    n606,
    n532,
    n421,
    n518,
    n484
  );


  nor
  g564
  (
    n590,
    n336,
    n524,
    n540,
    n344
  );


  nand
  g565
  (
    n576,
    n535,
    n545,
    n551,
    n508
  );


  xnor
  g566
  (
    n569,
    n543,
    n379,
    n391,
    n491
  );


  nand
  g567
  (
    n639,
    n436,
    n451,
    n548,
    n496
  );


  nand
  g568
  (
    n643,
    n519,
    n527,
    n518,
    n490
  );


  xnor
  g569
  (
    n586,
    n542,
    n527,
    n524,
    n529
  );


  or
  g570
  (
    n646,
    n347,
    n494,
    n521,
    n383
  );


  xnor
  g571
  (
    n616,
    n444,
    n522,
    n544,
    n454
  );


  nor
  g572
  (
    n580,
    n335,
    n427,
    n513,
    n538
  );


  or
  g573
  (
    n565,
    n352,
    n515,
    n507,
    n523
  );


  xor
  g574
  (
    n568,
    n354,
    n498,
    n333,
    n551
  );


  and
  g575
  (
    n605,
    n425,
    n489,
    n546,
    n364
  );


  or
  g576
  (
    n599,
    n417,
    n449,
    n534,
    n510
  );


  and
  g577
  (
    n572,
    n558,
    n460,
    n467,
    n539
  );


  xnor
  g578
  (
    n630,
    n525,
    n554,
    n388,
    n517
  );


  nor
  g579
  (
    n617,
    n537,
    n549,
    n356,
    n409
  );


  nand
  g580
  (
    n581,
    n523,
    n431,
    n390,
    n433
  );


  xor
  g581
  (
    n562,
    n546,
    n374,
    n495,
    n514
  );


  xnor
  g582
  (
    n655,
    n488,
    n488,
    n491,
    n357
  );


  nor
  g583
  (
    n594,
    n500,
    n492,
    n497,
    n452
  );


  xor
  g584
  (
    n585,
    n481,
    n369,
    n559,
    n526
  );


  xor
  g585
  (
    n644,
    n559,
    n506,
    n435,
    n496
  );


  xnor
  g586
  (
    n628,
    n499,
    n470,
    n473,
    n497
  );


  nor
  g587
  (
    n622,
    n461,
    n547,
    n346,
    n553
  );


  nor
  g588
  (
    n635,
    n526,
    n546,
    n397,
    n511
  );


  and
  g589
  (
    n652,
    n557,
    n555,
    n537,
    n513
  );


  or
  g590
  (
    n642,
    n504,
    n506,
    n520,
    n402
  );


  xor
  g591
  (
    n591,
    n445,
    n540,
    n504,
    n503
  );


  or
  g592
  (
    n649,
    n544,
    n378,
    n525,
    n334
  );


  and
  g593
  (
    n573,
    n525,
    n493,
    n533,
    n328
  );


  xor
  g594
  (
    n629,
    n373,
    n331,
    n540,
    n547
  );


  xnor
  g595
  (
    n637,
    n530,
    n501,
    n536,
    n498
  );


  nor
  g596
  (
    n648,
    n559,
    n536,
    n483,
    n553
  );


  nand
  g597
  (
    n608,
    n462,
    n550,
    n557,
    n432
  );


  nand
  g598
  (
    n647,
    n327,
    n561,
    n535,
    n441
  );


  and
  g599
  (
    n620,
    n468,
    n548,
    n517,
    n535
  );


  xnor
  g600
  (
    n597,
    n408,
    n446,
    n400,
    n519
  );


  or
  g601
  (
    n588,
    n486,
    n521,
    n511,
    n382
  );


  xnor
  g602
  (
    n624,
    n476,
    n513,
    n492,
    n475
  );


  nand
  g603
  (
    n634,
    n515,
    n499,
    n550,
    n542
  );


  xor
  g604
  (
    n651,
    n367,
    n365,
    n340,
    n501
  );


  nand
  g605
  (
    n595,
    n560,
    n453,
    n478,
    n504
  );


  xor
  g606
  (
    n566,
    n495,
    n360,
    n510,
    n386
  );


  xor
  g607
  (
    n645,
    n330,
    n370,
    n512,
    n557
  );


  xnor
  g608
  (
    n611,
    n549,
    n380,
    n405,
    n497
  );


  nor
  g609
  (
    n589,
    n531,
    n558,
    n556,
    n544
  );


  xnor
  g610
  (
    n563,
    n474,
    n561,
    n536,
    n458
  );


  xnor
  g611
  (
    n609,
    n520,
    n552,
    n371,
    n416
  );


  nand
  g612
  (
    n618,
    n507,
    n522,
    n545,
    n528
  );


  xnor
  g613
  (
    n607,
    n555,
    n526,
    n394,
    n552
  );


  nor
  g614
  (
    n601,
    n447,
    n560,
    n443,
    n479
  );


  xor
  g615
  (
    n575,
    n448,
    n489,
    n514,
    n498
  );


  nor
  g616
  (
    n633,
    n495,
    n381,
    n500,
    n502
  );


  nor
  g617
  (
    n577,
    n456,
    n492,
    n368,
    n442
  );


  and
  g618
  (
    n582,
    n332,
    n403,
    n494,
    n423
  );


  nand
  g619
  (
    n632,
    n518,
    n534,
    n551,
    n366
  );


  xnor
  g620
  (
    n619,
    n521,
    n326,
    n485,
    n530
  );


  xor
  g621
  (
    n657,
    n522,
    n560,
    n502,
    n538
  );


  xnor
  g622
  (
    n592,
    n358,
    n376,
    n509,
    n499
  );


  and
  g623
  (
    n571,
    n541,
    n516,
    n459,
    n520
  );


  or
  g624
  (
    n653,
    n412,
    n554,
    n457,
    n393
  );


  or
  g625
  (
    n612,
    n406,
    n438,
    n514,
    n411
  );


  xnor
  g626
  (
    n602,
    n387,
    n437,
    n362,
    n372
  );


  xnor
  g627
  (
    n654,
    n464,
    n419,
    n542,
    n547
  );


  xor
  g628
  (
    n610,
    n377,
    n337,
    n486,
    n485
  );


  nor
  g629
  (
    n574,
    n351,
    n532,
    n516,
    n501
  );


  nor
  g630
  (
    n638,
    n561,
    n500,
    n533,
    n350
  );


  nor
  g631
  (
    n681,
    n630,
    n648,
    n612,
    n640
  );


  or
  g632
  (
    n678,
    n590,
    n597,
    n592,
    n609
  );


  nand
  g633
  (
    n666,
    n654,
    n655,
    n633,
    n573
  );


  xnor
  g634
  (
    n667,
    n582,
    n577,
    n619,
    n599
  );


  and
  g635
  (
    n677,
    n626,
    n644,
    n580,
    n584
  );


  xor
  g636
  (
    n659,
    n574,
    n638,
    n576,
    n623
  );


  nor
  g637
  (
    n672,
    n646,
    n610,
    n650,
    n589
  );


  xor
  g638
  (
    n675,
    n656,
    n642,
    n570,
    n616
  );


  xnor
  g639
  (
    n673,
    n594,
    n637,
    n635,
    n583
  );


  or
  g640
  (
    n671,
    n604,
    n613,
    n563,
    n566
  );


  and
  g641
  (
    n668,
    n617,
    n595,
    n602,
    n657
  );


  nand
  g642
  (
    n662,
    n634,
    n627,
    n628,
    n629
  );


  or
  g643
  (
    n679,
    n631,
    n575,
    n622,
    n649
  );


  nor
  g644
  (
    n663,
    n586,
    n632,
    n591,
    n601
  );


  nand
  g645
  (
    n669,
    n614,
    n621,
    n588,
    n620
  );


  xor
  g646
  (
    n658,
    n568,
    n579,
    n569,
    n652
  );


  nand
  g647
  (
    n664,
    n567,
    n643,
    n600,
    n618
  );


  nand
  g648
  (
    n670,
    n607,
    n651,
    n605,
    n571
  );


  nand
  g649
  (
    n665,
    n598,
    n585,
    n603,
    n564
  );


  nand
  g650
  (
    n680,
    n639,
    n593,
    n578,
    n606
  );


  xnor
  g651
  (
    n660,
    n641,
    n647,
    n596,
    n562
  );


  nor
  g652
  (
    AntiSAT_key_wire,
    n565,
    n653,
    n572,
    n636
  );


  xor
  g653
  (
    n674,
    n645,
    n611,
    n624,
    n587
  );


  nor
  g654
  (
    n661,
    n608,
    n581,
    n615,
    n625
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_0,
    keyIn_0_26,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_1,
    keyIn_0_27,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_2,
    keyIn_0_28,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_3,
    keyIn_0_29,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_4,
    keyIn_0_30,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_5,
    keyIn_0_31,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_6,
    keyIn_0_32,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_7,
    keyIn_0_33,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_8,
    keyIn_0_34,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_9,
    keyIn_0_35,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_10,
    keyIn_0_36,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_11,
    keyIn_0_37,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_12,
    keyIn_0_38,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_13,
    keyIn_0_39,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_14,
    keyIn_0_40,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_15,
    keyIn_0_41,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_16,
    keyIn_0_42,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_17,
    keyIn_0_43,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_18,
    keyIn_0_44,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_19,
    keyIn_0_45,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_20,
    keyIn_0_46,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_21,
    keyIn_0_47,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_22,
    keyIn_0_48,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_23,
    keyIn_0_49,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_24,
    keyIn_0_50,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_25,
    keyIn_0_51,
    n26
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n676,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

