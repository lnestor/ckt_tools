

module Stat_100_56
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  nCHANGED,
  n105,
  n120,
  n101,
  n102,
  n104,
  n117,
  n122,
  n116,
  n123,
  n108,
  n99,
  n97,
  n121,
  n115,
  n95,
  n93,
  n107,
  n118,
  n98,
  n113,
  n106,
  n96,
  n109,
  n112,
  n114,
  n100,
  n128,
  n129,
  n130,
  n132,
  n131
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output nCHANGED;output n105;output n120;output n101;output n102;output n104;output n117;output n122;output n116;output n123;output n108;output n99;output n97;output n121;output n115;output n95;output n93;output n107;output n118;output n98;output n113;output n106;output n96;output n109;output n112;output n114;output n100;output n128;output n129;output n130;output n132;output n131;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n94;wire n103;wire n110;wire n111;wire n119;wire n124;wire n125;wire n126;wire n127;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    n52,
    n20
  );


  not
  g1
  (
    KeyWire_0_52,
    n28
  );


  not
  g2
  (
    KeyWire_0_30,
    n19
  );


  not
  g3
  (
    n60,
    n19
  );


  not
  g4
  (
    KeyWire_0_31,
    n12
  );


  not
  g5
  (
    n42,
    n18
  );


  buf
  g6
  (
    KeyWire_0_34,
    n25
  );


  not
  g7
  (
    KeyWire_0_48,
    n28
  );


  not
  g8
  (
    KeyWire_0_47,
    n25
  );


  not
  g9
  (
    n34,
    n17
  );


  buf
  g10
  (
    KeyWire_0_32,
    n6
  );


  buf
  g11
  (
    KeyWire_0_4,
    n22
  );


  not
  g12
  (
    n54,
    n23
  );


  not
  g13
  (
    KeyWire_0_29,
    n22
  );


  not
  g14
  (
    KeyWire_0_27,
    n16
  );


  not
  g15
  (
    n58,
    n20
  );


  not
  g16
  (
    KeyWire_0_11,
    n23
  );


  buf
  g17
  (
    KeyWire_0_26,
    n3
  );


  buf
  g18
  (
    KeyWire_0_33,
    n25
  );


  not
  g19
  (
    n33,
    n27
  );


  buf
  g20
  (
    KeyWire_0_8,
    n7
  );


  buf
  g21
  (
    KeyWire_0_10,
    n2
  );


  not
  g22
  (
    n63,
    n26
  );


  buf
  g23
  (
    KeyWire_0_23,
    n24
  );


  not
  g24
  (
    KeyWire_0_36,
    n13
  );


  not
  g25
  (
    KeyWire_0_44,
    n15
  );


  buf
  g26
  (
    KeyWire_0_1,
    n11
  );


  buf
  g27
  (
    n70,
    n22
  );


  buf
  g28
  (
    n48,
    n24
  );


  not
  g29
  (
    n37,
    n26
  );


  buf
  g30
  (
    KeyWire_0_42,
    n27
  );


  buf
  g31
  (
    n65,
    n24
  );


  buf
  g32
  (
    KeyWire_0_62,
    n18
  );


  buf
  g33
  (
    n41,
    n21
  );


  buf
  g34
  (
    n82,
    n21
  );


  buf
  g35
  (
    KeyWire_0_28,
    n4
  );


  buf
  g36
  (
    KeyWire_0_39,
    n9
  );


  not
  g37
  (
    KeyWire_0_43,
    n20
  );


  buf
  g38
  (
    KeyWire_0_19,
    n27
  );


  buf
  g39
  (
    n75,
    n21
  );


  not
  g40
  (
    KeyWire_0_22,
    n19
  );


  buf
  g41
  (
    KeyWire_0_0,
    n14
  );


  buf
  g42
  (
    KeyWire_0_7,
    n29
  );


  buf
  g43
  (
    n77,
    n10
  );


  buf
  g44
  (
    KeyWire_0_56,
    n29
  );


  buf
  g45
  (
    n62,
    n28
  );


  not
  g46
  (
    n53,
    n23
  );


  not
  g47
  (
    n73,
    n1
  );


  not
  g48
  (
    n45,
    n5
  );


  buf
  g49
  (
    KeyWire_0_49,
    n8
  );


  not
  g50
  (
    KeyWire_0_61,
    n26
  );


  not
  g51
  (
    KeyWire_0_9,
    n18
  );


  buf
  g52
  (
    n85,
    n35
  );


  buf
  g53
  (
    KeyWire_0_60,
    n34
  );


  not
  g54
  (
    n86,
    n36
  );


  buf
  g55
  (
    n87,
    n37
  );


  not
  g56
  (
    KeyWire_0_53,
    n33
  );


  buf
  g57
  (
    KeyWire_0_18,
    n38
  );


  not
  g58
  (
    n92,
    n39
  );


  buf
  g59
  (
    KeyWire_0_15,
    n40
  );


  xor
  g60
  (
    n121,
    n68,
    n82,
    n74,
    n85
  );


  nor
  g61
  (
    KeyWire_0_3,
    n57,
    n84,
    n75,
    n59
  );


  nor
  g62
  (
    n117,
    n75,
    n88,
    n83,
    n42
  );


  and
  g63
  (
    KeyWire_0_35,
    n86,
    n56,
    n46,
    n71
  );


  xor
  g64
  (
    KeyWire_0_51,
    n63,
    n86,
    n91,
    n62
  );


  nor
  g65
  (
    KeyWire_0_17,
    n73,
    n79,
    n67
  );


  xnor
  g66
  (
    KeyWire_0_38,
    n82,
    n83,
    n89,
    n81
  );


  nand
  g67
  (
    KeyWire_0_13,
    n90,
    n85,
    n92,
    n78
  );


  nand
  g68
  (
    KeyWire_0_46,
    n67,
    n70,
    n87,
    n78
  );


  xnor
  g69
  (
    KeyWire_0_40,
    n74,
    n84,
    n77,
    n91
  );


  or
  g70
  (
    KeyWire_0_21,
    n76,
    n61,
    n73,
    n79
  );


  xor
  g71
  (
    KeyWire_0_54,
    n53,
    n92,
    n65,
    n89
  );


  nand
  g72
  (
    KeyWire_0_57,
    n80,
    n72,
    n63
  );


  nand
  g73
  (
    KeyWire_0_55,
    n77,
    n69
  );


  nand
  g74
  (
    KeyWire_0_58,
    n75,
    n91,
    n86,
    n48
  );


  and
  g75
  (
    KeyWire_0_2,
    n89,
    n71,
    n77,
    n52
  );


  and
  g76
  (
    KeyWire_0_20,
    n91,
    n85,
    n54,
    n60
  );


  nand
  g77
  (
    KeyWire_0_24,
    n62,
    n61,
    n87
  );


  xnor
  g78
  (
    KeyWire_0_50,
    n71,
    n59,
    n50,
    n58
  );


  nor
  g79
  (
    n96,
    n72,
    n79,
    n51,
    n88
  );


  nor
  g80
  (
    n103,
    n65,
    n70,
    n76,
    n49
  );


  xnor
  g81
  (
    KeyWire_0_41,
    n84,
    n90,
    n62,
    n80
  );


  or
  g82
  (
    n118,
    n45,
    n66,
    n64,
    n90
  );


  nor
  g83
  (
    KeyWire_0_14,
    n66,
    n41,
    n47,
    n78
  );


  nor
  g84
  (
    KeyWire_0_45,
    n60,
    n43,
    n87,
    n89
  );


  and
  g85
  (
    KeyWire_0_37,
    n90,
    n61,
    n64,
    n83
  );


  or
  g86
  (
    KeyWire_0_59,
    n68,
    n55,
    n81,
    n72
  );


  or
  g87
  (
    KeyWire_0_6,
    n92,
    n73,
    n74,
    n85
  );


  xor
  g88
  (
    n115,
    n76,
    n82,
    n60,
    n59
  );


  or
  g89
  (
    KeyWire_0_16,
    n64,
    n70,
    n68,
    n80
  );


  xor
  g90
  (
    KeyWire_0_25,
    n44,
    n92,
    n86,
    n88
  );


  xnor
  g91
  (
    n120,
    n81,
    n66,
    n65,
    n88
  );


  not
  g92
  (
    n127,
    n121
  );


  not
  g93
  (
    KeyWire_0_12,
    n120
  );


  not
  g94
  (
    KeyWire_0_5,
    n119
  );


  xnor
  g95
  (
    n128,
    n123,
    n122,
    n127,
    n30
  );


  and
  g96
  (
    n131,
    n126,
    n29,
    n31
  );


  nor
  g97
  (
    n130,
    n125,
    n126,
    n30
  );


  nand
  g98
  (
    n129,
    n124,
    n32
  );


  and
  g99
  (
    KeyWire_0_63,
    n31,
    n127,
    n126
  );


  buf
  g100
  (
    nCHANGED,
    n10
  );


  xnor
  KeyGate_0_0
  (
    n43,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n66,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n116,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n104,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n35,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n125,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n119,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n84,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n46,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n50,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n67,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n80,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n126,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n111,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n95,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n91,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n93,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n107,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n89,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n74,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n124,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n122,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n38,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n56,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n94,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n106,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n51,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n69,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n61,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n81,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n36,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n64,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n47,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n59,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n44,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n99,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n78,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n100,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n110,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n49,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n108,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n97,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n72,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n83,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n40,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n102,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n113,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n68,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n71,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n39,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n101,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n98,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n76,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n90,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n112,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n123,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n79,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n105,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n109,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n114,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n88,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n55,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n57,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n132,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


