

module Stat_2000_204
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n401,
  n788,
  n758,
  n763,
  n796,
  n760,
  n795,
  n783,
  n779,
  n761,
  n771,
  n787,
  n764,
  n798,
  n767,
  n765,
  n791,
  n1288,
  n2023,
  n2020,
  n2027,
  n2032,
  n2031,
  n2028,
  n2019,
  n2029,
  n2022,
  n2030,
  n2024,
  n2021,
  n2026,
  n2025
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n401;output n788;output n758;output n763;output n796;output n760;output n795;output n783;output n779;output n761;output n771;output n787;output n764;output n798;output n767;output n765;output n791;output n1288;output n2023;output n2020;output n2027;output n2032;output n2031;output n2028;output n2019;output n2029;output n2022;output n2030;output n2024;output n2021;output n2026;output n2025;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n759;wire n762;wire n766;wire n768;wire n769;wire n770;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n780;wire n781;wire n782;wire n784;wire n785;wire n786;wire n789;wire n790;wire n792;wire n793;wire n794;wire n797;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    n69,
    n22
  );


  not
  g1
  (
    KeyWire_0_12,
    n15
  );


  not
  g2
  (
    n101,
    n29
  );


  not
  g3
  (
    n144,
    n25
  );


  buf
  g4
  (
    n55,
    n14
  );


  not
  g5
  (
    n65,
    n9
  );


  buf
  g6
  (
    n135,
    n12
  );


  buf
  g7
  (
    n136,
    n5
  );


  not
  g8
  (
    n59,
    n16
  );


  not
  g9
  (
    n109,
    n8
  );


  not
  g10
  (
    n130,
    n14
  );


  not
  g11
  (
    n71,
    n17
  );


  buf
  g12
  (
    n94,
    n20
  );


  buf
  g13
  (
    n60,
    n1
  );


  not
  g14
  (
    n97,
    n24
  );


  not
  g15
  (
    n99,
    n22
  );


  buf
  g16
  (
    n124,
    n28
  );


  not
  g17
  (
    n98,
    n10
  );


  not
  g18
  (
    n146,
    n3
  );


  buf
  g19
  (
    n41,
    n21
  );


  buf
  g20
  (
    n148,
    n25
  );


  not
  g21
  (
    n64,
    n11
  );


  buf
  g22
  (
    n77,
    n7
  );


  not
  g23
  (
    n139,
    n9
  );


  not
  g24
  (
    n68,
    n18
  );


  buf
  g25
  (
    n145,
    n23
  );


  not
  g26
  (
    n104,
    n6
  );


  buf
  g27
  (
    n83,
    n16
  );


  not
  g28
  (
    n47,
    n20
  );


  buf
  g29
  (
    n103,
    n19
  );


  buf
  g30
  (
    n96,
    n26
  );


  not
  g31
  (
    n108,
    n26
  );


  not
  g32
  (
    n56,
    n19
  );


  not
  g33
  (
    n50,
    n10
  );


  buf
  g34
  (
    n53,
    n2
  );


  not
  g35
  (
    n63,
    n5
  );


  buf
  g36
  (
    n76,
    n1
  );


  buf
  g37
  (
    n79,
    n15
  );


  buf
  g38
  (
    n52,
    n3
  );


  not
  g39
  (
    n46,
    n9
  );


  not
  g40
  (
    n92,
    n18
  );


  buf
  g41
  (
    n116,
    n5
  );


  buf
  g42
  (
    n80,
    n27
  );


  not
  g43
  (
    n82,
    n9
  );


  not
  g44
  (
    n62,
    n22
  );


  not
  g45
  (
    n102,
    n23
  );


  not
  g46
  (
    n72,
    n20
  );


  buf
  g47
  (
    n114,
    n4
  );


  not
  g48
  (
    n143,
    n24
  );


  not
  g49
  (
    n87,
    n30
  );


  buf
  g50
  (
    n89,
    n19
  );


  buf
  g51
  (
    n127,
    n11
  );


  not
  g52
  (
    n118,
    n11
  );


  not
  g53
  (
    n58,
    n13
  );


  buf
  g54
  (
    n54,
    n30
  );


  not
  g55
  (
    n73,
    n27
  );


  buf
  g56
  (
    n107,
    n21
  );


  not
  g57
  (
    n128,
    n24
  );


  buf
  g58
  (
    n141,
    n17
  );


  buf
  g59
  (
    n121,
    n7
  );


  not
  g60
  (
    n34,
    n12
  );


  not
  g61
  (
    n132,
    n22
  );


  buf
  g62
  (
    n86,
    n25
  );


  buf
  g63
  (
    n110,
    n15
  );


  not
  g64
  (
    n61,
    n31
  );


  not
  g65
  (
    n74,
    n24
  );


  not
  g66
  (
    n78,
    n29
  );


  buf
  g67
  (
    n90,
    n25
  );


  not
  g68
  (
    n93,
    n14
  );


  buf
  g69
  (
    n81,
    n8
  );


  buf
  g70
  (
    n35,
    n30
  );


  buf
  g71
  (
    n122,
    n27
  );


  buf
  g72
  (
    n112,
    n4
  );


  buf
  g73
  (
    n113,
    n14
  );


  not
  g74
  (
    n137,
    n12
  );


  not
  g75
  (
    n138,
    n18
  );


  buf
  g76
  (
    n131,
    n31
  );


  not
  g77
  (
    n51,
    n28
  );


  not
  g78
  (
    n142,
    n6
  );


  not
  g79
  (
    n95,
    n7
  );


  not
  g80
  (
    n66,
    n18
  );


  buf
  g81
  (
    n67,
    n2
  );


  not
  g82
  (
    n105,
    n13
  );


  buf
  g83
  (
    n147,
    n16
  );


  buf
  g84
  (
    n133,
    n16
  );


  buf
  g85
  (
    n37,
    n3
  );


  buf
  g86
  (
    n119,
    n4
  );


  not
  g87
  (
    KeyWire_0_33,
    n13
  );


  buf
  g88
  (
    KeyWire_0_11,
    n17
  );


  buf
  g89
  (
    n123,
    n19
  );


  buf
  g90
  (
    n115,
    n6
  );


  buf
  g91
  (
    n117,
    n26
  );


  buf
  g92
  (
    n140,
    n2
  );


  buf
  g93
  (
    n129,
    n29
  );


  not
  g94
  (
    n44,
    n13
  );


  not
  g95
  (
    n43,
    n11
  );


  buf
  g96
  (
    n36,
    n29
  );


  not
  g97
  (
    n70,
    n30
  );


  buf
  g98
  (
    n100,
    n17
  );


  buf
  g99
  (
    n42,
    n10
  );


  not
  g100
  (
    n38,
    n23
  );


  not
  g101
  (
    n125,
    n8
  );


  not
  g102
  (
    n33,
    n12
  );


  buf
  g103
  (
    n84,
    n8
  );


  not
  g104
  (
    n88,
    n21
  );


  not
  g105
  (
    n111,
    n27
  );


  not
  g106
  (
    n57,
    n15
  );


  buf
  g107
  (
    n48,
    n20
  );


  not
  g108
  (
    n106,
    n23
  );


  buf
  g109
  (
    n45,
    n31
  );


  buf
  g110
  (
    n134,
    n28
  );


  not
  g111
  (
    n85,
    n28
  );


  not
  g112
  (
    n149,
    n26
  );


  not
  g113
  (
    n75,
    n10
  );


  not
  g114
  (
    n39,
    n1
  );


  not
  g115
  (
    n120,
    n21
  );


  buf
  g116
  (
    n49,
    n7
  );


  xor
  g117
  (
    n254,
    n113,
    n87
  );


  nand
  g118
  (
    n253,
    n52,
    n68
  );


  xnor
  g119
  (
    n286,
    n127,
    n67
  );


  or
  g120
  (
    n263,
    n75,
    n89
  );


  nor
  g121
  (
    n191,
    n81,
    n36
  );


  nor
  g122
  (
    n192,
    n80,
    n148
  );


  or
  g123
  (
    n203,
    n131,
    n67
  );


  and
  g124
  (
    n228,
    n130,
    n136
  );


  buf
  g125
  (
    n256,
    n68
  );


  and
  g126
  (
    n268,
    n114,
    n94
  );


  xnor
  g127
  (
    n164,
    n116,
    n141
  );


  xnor
  g128
  (
    n187,
    n40,
    n34
  );


  nand
  g129
  (
    n311,
    n120,
    n81
  );


  nand
  g130
  (
    n283,
    n72,
    n117
  );


  nor
  g131
  (
    n237,
    n104,
    n63
  );


  xnor
  g132
  (
    n292,
    n45,
    n79
  );


  or
  g133
  (
    n333,
    n56,
    n133
  );


  xnor
  g134
  (
    n209,
    n87,
    n50
  );


  xor
  g135
  (
    n193,
    n47,
    n57
  );


  xnor
  g136
  (
    n273,
    n126,
    n74
  );


  nand
  g137
  (
    n165,
    n142,
    n97
  );


  xor
  g138
  (
    n173,
    n121,
    n41
  );


  or
  g139
  (
    n304,
    n97,
    n80
  );


  xor
  g140
  (
    n274,
    n127,
    n113
  );


  nand
  g141
  (
    n244,
    n119,
    n49
  );


  and
  g142
  (
    n294,
    n38,
    n145
  );


  and
  g143
  (
    n227,
    n44,
    n100
  );


  and
  g144
  (
    KeyWire_0_44,
    n53,
    n108
  );


  or
  g145
  (
    n305,
    n105,
    n97
  );


  nor
  g146
  (
    n277,
    n55,
    n145
  );


  nand
  g147
  (
    n151,
    n50,
    n70
  );


  nor
  g148
  (
    n177,
    n36,
    n43
  );


  nor
  g149
  (
    n334,
    n92,
    n83
  );


  nor
  g150
  (
    n276,
    n84,
    n83
  );


  or
  g151
  (
    n229,
    n111,
    n115
  );


  or
  g152
  (
    KeyWire_0_4,
    n78,
    n33
  );


  and
  g153
  (
    n196,
    n106,
    n64
  );


  xnor
  g154
  (
    n302,
    n35,
    n118
  );


  nor
  g155
  (
    n329,
    n134,
    n66
  );


  xor
  g156
  (
    n299,
    n33,
    n108
  );


  xnor
  g157
  (
    n295,
    n109,
    n54
  );


  or
  g158
  (
    n284,
    n45,
    n75
  );


  xnor
  g159
  (
    n331,
    n132,
    n137
  );


  and
  g160
  (
    n324,
    n71,
    n56
  );


  nor
  g161
  (
    n234,
    n117,
    n88
  );


  xnor
  g162
  (
    n330,
    n72,
    n93
  );


  xor
  g163
  (
    n188,
    n57,
    n99
  );


  xnor
  g164
  (
    n251,
    n143,
    n102
  );


  nor
  g165
  (
    KeyWire_0_51,
    n145,
    n102
  );


  xnor
  g166
  (
    n179,
    n112,
    n42
  );


  nor
  g167
  (
    n221,
    n136,
    n58
  );


  nor
  g168
  (
    n214,
    n75,
    n44
  );


  and
  g169
  (
    n326,
    n65,
    n102
  );


  xor
  g170
  (
    n303,
    n123,
    n77
  );


  buf
  g171
  (
    n325,
    n113
  );


  xnor
  g172
  (
    n181,
    n37,
    n133
  );


  xor
  g173
  (
    n172,
    n101,
    n97
  );


  or
  g174
  (
    n157,
    n84,
    n77
  );


  xor
  g175
  (
    n266,
    n123,
    n117
  );


  and
  g176
  (
    n150,
    n139,
    n55
  );


  xnor
  g177
  (
    n225,
    n141,
    n89
  );


  and
  g178
  (
    n242,
    n89,
    n36
  );


  xnor
  g179
  (
    n280,
    n67,
    n49
  );


  xnor
  g180
  (
    n269,
    n46,
    n147
  );


  nor
  g181
  (
    n185,
    n82,
    n112
  );


  nor
  g182
  (
    n322,
    n78,
    n133
  );


  and
  g183
  (
    n246,
    n102,
    n91
  );


  nor
  g184
  (
    n171,
    n35,
    n125
  );


  nor
  g185
  (
    n289,
    n110,
    n114
  );


  xnor
  g186
  (
    n211,
    n86,
    n71
  );


  xor
  g187
  (
    n261,
    n125,
    n105
  );


  xnor
  g188
  (
    n167,
    n37,
    n79
  );


  xnor
  g189
  (
    n252,
    n42,
    n138
  );


  and
  g190
  (
    n265,
    n103,
    n73
  );


  or
  g191
  (
    n160,
    n147,
    n121
  );


  and
  g192
  (
    n314,
    n143,
    n94
  );


  nor
  g193
  (
    n190,
    n74,
    n135
  );


  or
  g194
  (
    n180,
    n108,
    n91
  );


  xor
  g195
  (
    n220,
    n115,
    n88
  );


  nor
  g196
  (
    n236,
    n121,
    n92
  );


  xor
  g197
  (
    n258,
    n124,
    n96
  );


  xnor
  g198
  (
    n176,
    n138,
    n95
  );


  and
  g199
  (
    n257,
    n147,
    n85
  );


  and
  g200
  (
    n158,
    n145,
    n127
  );


  nor
  g201
  (
    n279,
    n128,
    n40
  );


  and
  g202
  (
    n186,
    n87,
    n136
  );


  nand
  g203
  (
    n247,
    n107,
    n100
  );


  nor
  g204
  (
    n243,
    n109,
    n42
  );


  xor
  g205
  (
    KeyWire_0_10,
    n40,
    n57
  );


  nand
  g206
  (
    n204,
    n149,
    n66
  );


  xnor
  g207
  (
    n259,
    n93,
    n84
  );


  nor
  g208
  (
    n208,
    n76,
    n73
  );


  nand
  g209
  (
    n332,
    n140,
    n139
  );


  nand
  g210
  (
    n278,
    n33,
    n76
  );


  nor
  g211
  (
    n189,
    n116,
    n92
  );


  or
  g212
  (
    n307,
    n57,
    n107
  );


  xnor
  g213
  (
    n308,
    n46,
    n86
  );


  nor
  g214
  (
    n178,
    n38,
    n90
  );


  xor
  g215
  (
    n312,
    n69,
    n68
  );


  and
  g216
  (
    n210,
    n142,
    n91
  );


  nand
  g217
  (
    n238,
    n80,
    n46
  );


  xor
  g218
  (
    n301,
    n134,
    n148
  );


  xnor
  g219
  (
    n161,
    n79,
    n114
  );


  nor
  g220
  (
    n262,
    n111,
    n87
  );


  xnor
  g221
  (
    n300,
    n140,
    n74
  );


  or
  g222
  (
    n313,
    n48,
    n118
  );


  and
  g223
  (
    n288,
    n135,
    n78
  );


  and
  g224
  (
    n282,
    n126,
    n148
  );


  nor
  g225
  (
    n213,
    n83,
    n88
  );


  nand
  g226
  (
    n182,
    n46,
    n90
  );


  nand
  g227
  (
    n152,
    n128,
    n122
  );


  xor
  g228
  (
    n169,
    n60,
    n82
  );


  and
  g229
  (
    n249,
    n141,
    n144
  );


  or
  g230
  (
    n223,
    n48,
    n76
  );


  xor
  g231
  (
    n216,
    n103,
    n105
  );


  or
  g232
  (
    n154,
    n115,
    n80
  );


  xor
  g233
  (
    n200,
    n62,
    n43
  );


  nor
  g234
  (
    n195,
    n146,
    n100
  );


  or
  g235
  (
    n297,
    n146,
    n117
  );


  nand
  g236
  (
    KeyWire_0_62,
    n60,
    n48
  );


  nand
  g237
  (
    n335,
    n118,
    n37
  );


  xnor
  g238
  (
    n235,
    n55,
    n65
  );


  xor
  g239
  (
    n202,
    n47,
    n112
  );


  nand
  g240
  (
    n260,
    n53,
    n81
  );


  xor
  g241
  (
    n270,
    n63,
    n143
  );


  nand
  g242
  (
    n281,
    n51,
    n137
  );


  and
  g243
  (
    n217,
    n64,
    n39
  );


  nand
  g244
  (
    n318,
    n106,
    n99
  );


  xor
  g245
  (
    n184,
    n119,
    n56
  );


  nand
  g246
  (
    n175,
    n58,
    n66
  );


  xor
  g247
  (
    n287,
    n139,
    n82
  );


  xor
  g248
  (
    n309,
    n38,
    n131
  );


  or
  g249
  (
    n298,
    n78,
    n55
  );


  nor
  g250
  (
    n290,
    n89,
    n34
  );


  nor
  g251
  (
    n255,
    n141,
    n115
  );


  or
  g252
  (
    n316,
    n48,
    n54
  );


  xor
  g253
  (
    n219,
    n138,
    n85
  );


  or
  g254
  (
    n275,
    n129,
    n109
  );


  and
  g255
  (
    n317,
    n122,
    n111,
    n86
  );


  and
  g256
  (
    n215,
    n61,
    n111,
    n101,
    n66
  );


  xor
  g257
  (
    n230,
    n126,
    n60,
    n129,
    n149
  );


  xor
  g258
  (
    n201,
    n130,
    n40,
    n79,
    n54
  );


  xor
  g259
  (
    n328,
    n72,
    n124,
    n47,
    n130
  );


  or
  g260
  (
    n207,
    n45,
    n103,
    n104
  );


  xor
  g261
  (
    n264,
    n104,
    n77,
    n98,
    n51
  );


  or
  g262
  (
    n224,
    n122,
    n64,
    n140,
    n76
  );


  nor
  g263
  (
    n159,
    n82,
    n138,
    n96,
    n72
  );


  xor
  g264
  (
    n174,
    n99,
    n95,
    n34,
    n129
  );


  xnor
  g265
  (
    n319,
    n83,
    n44,
    n135,
    n47
  );


  and
  g266
  (
    n267,
    n126,
    n39,
    n85,
    n147
  );


  nand
  g267
  (
    n321,
    n119,
    n44,
    n59,
    n62
  );


  nor
  g268
  (
    n296,
    n137,
    n104,
    n41,
    n110
  );


  nand
  g269
  (
    n153,
    n36,
    n61,
    n84,
    n136
  );


  and
  g270
  (
    n245,
    n61,
    n122,
    n69,
    n49
  );


  xor
  g271
  (
    n233,
    n101,
    n73,
    n59,
    n81
  );


  xnor
  g272
  (
    n183,
    n107,
    n51,
    n75,
    n131
  );


  nor
  g273
  (
    n248,
    n146,
    n110,
    n50,
    n90
  );


  xor
  g274
  (
    n162,
    n106,
    n85,
    n43,
    n59
  );


  or
  g275
  (
    n163,
    n52,
    n34,
    n35
  );


  nor
  g276
  (
    n250,
    n142,
    n69,
    n74,
    n120
  );


  or
  g277
  (
    n310,
    n58,
    n98,
    n125,
    n116
  );


  nand
  g278
  (
    n231,
    n98,
    n107,
    n129,
    n112
  );


  and
  g279
  (
    n166,
    n58,
    n135,
    n51,
    n120
  );


  or
  g280
  (
    n291,
    n144,
    n125,
    n94,
    n109
  );


  and
  g281
  (
    n198,
    n70,
    n146,
    n65,
    n92
  );


  or
  g282
  (
    KeyWire_0_15,
    n148,
    n42,
    n100,
    n63
  );


  xnor
  g283
  (
    n293,
    n132,
    n70,
    n52,
    n64
  );


  xor
  g284
  (
    n155,
    n95,
    n65,
    n143,
    n130
  );


  nor
  g285
  (
    n205,
    n149,
    n121,
    n62
  );


  or
  g286
  (
    n197,
    n132,
    n38,
    n118,
    n33
  );


  or
  g287
  (
    n226,
    n101,
    n108,
    n77,
    n96
  );


  and
  g288
  (
    n240,
    n41,
    n69,
    n142,
    n50
  );


  nand
  g289
  (
    n323,
    n133,
    n99,
    n110,
    n123
  );


  nor
  g290
  (
    n272,
    n95,
    n91,
    n127,
    n128
  );


  xnor
  g291
  (
    n327,
    n94,
    n98,
    n134,
    n39
  );


  and
  g292
  (
    n199,
    n144,
    n114,
    n53,
    n134
  );


  xnor
  g293
  (
    n271,
    n86,
    n131,
    n71,
    n105
  );


  and
  g294
  (
    n212,
    n61,
    n45,
    n39,
    n144
  );


  nand
  g295
  (
    n232,
    n93,
    n73,
    n139,
    n43
  );


  nor
  g296
  (
    n156,
    n132,
    n119,
    n123,
    n137
  );


  xor
  g297
  (
    KeyWire_0_17,
    n71,
    n116,
    n54,
    n49
  );


  or
  g298
  (
    n168,
    n88,
    n124,
    n52,
    n53
  );


  nand
  g299
  (
    n218,
    n63,
    n41,
    n124,
    n128
  );


  xor
  g300
  (
    n320,
    n37,
    n96,
    n67,
    n106
  );


  xor
  g301
  (
    n206,
    n140,
    n59,
    n120,
    n93
  );


  and
  g302
  (
    n306,
    n60,
    n90,
    n56,
    n70
  );


  and
  g303
  (
    n406,
    n328,
    n235,
    n230
  );


  nand
  g304
  (
    n351,
    n246,
    n284,
    n166,
    n234
  );


  nor
  g305
  (
    n430,
    n265,
    n298,
    n264,
    n331
  );


  and
  g306
  (
    n436,
    n174,
    n183,
    n333,
    n250
  );


  or
  g307
  (
    n451,
    n250,
    n177,
    n319,
    n323
  );


  and
  g308
  (
    n374,
    n249,
    n215,
    n315,
    n260
  );


  nand
  g309
  (
    n453,
    n329,
    n229,
    n271,
    n300
  );


  xor
  g310
  (
    n395,
    n249,
    n245,
    n252,
    n181
  );


  xor
  g311
  (
    n409,
    n199,
    n220,
    n225,
    n277
  );


  and
  g312
  (
    n461,
    n272,
    n211,
    n184,
    n232
  );


  nor
  g313
  (
    n364,
    n173,
    n181,
    n175,
    n268
  );


  or
  g314
  (
    n355,
    n237,
    n304,
    n257,
    n233
  );


  nand
  g315
  (
    n357,
    n272,
    n177,
    n248,
    n320
  );


  or
  g316
  (
    n435,
    n293,
    n305,
    n243,
    n208
  );


  xor
  g317
  (
    n399,
    n289,
    n291,
    n257,
    n274
  );


  or
  g318
  (
    n428,
    n191,
    n292,
    n267,
    n228
  );


  xnor
  g319
  (
    n337,
    n181,
    n312,
    n207,
    n259
  );


  nor
  g320
  (
    n367,
    n279,
    n219,
    n285,
    n209
  );


  nor
  g321
  (
    n443,
    n280,
    n288,
    n180,
    n227
  );


  xor
  g322
  (
    n347,
    n253,
    n283,
    n239,
    n190
  );


  nor
  g323
  (
    n343,
    n160,
    n254,
    n258,
    n280
  );


  xnor
  g324
  (
    n441,
    n157,
    n285,
    n251,
    n322
  );


  nor
  g325
  (
    n446,
    n318,
    n317,
    n266,
    n270
  );


  nand
  g326
  (
    n372,
    n296,
    n167,
    n212,
    n236
  );


  xnor
  g327
  (
    n348,
    n332,
    n206,
    n214,
    n331
  );


  nand
  g328
  (
    n417,
    n255,
    n251,
    n229,
    n310
  );


  or
  g329
  (
    n464,
    n228,
    n243,
    n242,
    n333
  );


  nor
  g330
  (
    KeyWire_0_56,
    n161,
    n237,
    n240
  );


  xor
  g331
  (
    n339,
    n155,
    n185,
    n253,
    n221
  );


  nor
  g332
  (
    n437,
    n189,
    n153,
    n292,
    n210
  );


  xnor
  g333
  (
    n456,
    n234,
    n169,
    n327,
    n307
  );


  and
  g334
  (
    n394,
    n244,
    n165,
    n311,
    n276
  );


  xnor
  g335
  (
    n360,
    n159,
    n196,
    n167,
    n264
  );


  xnor
  g336
  (
    n392,
    n297,
    n203,
    n315,
    n187
  );


  xnor
  g337
  (
    n376,
    n321,
    n280,
    n188,
    n250
  );


  xnor
  g338
  (
    n359,
    n196,
    n294,
    n275,
    n334
  );


  or
  g339
  (
    n401,
    n242,
    n316,
    n265,
    n227
  );


  nand
  g340
  (
    n466,
    n325,
    n300,
    n172,
    n295
  );


  xor
  g341
  (
    n362,
    n239,
    n308,
    n326,
    n327
  );


  nand
  g342
  (
    n391,
    n211,
    n238,
    n203,
    n205
  );


  xor
  g343
  (
    n455,
    n204,
    n180,
    n283,
    n245
  );


  xnor
  g344
  (
    n373,
    n210,
    n301,
    n241,
    n287
  );


  xnor
  g345
  (
    n440,
    n199,
    n186,
    n190,
    n303
  );


  or
  g346
  (
    n387,
    n271,
    n258,
    n303,
    n214
  );


  nand
  g347
  (
    n452,
    n311,
    n238,
    n281,
    n195
  );


  nand
  g348
  (
    n340,
    n229,
    n266,
    n281,
    n325
  );


  xnor
  g349
  (
    n410,
    n314,
    n178,
    n194,
    n312
  );


  and
  g350
  (
    n434,
    n307,
    n316,
    n299,
    n286
  );


  nor
  g351
  (
    n336,
    n268,
    n251,
    n158,
    n278
  );


  xor
  g352
  (
    n465,
    n208,
    n326,
    n291,
    n168
  );


  and
  g353
  (
    n458,
    n219,
    n224,
    n270,
    n218
  );


  and
  g354
  (
    n414,
    n330,
    n168,
    n243,
    n309
  );


  xor
  g355
  (
    n349,
    n311,
    n252,
    n191,
    n320
  );


  xnor
  g356
  (
    n344,
    n171,
    n266,
    n224,
    n201
  );


  nor
  g357
  (
    n378,
    n201,
    n210,
    n297,
    n151
  );


  xor
  g358
  (
    n382,
    n175,
    n202,
    n320,
    n217
  );


  xor
  g359
  (
    n413,
    n286,
    n190,
    n329,
    n192
  );


  nand
  g360
  (
    n462,
    n192,
    n333,
    n308,
    n272
  );


  xor
  g361
  (
    n352,
    n224,
    n294,
    n218,
    n222
  );


  and
  g362
  (
    n370,
    n169,
    n192,
    n197,
    n202
  );


  xnor
  g363
  (
    n368,
    n275,
    n230,
    n277,
    n310
  );


  or
  g364
  (
    n420,
    n291,
    n314,
    n182,
    n207
  );


  nor
  g365
  (
    n442,
    n254,
    n271,
    n292,
    n205
  );


  and
  g366
  (
    n363,
    n154,
    n240,
    n199,
    n263
  );


  xnor
  g367
  (
    n380,
    n188,
    n216,
    n232,
    n179
  );


  xnor
  g368
  (
    n386,
    n267,
    n207,
    n259,
    n217
  );


  and
  g369
  (
    n422,
    n306,
    n215,
    n209,
    n216
  );


  nand
  g370
  (
    n402,
    n302,
    n261,
    n212
  );


  and
  g371
  (
    n384,
    n220,
    n273,
    n282,
    n334
  );


  xnor
  g372
  (
    n412,
    n184,
    n227,
    n216,
    n201
  );


  nor
  g373
  (
    n385,
    n220,
    n282,
    n214,
    n168
  );


  and
  g374
  (
    n425,
    n294,
    n156,
    n178,
    n293
  );


  or
  g375
  (
    n365,
    n174,
    n188,
    n193,
    n327
  );


  xnor
  g376
  (
    n346,
    n183,
    n187,
    n197,
    n182
  );


  xnor
  g377
  (
    n375,
    n262,
    n262,
    n264,
    n171
  );


  xnor
  g378
  (
    n369,
    n267,
    n194,
    n317,
    n326
  );


  or
  g379
  (
    n381,
    n206,
    n325,
    n329,
    n178
  );


  and
  g380
  (
    n354,
    n173,
    n302,
    n189,
    n247
  );


  nand
  g381
  (
    n459,
    n313,
    n274,
    n186,
    n223
  );


  xnor
  g382
  (
    n439,
    n198,
    n328,
    n260,
    n191
  );


  and
  g383
  (
    n450,
    n301,
    n304,
    n323,
    n176
  );


  and
  g384
  (
    n398,
    n262,
    n166,
    n170,
    n226
  );


  xor
  g385
  (
    n388,
    n172,
    n189,
    n242,
    n296
  );


  nor
  g386
  (
    n438,
    n166,
    n164,
    n185,
    n295
  );


  nand
  g387
  (
    n397,
    n306,
    n305,
    n328,
    n179
  );


  nand
  g388
  (
    n383,
    n330,
    n246,
    n231,
    n200
  );


  and
  g389
  (
    n419,
    n287,
    n284,
    n286,
    n241
  );


  or
  g390
  (
    n463,
    n184,
    n303,
    n319,
    n322
  );


  xor
  g391
  (
    n405,
    n223,
    n269,
    n310,
    n233
  );


  nand
  g392
  (
    n371,
    n203,
    n183,
    n295,
    n259
  );


  nand
  g393
  (
    n379,
    n330,
    n176,
    n313,
    n324
  );


  and
  g394
  (
    n444,
    n206,
    n315,
    n278,
    n300
  );


  nor
  g395
  (
    n408,
    n235,
    n301,
    n177,
    n257
  );


  xnor
  g396
  (
    n460,
    n204,
    n231,
    n334,
    n234
  );


  or
  g397
  (
    n400,
    n274,
    n163,
    n236,
    n194
  );


  xnor
  g398
  (
    n432,
    n290,
    n255,
    n283,
    n256
  );


  xor
  g399
  (
    n411,
    n215,
    n232,
    n299,
    n279
  );


  or
  g400
  (
    n345,
    n287,
    n172,
    n321,
    n244
  );


  nand
  g401
  (
    n390,
    n304,
    n273,
    n219,
    n314
  );


  nor
  g402
  (
    n350,
    n213,
    n324,
    n276,
    n240
  );


  xor
  g403
  (
    n448,
    n255,
    n306,
    n200,
    n313
  );


  nand
  g404
  (
    n353,
    n179,
    n175,
    n263,
    n222
  );


  nor
  g405
  (
    n366,
    n169,
    n309,
    n182,
    n285
  );


  nand
  g406
  (
    KeyWire_0_2,
    n223,
    n180,
    n278,
    n308
  );


  or
  g407
  (
    n338,
    n247,
    n202,
    n261,
    n296
  );


  nand
  g408
  (
    n358,
    n239,
    n171,
    n218,
    n204
  );


  xnor
  g409
  (
    n429,
    n195,
    n230,
    n225,
    n253
  );


  and
  g410
  (
    n445,
    n284,
    n332,
    n289,
    n324
  );


  xor
  g411
  (
    n454,
    n221,
    n225,
    n236,
    n307
  );


  nand
  g412
  (
    n423,
    n198,
    n197,
    n195,
    n193
  );


  nor
  g413
  (
    n341,
    n212,
    n167,
    n279,
    n269
  );


  and
  g414
  (
    n342,
    n322,
    n187,
    n319,
    n198
  );


  nand
  g415
  (
    n449,
    n162,
    n273,
    n185,
    n200
  );


  xor
  g416
  (
    n457,
    n150,
    n312,
    n245,
    n265
  );


  nor
  g417
  (
    n418,
    n289,
    n282,
    n252,
    n318
  );


  nand
  g418
  (
    n389,
    n270,
    n213,
    n233,
    n222
  );


  xor
  g419
  (
    n393,
    n254,
    n196,
    n248,
    n331
  );


  nand
  g420
  (
    n361,
    n256,
    n318,
    n263,
    n298
  );


  and
  g421
  (
    n431,
    n302,
    n238,
    n277,
    n317
  );


  nor
  g422
  (
    n433,
    n170,
    n235,
    n221,
    n288
  );


  or
  g423
  (
    n416,
    n174,
    n332,
    n258,
    n152
  );


  nand
  g424
  (
    n415,
    n193,
    n226,
    n246,
    n269
  );


  and
  g425
  (
    n377,
    n275,
    n293,
    n290,
    n305
  );


  xor
  g426
  (
    n396,
    n209,
    n186,
    n249,
    n290
  );


  and
  g427
  (
    n427,
    n205,
    n321,
    n176,
    n226
  );


  and
  g428
  (
    n447,
    n241,
    n323,
    n268,
    n244
  );


  or
  g429
  (
    n426,
    n228,
    n298,
    n248,
    n213
  );


  nor
  g430
  (
    n421,
    n173,
    n211,
    n208,
    n247
  );


  nand
  g431
  (
    n407,
    n260,
    n276,
    n170,
    n309
  );


  or
  g432
  (
    n356,
    n316,
    n288,
    n299,
    n231
  );


  xnor
  g433
  (
    n403,
    n256,
    n217,
    n281,
    n297
  );


  not
  g434
  (
    n615,
    n364
  );


  buf
  g435
  (
    n534,
    n442
  );


  buf
  g436
  (
    n593,
    n442
  );


  buf
  g437
  (
    n588,
    n435
  );


  not
  g438
  (
    n527,
    n360
  );


  buf
  g439
  (
    n565,
    n399
  );


  not
  g440
  (
    n591,
    n408
  );


  not
  g441
  (
    n499,
    n413
  );


  buf
  g442
  (
    n523,
    n370
  );


  buf
  g443
  (
    n516,
    n436
  );


  not
  g444
  (
    n554,
    n417
  );


  buf
  g445
  (
    KeyWire_0_47,
    n405
  );


  buf
  g446
  (
    n555,
    n394
  );


  not
  g447
  (
    n528,
    n363
  );


  not
  g448
  (
    n542,
    n437
  );


  not
  g449
  (
    n473,
    n359
  );


  buf
  g450
  (
    n530,
    n371
  );


  not
  g451
  (
    n572,
    n428
  );


  buf
  g452
  (
    n569,
    n427
  );


  buf
  g453
  (
    n561,
    n409
  );


  buf
  g454
  (
    n510,
    n368
  );


  not
  g455
  (
    KeyWire_0_35,
    n367
  );


  buf
  g456
  (
    n574,
    n422
  );


  not
  g457
  (
    KeyWire_0_30,
    n441
  );


  not
  g458
  (
    n557,
    n425
  );


  not
  g459
  (
    n536,
    n424
  );


  not
  g460
  (
    n540,
    n395
  );


  not
  g461
  (
    n623,
    n393
  );


  buf
  g462
  (
    n525,
    n420
  );


  buf
  g463
  (
    n550,
    n362
  );


  not
  g464
  (
    n511,
    n337
  );


  buf
  g465
  (
    n594,
    n348
  );


  buf
  g466
  (
    n468,
    n401
  );


  buf
  g467
  (
    n496,
    n361
  );


  not
  g468
  (
    n486,
    n416
  );


  not
  g469
  (
    n548,
    n375
  );


  not
  g470
  (
    n607,
    n398
  );


  not
  g471
  (
    n590,
    n433
  );


  buf
  g472
  (
    n610,
    n437
  );


  not
  g473
  (
    n531,
    n430
  );


  buf
  g474
  (
    n620,
    n419
  );


  buf
  g475
  (
    n599,
    n347
  );


  buf
  g476
  (
    n503,
    n438
  );


  buf
  g477
  (
    n609,
    n442
  );


  buf
  g478
  (
    n582,
    n431
  );


  not
  g479
  (
    n492,
    n419
  );


  not
  g480
  (
    n489,
    n374
  );


  buf
  g481
  (
    n549,
    n427
  );


  not
  g482
  (
    n533,
    n441
  );


  not
  g483
  (
    n537,
    n357
  );


  not
  g484
  (
    n556,
    n438
  );


  not
  g485
  (
    n475,
    n432
  );


  not
  g486
  (
    n621,
    n406
  );


  not
  g487
  (
    n513,
    n440
  );


  not
  g488
  (
    n545,
    n435
  );


  not
  g489
  (
    n471,
    n407
  );


  not
  g490
  (
    n584,
    n439
  );


  buf
  g491
  (
    n587,
    n426
  );


  not
  g492
  (
    n477,
    n380
  );


  buf
  g493
  (
    n570,
    n391
  );


  not
  g494
  (
    n551,
    n422
  );


  buf
  g495
  (
    n539,
    n340
  );


  not
  g496
  (
    n566,
    n378
  );


  not
  g497
  (
    n470,
    n425
  );


  not
  g498
  (
    n543,
    n373
  );


  not
  g499
  (
    n597,
    n431
  );


  buf
  g500
  (
    n508,
    n377
  );


  not
  g501
  (
    n515,
    n392
  );


  buf
  g502
  (
    n577,
    n381
  );


  buf
  g503
  (
    n541,
    n403
  );


  not
  g504
  (
    n506,
    n429
  );


  not
  g505
  (
    n618,
    n387
  );


  buf
  g506
  (
    KeyWire_0_55,
    n410
  );


  buf
  g507
  (
    n512,
    n436
  );


  not
  g508
  (
    n480,
    n438
  );


  buf
  g509
  (
    n529,
    n388
  );


  not
  g510
  (
    n553,
    n354
  );


  not
  g511
  (
    n520,
    n434
  );


  not
  g512
  (
    n576,
    n345
  );


  not
  g513
  (
    n589,
    n424
  );


  not
  g514
  (
    n521,
    n443
  );


  not
  g515
  (
    n564,
    n351
  );


  buf
  g516
  (
    n573,
    n423
  );


  not
  g517
  (
    n559,
    n396
  );


  buf
  g518
  (
    n494,
    n432
  );


  not
  g519
  (
    n600,
    n417
  );


  buf
  g520
  (
    n580,
    n434
  );


  buf
  g521
  (
    n507,
    n421
  );


  buf
  g522
  (
    n481,
    n413
  );


  buf
  g523
  (
    n505,
    n355
  );


  not
  g524
  (
    n622,
    n440
  );


  not
  g525
  (
    n614,
    n342
  );


  not
  g526
  (
    n560,
    n431
  );


  not
  g527
  (
    n586,
    n412
  );


  buf
  g528
  (
    n578,
    n365
  );


  buf
  g529
  (
    n474,
    n379
  );


  buf
  g530
  (
    n571,
    n336
  );


  not
  g531
  (
    n524,
    n432
  );


  buf
  g532
  (
    n518,
    n356
  );


  buf
  g533
  (
    n485,
    n411
  );


  buf
  g534
  (
    n526,
    n435
  );


  not
  g535
  (
    KeyWire_0_21,
    n443
  );


  buf
  g536
  (
    n579,
    n429
  );


  buf
  g537
  (
    n472,
    n429
  );


  buf
  g538
  (
    n535,
    n439
  );


  not
  g539
  (
    n603,
    n423
  );


  not
  g540
  (
    n568,
    n366
  );


  not
  g541
  (
    n493,
    n428
  );


  not
  g542
  (
    n575,
    n390
  );


  not
  g543
  (
    n501,
    n433
  );


  not
  g544
  (
    n604,
    n384
  );


  buf
  g545
  (
    n619,
    n420
  );


  not
  g546
  (
    n483,
    n415
  );


  buf
  g547
  (
    n601,
    n397
  );


  buf
  g548
  (
    n612,
    n426
  );


  buf
  g549
  (
    n562,
    n414
  );


  not
  g550
  (
    n478,
    n386
  );


  not
  g551
  (
    n567,
    n383
  );


  buf
  g552
  (
    n487,
    n436
  );


  buf
  g553
  (
    n596,
    n404
  );


  not
  g554
  (
    n484,
    n421
  );


  buf
  g555
  (
    n514,
    n411
  );


  not
  g556
  (
    n544,
    n410
  );


  buf
  g557
  (
    n581,
    n418
  );


  not
  g558
  (
    n495,
    n441
  );


  buf
  g559
  (
    n498,
    n430
  );


  not
  g560
  (
    n509,
    n352
  );


  buf
  g561
  (
    n585,
    n412
  );


  not
  g562
  (
    n488,
    n350
  );


  not
  g563
  (
    n490,
    n434
  );


  buf
  g564
  (
    n592,
    n428
  );


  buf
  g565
  (
    n611,
    n382
  );


  not
  g566
  (
    n595,
    n344
  );


  not
  g567
  (
    n552,
    n389
  );


  buf
  g568
  (
    n617,
    n400
  );


  not
  g569
  (
    n517,
    n415
  );


  buf
  g570
  (
    n482,
    n341
  );


  buf
  g571
  (
    n606,
    n339
  );


  buf
  g572
  (
    KeyWire_0_26,
    n418
  );


  not
  g573
  (
    n613,
    n433
  );


  buf
  g574
  (
    n497,
    n439
  );


  buf
  g575
  (
    n504,
    n385
  );


  not
  g576
  (
    n502,
    n338
  );


  not
  g577
  (
    n608,
    n343
  );


  not
  g578
  (
    n546,
    n414
  );


  not
  g579
  (
    n583,
    n369
  );


  not
  g580
  (
    n547,
    n372
  );


  buf
  g581
  (
    n532,
    n440
  );


  buf
  g582
  (
    n500,
    n346
  );


  buf
  g583
  (
    n605,
    n430
  );


  buf
  g584
  (
    n522,
    n402
  );


  buf
  g585
  (
    n469,
    n376
  );


  not
  g586
  (
    n479,
    n353
  );


  buf
  g587
  (
    n558,
    n437
  );


  not
  g588
  (
    n467,
    n349
  );


  not
  g589
  (
    n519,
    n416
  );


  not
  g590
  (
    n598,
    n358
  );


  or
  g591
  (
    n724,
    n508,
    n555,
    n497,
    n580
  );


  nand
  g592
  (
    n631,
    n491,
    n476,
    n527,
    n584
  );


  nand
  g593
  (
    n657,
    n542,
    n507,
    n500,
    n581
  );


  nand
  g594
  (
    n721,
    n585,
    n542,
    n524,
    n541
  );


  xor
  g595
  (
    n746,
    n532,
    n555,
    n475,
    n543
  );


  nor
  g596
  (
    n691,
    n552,
    n581,
    n525,
    n486
  );


  and
  g597
  (
    n661,
    n529,
    n585,
    n574,
    n570
  );


  xor
  g598
  (
    n737,
    n535,
    n492,
    n542,
    n478
  );


  and
  g599
  (
    KeyWire_0_52,
    n505,
    n494,
    n558,
    n499
  );


  xor
  g600
  (
    n649,
    n525,
    n574,
    n531,
    n485
  );


  xor
  g601
  (
    n738,
    n512,
    n570,
    n528,
    n471
  );


  nor
  g602
  (
    n723,
    n498,
    n588,
    n513
  );


  xor
  g603
  (
    n702,
    n493,
    n498,
    n568,
    n539
  );


  or
  g604
  (
    n638,
    n499,
    n488,
    n475,
    n527
  );


  nand
  g605
  (
    n630,
    n540,
    n591,
    n545,
    n495
  );


  or
  g606
  (
    n728,
    n533,
    n547,
    n577,
    n515
  );


  xor
  g607
  (
    n665,
    n492,
    n502,
    n480,
    n584
  );


  nand
  g608
  (
    n643,
    n553,
    n587,
    n564,
    n495
  );


  nor
  g609
  (
    n686,
    n478,
    n570,
    n489,
    n488
  );


  or
  g610
  (
    n624,
    n554,
    n530,
    n513,
    n591
  );


  nand
  g611
  (
    n708,
    n550,
    n589,
    n536,
    n567
  );


  xnor
  g612
  (
    n729,
    n580,
    n590,
    n471,
    n555
  );


  and
  g613
  (
    n651,
    n565,
    n508,
    n510,
    n534
  );


  or
  g614
  (
    n732,
    n474,
    n557,
    n580,
    n561
  );


  xor
  g615
  (
    n694,
    n517,
    n545,
    n487,
    n585
  );


  or
  g616
  (
    n662,
    n535,
    n501,
    n487,
    n497
  );


  nor
  g617
  (
    n712,
    n524,
    n483,
    n582,
    n535
  );


  nand
  g618
  (
    n650,
    n526,
    n479,
    n519,
    n473
  );


  or
  g619
  (
    n625,
    n471,
    n468,
    n532,
    n559
  );


  nand
  g620
  (
    n684,
    n490,
    n576,
    n562,
    n542
  );


  xor
  g621
  (
    n741,
    n502,
    n524,
    n507,
    n494
  );


  or
  g622
  (
    n666,
    n566,
    n491,
    n574,
    n582
  );


  and
  g623
  (
    n711,
    n468,
    n575,
    n571,
    n519
  );


  xor
  g624
  (
    n727,
    n496,
    n564,
    n512,
    n481
  );


  xnor
  g625
  (
    n656,
    n509,
    n513,
    n489,
    n491
  );


  nand
  g626
  (
    n640,
    n482,
    n556,
    n509,
    n505
  );


  or
  g627
  (
    n710,
    n486,
    n582,
    n576,
    n557
  );


  and
  g628
  (
    n736,
    n588,
    n521,
    n578,
    n519
  );


  or
  g629
  (
    n716,
    n476,
    n483,
    n484,
    n511
  );


  xnor
  g630
  (
    n648,
    n493,
    n583,
    n541,
    n540
  );


  xnor
  g631
  (
    n720,
    n538,
    n482,
    n525,
    n518
  );


  xnor
  g632
  (
    n670,
    n517,
    n504,
    n587,
    n529
  );


  nand
  g633
  (
    n730,
    n527,
    n477,
    n474,
    n538
  );


  xor
  g634
  (
    n726,
    n511,
    n510,
    n566,
    n520
  );


  or
  g635
  (
    n654,
    n566,
    n534,
    n562,
    n543
  );


  nand
  g636
  (
    n725,
    n483,
    n544,
    n501,
    n553
  );


  nand
  g637
  (
    n641,
    n494,
    n521,
    n506,
    n532
  );


  xor
  g638
  (
    n669,
    n537,
    n568,
    n552,
    n585
  );


  nand
  g639
  (
    n699,
    n546,
    n530,
    n498,
    n559
  );


  xnor
  g640
  (
    n700,
    n497,
    n473,
    n558,
    n480
  );


  and
  g641
  (
    n733,
    n575,
    n549,
    n584,
    n534
  );


  xnor
  g642
  (
    n645,
    n514,
    n529,
    n490,
    n592
  );


  nand
  g643
  (
    n663,
    n482,
    n531,
    n473,
    n492
  );


  xnor
  g644
  (
    n689,
    n539,
    n569,
    n556,
    n566
  );


  xnor
  g645
  (
    n677,
    n588,
    n470,
    n513,
    n549
  );


  nor
  g646
  (
    n706,
    n479,
    n552,
    n509,
    n495
  );


  and
  g647
  (
    n671,
    n577,
    n556,
    n584,
    n572
  );


  nor
  g648
  (
    KeyWire_0_50,
    n480,
    n541,
    n504,
    n469
  );


  nand
  g649
  (
    n688,
    n579,
    n518,
    n553,
    n496
  );


  and
  g650
  (
    n642,
    n567,
    n544,
    n504,
    n589
  );


  nor
  g651
  (
    n674,
    n553,
    n591,
    n485,
    n580
  );


  nor
  g652
  (
    n637,
    n573,
    n545,
    n522,
    n521
  );


  nand
  g653
  (
    n719,
    n491,
    n545,
    n551,
    n503
  );


  or
  g654
  (
    n635,
    n560,
    n531,
    n541,
    n507
  );


  nor
  g655
  (
    n739,
    n490,
    n492,
    n515,
    n561
  );


  xnor
  g656
  (
    n646,
    n511,
    n505,
    n536,
    n534
  );


  xor
  g657
  (
    n696,
    n573,
    n526,
    n502,
    n536
  );


  nor
  g658
  (
    n713,
    n468,
    n526,
    n537,
    n568
  );


  and
  g659
  (
    n714,
    n564,
    n563,
    n569,
    n482
  );


  xor
  g660
  (
    n679,
    n530,
    n493,
    n578,
    n528
  );


  nand
  g661
  (
    n628,
    n489,
    n570,
    n569,
    n587
  );


  xor
  g662
  (
    n639,
    n496,
    n490,
    n583,
    n483
  );


  nand
  g663
  (
    n632,
    n543,
    n503,
    n476,
    n590
  );


  xnor
  g664
  (
    n676,
    n575,
    n515,
    n525,
    n536
  );


  nand
  g665
  (
    n658,
    n527,
    n554,
    n516,
    n510
  );


  and
  g666
  (
    n707,
    n488,
    n509,
    n470,
    n579
  );


  xnor
  g667
  (
    n745,
    n548,
    n551,
    n520,
    n484
  );


  nand
  g668
  (
    n680,
    n539,
    n498,
    n533,
    n572
  );


  xor
  g669
  (
    n692,
    n505,
    n583,
    n546,
    n488
  );


  or
  g670
  (
    n682,
    n574,
    n499,
    n518,
    n577
  );


  nor
  g671
  (
    n678,
    n494,
    n496,
    n480,
    n508
  );


  xor
  g672
  (
    n653,
    n506,
    n554,
    n467,
    n562
  );


  nor
  g673
  (
    n636,
    n577,
    n469,
    n558,
    n568
  );


  or
  g674
  (
    n717,
    n489,
    n551,
    n548,
    n589
  );


  xor
  g675
  (
    n698,
    n520,
    n535,
    n526,
    n557
  );


  or
  g676
  (
    n740,
    n511,
    n484,
    n495,
    n563
  );


  nand
  g677
  (
    n722,
    n552,
    n493,
    n591,
    n567
  );


  nand
  g678
  (
    n705,
    n474,
    n516,
    n563,
    n582
  );


  and
  g679
  (
    n731,
    n571,
    n550,
    n547,
    n537
  );


  nor
  g680
  (
    n744,
    n571,
    n586,
    n549,
    n504
  );


  and
  g681
  (
    n681,
    n579,
    n560,
    n548
  );


  xnor
  g682
  (
    n644,
    n486,
    n487,
    n561,
    n517
  );


  xor
  g683
  (
    n685,
    n572,
    n514,
    n524,
    n550
  );


  nand
  g684
  (
    n701,
    n551,
    n470,
    n569,
    n523
  );


  nand
  g685
  (
    n647,
    n589,
    n555,
    n517,
    n519
  );


  nand
  g686
  (
    n627,
    n567,
    n479,
    n538,
    n547
  );


  or
  g687
  (
    n743,
    n510,
    n472,
    n516,
    n487
  );


  or
  g688
  (
    n715,
    n467,
    n467,
    n539,
    n499
  );


  nor
  g689
  (
    n695,
    n531,
    n479,
    n522,
    n558
  );


  nor
  g690
  (
    n652,
    n572,
    n514,
    n587,
    n537
  );


  or
  g691
  (
    n718,
    n518,
    n564,
    n561,
    n547
  );


  and
  g692
  (
    n709,
    n550,
    n485,
    n506,
    n575
  );


  or
  g693
  (
    n683,
    n478,
    n512,
    n485,
    n586
  );


  xnor
  g694
  (
    n664,
    n538,
    n565,
    n578,
    n559
  );


  or
  g695
  (
    n704,
    n522,
    n523,
    n563,
    n469
  );


  xor
  g696
  (
    n675,
    n500,
    n559,
    n507,
    n530
  );


  or
  g697
  (
    n626,
    n481,
    n472,
    n529,
    n528
  );


  nand
  g698
  (
    n690,
    n508,
    n573,
    n481,
    n506
  );


  and
  g699
  (
    n687,
    n522,
    n543,
    n486,
    n523
  );


  xor
  g700
  (
    n667,
    n576,
    n554,
    n501,
    n571
  );


  nand
  g701
  (
    n735,
    n532,
    n581,
    n583,
    n516
  );


  or
  g702
  (
    n703,
    n549,
    n533,
    n523,
    n540
  );


  and
  g703
  (
    n629,
    n546,
    n503,
    n590,
    n520
  );


  nand
  g704
  (
    n633,
    n484,
    n556,
    n560,
    n512
  );


  nor
  g705
  (
    n734,
    n514,
    n528,
    n472,
    n477
  );


  nand
  g706
  (
    n673,
    n557,
    n565,
    n501,
    n503
  );


  and
  g707
  (
    n660,
    n500,
    n478,
    n533,
    n515
  );


  or
  g708
  (
    n655,
    n592,
    n497,
    n581,
    n540
  );


  xor
  g709
  (
    n693,
    n586,
    n477,
    n475,
    n500
  );


  xor
  g710
  (
    n668,
    n586,
    n592,
    n578,
    n502
  );


  or
  g711
  (
    n634,
    n565,
    n579,
    n590,
    n544
  );


  and
  g712
  (
    n659,
    n546,
    n573,
    n544,
    n481
  );


  xor
  g713
  (
    n742,
    n576,
    n548,
    n521,
    n562
  );


  not
  g714
  (
    n749,
    n630
  );


  not
  g715
  (
    n754,
    n633
  );


  buf
  g716
  (
    n752,
    n628
  );


  not
  g717
  (
    n757,
    n632
  );


  buf
  g718
  (
    n753,
    n629
  );


  not
  g719
  (
    n756,
    n624
  );


  buf
  g720
  (
    n751,
    n625
  );


  not
  g721
  (
    n755,
    n627
  );


  not
  g722
  (
    n747,
    n626
  );


  buf
  g723
  (
    n748,
    n634
  );


  buf
  g724
  (
    n750,
    n631
  );


  xor
  g725
  (
    n773,
    n465,
    n757,
    n601,
    n603
  );


  xor
  g726
  (
    n789,
    n749,
    n595,
    n458,
    n448
  );


  or
  g727
  (
    n769,
    n757,
    n602,
    n599,
    n750
  );


  xnor
  g728
  (
    n780,
    n444,
    n752,
    n598,
    n754
  );


  and
  g729
  (
    n785,
    n747,
    n459,
    n444,
    n149
  );


  xnor
  g730
  (
    n771,
    n453,
    n454,
    n756
  );


  xnor
  g731
  (
    n783,
    n458,
    n455,
    n463,
    n753
  );


  xor
  g732
  (
    n792,
    n465,
    n462,
    n755
  );


  nor
  g733
  (
    n770,
    n448,
    n747,
    n601,
    n455
  );


  nor
  g734
  (
    n781,
    n464,
    n751,
    n460,
    n463
  );


  and
  g735
  (
    n787,
    n752,
    n600,
    n447,
    n755
  );


  and
  g736
  (
    n765,
    n748,
    n604,
    n449,
    n751
  );


  xnor
  g737
  (
    n796,
    n595,
    n594,
    n465,
    n461
  );


  xnor
  g738
  (
    n778,
    n460,
    n453,
    n597,
    n598
  );


  xor
  g739
  (
    n760,
    n444,
    n599,
    n601,
    n460
  );


  or
  g740
  (
    n758,
    n452,
    n446,
    n754,
    n449
  );


  nor
  g741
  (
    n793,
    n748,
    n755,
    n597
  );


  or
  g742
  (
    n774,
    n601,
    n604,
    n445,
    n756
  );


  nor
  g743
  (
    n799,
    n447,
    n596,
    n335,
    n456
  );


  xnor
  g744
  (
    n763,
    n32,
    n603,
    n443,
    n450
  );


  xor
  g745
  (
    n777,
    n450,
    n750,
    n598,
    n593
  );


  nand
  g746
  (
    n795,
    n449,
    n451,
    n754,
    n600
  );


  nand
  g747
  (
    n766,
    n463,
    n461,
    n596,
    n451
  );


  xor
  g748
  (
    n772,
    n32,
    n599,
    n757,
    n445
  );


  nor
  g749
  (
    n768,
    n751,
    n454,
    n602,
    n31
  );


  nor
  g750
  (
    n790,
    n600,
    n603,
    n593,
    n466
  );


  xnor
  g751
  (
    n767,
    n448,
    n447,
    n595,
    n594
  );


  xnor
  g752
  (
    n791,
    n466,
    n446,
    n462,
    n756
  );


  nand
  g753
  (
    n764,
    n602,
    n466,
    n750,
    n456
  );


  or
  g754
  (
    n794,
    n597,
    n593,
    n464,
    n456
  );


  xor
  g755
  (
    n775,
    n593,
    n457,
    n749,
    n458
  );


  or
  g756
  (
    n786,
    n453,
    n753,
    n749
  );


  xor
  g757
  (
    n788,
    n459,
    n335,
    n752,
    n596
  );


  or
  g758
  (
    n761,
    n748,
    n594,
    n451,
    n597
  );


  nor
  g759
  (
    n776,
    n450,
    n600,
    n756,
    n32
  );


  and
  g760
  (
    n762,
    n459,
    n747,
    n752,
    n595
  );


  nor
  g761
  (
    n759,
    n604,
    n753,
    n751,
    n599
  );


  nand
  g762
  (
    n798,
    n754,
    n464,
    n592,
    n457
  );


  or
  g763
  (
    n782,
    n750,
    n455,
    n457,
    n452
  );


  nor
  g764
  (
    n797,
    n596,
    n753,
    n445,
    n602
  );


  nor
  g765
  (
    n784,
    n598,
    n452,
    n446,
    n594
  );


  and
  g766
  (
    n779,
    n335,
    n757,
    n603,
    n461
  );


  xnor
  g767
  (
    n812,
    n615,
    n774,
    n608
  );


  and
  g768
  (
    n823,
    n615,
    n606,
    n605
  );


  nor
  g769
  (
    n819,
    n781,
    n798,
    n611
  );


  or
  g770
  (
    n816,
    n604,
    n787,
    n614
  );


  nand
  g771
  (
    n803,
    n607,
    n609
  );


  and
  g772
  (
    n805,
    n616,
    n795,
    n613
  );


  or
  g773
  (
    n820,
    n793,
    n614
  );


  nand
  g774
  (
    n817,
    n606,
    n617
  );


  nor
  g775
  (
    n818,
    n784,
    n791,
    n796
  );


  and
  g776
  (
    n821,
    n609,
    n608,
    n610
  );


  xnor
  g777
  (
    n814,
    n782,
    n607,
    n605
  );


  and
  g778
  (
    n813,
    n783,
    n613,
    n610
  );


  or
  g779
  (
    n807,
    n611,
    n790,
    n780
  );


  or
  g780
  (
    n808,
    n788,
    n776,
    n612
  );


  nand
  g781
  (
    n800,
    n608,
    n611,
    n609
  );


  nor
  g782
  (
    n801,
    n613,
    n777,
    n775
  );


  and
  g783
  (
    n806,
    n606,
    n605,
    n789,
    n616
  );


  and
  g784
  (
    n809,
    n617,
    n785,
    n615,
    n778
  );


  nor
  g785
  (
    n810,
    n610,
    n617,
    n792,
    n615
  );


  and
  g786
  (
    n804,
    n794,
    n612,
    n786,
    n605
  );


  xnor
  g787
  (
    n815,
    n614,
    n606,
    n611,
    n607
  );


  nor
  g788
  (
    n802,
    n616,
    n616,
    n797,
    n608
  );


  xnor
  g789
  (
    KeyWire_0_59,
    n613,
    n610,
    n612
  );


  nor
  g790
  (
    n822,
    n618,
    n799,
    n779,
    n607
  );


  not
  g791
  (
    n900,
    n642
  );


  buf
  g792
  (
    n886,
    n816
  );


  buf
  g793
  (
    n833,
    n726
  );


  not
  g794
  (
    n899,
    n663
  );


  buf
  g795
  (
    n898,
    n819
  );


  not
  g796
  (
    n849,
    n820
  );


  buf
  g797
  (
    n887,
    n802
  );


  not
  g798
  (
    n826,
    n809
  );


  not
  g799
  (
    n830,
    n661
  );


  buf
  g800
  (
    n892,
    n814
  );


  not
  g801
  (
    n860,
    n666
  );


  not
  g802
  (
    n878,
    n800
  );


  not
  g803
  (
    n840,
    n815
  );


  buf
  g804
  (
    n879,
    n685
  );


  not
  g805
  (
    n850,
    n706
  );


  not
  g806
  (
    n846,
    n712
  );


  not
  g807
  (
    n896,
    n811
  );


  not
  g808
  (
    n842,
    n669
  );


  buf
  g809
  (
    n883,
    n822
  );


  not
  g810
  (
    n847,
    n817
  );


  not
  g811
  (
    n880,
    n674
  );


  not
  g812
  (
    n889,
    n671
  );


  not
  g813
  (
    n858,
    n636
  );


  buf
  g814
  (
    n863,
    n808
  );


  not
  g815
  (
    n851,
    n716
  );


  buf
  g816
  (
    n864,
    n820
  );


  buf
  g817
  (
    n877,
    n744
  );


  not
  g818
  (
    n825,
    n700
  );


  not
  g819
  (
    n866,
    n822
  );


  buf
  g820
  (
    n869,
    n815
  );


  not
  g821
  (
    n884,
    n646
  );


  buf
  g822
  (
    n873,
    n820
  );


  buf
  g823
  (
    n875,
    n668
  );


  buf
  g824
  (
    n843,
    n692
  );


  buf
  g825
  (
    n861,
    n821
  );


  buf
  g826
  (
    n868,
    n724
  );


  buf
  g827
  (
    n834,
    n819
  );


  buf
  g828
  (
    n836,
    n660
  );


  buf
  g829
  (
    n871,
    n697
  );


  nand
  g830
  (
    n876,
    n688,
    n714
  );


  and
  g831
  (
    n852,
    n664,
    n810,
    n808,
    n732
  );


  xnor
  g832
  (
    n870,
    n821,
    n641,
    n807,
    n649
  );


  xor
  g833
  (
    n827,
    n819,
    n731,
    n643,
    n676
  );


  nor
  g834
  (
    n837,
    n659,
    n677,
    n696,
    n667
  );


  xnor
  g835
  (
    n882,
    n698,
    n823,
    n810
  );


  xnor
  g836
  (
    n893,
    n717,
    n812,
    n739,
    n662
  );


  or
  g837
  (
    n859,
    n822,
    n679,
    n802,
    n687
  );


  nand
  g838
  (
    n872,
    n811,
    n719,
    n742,
    n745
  );


  xor
  g839
  (
    n854,
    n684,
    n822,
    n699,
    n819
  );


  nand
  g840
  (
    n856,
    n727,
    n812,
    n728,
    n715
  );


  nor
  g841
  (
    n891,
    n808,
    n811,
    n823,
    n740
  );


  or
  g842
  (
    n832,
    n803,
    n816,
    n813,
    n673
  );


  nand
  g843
  (
    n895,
    n816,
    n713,
    n818,
    n683
  );


  or
  g844
  (
    n897,
    n820,
    n705,
    n813,
    n665
  );


  nor
  g845
  (
    n845,
    n645,
    n805,
    n658,
    n723
  );


  or
  g846
  (
    n865,
    n701,
    n735,
    n736,
    n814
  );


  nand
  g847
  (
    n888,
    n707,
    n722,
    n809,
    n710
  );


  xor
  g848
  (
    n862,
    n694,
    n809,
    n704,
    n695
  );


  xor
  g849
  (
    n824,
    n804,
    n741,
    n702,
    n821
  );


  nor
  g850
  (
    n885,
    n806,
    n805,
    n818,
    n738
  );


  or
  g851
  (
    n828,
    n678,
    n721,
    n807
  );


  nor
  g852
  (
    n894,
    n815,
    n800,
    n801,
    n803
  );


  nor
  g853
  (
    n844,
    n672,
    n689,
    n817,
    n729
  );


  xnor
  g854
  (
    n874,
    n670,
    n644,
    n640,
    n651
  );


  xor
  g855
  (
    n890,
    n823,
    n805,
    n817,
    n709
  );


  xnor
  g856
  (
    n855,
    n686,
    n818,
    n675,
    n708
  );


  nand
  g857
  (
    n831,
    n654,
    n703,
    n806,
    n804
  );


  xor
  g858
  (
    n848,
    n637,
    n693,
    n734,
    n802
  );


  xnor
  g859
  (
    n841,
    n682,
    n655,
    n804,
    n725
  );


  xnor
  g860
  (
    n835,
    n800,
    n647,
    n801,
    n639
  );


  xnor
  g861
  (
    n839,
    n657,
    n803,
    n635,
    n810
  );


  or
  g862
  (
    n881,
    n814,
    n680,
    n656,
    n801
  );


  nand
  g863
  (
    n867,
    n746,
    n737,
    n690,
    n821
  );


  nand
  g864
  (
    n838,
    n812,
    n730,
    n711,
    n650
  );


  or
  g865
  (
    n853,
    n681,
    n733,
    n648,
    n653
  );


  or
  g866
  (
    n857,
    n806,
    n720,
    n743,
    n718
  );


  xnor
  g867
  (
    n829,
    n652,
    n638,
    n691,
    n813
  );


  buf
  g868
  (
    n948,
    n844
  );


  buf
  g869
  (
    n945,
    n849
  );


  buf
  g870
  (
    n1036,
    n875
  );


  buf
  g871
  (
    n976,
    n844
  );


  buf
  g872
  (
    n941,
    n894
  );


  not
  g873
  (
    n1001,
    n837
  );


  buf
  g874
  (
    n1053,
    n856
  );


  not
  g875
  (
    n1049,
    n869
  );


  buf
  g876
  (
    n1011,
    n878
  );


  not
  g877
  (
    KeyWire_0_22,
    n890
  );


  buf
  g878
  (
    n1075,
    n889
  );


  buf
  g879
  (
    n959,
    n826
  );


  not
  g880
  (
    n989,
    n851
  );


  not
  g881
  (
    n1103,
    n828
  );


  buf
  g882
  (
    n1045,
    n869
  );


  buf
  g883
  (
    n914,
    n876
  );


  not
  g884
  (
    n1030,
    n886
  );


  buf
  g885
  (
    n942,
    n850
  );


  not
  g886
  (
    n1048,
    n831
  );


  buf
  g887
  (
    n1077,
    n875
  );


  not
  g888
  (
    n1102,
    n827
  );


  buf
  g889
  (
    n917,
    n831
  );


  buf
  g890
  (
    n980,
    n870
  );


  buf
  g891
  (
    n1004,
    n870
  );


  not
  g892
  (
    n964,
    n899
  );


  not
  g893
  (
    n953,
    n883
  );


  buf
  g894
  (
    n1104,
    n833
  );


  buf
  g895
  (
    n936,
    n852
  );


  buf
  g896
  (
    n934,
    n874
  );


  not
  g897
  (
    n1134,
    n836
  );


  not
  g898
  (
    n937,
    n837
  );


  buf
  g899
  (
    n935,
    n891
  );


  buf
  g900
  (
    n1044,
    n832
  );


  not
  g901
  (
    n1046,
    n849
  );


  not
  g902
  (
    n1023,
    n854
  );


  buf
  g903
  (
    n921,
    n884
  );


  buf
  g904
  (
    n1121,
    n830
  );


  not
  g905
  (
    n1109,
    n881
  );


  not
  g906
  (
    n927,
    n875
  );


  not
  g907
  (
    n1013,
    n859
  );


  buf
  g908
  (
    n1024,
    n874
  );


  not
  g909
  (
    n1073,
    n875
  );


  buf
  g910
  (
    n965,
    n898
  );


  buf
  g911
  (
    n975,
    n891
  );


  buf
  g912
  (
    n1116,
    n845
  );


  not
  g913
  (
    n926,
    n835
  );


  buf
  g914
  (
    n905,
    n885
  );


  buf
  g915
  (
    n1101,
    n829
  );


  buf
  g916
  (
    n990,
    n893
  );


  buf
  g917
  (
    n916,
    n874
  );


  buf
  g918
  (
    n955,
    n855
  );


  not
  g919
  (
    n946,
    n858
  );


  buf
  g920
  (
    n1113,
    n886
  );


  buf
  g921
  (
    n974,
    n863
  );


  buf
  g922
  (
    n987,
    n829
  );


  buf
  g923
  (
    n1087,
    n900
  );


  not
  g924
  (
    n1063,
    n899
  );


  not
  g925
  (
    n1090,
    n882
  );


  buf
  g926
  (
    n1043,
    n864
  );


  not
  g927
  (
    n1136,
    n827
  );


  not
  g928
  (
    n1095,
    n871
  );


  not
  g929
  (
    n910,
    n853
  );


  buf
  g930
  (
    n909,
    n882
  );


  not
  g931
  (
    n1032,
    n900
  );


  buf
  g932
  (
    n1082,
    n825
  );


  not
  g933
  (
    n991,
    n865
  );


  not
  g934
  (
    n1108,
    n880
  );


  not
  g935
  (
    n1000,
    n847
  );


  buf
  g936
  (
    n1100,
    n893
  );


  buf
  g937
  (
    n988,
    n848
  );


  not
  g938
  (
    n1010,
    n831
  );


  not
  g939
  (
    KeyWire_0_45,
    n894
  );


  not
  g940
  (
    n1006,
    n847
  );


  not
  g941
  (
    n1062,
    n840
  );


  not
  g942
  (
    n960,
    n879
  );


  not
  g943
  (
    n1114,
    n882
  );


  not
  g944
  (
    n985,
    n842
  );


  not
  g945
  (
    n1017,
    n853
  );


  not
  g946
  (
    n1015,
    n884
  );


  buf
  g947
  (
    n1098,
    n883
  );


  not
  g948
  (
    n1034,
    n843
  );


  not
  g949
  (
    n1089,
    n898
  );


  buf
  g950
  (
    n923,
    n861
  );


  not
  g951
  (
    n1022,
    n847
  );


  not
  g952
  (
    n996,
    n854
  );


  buf
  g953
  (
    n918,
    n895
  );


  buf
  g954
  (
    n1107,
    n856
  );


  not
  g955
  (
    n932,
    n840
  );


  buf
  g956
  (
    n939,
    n858
  );


  buf
  g957
  (
    n924,
    n866
  );


  not
  g958
  (
    n1132,
    n824
  );


  not
  g959
  (
    n1084,
    n892
  );


  not
  g960
  (
    n995,
    n872
  );


  buf
  g961
  (
    n994,
    n888
  );


  not
  g962
  (
    n969,
    n834
  );


  buf
  g963
  (
    n922,
    n886
  );


  not
  g964
  (
    n1038,
    n827
  );


  not
  g965
  (
    n1068,
    n847
  );


  not
  g966
  (
    n1129,
    n838
  );


  buf
  g967
  (
    n1092,
    n900
  );


  not
  g968
  (
    n954,
    n878
  );


  not
  g969
  (
    n1076,
    n854
  );


  buf
  g970
  (
    n1009,
    n880
  );


  buf
  g971
  (
    n1037,
    n834
  );


  not
  g972
  (
    n1067,
    n838
  );


  buf
  g973
  (
    n1131,
    n841
  );


  not
  g974
  (
    n1039,
    n888
  );


  not
  g975
  (
    KeyWire_0_0,
    n896
  );


  buf
  g976
  (
    n1056,
    n866
  );


  not
  g977
  (
    n1065,
    n860
  );


  buf
  g978
  (
    n943,
    n869
  );


  buf
  g979
  (
    n949,
    n876
  );


  buf
  g980
  (
    n1091,
    n825
  );


  not
  g981
  (
    n1083,
    n834
  );


  buf
  g982
  (
    n1072,
    n866
  );


  not
  g983
  (
    n1081,
    n857
  );


  not
  g984
  (
    n1016,
    n864
  );


  buf
  g985
  (
    KeyWire_0_13,
    n881
  );


  not
  g986
  (
    n1020,
    n872
  );


  not
  g987
  (
    n940,
    n884
  );


  buf
  g988
  (
    n1099,
    n867
  );


  not
  g989
  (
    n1019,
    n843
  );


  buf
  g990
  (
    n970,
    n860
  );


  buf
  g991
  (
    n1078,
    n858
  );


  buf
  g992
  (
    n1110,
    n835
  );


  not
  g993
  (
    n1025,
    n863
  );


  not
  g994
  (
    n956,
    n870
  );


  not
  g995
  (
    n915,
    n839
  );


  not
  g996
  (
    n1012,
    n849
  );


  buf
  g997
  (
    n1086,
    n855
  );


  not
  g998
  (
    n1050,
    n857
  );


  buf
  g999
  (
    KeyWire_0_60,
    n828
  );


  buf
  g1000
  (
    n930,
    n888
  );


  not
  g1001
  (
    n967,
    n841
  );


  not
  g1002
  (
    n1014,
    n839
  );


  buf
  g1003
  (
    n977,
    n885
  );


  buf
  g1004
  (
    n944,
    n869
  );


  buf
  g1005
  (
    n1120,
    n842
  );


  not
  g1006
  (
    n1027,
    n851
  );


  buf
  g1007
  (
    n1054,
    n857
  );


  not
  g1008
  (
    n925,
    n863
  );


  buf
  g1009
  (
    n973,
    n844
  );


  buf
  g1010
  (
    n1088,
    n892
  );


  buf
  g1011
  (
    n1031,
    n887
  );


  buf
  g1012
  (
    n1135,
    n889
  );


  not
  g1013
  (
    n1071,
    n896
  );


  not
  g1014
  (
    n1005,
    n892
  );


  not
  g1015
  (
    n1051,
    n826
  );


  buf
  g1016
  (
    n986,
    n862
  );


  not
  g1017
  (
    n1057,
    n825
  );


  buf
  g1018
  (
    n1026,
    n864
  );


  buf
  g1019
  (
    n962,
    n888
  );


  buf
  g1020
  (
    n904,
    n836
  );


  buf
  g1021
  (
    n913,
    n883
  );


  not
  g1022
  (
    n1128,
    n862
  );


  not
  g1023
  (
    n908,
    n862
  );


  not
  g1024
  (
    n1112,
    n894
  );


  not
  g1025
  (
    n1021,
    n881
  );


  not
  g1026
  (
    n1059,
    n880
  );


  buf
  g1027
  (
    n950,
    n890
  );


  not
  g1028
  (
    n1070,
    n828
  );


  buf
  g1029
  (
    n1061,
    n852
  );


  not
  g1030
  (
    n1003,
    n861
  );


  buf
  g1031
  (
    n1133,
    n851
  );


  not
  g1032
  (
    n1122,
    n855
  );


  buf
  g1033
  (
    n1058,
    n832
  );


  not
  g1034
  (
    n982,
    n881
  );


  not
  g1035
  (
    n1066,
    n846
  );


  not
  g1036
  (
    KeyWire_0_28,
    n860
  );


  buf
  g1037
  (
    n1130,
    n863
  );


  buf
  g1038
  (
    n1029,
    n832
  );


  not
  g1039
  (
    n966,
    n842
  );


  not
  g1040
  (
    n1096,
    n858
  );


  buf
  g1041
  (
    n1040,
    n830
  );


  buf
  g1042
  (
    n1125,
    n825
  );


  buf
  g1043
  (
    n1007,
    n845
  );


  not
  g1044
  (
    KeyWire_0_19,
    n828
  );


  not
  g1045
  (
    n1035,
    n831
  );


  buf
  g1046
  (
    n1047,
    n833
  );


  buf
  g1047
  (
    n938,
    n827
  );


  not
  g1048
  (
    n971,
    n845
  );


  buf
  g1049
  (
    n1097,
    n868
  );


  buf
  g1050
  (
    n947,
    n859
  );


  not
  g1051
  (
    n998,
    n878
  );


  buf
  g1052
  (
    KeyWire_0_24,
    n841
  );


  buf
  g1053
  (
    n931,
    n871
  );


  buf
  g1054
  (
    n963,
    n883
  );


  buf
  g1055
  (
    n929,
    n861
  );


  not
  g1056
  (
    n1085,
    n880
  );


  buf
  g1057
  (
    n928,
    n876
  );


  buf
  g1058
  (
    n1018,
    n879
  );


  buf
  g1059
  (
    n992,
    n829
  );


  buf
  g1060
  (
    n911,
    n865
  );


  buf
  g1061
  (
    n1002,
    n840
  );


  buf
  g1062
  (
    n983,
    n886
  );


  buf
  g1063
  (
    n1080,
    n870
  );


  not
  g1064
  (
    n902,
    n854
  );


  buf
  g1065
  (
    n957,
    n837
  );


  buf
  g1066
  (
    n1052,
    n877
  );


  not
  g1067
  (
    n1064,
    n887
  );


  or
  g1068
  (
    n1028,
    n832,
    n897,
    n873
  );


  and
  g1069
  (
    n1124,
    n879,
    n845,
    n868
  );


  nand
  g1070
  (
    n1117,
    n892,
    n850,
    n859
  );


  nand
  g1071
  (
    n1115,
    n853,
    n868,
    n890
  );


  or
  g1072
  (
    n1127,
    n885,
    n899,
    n830
  );


  xnor
  g1073
  (
    n1126,
    n876,
    n841,
    n871
  );


  xnor
  g1074
  (
    n1042,
    n871,
    n824,
    n855
  );


  nor
  g1075
  (
    KeyWire_0_18,
    n826,
    n866,
    n882
  );


  xnor
  g1076
  (
    n1093,
    n897,
    n838,
    n895
  );


  or
  g1077
  (
    n912,
    n872,
    n850,
    n826
  );


  nor
  g1078
  (
    n1055,
    n867,
    n824,
    n885
  );


  xnor
  g1079
  (
    n920,
    n838,
    n864,
    n891
  );


  xnor
  g1080
  (
    n903,
    n889,
    n853,
    n824
  );


  nand
  g1081
  (
    n958,
    n894,
    n896,
    n867
  );


  and
  g1082
  (
    n997,
    n835,
    n898,
    n851
  );


  nor
  g1083
  (
    n1123,
    n900,
    n873,
    n846
  );


  and
  g1084
  (
    n968,
    n893,
    n861,
    n844
  );


  nor
  g1085
  (
    n906,
    n830,
    n857,
    n867
  );


  xnor
  g1086
  (
    n1008,
    n856,
    n829,
    n891
  );


  and
  g1087
  (
    n1105,
    n865,
    n840,
    n899
  );


  nand
  g1088
  (
    n981,
    n842,
    n872,
    n833
  );


  nand
  g1089
  (
    n933,
    n898,
    n895,
    n890
  );


  xnor
  g1090
  (
    n993,
    n848,
    n879,
    n859
  );


  nor
  g1091
  (
    n1060,
    n865,
    n836,
    n896
  );


  xnor
  g1092
  (
    n952,
    n848,
    n837,
    n849
  );


  xor
  g1093
  (
    n979,
    n874,
    n856,
    n893
  );


  nand
  g1094
  (
    n1119,
    n839,
    n846,
    n843
  );


  nor
  g1095
  (
    n1094,
    n895,
    n887,
    n843
  );


  and
  g1096
  (
    n951,
    n862,
    n873
  );


  xnor
  g1097
  (
    n1079,
    n850,
    n836,
    n839
  );


  or
  g1098
  (
    n1111,
    n897,
    n884,
    n833
  );


  xor
  g1099
  (
    n901,
    n877,
    n889,
    n897
  );


  xor
  g1100
  (
    n984,
    n834,
    n852,
    n877
  );


  xnor
  g1101
  (
    n961,
    n848,
    n846,
    n887
  );


  and
  g1102
  (
    n1069,
    n868,
    n835,
    n860
  );


  or
  g1103
  (
    n978,
    n877,
    n852,
    n878
  );


  buf
  g1104
  (
    n1161,
    n1002
  );


  buf
  g1105
  (
    n1313,
    n954
  );


  not
  g1106
  (
    n1200,
    n925
  );


  buf
  g1107
  (
    n1269,
    n1008
  );


  buf
  g1108
  (
    n1204,
    n957
  );


  buf
  g1109
  (
    n1210,
    n916
  );


  buf
  g1110
  (
    n1265,
    n1024
  );


  buf
  g1111
  (
    n1159,
    n949
  );


  not
  g1112
  (
    n1237,
    n1004
  );


  not
  g1113
  (
    n1244,
    n901
  );


  not
  g1114
  (
    n1256,
    n1015
  );


  not
  g1115
  (
    n1199,
    n965
  );


  not
  g1116
  (
    n1271,
    n999
  );


  not
  g1117
  (
    n1208,
    n920
  );


  not
  g1118
  (
    n1314,
    n987
  );


  buf
  g1119
  (
    n1287,
    n994
  );


  buf
  g1120
  (
    n1299,
    n950
  );


  buf
  g1121
  (
    n1290,
    n1015
  );


  not
  g1122
  (
    n1266,
    n948
  );


  not
  g1123
  (
    n1267,
    n1020
  );


  buf
  g1124
  (
    n1203,
    n972
  );


  buf
  g1125
  (
    n1138,
    n956
  );


  buf
  g1126
  (
    n1273,
    n944
  );


  buf
  g1127
  (
    n1140,
    n1027
  );


  not
  g1128
  (
    n1195,
    n951
  );


  buf
  g1129
  (
    n1181,
    n970
  );


  not
  g1130
  (
    n1320,
    n990
  );


  not
  g1131
  (
    n1231,
    n955
  );


  buf
  g1132
  (
    n1205,
    n999
  );


  buf
  g1133
  (
    n1250,
    n1022
  );


  buf
  g1134
  (
    n1167,
    n1010
  );


  buf
  g1135
  (
    n1225,
    n921
  );


  buf
  g1136
  (
    n1221,
    n924
  );


  buf
  g1137
  (
    n1189,
    n1026
  );


  buf
  g1138
  (
    n1169,
    n1025
  );


  not
  g1139
  (
    n1139,
    n917
  );


  not
  g1140
  (
    n1170,
    n1016
  );


  buf
  g1141
  (
    KeyWire_0_53,
    n984
  );


  buf
  g1142
  (
    n1303,
    n1006
  );


  not
  g1143
  (
    n1247,
    n1021
  );


  not
  g1144
  (
    n1270,
    n1007
  );


  buf
  g1145
  (
    n1274,
    n950
  );


  not
  g1146
  (
    n1281,
    n941
  );


  not
  g1147
  (
    n1277,
    n1005
  );


  not
  g1148
  (
    n1318,
    n977
  );


  buf
  g1149
  (
    n1248,
    n972
  );


  buf
  g1150
  (
    n1178,
    n964
  );


  not
  g1151
  (
    n1311,
    n1014
  );


  not
  g1152
  (
    n1147,
    n974
  );


  not
  g1153
  (
    n1211,
    n976
  );


  not
  g1154
  (
    n1259,
    n1019
  );


  buf
  g1155
  (
    n1152,
    n958
  );


  not
  g1156
  (
    n1184,
    n996
  );


  buf
  g1157
  (
    n1307,
    n982
  );


  buf
  g1158
  (
    n1213,
    n988
  );


  buf
  g1159
  (
    n1230,
    n959
  );


  not
  g1160
  (
    n1218,
    n1015
  );


  not
  g1161
  (
    n1212,
    n937
  );


  not
  g1162
  (
    n1272,
    n989
  );


  buf
  g1163
  (
    n1235,
    n1002
  );


  not
  g1164
  (
    n1193,
    n967
  );


  not
  g1165
  (
    KeyWire_0_31,
    n997
  );


  buf
  g1166
  (
    n1188,
    n970
  );


  not
  g1167
  (
    n1260,
    n996
  );


  not
  g1168
  (
    n1223,
    n986
  );


  not
  g1169
  (
    n1162,
    n974
  );


  buf
  g1170
  (
    n1252,
    n982
  );


  not
  g1171
  (
    n1308,
    n966
  );


  not
  g1172
  (
    n1141,
    n1003
  );


  buf
  g1173
  (
    n1217,
    n980
  );


  buf
  g1174
  (
    n1191,
    n994
  );


  not
  g1175
  (
    n1295,
    n1014
  );


  not
  g1176
  (
    n1183,
    n978
  );


  not
  g1177
  (
    n1192,
    n980
  );


  not
  g1178
  (
    n1306,
    n968
  );


  not
  g1179
  (
    n1196,
    n1013
  );


  not
  g1180
  (
    n1245,
    n968
  );


  buf
  g1181
  (
    n1209,
    n974
  );


  buf
  g1182
  (
    n1142,
    n981
  );


  not
  g1183
  (
    n1317,
    n977
  );


  not
  g1184
  (
    n1278,
    n906
  );


  buf
  g1185
  (
    n1238,
    n950
  );


  buf
  g1186
  (
    n1155,
    n971
  );


  buf
  g1187
  (
    n1156,
    n969
  );


  not
  g1188
  (
    n1175,
    n965
  );


  not
  g1189
  (
    n1243,
    n1028
  );


  not
  g1190
  (
    n1216,
    n904
  );


  buf
  g1191
  (
    n1309,
    n960
  );


  not
  g1192
  (
    n1282,
    n984
  );


  not
  g1193
  (
    n1145,
    n982
  );


  buf
  g1194
  (
    n1240,
    n967
  );


  buf
  g1195
  (
    KeyWire_0_5,
    n1011
  );


  buf
  g1196
  (
    n1286,
    n910
  );


  buf
  g1197
  (
    KeyWire_0_37,
    n962
  );


  buf
  g1198
  (
    n1284,
    n949
  );


  not
  g1199
  (
    n1239,
    n965
  );


  buf
  g1200
  (
    n1214,
    n960
  );


  buf
  g1201
  (
    n1215,
    n964
  );


  buf
  g1202
  (
    n1293,
    n1009
  );


  not
  g1203
  (
    n1224,
    n1024
  );


  not
  g1204
  (
    n1319,
    n973
  );


  not
  g1205
  (
    n1268,
    n1004
  );


  buf
  g1206
  (
    n1279,
    n995
  );


  not
  g1207
  (
    n1264,
    n983
  );


  buf
  g1208
  (
    n1174,
    n940
  );


  not
  g1209
  (
    n1297,
    n955
  );


  not
  g1210
  (
    n1305,
    n1028
  );


  buf
  g1211
  (
    n1202,
    n1008
  );


  not
  g1212
  (
    n1197,
    n934
  );


  not
  g1213
  (
    n1187,
    n918
  );


  buf
  g1214
  (
    n1190,
    n1009
  );


  buf
  g1215
  (
    n1226,
    n1012
  );


  not
  g1216
  (
    n1146,
    n993
  );


  buf
  g1217
  (
    n1285,
    n1013
  );


  not
  g1218
  (
    n1166,
    n963
  );


  buf
  g1219
  (
    n1158,
    n1000
  );


  not
  g1220
  (
    n1144,
    n939
  );


  buf
  g1221
  (
    KeyWire_0_40,
    n973
  );


  buf
  g1222
  (
    KeyWire_0_36,
    n948
  );


  not
  g1223
  (
    n1227,
    n936
  );


  not
  g1224
  (
    n1219,
    n952
  );


  buf
  g1225
  (
    n1257,
    n1001
  );


  buf
  g1226
  (
    n1310,
    n955
  );


  not
  g1227
  (
    n1291,
    n1022
  );


  buf
  g1228
  (
    n1229,
    n960
  );


  buf
  g1229
  (
    n1241,
    n947
  );


  not
  g1230
  (
    n1300,
    n962
  );


  not
  g1231
  (
    n1164,
    n1019
  );


  buf
  g1232
  (
    n1173,
    n972
  );


  not
  g1233
  (
    n1312,
    n945
  );


  buf
  g1234
  (
    n1228,
    n979
  );


  not
  g1235
  (
    n1176,
    n946
  );


  not
  g1236
  (
    n1222,
    n966
  );


  buf
  g1237
  (
    n1283,
    n964
  );


  not
  g1238
  (
    n1302,
    n923
  );


  not
  g1239
  (
    n1246,
    n971
  );


  buf
  g1240
  (
    n1316,
    n975
  );


  buf
  g1241
  (
    n1179,
    n913
  );


  not
  g1242
  (
    n1149,
    n952
  );


  buf
  g1243
  (
    n1255,
    n1028
  );


  buf
  g1244
  (
    n1153,
    n1001
  );


  not
  g1245
  (
    n1150,
    n1018
  );


  not
  g1246
  (
    n1165,
    n922
  );


  not
  g1247
  (
    n1160,
    n1006
  );


  buf
  g1248
  (
    n1180,
    n987
  );


  buf
  g1249
  (
    n1163,
    n1012
  );


  buf
  g1250
  (
    KeyWire_0_1,
    n988
  );


  buf
  g1251
  (
    n1198,
    n958
  );


  xnor
  g1252
  (
    n1233,
    n1002,
    n980,
    n958,
    n1011
  );


  nand
  g1253
  (
    n1206,
    n1016,
    n938,
    n930,
    n990
  );


  and
  g1254
  (
    n1171,
    n992,
    n951,
    n966,
    n942
  );


  xnor
  g1255
  (
    n1294,
    n1027,
    n1025,
    n967,
    n951
  );


  nand
  g1256
  (
    n1185,
    n932,
    n970,
    n1026,
    n973
  );


  nor
  g1257
  (
    n1143,
    n997,
    n949,
    n1007,
    n911
  );


  xor
  g1258
  (
    n1232,
    n1000,
    n909,
    n962,
    n1020
  );


  and
  g1259
  (
    KeyWire_0_34,
    n943,
    n985,
    n1010
  );


  or
  g1260
  (
    n1194,
    n902,
    n1004,
    n931,
    n998
  );


  nor
  g1261
  (
    n1148,
    n991,
    n971,
    n975,
    n978
  );


  nor
  g1262
  (
    n1263,
    n956,
    n1012,
    n912,
    n1014
  );


  or
  g1263
  (
    n1220,
    n1020,
    n991,
    n915,
    n1024
  );


  nor
  g1264
  (
    n1151,
    n1005,
    n984,
    n954,
    n1021
  );


  xor
  g1265
  (
    n1280,
    n978,
    n983,
    n995,
    n908
  );


  xor
  g1266
  (
    n1292,
    n1017,
    n981,
    n1023,
    n992
  );


  or
  g1267
  (
    n1234,
    n1011,
    n919,
    n1013,
    n947
  );


  xor
  g1268
  (
    n1288,
    n1027,
    n990,
    n986,
    n963
  );


  or
  g1269
  (
    n1172,
    n1025,
    n963,
    n1021,
    n988
  );


  nand
  g1270
  (
    n1186,
    n969,
    n985,
    n1001,
    n959
  );


  xor
  g1271
  (
    n1242,
    n979,
    n1023,
    n989,
    n986
  );


  xor
  g1272
  (
    n1251,
    n1018,
    n935,
    n961,
    n1017
  );


  nand
  g1273
  (
    n1207,
    n953,
    n1008,
    n961,
    n903
  );


  xnor
  g1274
  (
    n1201,
    n928,
    n959,
    n1003,
    n969
  );


  xor
  g1275
  (
    n1258,
    n961,
    n948,
    n927,
    n933
  );


  and
  g1276
  (
    n1296,
    n1009,
    n987,
    n1010,
    n1017
  );


  xor
  g1277
  (
    n1254,
    n953,
    n956,
    n977,
    n1007
  );


  nor
  g1278
  (
    n1177,
    n905,
    n993,
    n996,
    n976
  );


  xor
  g1279
  (
    n1182,
    n991,
    n1019,
    n1006,
    n995
  );


  or
  g1280
  (
    n1289,
    n914,
    n979,
    n954,
    n953
  );


  and
  g1281
  (
    n1236,
    n993,
    n997,
    n968,
    n976
  );


  nor
  g1282
  (
    n1315,
    n1026,
    n957,
    n981,
    n998
  );


  and
  g1283
  (
    n1168,
    n1005,
    n999,
    n1023,
    n1016
  );


  or
  g1284
  (
    n1154,
    n1022,
    n907,
    n992,
    n998
  );


  xor
  g1285
  (
    n1276,
    n957,
    n989,
    n926,
    n947
  );


  nand
  g1286
  (
    KeyWire_0_9,
    n1000,
    n952,
    n929,
    n975
  );


  xnor
  g1287
  (
    n1262,
    n983,
    n1018,
    n994,
    n1003
  );


  xor
  g1288
  (
    n1327,
    n1144,
    n1137
  );


  nand
  g1289
  (
    n1330,
    n618,
    n1141,
    n619,
    n1144
  );


  nor
  g1290
  (
    n1324,
    n1144,
    n618,
    n1140
  );


  and
  g1291
  (
    n1326,
    n1137,
    n619,
    n1138,
    n1139
  );


  xor
  g1292
  (
    n1325,
    n618,
    n1141,
    n1139,
    n1143
  );


  xor
  g1293
  (
    n1323,
    n1142,
    n1138,
    n1137
  );


  xor
  g1294
  (
    n1321,
    n1140,
    n1142,
    n1143
  );


  xor
  g1295
  (
    n1322,
    n1139,
    n619,
    n1140
  );


  and
  g1296
  (
    n1329,
    n1144,
    n1143,
    n1138
  );


  and
  g1297
  (
    n1328,
    n1139,
    n1142,
    n1141
  );


  not
  g1298
  (
    n1355,
    n1329
  );


  not
  g1299
  (
    n1347,
    n1321
  );


  not
  g1300
  (
    n1340,
    n622
  );


  not
  g1301
  (
    n1341,
    n1329
  );


  not
  g1302
  (
    n1337,
    n621
  );


  not
  g1303
  (
    n1351,
    n1322
  );


  not
  g1304
  (
    n1354,
    n620
  );


  not
  g1305
  (
    n1336,
    n1329
  );


  not
  g1306
  (
    n1333,
    n1324
  );


  not
  g1307
  (
    n1343,
    n1326
  );


  not
  g1308
  (
    n1353,
    n1324
  );


  nor
  g1309
  (
    n1335,
    n621,
    n620
  );


  or
  g1310
  (
    n1349,
    n1327,
    n1330
  );


  xor
  g1311
  (
    n1334,
    n1325,
    n621
  );


  xnor
  g1312
  (
    n1346,
    n1326,
    n1323
  );


  nor
  g1313
  (
    KeyWire_0_25,
    n1323,
    n623
  );


  xor
  g1314
  (
    n1350,
    n1324,
    n620
  );


  not
  g1315
  (
    n1348,
    n1328
  );


  nand
  g1316
  (
    n1357,
    n1322,
    n622
  );


  or
  g1317
  (
    n1356,
    n1330,
    n622
  );


  and
  g1318
  (
    n1352,
    n623,
    n1323
  );


  and
  g1319
  (
    n1342,
    n622,
    n1327
  );


  nand
  g1320
  (
    n1345,
    n620,
    n623
  );


  not
  g1321
  (
    n1339,
    n1325
  );


  nor
  g1322
  (
    n1344,
    n1327,
    n1330
  );


  and
  g1323
  (
    n1332,
    n1326,
    n1328
  );


  xnor
  g1324
  (
    n1338,
    n621,
    n623
  );


  or
  g1325
  (
    n1407,
    n1031,
    n1046,
    n1089,
    n1349
  );


  nand
  g1326
  (
    n1413,
    n1352,
    n1118,
    n1338,
    n1111
  );


  nand
  g1327
  (
    n1417,
    n1115,
    n1133,
    n1124,
    n1331
  );


  xnor
  g1328
  (
    n1370,
    n1077,
    n1033,
    n1078,
    n1350
  );


  xnor
  g1329
  (
    n1458,
    n1119,
    n1122,
    n1332,
    n1045
  );


  xnor
  g1330
  (
    n1420,
    n1030,
    n1091,
    n1349,
    n1081
  );


  nor
  g1331
  (
    n1406,
    n1052,
    n1029,
    n1104,
    n1091
  );


  xnor
  g1332
  (
    n1388,
    n1045,
    n1114,
    n1355,
    n1034
  );


  or
  g1333
  (
    n1375,
    n1047,
    n1352,
    n1335,
    n1046
  );


  xnor
  g1334
  (
    n1429,
    n1047,
    n1050,
    n1065,
    n1097
  );


  xor
  g1335
  (
    n1409,
    n1096,
    n1094,
    n1069,
    n1334
  );


  xor
  g1336
  (
    n1428,
    n1135,
    n1333,
    n1105,
    n1115
  );


  xor
  g1337
  (
    n1399,
    n1029,
    n1031,
    n1354,
    n1037
  );


  nor
  g1338
  (
    n1426,
    n1051,
    n1039,
    n1065,
    n1083
  );


  or
  g1339
  (
    n1461,
    n1340,
    n1055,
    n1088,
    n1080
  );


  or
  g1340
  (
    n1395,
    n1341,
    n1096,
    n1042,
    n1052
  );


  xor
  g1341
  (
    n1460,
    n1034,
    n1095,
    n1111,
    n1042
  );


  or
  g1342
  (
    n1425,
    n1341,
    n1115,
    n1036,
    n1351
  );


  nand
  g1343
  (
    KeyWire_0_48,
    n1133,
    n1039,
    n1355,
    n1057
  );


  or
  g1344
  (
    n1361,
    n1077,
    n1342,
    n1356,
    n1099
  );


  and
  g1345
  (
    n1368,
    n1067,
    n1353,
    n1076,
    n1113
  );


  nand
  g1346
  (
    n1359,
    n1095,
    n1030,
    n1337,
    n1097
  );


  xnor
  g1347
  (
    n1394,
    n1051,
    n1057,
    n1100,
    n1331
  );


  nor
  g1348
  (
    n1367,
    n1036,
    n1357,
    n1092,
    n1106
  );


  and
  g1349
  (
    n1442,
    n1032,
    n1041,
    n1117,
    n1100
  );


  nor
  g1350
  (
    n1435,
    n1073,
    n1043,
    n1072,
    n1081
  );


  or
  g1351
  (
    n1463,
    n1064,
    n1074,
    n1129,
    n1132
  );


  xor
  g1352
  (
    n1404,
    n1113,
    n1342,
    n1056,
    n1345
  );


  nor
  g1353
  (
    n1389,
    n1054,
    n1134,
    n1118,
    n1086
  );


  and
  g1354
  (
    n1424,
    n1340,
    n1056,
    n1051,
    n1071
  );


  xnor
  g1355
  (
    n1465,
    n1112,
    n1053,
    n1049,
    n1069
  );


  xor
  g1356
  (
    n1434,
    n1338,
    n1087,
    n1075,
    n1062
  );


  and
  g1357
  (
    n1448,
    n1107,
    n1356,
    n1063,
    n1072
  );


  nand
  g1358
  (
    n1363,
    n1092,
    n1107,
    n1354,
    n1112
  );


  and
  g1359
  (
    n1390,
    n1355,
    n1354,
    n1098,
    n1333
  );


  xnor
  g1360
  (
    n1439,
    n1339,
    n1356,
    n1073,
    n1113
  );


  and
  g1361
  (
    n1455,
    n1352,
    n1120,
    n1049,
    n1080
  );


  nand
  g1362
  (
    n1400,
    n1130,
    n1053,
    n1126,
    n1111
  );


  and
  g1363
  (
    n1438,
    n1333,
    n1343,
    n1074,
    n1126
  );


  or
  g1364
  (
    n1408,
    n1039,
    n1345,
    n1081,
    n1066
  );


  xor
  g1365
  (
    n1436,
    n1101,
    n1357,
    n1114,
    n1035
  );


  xor
  g1366
  (
    n1402,
    n1339,
    n1106,
    n1105,
    n1341
  );


  and
  g1367
  (
    n1380,
    n1344,
    n1082,
    n1129,
    n1078
  );


  nor
  g1368
  (
    n1393,
    n1063,
    n1088,
    n1060,
    n1135
  );


  nand
  g1369
  (
    n1373,
    n1342,
    n1128,
    n1134,
    n1083
  );


  nor
  g1370
  (
    n1358,
    n1066,
    n1336,
    n1350,
    n1123
  );


  nor
  g1371
  (
    n1385,
    n1037,
    n1048,
    n1102,
    n1333
  );


  or
  g1372
  (
    n1397,
    n1357,
    n1059,
    n1101,
    n1104
  );


  nor
  g1373
  (
    n1437,
    n1122,
    n1121,
    n1336,
    n1110
  );


  xnor
  g1374
  (
    n1376,
    n1353,
    n1132,
    n1053,
    n1352
  );


  xor
  g1375
  (
    n1410,
    n1110,
    n1079,
    n1106,
    n1088
  );


  nand
  g1376
  (
    n1382,
    n1045,
    n1033,
    n1334,
    n1340
  );


  xnor
  g1377
  (
    KeyWire_0_6,
    n1085,
    n1048,
    n1092,
    n1063
  );


  xnor
  g1378
  (
    n1365,
    n1084,
    n1054,
    n1133,
    n1046
  );


  xor
  g1379
  (
    n1430,
    n1055,
    n1054,
    n1061,
    n1337
  );


  and
  g1380
  (
    n1418,
    n1040,
    n1131,
    n1348,
    n1071
  );


  or
  g1381
  (
    n1432,
    n1125,
    n1072,
    n1136,
    n1047
  );


  nor
  g1382
  (
    n1415,
    n1085,
    n1343,
    n1079,
    n1044
  );


  nor
  g1383
  (
    n1423,
    n1351,
    n1077,
    n1061,
    n1108
  );


  xnor
  g1384
  (
    KeyWire_0_54,
    n1043,
    n1127,
    n1056,
    n1068
  );


  nor
  g1385
  (
    n1391,
    n1120,
    n1075,
    n1347,
    n1087
  );


  xor
  g1386
  (
    n1371,
    n1031,
    n1094,
    n1059,
    n1357
  );


  or
  g1387
  (
    n1366,
    n1084,
    n1070,
    n1030,
    n1110
  );


  nand
  g1388
  (
    n1459,
    n1058,
    n1345,
    n1082,
    n1071
  );


  or
  g1389
  (
    n1405,
    n1335,
    n1349,
    n1093,
    n1044
  );


  and
  g1390
  (
    n1362,
    n1347,
    n1351,
    n1040,
    n1038
  );


  and
  g1391
  (
    n1384,
    n1344,
    n1350,
    n1346,
    n1332
  );


  nand
  g1392
  (
    n1447,
    n1065,
    n1109,
    n1100,
    n1080
  );


  xor
  g1393
  (
    n1414,
    n1089,
    n1086,
    n1331
  );


  nor
  g1394
  (
    n1422,
    n1085,
    n1116,
    n1124,
    n1332
  );


  xnor
  g1395
  (
    n1457,
    n1097,
    n1340,
    n1339,
    n1347
  );


  or
  g1396
  (
    n1374,
    n1076,
    n1116,
    n1135,
    n1049
  );


  xor
  g1397
  (
    n1450,
    n1339,
    n1108,
    n1082,
    n1037
  );


  xor
  g1398
  (
    n1427,
    n1074,
    n1120,
    n1123,
    n1132
  );


  and
  g1399
  (
    n1387,
    n1067,
    n1079,
    n1032,
    n1344
  );


  xnor
  g1400
  (
    n1445,
    n1035,
    n1338,
    n1335,
    n1036
  );


  nor
  g1401
  (
    n1360,
    n1337,
    n1058,
    n1109,
    n1348
  );


  nor
  g1402
  (
    n1377,
    n1107,
    n1032,
    n1353,
    n1351
  );


  and
  g1403
  (
    n1378,
    n1114,
    n1091,
    n1078,
    n1112
  );


  and
  g1404
  (
    n1443,
    n1346,
    n1338,
    n1042,
    n1127
  );


  or
  g1405
  (
    n1398,
    n1069,
    n1104,
    n1126,
    n1064
  );


  or
  g1406
  (
    n1383,
    n1098,
    n1093,
    n1128,
    n1050
  );


  nor
  g1407
  (
    n1396,
    n1062,
    n1070,
    n1068,
    n1103
  );


  nor
  g1408
  (
    n1386,
    n1073,
    n1130,
    n1127,
    n1060
  );


  nand
  g1409
  (
    n1419,
    n1117,
    n1109,
    n1119,
    n1343
  );


  nand
  g1410
  (
    n1454,
    n1070,
    n1125,
    n1343,
    n1121
  );


  and
  g1411
  (
    n1431,
    n1044,
    n1076,
    n1347,
    n1061
  );


  nor
  g1412
  (
    n1421,
    n1336,
    n1119,
    n1108,
    n1349
  );


  nand
  g1413
  (
    n1369,
    n1087,
    n1346,
    n1355,
    n1066
  );


  nor
  g1414
  (
    n1392,
    n1062,
    n1083,
    n1121,
    n1034
  );


  nor
  g1415
  (
    n1444,
    n1332,
    n1089,
    n1353,
    n1341
  );


  xnor
  g1416
  (
    n1449,
    n1094,
    n1356,
    n1090,
    n1103
  );


  xnor
  g1417
  (
    n1412,
    n1075,
    n1090,
    n1342,
    n1348
  );


  or
  g1418
  (
    n1411,
    n1344,
    n1334,
    n1043,
    n1093
  );


  xor
  g1419
  (
    n1452,
    n1099,
    n1116,
    n1334,
    n1038
  );


  nor
  g1420
  (
    n1446,
    n1348,
    n1122,
    n1128,
    n1068
  );


  nand
  g1421
  (
    n1364,
    n1331,
    n1131,
    n1059,
    n1124
  );


  and
  g1422
  (
    n1441,
    n1134,
    n1337,
    n1048,
    n1102
  );


  nor
  g1423
  (
    n1379,
    n1350,
    n1095,
    n1029,
    n1354
  );


  nand
  g1424
  (
    n1403,
    n1058,
    n1057,
    n1035,
    n1336
  );


  nor
  g1425
  (
    KeyWire_0_58,
    n1130,
    n1090,
    n1038,
    n1136
  );


  or
  g1426
  (
    n1451,
    n1345,
    n1067,
    n1052,
    n1117
  );


  or
  g1427
  (
    n1372,
    n1040,
    n1041,
    n1098,
    n1102
  );


  or
  g1428
  (
    n1401,
    n1064,
    n1125,
    n1033,
    n1105
  );


  or
  g1429
  (
    n1433,
    n1123,
    n1041,
    n1055,
    n1060
  );


  nor
  g1430
  (
    n1453,
    n1099,
    n1096,
    n1101,
    n1050
  );


  nand
  g1431
  (
    n1456,
    n1136,
    n1103,
    n1118,
    n1346
  );


  xor
  g1432
  (
    n1381,
    n1131,
    n1084,
    n1335,
    n1129
  );


  xor
  g1433
  (
    n1492,
    n1309,
    n1386,
    n1176,
    n1368
  );


  and
  g1434
  (
    n1635,
    n1243,
    n1156,
    n1405,
    n1225
  );


  nor
  g1435
  (
    n1674,
    n1269,
    n1165,
    n1389,
    n1300
  );


  xor
  g1436
  (
    n1606,
    n1410,
    n1188,
    n1183,
    n1320
  );


  xor
  g1437
  (
    KeyWire_0_39,
    n1412,
    n1158,
    n1408,
    n1162
  );


  nor
  g1438
  (
    n1569,
    n1388,
    n1208,
    n1166,
    n1191
  );


  xnor
  g1439
  (
    n1658,
    n1164,
    n1396,
    n1408,
    n1233
  );


  and
  g1440
  (
    n1732,
    n1446,
    n1419,
    n1364,
    n1173
  );


  nand
  g1441
  (
    n1709,
    n1371,
    n1387,
    n1456,
    n1214
  );


  nor
  g1442
  (
    n1718,
    n1421,
    n1377,
    n1428,
    n1396
  );


  xor
  g1443
  (
    n1708,
    n1427,
    n1299,
    n1435,
    n1159
  );


  and
  g1444
  (
    n1679,
    n1283,
    n1165,
    n1213,
    n1223
  );


  xnor
  g1445
  (
    n1628,
    n1207,
    n1225,
    n1193,
    n1295
  );


  or
  g1446
  (
    n1530,
    n1254,
    n1278,
    n1184,
    n1221
  );


  nor
  g1447
  (
    n1731,
    n1229,
    n1221,
    n1191,
    n1403
  );


  xor
  g1448
  (
    n1644,
    n1284,
    n1196,
    n1364,
    n1269
  );


  nand
  g1449
  (
    n1643,
    n1392,
    n1393,
    n1219,
    n1367
  );


  nor
  g1450
  (
    n1648,
    n1452,
    n1263,
    n1284,
    n1174
  );


  xor
  g1451
  (
    n1553,
    n1155,
    n1275,
    n1378,
    n1460
  );


  nor
  g1452
  (
    n1476,
    n1282,
    n1414,
    n1251,
    n1227
  );


  xor
  g1453
  (
    n1595,
    n1205,
    n1189,
    n1217,
    n1230
  );


  nand
  g1454
  (
    n1626,
    n1405,
    n1275,
    n1433,
    n1461
  );


  or
  g1455
  (
    n1676,
    n1223,
    n1306,
    n1457,
    n1280
  );


  nor
  g1456
  (
    KeyWire_0_38,
    n1448,
    n1398,
    n1232,
    n1443
  );


  or
  g1457
  (
    n1474,
    n1203,
    n1287,
    n1210,
    n1265
  );


  and
  g1458
  (
    n1570,
    n1161,
    n1237,
    n1163,
    n1288
  );


  and
  g1459
  (
    n1488,
    n1215,
    n1315,
    n1159,
    n1177
  );


  or
  g1460
  (
    n1480,
    n1313,
    n1423,
    n1372,
    n1259
  );


  xnor
  g1461
  (
    n1712,
    n1434,
    n1222,
    n1408
  );


  nor
  g1462
  (
    KeyWire_0_27,
    n1152,
    n1160,
    n1239,
    n1434
  );


  nand
  g1463
  (
    n1498,
    n1213,
    n1418,
    n1280,
    n1463
  );


  and
  g1464
  (
    n1733,
    n1264,
    n1238,
    n1302,
    n1396
  );


  xnor
  g1465
  (
    n1526,
    n1366,
    n1365,
    n1371,
    n1190
  );


  nand
  g1466
  (
    n1486,
    n1269,
    n1273,
    n1169,
    n1221
  );


  or
  g1467
  (
    n1680,
    n1267,
    n1445,
    n1255,
    n1270
  );


  xnor
  g1468
  (
    KeyWire_0_8,
    n1171,
    n1305,
    n1169,
    n1365
  );


  xnor
  g1469
  (
    n1605,
    n1436,
    n1149,
    n1258,
    n1264
  );


  xnor
  g1470
  (
    n1616,
    n1438,
    n1432,
    n1213,
    n1274
  );


  or
  g1471
  (
    n1721,
    n1242,
    n1206,
    n1170,
    n1260
  );


  xnor
  g1472
  (
    n1537,
    n1370,
    n1226,
    n1395,
    n1425
  );


  xor
  g1473
  (
    n1525,
    n1229,
    n1279,
    n1305,
    n1307
  );


  or
  g1474
  (
    n1522,
    n1383,
    n1178,
    n1308,
    n1365
  );


  and
  g1475
  (
    n1466,
    n1463,
    n1146,
    n1410,
    n1171
  );


  xnor
  g1476
  (
    n1631,
    n1172,
    n1194,
    n1294,
    n1367
  );


  xor
  g1477
  (
    n1617,
    n1450,
    n1256,
    n1184,
    n1230
  );


  or
  g1478
  (
    n1566,
    n1294,
    n1317,
    n1179,
    n1235
  );


  or
  g1479
  (
    n1707,
    n1271,
    n1154,
    n1204,
    n1421
  );


  nand
  g1480
  (
    n1582,
    n1298,
    n1307,
    n1391,
    n1458
  );


  nand
  g1481
  (
    n1729,
    n1385,
    n1193,
    n1219,
    n1303
  );


  and
  g1482
  (
    n1510,
    n1422,
    n1389,
    n1415,
    n1236
  );


  or
  g1483
  (
    n1573,
    n1228,
    n1406,
    n1385,
    n1367
  );


  and
  g1484
  (
    n1501,
    n1370,
    n1219,
    n1249,
    n1463
  );


  xnor
  g1485
  (
    n1654,
    n1151,
    n1218,
    n1254,
    n1287
  );


  and
  g1486
  (
    n1613,
    n1286,
    n1284,
    n1262,
    n1186
  );


  nor
  g1487
  (
    n1650,
    n1261,
    n1178,
    n1364,
    n1215
  );


  xnor
  g1488
  (
    n1506,
    n1387,
    n1411,
    n1442,
    n1214
  );


  nand
  g1489
  (
    n1653,
    n1314,
    n1316,
    n1285,
    n1290
  );


  xor
  g1490
  (
    n1604,
    n1288,
    n1232,
    n1462,
    n1464
  );


  xor
  g1491
  (
    n1568,
    n1292,
    n1456,
    n1305,
    n1359
  );


  or
  g1492
  (
    n1663,
    n1295,
    n1234,
    n1210,
    n1374
  );


  xor
  g1493
  (
    n1693,
    n1285,
    n1206,
    n1209,
    n1369
  );


  nor
  g1494
  (
    n1503,
    n1265,
    n1311,
    n1159,
    n1361
  );


  xor
  g1495
  (
    n1695,
    n1382,
    n1151,
    n1420,
    n1215
  );


  and
  g1496
  (
    n1562,
    n1269,
    n1267,
    n1191,
    n1455
  );


  nand
  g1497
  (
    n1584,
    n1412,
    n1390,
    n1152,
    n1403
  );


  or
  g1498
  (
    n1642,
    n1245,
    n1157,
    n1224,
    n1412
  );


  xor
  g1499
  (
    n1580,
    n1313,
    n1263,
    n1243,
    n1418
  );


  nand
  g1500
  (
    n1741,
    n1411,
    n1459,
    n1448,
    n1180
  );


  xor
  g1501
  (
    n1728,
    n1267,
    n1306,
    n1423,
    n1261
  );


  nand
  g1502
  (
    n1598,
    n1416,
    n1310,
    n1237,
    n1432
  );


  xnor
  g1503
  (
    n1597,
    n1319,
    n1409,
    n1196,
    n1173
  );


  or
  g1504
  (
    n1711,
    n1158,
    n1379,
    n1254,
    n1207
  );


  and
  g1505
  (
    n1565,
    n1318,
    n1194,
    n1465,
    n1175
  );


  xor
  g1506
  (
    n1685,
    n1451,
    n1277,
    n1177,
    n1402
  );


  and
  g1507
  (
    n1502,
    n1443,
    n1274,
    n1198,
    n1176
  );


  or
  g1508
  (
    n1509,
    n1309,
    n1247,
    n1196,
    n1448
  );


  xor
  g1509
  (
    n1484,
    n1435,
    n1282,
    n1259
  );


  xor
  g1510
  (
    n1673,
    n1449,
    n1414,
    n1233,
    n1444
  );


  or
  g1511
  (
    n1657,
    n1164,
    n1223,
    n1256,
    n1371
  );


  nor
  g1512
  (
    n1725,
    n1234,
    n1410,
    n1192,
    n1200
  );


  nor
  g1513
  (
    n1587,
    n1168,
    n1372,
    n1300,
    n1315
  );


  and
  g1514
  (
    n1527,
    n1266,
    n1195,
    n1226,
    n1394
  );


  and
  g1515
  (
    n1547,
    n1316,
    n1235,
    n1453,
    n1363
  );


  xor
  g1516
  (
    n1490,
    n1225,
    n1278,
    n1394,
    n1166
  );


  or
  g1517
  (
    n1646,
    n1378,
    n1202,
    n1199,
    n1175
  );


  nand
  g1518
  (
    n1575,
    n1260,
    n1456,
    n1380,
    n1397
  );


  nand
  g1519
  (
    n1551,
    n1167,
    n1438,
    n1359,
    n1371
  );


  or
  g1520
  (
    n1719,
    n1401,
    n1358,
    n1172,
    n1304
  );


  nor
  g1521
  (
    KeyWire_0_3,
    n1443,
    n1439,
    n1391,
    n1278
  );


  or
  g1522
  (
    n1585,
    n1166,
    n1392,
    n1202,
    n1317
  );


  nor
  g1523
  (
    n1491,
    n1462,
    n1375,
    n1460,
    n1185
  );


  nand
  g1524
  (
    n1543,
    n1380,
    n1203,
    n1262,
    n1146
  );


  xnor
  g1525
  (
    n1538,
    n1163,
    n1286,
    n1230,
    n1416
  );


  xnor
  g1526
  (
    n1610,
    n1167,
    n1417,
    n1173,
    n1317
  );


  nand
  g1527
  (
    n1529,
    n1241,
    n1299,
    n1406,
    n1431
  );


  nand
  g1528
  (
    n1714,
    n1207,
    n1393,
    n1385,
    n1154
  );


  or
  g1529
  (
    n1475,
    n1379,
    n1286,
    n1358,
    n1425
  );


  xor
  g1530
  (
    n1629,
    n1283,
    n1439,
    n1399,
    n1226
  );


  and
  g1531
  (
    n1500,
    n1449,
    n1251,
    n1410,
    n1312
  );


  and
  g1532
  (
    n1713,
    n1377,
    n1152,
    n1149,
    n1168
  );


  or
  g1533
  (
    n1636,
    n1423,
    n1393,
    n1263,
    n1228
  );


  xor
  g1534
  (
    n1469,
    n1220,
    n1412,
    n1452,
    n1314
  );


  xnor
  g1535
  (
    n1513,
    n1179,
    n1444,
    n1450,
    n1442
  );


  nand
  g1536
  (
    n1669,
    n1183,
    n1280,
    n1450,
    n1383
  );


  xnor
  g1537
  (
    n1523,
    n1181,
    n1238,
    n1197,
    n1185
  );


  xor
  g1538
  (
    n1517,
    n1441,
    n1272,
    n1402,
    n1400
  );


  or
  g1539
  (
    n1560,
    n1211,
    n1381,
    n1145,
    n1255
  );


  and
  g1540
  (
    n1633,
    n1396,
    n1145,
    n1217,
    n1190
  );


  xnor
  g1541
  (
    n1715,
    n1362,
    n1289,
    n1460,
    n1391
  );


  nand
  g1542
  (
    n1495,
    n1145,
    n1465,
    n1310,
    n1451
  );


  xor
  g1543
  (
    n1520,
    n1191,
    n1238,
    n1425,
    n1362
  );


  nand
  g1544
  (
    KeyWire_0_29,
    n1220,
    n1429,
    n1301,
    n1395
  );


  nand
  g1545
  (
    n1554,
    n1208,
    n1250,
    n1291,
    n1237
  );


  nor
  g1546
  (
    n1744,
    n1307,
    n1397,
    n1291,
    n1172
  );


  or
  g1547
  (
    n1666,
    n1180,
    n1239,
    n1197,
    n1270
  );


  and
  g1548
  (
    n1619,
    n1224,
    n1290,
    n1179,
    n1375
  );


  nand
  g1549
  (
    n1514,
    n1294,
    n1393,
    n1306,
    n1268
  );


  or
  g1550
  (
    KeyWire_0_41,
    n1188,
    n1147,
    n1399,
    n1299
  );


  or
  g1551
  (
    n1535,
    n1275,
    n1454,
    n1395,
    n1459
  );


  xor
  g1552
  (
    n1485,
    n1461,
    n1363,
    n1241,
    n1246
  );


  and
  g1553
  (
    n1528,
    n1204,
    n1411,
    n1233,
    n1433
  );


  nor
  g1554
  (
    n1662,
    n1247,
    n1318,
    n1417,
    n1205
  );


  and
  g1555
  (
    n1625,
    n1411,
    n1392,
    n1435,
    n1319
  );


  and
  g1556
  (
    n1655,
    n1183,
    n1407,
    n1362,
    n1461
  );


  nand
  g1557
  (
    n1637,
    n1434,
    n1433,
    n1363,
    n1240
  );


  and
  g1558
  (
    n1627,
    n1270,
    n1148,
    n1291,
    n1276
  );


  or
  g1559
  (
    n1603,
    n1277,
    n1200,
    n1158,
    n1302
  );


  and
  g1560
  (
    n1532,
    n1193,
    n1366,
    n1416,
    n1251
  );


  nand
  g1561
  (
    KeyWire_0_7,
    n1292,
    n1235,
    n1382,
    n1401
  );


  xor
  g1562
  (
    n1499,
    n1185,
    n1199,
    n1189,
    n1404
  );


  or
  g1563
  (
    n1722,
    n1150,
    n1223,
    n1268,
    n1381
  );


  nor
  g1564
  (
    n1577,
    n1212,
    n1362,
    n1229,
    n1436
  );


  nor
  g1565
  (
    n1586,
    n1147,
    n1415,
    n1458,
    n1150
  );


  nor
  g1566
  (
    n1645,
    n1193,
    n1368,
    n1296,
    n1453
  );


  and
  g1567
  (
    n1700,
    n1271,
    n1289,
    n1308,
    n1247
  );


  nand
  g1568
  (
    n1533,
    n1438,
    n1418,
    n1166,
    n1192
  );


  xnor
  g1569
  (
    n1477,
    n1382,
    n1405,
    n1185,
    n1243
  );


  and
  g1570
  (
    n1467,
    n1363,
    n1459,
    n1453,
    n1426
  );


  nor
  g1571
  (
    n1524,
    n1387,
    n1251,
    n1304,
    n1435
  );


  xor
  g1572
  (
    n1738,
    n1225,
    n1189,
    n1248,
    n1208
  );


  or
  g1573
  (
    n1688,
    n1161,
    n1442,
    n1195,
    n1449
  );


  xnor
  g1574
  (
    n1660,
    n1390,
    n1160,
    n1246
  );


  xnor
  g1575
  (
    n1640,
    n1210,
    n1234,
    n1163,
    n1218
  );


  or
  g1576
  (
    n1614,
    n1256,
    n1424,
    n1316,
    n1373
  );


  or
  g1577
  (
    n1727,
    n1430,
    n1372,
    n1156,
    n1266
  );


  xor
  g1578
  (
    n1683,
    n1424,
    n1444,
    n1448,
    n1370
  );


  and
  g1579
  (
    n1489,
    n1240,
    n1195,
    n1384,
    n1458
  );


  and
  g1580
  (
    n1682,
    n1273,
    n1231,
    n1168,
    n1422
  );


  nand
  g1581
  (
    n1483,
    n1302,
    n1419,
    n1405,
    n1232
  );


  and
  g1582
  (
    n1622,
    n1255,
    n1167,
    n1177,
    n1266
  );


  or
  g1583
  (
    n1544,
    n1394,
    n1413,
    n1187,
    n1290
  );


  xor
  g1584
  (
    n1567,
    n1279,
    n1292,
    n1437,
    n1159
  );


  nor
  g1585
  (
    n1564,
    n1162,
    n1313,
    n1302,
    n1389
  );


  or
  g1586
  (
    n1668,
    n1388,
    n1257,
    n1188,
    n1160
  );


  or
  g1587
  (
    n1540,
    n1271,
    n1431,
    n1154,
    n1442
  );


  nor
  g1588
  (
    n1596,
    n1426,
    n1150,
    n1192,
    n1258
  );


  xnor
  g1589
  (
    n1493,
    n1244,
    n1171,
    n1308,
    n1279
  );


  nor
  g1590
  (
    n1591,
    n1432,
    n1260,
    n1400,
    n1440
  );


  or
  g1591
  (
    n1612,
    n1286,
    n1274,
    n1214,
    n1175
  );


  nand
  g1592
  (
    n1689,
    n1426,
    n1276,
    n1390,
    n1429
  );


  xor
  g1593
  (
    n1630,
    n1275,
    n1409,
    n1364,
    n1457
  );


  xnor
  g1594
  (
    n1740,
    n1155,
    n1190,
    n1255,
    n1176
  );


  or
  g1595
  (
    n1703,
    n1418,
    n1446,
    n1187,
    n1184
  );


  xnor
  g1596
  (
    n1608,
    n1437,
    n1182,
    n1242,
    n1287
  );


  xor
  g1597
  (
    n1702,
    n1233,
    n1198,
    n1216,
    n1153
  );


  nand
  g1598
  (
    n1601,
    n1205,
    n1250,
    n1156,
    n1192
  );


  or
  g1599
  (
    n1748,
    n1183,
    n1319,
    n1279,
    n1164
  );


  or
  g1600
  (
    n1611,
    n1264,
    n1296,
    n1297,
    n1253
  );


  nor
  g1601
  (
    n1518,
    n1224,
    n1437,
    n1266,
    n1455
  );


  nand
  g1602
  (
    n1634,
    n1167,
    n1202,
    n1248,
    n1317
  );


  and
  g1603
  (
    n1670,
    n1247,
    n1209,
    n1381,
    n1454
  );


  or
  g1604
  (
    n1720,
    n1219,
    n1464,
    n1291,
    n1290
  );


  nand
  g1605
  (
    n1672,
    n1281,
    n1440,
    n1409,
    n1145
  );


  and
  g1606
  (
    n1472,
    n1258,
    n1397,
    n1383,
    n1272
  );


  nor
  g1607
  (
    n1494,
    n1216,
    n1243,
    n1394,
    n1224
  );


  or
  g1608
  (
    n1698,
    n1274,
    n1271,
    n1401,
    n1186
  );


  xor
  g1609
  (
    n1716,
    n1404,
    n1455,
    n1231,
    n1170
  );


  nor
  g1610
  (
    n1496,
    n1439,
    n1278,
    n1406,
    n1188
  );


  nand
  g1611
  (
    n1600,
    n1236,
    n1240,
    n1268,
    n1257
  );


  nor
  g1612
  (
    n1473,
    n1359,
    n1381,
    n1421,
    n1413
  );


  xor
  g1613
  (
    n1507,
    n1440,
    n1248,
    n1308,
    n1360
  );


  xor
  g1614
  (
    KeyWire_0_49,
    n1231,
    n1427,
    n1376,
    n1177
  );


  xnor
  g1615
  (
    n1552,
    n1298,
    n1273,
    n1208,
    n1417
  );


  xnor
  g1616
  (
    n1638,
    n1236,
    n1240,
    n1403,
    n1272
  );


  nor
  g1617
  (
    n1701,
    n1441,
    n1283,
    n1373,
    n1179
  );


  or
  g1618
  (
    n1534,
    n1182,
    n1284,
    n1181,
    n1299
  );


  nand
  g1619
  (
    n1561,
    n1382,
    n1220,
    n1446,
    n1261
  );


  and
  g1620
  (
    n1620,
    n1170,
    n1268,
    n1287,
    n1239
  );


  or
  g1621
  (
    n1632,
    n1420,
    n1427,
    n1270,
    n1277
  );


  nand
  g1622
  (
    n1692,
    n1305,
    n1404,
    n1253,
    n1460
  );


  xnor
  g1623
  (
    n1724,
    n1147,
    n1441,
    n1252,
    n1203
  );


  xor
  g1624
  (
    n1557,
    n1147,
    n1230,
    n1430,
    n1207
  );


  or
  g1625
  (
    n1588,
    n1262,
    n1180,
    n1319,
    n1249
  );


  xor
  g1626
  (
    n1735,
    n1458,
    n1419,
    n1174,
    n1200
  );


  nor
  g1627
  (
    n1747,
    n1386,
    n1184,
    n1424,
    n1374
  );


  nand
  g1628
  (
    n1508,
    n1407,
    n1379,
    n1260,
    n1403
  );


  and
  g1629
  (
    n1665,
    n1237,
    n1242,
    n1369,
    n1250
  );


  and
  g1630
  (
    n1556,
    n1280,
    n1216,
    n1298,
    n1281
  );


  xor
  g1631
  (
    n1504,
    n1199,
    n1397,
    n1296,
    n1309
  );


  xnor
  g1632
  (
    n1623,
    n1289,
    n1449,
    n1261,
    n1400
  );


  nor
  g1633
  (
    n1699,
    n1447,
    n1310,
    n1174,
    n1201
  );


  and
  g1634
  (
    n1677,
    n1420,
    n1257,
    n1388,
    n1265
  );


  and
  g1635
  (
    n1730,
    n1423,
    n1165,
    n1148,
    n1404
  );


  xnor
  g1636
  (
    KeyWire_0_46,
    n1439,
    n1300,
    n1406,
    n1432
  );


  xor
  g1637
  (
    n1736,
    n1399,
    n1189,
    n1366,
    n1414
  );


  or
  g1638
  (
    n1746,
    n1313,
    n1378,
    n1399,
    n1315
  );


  or
  g1639
  (
    n1686,
    n1386,
    n1402,
    n1395,
    n1370
  );


  and
  g1640
  (
    n1559,
    n1214,
    n1408,
    n1428,
    n1303
  );


  nor
  g1641
  (
    n1742,
    n1358,
    n1391,
    n1154,
    n1152
  );


  and
  g1642
  (
    n1516,
    n1267,
    n1297,
    n1197,
    n1238
  );


  nor
  g1643
  (
    n1479,
    n1398,
    n1200,
    n1376,
    n1303
  );


  or
  g1644
  (
    n1717,
    n1153,
    n1164,
    n1246,
    n1178
  );


  xnor
  g1645
  (
    n1687,
    n1264,
    n1218,
    n1293,
    n1265
  );


  xnor
  g1646
  (
    n1652,
    n1165,
    n1235,
    n1156,
    n1420
  );


  xnor
  g1647
  (
    n1618,
    n1301,
    n1228,
    n1281,
    n1380
  );


  and
  g1648
  (
    n1574,
    n1163,
    n1172,
    n1149,
    n1212
  );


  nand
  g1649
  (
    n1471,
    n1407,
    n1430,
    n1176,
    n1368
  );


  nor
  g1650
  (
    n1555,
    n1456,
    n1417,
    n1441,
    n1392
  );


  xnor
  g1651
  (
    n1578,
    n1358,
    n1451,
    n1272,
    n1197
  );


  xor
  g1652
  (
    n1726,
    n1289,
    n1384,
    n1186,
    n1293
  );


  xnor
  g1653
  (
    n1549,
    n1194,
    n1222,
    n1190,
    n1360
  );


  xnor
  g1654
  (
    n1734,
    n1462,
    n1306,
    n1259,
    n1196
  );


  xnor
  g1655
  (
    n1572,
    n1285,
    n1201,
    n1431,
    n1153
  );


  nand
  g1656
  (
    n1705,
    n1433,
    n1293,
    n1445,
    n1316
  );


  xor
  g1657
  (
    KeyWire_0_42,
    n1244,
    n1454,
    n1151,
    n1210
  );


  and
  g1658
  (
    n1678,
    n1315,
    n1361,
    n1369,
    n1379
  );


  xnor
  g1659
  (
    n1589,
    n1252,
    n1366,
    n1307,
    n1427
  );


  or
  g1660
  (
    n1743,
    n1155,
    n1459,
    n1252,
    n1359
  );


  or
  g1661
  (
    n1536,
    n1202,
    n1174,
    n1436,
    n1257
  );


  nor
  g1662
  (
    n1550,
    n1378,
    n1310,
    n1241,
    n1157
  );


  xnor
  g1663
  (
    n1697,
    n1311,
    n1450,
    n1443,
    n1440
  );


  xnor
  g1664
  (
    n1482,
    n1389,
    n1203,
    n1424,
    n1409
  );


  nor
  g1665
  (
    n1615,
    n1178,
    n1303,
    n1198,
    n1180
  );


  and
  g1666
  (
    n1576,
    n1249,
    n1258,
    n1430,
    n1462
  );


  nor
  g1667
  (
    n1706,
    n1311,
    n1452,
    n1447,
    n1151
  );


  xnor
  g1668
  (
    n1590,
    n1245,
    n1211,
    n1244,
    n1228
  );


  and
  g1669
  (
    n1546,
    n1312,
    n1298,
    n1253,
    n1249
  );


  nand
  g1670
  (
    n1675,
    n1375,
    n1301,
    n1236,
    n1463
  );


  xnor
  g1671
  (
    n1571,
    n1148,
    n1181,
    n1421,
    n1256
  );


  or
  g1672
  (
    n1481,
    n1146,
    n1416,
    n1311,
    n1276
  );


  xor
  g1673
  (
    n1690,
    n1285,
    n1182,
    n1374,
    n1415
  );


  or
  g1674
  (
    n1723,
    n1201,
    n1209,
    n1212,
    n1465
  );


  or
  g1675
  (
    n1667,
    n1171,
    n1294,
    n1158,
    n1445
  );


  xnor
  g1676
  (
    KeyWire_0_61,
    n1386,
    n1242,
    n1312,
    n1220
  );


  nand
  g1677
  (
    n1583,
    n1384,
    n1157,
    n1173,
    n1297
  );


  xor
  g1678
  (
    n1521,
    n1376,
    n1457,
    n1216
  );


  xnor
  g1679
  (
    n1593,
    n1199,
    n1245,
    n1438,
    n1387
  );


  or
  g1680
  (
    n1659,
    n1413,
    n1181,
    n1320,
    n1375
  );


  nand
  g1681
  (
    n1468,
    n1380,
    n1436,
    n1263,
    n1222
  );


  xor
  g1682
  (
    n1656,
    n1413,
    n1227,
    n1428,
    n1446
  );


  xor
  g1683
  (
    n1542,
    n1231,
    n1384,
    n1162,
    n1218
  );


  nor
  g1684
  (
    n1624,
    n1244,
    n1422,
    n1283,
    n1215
  );


  nor
  g1685
  (
    n1545,
    n1169,
    n1373,
    n1175,
    n1415
  );


  xor
  g1686
  (
    n1749,
    n1162,
    n1187,
    n1169,
    n1296
  );


  xnor
  g1687
  (
    n1691,
    n1367,
    n1398,
    n1374,
    n1186
  );


  or
  g1688
  (
    n1647,
    n1155,
    n1383,
    n1452,
    n1373
  );


  xnor
  g1689
  (
    n1592,
    n1301,
    n1444,
    n1314,
    n1206
  );


  or
  g1690
  (
    n1737,
    n1320,
    n1447,
    n1239,
    n1398
  );


  xnor
  g1691
  (
    n1739,
    n1465,
    n1204,
    n1211,
    n1182
  );


  xnor
  g1692
  (
    n1478,
    n1402,
    n1390,
    n1360,
    n1288
  );


  xnor
  g1693
  (
    n1684,
    n1217,
    n1157,
    n1221,
    n1150
  );


  and
  g1694
  (
    n1541,
    n1320,
    n1318,
    n1372,
    n1254
  );


  and
  g1695
  (
    n1548,
    n1206,
    n1297,
    n1234,
    n1414
  );


  xnor
  g1696
  (
    n1470,
    n1447,
    n1431,
    n1187,
    n1245
  );


  nor
  g1697
  (
    n1511,
    n1461,
    n1204,
    n1232,
    n1437
  );


  xnor
  g1698
  (
    n1581,
    n1217,
    n1211,
    n1453,
    n1161
  );


  or
  g1699
  (
    n1661,
    n1282,
    n1361,
    n1400,
    n1295
  );


  xnor
  g1700
  (
    n1594,
    n1454,
    n1205,
    n1425,
    n1376
  );


  xor
  g1701
  (
    n1519,
    n1288,
    n1434,
    n1419,
    n1262
  );


  or
  g1702
  (
    n1681,
    n1282,
    n1229,
    n1148,
    n1281
  );


  and
  g1703
  (
    n1558,
    n1253,
    n1385,
    n1455,
    n1277
  );


  or
  g1704
  (
    n1671,
    n1252,
    n1312,
    n1226,
    n1401
  );


  nand
  g1705
  (
    KeyWire_0_16,
    n1250,
    n1209,
    n1241,
    n1369
  );


  nor
  g1706
  (
    n1505,
    n1300,
    n1429,
    n1422,
    n1388
  );


  and
  g1707
  (
    n1641,
    n1195,
    n1201,
    n1153,
    n1146
  );


  xor
  g1708
  (
    n1599,
    n1428,
    n1273,
    n1213,
    n1464
  );


  xnor
  g1709
  (
    n1651,
    n1314,
    n1168,
    n1212,
    n1304
  );


  and
  g1710
  (
    n1515,
    n1365,
    n1429,
    n1377,
    n1426
  );


  xor
  g1711
  (
    n1710,
    n1451,
    n1227,
    n1248,
    n1361
  );


  nand
  g1712
  (
    n1497,
    n1246,
    n1161,
    n1377,
    n1407
  );


  or
  g1713
  (
    n1639,
    n1170,
    n1149,
    n1368,
    n1293
  );


  nand
  g1714
  (
    n1745,
    n1198,
    n1318,
    n1445,
    n1227
  );


  nand
  g1715
  (
    n1531,
    n1309,
    n1276,
    n1464,
    n1295
  );


  nor
  g1716
  (
    n1512,
    n1304,
    n1360,
    n1194,
    n1292
  );


  or
  g1717
  (
    n1799,
    n1566,
    n1476,
    n1721,
    n1473
  );


  or
  g1718
  (
    n1808,
    n1620,
    n1697,
    n1691,
    n1669
  );


  nor
  g1719
  (
    n1791,
    n1714,
    n1734,
    n1600,
    n1526
  );


  or
  g1720
  (
    n1832,
    n1674,
    n1653,
    n1722,
    n1727
  );


  nand
  g1721
  (
    n1756,
    n1675,
    n1712,
    n1497,
    n1717
  );


  nand
  g1722
  (
    n1817,
    n1468,
    n1606,
    n1702,
    n1715
  );


  or
  g1723
  (
    n1779,
    n1518,
    n1745,
    n1719,
    n1747
  );


  nor
  g1724
  (
    n1780,
    n1555,
    n1642,
    n1582,
    n1718
  );


  and
  g1725
  (
    n1837,
    n1517,
    n1571,
    n1646,
    n1688
  );


  xor
  g1726
  (
    n1859,
    n1654,
    n1535,
    n1677,
    n1632
  );


  xor
  g1727
  (
    n1842,
    n1564,
    n1704,
    n1622,
    n1602
  );


  nor
  g1728
  (
    n1850,
    n1730,
    n1586,
    n1736,
    n1737
  );


  nor
  g1729
  (
    n1852,
    n1724,
    n1696,
    n1698,
    n1482
  );


  xnor
  g1730
  (
    n1750,
    n1702,
    n1742,
    n1713,
    n1480
  );


  xnor
  g1731
  (
    n1769,
    n1672,
    n1494,
    n1710,
    n1590
  );


  nor
  g1732
  (
    n1797,
    n1638,
    n1617,
    n1619,
    n1682
  );


  and
  g1733
  (
    n1845,
    n1495,
    n1711,
    n1596,
    n1651
  );


  xor
  g1734
  (
    n1854,
    n1696,
    n1498,
    n1679,
    n1705
  );


  xnor
  g1735
  (
    n1861,
    n1492,
    n1707,
    n1516,
    n1722
  );


  nor
  g1736
  (
    n1829,
    n1677,
    n1692,
    n1686,
    n1631
  );


  xnor
  g1737
  (
    n1803,
    n1501,
    n1739,
    n1489,
    n1668
  );


  nand
  g1738
  (
    n1762,
    n1676,
    n1717,
    n1486,
    n1682
  );


  and
  g1739
  (
    n1789,
    n1592,
    n1715,
    n1519,
    n1745
  );


  xnor
  g1740
  (
    n1805,
    n1578,
    n1543,
    n1681,
    n1591
  );


  xnor
  g1741
  (
    n1800,
    n1747,
    n1569,
    n1595,
    n1528
  );


  xnor
  g1742
  (
    n1770,
    n1727,
    n1467,
    n1562,
    n1540
  );


  xor
  g1743
  (
    n1766,
    n1706,
    n1699,
    n1558,
    n1694
  );


  or
  g1744
  (
    n1807,
    n1510,
    n1479,
    n1683,
    n1522
  );


  or
  g1745
  (
    n1768,
    n1670,
    n1694,
    n1698,
    n1671
  );


  or
  g1746
  (
    n1821,
    n1554,
    n1704,
    n1659,
    n1703
  );


  xnor
  g1747
  (
    n1757,
    n1471,
    n1712,
    n1743,
    n1594
  );


  nand
  g1748
  (
    n1815,
    n1675,
    n1699,
    n1731,
    n1469
  );


  or
  g1749
  (
    n1796,
    n1530,
    n1673,
    n1639,
    n1747
  );


  and
  g1750
  (
    n1806,
    n1615,
    n1705,
    n1725,
    n1688
  );


  or
  g1751
  (
    n1822,
    n1722,
    n1741,
    n1664,
    n1710
  );


  nand
  g1752
  (
    n1860,
    n1478,
    n1727,
    n1618,
    n1736
  );


  xnor
  g1753
  (
    n1840,
    n1740,
    n1684,
    n1739,
    n1695
  );


  nand
  g1754
  (
    n1813,
    n1711,
    n1514,
    n1700
  );


  xnor
  g1755
  (
    n1763,
    n1521,
    n1680,
    n1504,
    n1674
  );


  nand
  g1756
  (
    n1753,
    n1539,
    n1561,
    n1601,
    n1644
  );


  nor
  g1757
  (
    n1774,
    n1732,
    n1506,
    n1742,
    n1678
  );


  or
  g1758
  (
    n1776,
    n1723,
    n1714,
    n1730,
    n1529
  );


  and
  g1759
  (
    n1783,
    n1679,
    n1705,
    n1691,
    n1474
  );


  and
  g1760
  (
    n1834,
    n1724,
    n1707,
    n1725,
    n1546
  );


  xor
  g1761
  (
    n1855,
    n1685,
    n1610,
    n1741,
    n1713
  );


  nand
  g1762
  (
    n1825,
    n1534,
    n1708,
    n1729,
    n1556
  );


  and
  g1763
  (
    n1771,
    n1598,
    n1718,
    n1726,
    n1701
  );


  xor
  g1764
  (
    n1765,
    n1719,
    n1708,
    n1728,
    n1608
  );


  xnor
  g1765
  (
    n1828,
    n1697,
    n1484,
    n1648,
    n1509
  );


  nor
  g1766
  (
    n1848,
    n1493,
    n1667,
    n1674,
    n1672
  );


  xor
  g1767
  (
    n1773,
    n1656,
    n1605,
    n1533,
    n1570
  );


  xor
  g1768
  (
    n1790,
    n1589,
    n1676,
    n1490,
    n1581
  );


  or
  g1769
  (
    n1841,
    n1637,
    n1574,
    n1748,
    n1704
  );


  xor
  g1770
  (
    n1856,
    n1669,
    n1613,
    n1732,
    n1665
  );


  xor
  g1771
  (
    n1759,
    n1548,
    n1593,
    n1496,
    n1731
  );


  or
  g1772
  (
    n1764,
    n1697,
    n1502,
    n1716,
    n1745
  );


  nand
  g1773
  (
    n1838,
    n1567,
    n1715,
    n1725,
    n1576
  );


  nand
  g1774
  (
    n1818,
    n1623,
    n1597,
    n1672,
    n1542
  );


  or
  g1775
  (
    n1760,
    n1655,
    n1692,
    n1621,
    n1527
  );


  nand
  g1776
  (
    n1802,
    n1573,
    n1604,
    n1662,
    n1660
  );


  or
  g1777
  (
    n1793,
    n1723,
    n1511,
    n1738,
    n1726
  );


  xnor
  g1778
  (
    KeyWire_0_57,
    n1579,
    n1658,
    n1627,
    n1686
  );


  xor
  g1779
  (
    n1835,
    n1736,
    n1729,
    n1701,
    n1741
  );


  or
  g1780
  (
    KeyWire_0_43,
    n1684,
    n1577,
    n1500,
    n1737
  );


  nand
  g1781
  (
    n1857,
    n1690,
    n1711,
    n1575,
    n1696
  );


  xor
  g1782
  (
    n1826,
    n1675,
    n1544,
    n1746,
    n1691
  );


  and
  g1783
  (
    n1827,
    n1536,
    n1738,
    n1483,
    n1634
  );


  nor
  g1784
  (
    n1781,
    n1609,
    n1666,
    n1702,
    n1680
  );


  and
  g1785
  (
    n1794,
    n1718,
    n1724,
    n1669,
    n1694
  );


  xor
  g1786
  (
    n1849,
    n1678,
    n1491,
    n1565,
    n1508
  );


  and
  g1787
  (
    n1839,
    n1701,
    n1481,
    n1532,
    n1710
  );


  and
  g1788
  (
    n1798,
    n1686,
    n1538,
    n1698,
    n1743
  );


  xnor
  g1789
  (
    n1814,
    n1475,
    n1734,
    n1488,
    n1641
  );


  or
  g1790
  (
    n1811,
    n1735,
    n1733,
    n1706,
    n1734
  );


  nor
  g1791
  (
    n1801,
    n1524,
    n1583,
    n1551,
    n1633
  );


  xor
  g1792
  (
    n1788,
    n1740,
    n1466,
    n1742,
    n1611
  );


  xor
  g1793
  (
    n1843,
    n1748,
    n1746,
    n1505,
    n1685
  );


  nor
  g1794
  (
    n1833,
    n1721,
    n1673,
    n1507,
    n1726
  );


  nor
  g1795
  (
    KeyWire_0_63,
    n1682,
    n1537,
    n1703,
    n1749
  );


  nand
  g1796
  (
    n1831,
    n1679,
    n1681,
    n1730,
    n1547
  );


  xnor
  g1797
  (
    n1836,
    n1728,
    n1477,
    n1689,
    n1643
  );


  nor
  g1798
  (
    n1804,
    n1748,
    n1716,
    n1735,
    n1720
  );


  and
  g1799
  (
    n1816,
    n1684,
    n1515,
    n1588,
    n1541
  );


  nand
  g1800
  (
    n1820,
    n1640,
    n1607,
    n1630,
    n1676
  );


  or
  g1801
  (
    n1824,
    n1650,
    n1709,
    n1563,
    n1513
  );


  and
  g1802
  (
    n1819,
    n1693,
    n1560,
    n1706,
    n1709
  );


  or
  g1803
  (
    n1786,
    n1731,
    n1557,
    n1744,
    n1720
  );


  nand
  g1804
  (
    n1830,
    n1717,
    n1728,
    n1714,
    n1628
  );


  xor
  g1805
  (
    n1851,
    n1668,
    n1689,
    n1692,
    n1733
  );


  and
  g1806
  (
    n1767,
    n1624,
    n1487,
    n1614,
    n1661
  );


  or
  g1807
  (
    n1761,
    n1470,
    n1712,
    n1683,
    n1599
  );


  xor
  g1808
  (
    n1792,
    n1647,
    n1616,
    n1743,
    n1700
  );


  nand
  g1809
  (
    n1858,
    n1740,
    n1549,
    n1670,
    n1550
  );


  nand
  g1810
  (
    n1853,
    n1531,
    n1523,
    n1503,
    n1645
  );


  xnor
  g1811
  (
    KeyWire_0_23,
    n1699,
    n1690,
    n1744,
    n1687
  );


  nor
  g1812
  (
    n1810,
    n1678,
    n1652,
    n1708,
    n1737
  );


  xnor
  g1813
  (
    n1785,
    n1707,
    n1720,
    n1729,
    n1749
  );


  or
  g1814
  (
    n1787,
    n1668,
    n1525,
    n1685,
    n1568
  );


  xor
  g1815
  (
    n1752,
    n1580,
    n1559,
    n1693,
    n1485
  );


  and
  g1816
  (
    n1784,
    n1545,
    n1687,
    n1512,
    n1635
  );


  nand
  g1817
  (
    n1772,
    n1649,
    n1690,
    n1657,
    n1738
  );


  and
  g1818
  (
    n1782,
    n1746,
    n1584,
    n1683,
    n1499
  );


  xor
  g1819
  (
    n1754,
    n1612,
    n1472,
    n1629,
    n1744
  );


  and
  g1820
  (
    n1844,
    n1626,
    n1689,
    n1681,
    n1695
  );


  xnor
  g1821
  (
    n1751,
    n1553,
    n1572,
    n1688,
    n1749
  );


  and
  g1822
  (
    n1755,
    n1695,
    n1687,
    n1680,
    n1732
  );


  xor
  g1823
  (
    n1812,
    n1733,
    n1663,
    n1739,
    n1703
  );


  xnor
  g1824
  (
    n1847,
    n1625,
    n1671,
    n1677,
    n1719
  );


  or
  g1825
  (
    n1758,
    n1673,
    n1693,
    n1716,
    n1713
  );


  and
  g1826
  (
    n1846,
    n1552,
    n1671,
    n1709,
    n1735
  );


  nand
  g1827
  (
    n1778,
    n1587,
    n1603,
    n1520,
    n1585
  );


  xnor
  g1828
  (
    n1777,
    n1670,
    n1723,
    n1721,
    n1636
  );


  not
  g1829
  (
    n1874,
    n1770
  );


  buf
  g1830
  (
    n1887,
    n1757
  );


  not
  g1831
  (
    KeyWire_0_14,
    n1780
  );


  buf
  g1832
  (
    n1870,
    n1776
  );


  xor
  g1833
  (
    n1886,
    n1773,
    n1750,
    n1775,
    n1751
  );


  xor
  g1834
  (
    n1888,
    n1754,
    n1763,
    n1762,
    n1759
  );


  or
  g1835
  (
    n1890,
    n1763,
    n1761,
    n1762,
    n1758
  );


  and
  g1836
  (
    n1863,
    n1755,
    n1768,
    n1769,
    n1758
  );


  and
  g1837
  (
    n1877,
    n1750,
    n1766,
    n1765,
    n1761
  );


  xor
  g1838
  (
    n1869,
    n1766,
    n1756,
    n1751,
    n1782
  );


  and
  g1839
  (
    n1867,
    n1779,
    n1758,
    n1757,
    n1753
  );


  nand
  g1840
  (
    n1871,
    n1770,
    n1777,
    n1760
  );


  nand
  g1841
  (
    n1882,
    n1773,
    n1767,
    n1750,
    n1764
  );


  nand
  g1842
  (
    n1896,
    n1751,
    n1763,
    n1758,
    n1760
  );


  xnor
  g1843
  (
    n1872,
    n1778,
    n1779,
    n1765,
    n1769
  );


  xnor
  g1844
  (
    n1865,
    n1753,
    n1776,
    n1764,
    n1771
  );


  xor
  g1845
  (
    n1881,
    n1767,
    n1771,
    n1780,
    n1752
  );


  and
  g1846
  (
    n1885,
    n1769,
    n1755,
    n1761,
    n1764
  );


  nand
  g1847
  (
    n1866,
    n1768,
    n1773,
    n1761,
    n1767
  );


  or
  g1848
  (
    n1893,
    n1768,
    n1772,
    n1755,
    n1770
  );


  or
  g1849
  (
    n1868,
    n1756,
    n1782,
    n1778,
    n1753
  );


  nor
  g1850
  (
    n1897,
    n1769,
    n1782,
    n1764,
    n1772
  );


  or
  g1851
  (
    n1880,
    n1759,
    n1766,
    n1750,
    n1775
  );


  xor
  g1852
  (
    n1891,
    n1775,
    n1779,
    n1781
  );


  and
  g1853
  (
    n1875,
    n1765,
    n1753,
    n1763,
    n1768
  );


  xor
  g1854
  (
    n1864,
    n1770,
    n1754,
    n1775,
    n1781
  );


  or
  g1855
  (
    n1883,
    n1754,
    n1759,
    n1781,
    n1771
  );


  and
  g1856
  (
    n1876,
    n1776,
    n1774,
    n1771,
    n1778
  );


  or
  g1857
  (
    n1879,
    n1774,
    n1757,
    n1762
  );


  nor
  g1858
  (
    n1862,
    n1752,
    n1773,
    n1760,
    n1751
  );


  xor
  g1859
  (
    n1873,
    n1759,
    n1754,
    n1756,
    n1780
  );


  nor
  g1860
  (
    n1889,
    n1752,
    n1772,
    n1774
  );


  and
  g1861
  (
    n1878,
    n1760,
    n1778,
    n1757,
    n1782
  );


  nor
  g1862
  (
    n1892,
    n1752,
    n1781,
    n1756,
    n1766
  );


  nand
  g1863
  (
    n1884,
    n1776,
    n1767,
    n1780,
    n1765
  );


  xor
  g1864
  (
    n1894,
    n1772,
    n1755,
    n1777
  );


  nor
  g1865
  (
    n1978,
    n1808,
    n1805,
    n1842,
    n1815
  );


  nor
  g1866
  (
    n1976,
    n1804,
    n1812,
    n1840,
    n1875
  );


  or
  g1867
  (
    n1931,
    n1831,
    n1882,
    n1797,
    n1809
  );


  and
  g1868
  (
    n1966,
    n1793,
    n1783,
    n1895,
    n1843
  );


  nor
  g1869
  (
    n1983,
    n1828,
    n1792,
    n1866,
    n1881
  );


  nor
  g1870
  (
    n1970,
    n1825,
    n1884,
    n1800,
    n1818
  );


  nand
  g1871
  (
    n1922,
    n1871,
    n1892,
    n1807,
    n1828
  );


  or
  g1872
  (
    n1942,
    n1870,
    n1792,
    n1820,
    n1831
  );


  or
  g1873
  (
    n1925,
    n1879,
    n1837,
    n1864,
    n1888
  );


  or
  g1874
  (
    n1973,
    n1829,
    n1883,
    n1819,
    n1890
  );


  xor
  g1875
  (
    n1926,
    n1841,
    n1893,
    n1838,
    n1882
  );


  nand
  g1876
  (
    n1940,
    n1800,
    n1892,
    n1807,
    n1795
  );


  nor
  g1877
  (
    n1957,
    n1815,
    n1830,
    n1825,
    n1834
  );


  xor
  g1878
  (
    n1971,
    n1802,
    n1883,
    n1889,
    n1831
  );


  nor
  g1879
  (
    n1924,
    n1830,
    n1785,
    n1827,
    n1882
  );


  or
  g1880
  (
    n1972,
    n1826,
    n1817,
    n1821,
    n1841
  );


  or
  g1881
  (
    n1963,
    n1795,
    n1873,
    n1874,
    n1894
  );


  nor
  g1882
  (
    n1949,
    n1789,
    n1822,
    n1895,
    n1814
  );


  xnor
  g1883
  (
    n1916,
    n1786,
    n1789,
    n1888,
    n1807
  );


  and
  g1884
  (
    n1907,
    n1883,
    n1821,
    n1872,
    n1811
  );


  and
  g1885
  (
    n1932,
    n1897,
    n1836,
    n1789,
    n1792
  );


  xnor
  g1886
  (
    n1953,
    n1808,
    n1791,
    n1837,
    n1790
  );


  and
  g1887
  (
    n1903,
    n1827,
    n1896,
    n1784,
    n1865
  );


  xor
  g1888
  (
    n1964,
    n1881,
    n1783,
    n1810,
    n1893
  );


  nor
  g1889
  (
    n1969,
    n1840,
    n1835,
    n1821,
    n1801
  );


  and
  g1890
  (
    n1950,
    n1793,
    n1822,
    n1840,
    n1832
  );


  xnor
  g1891
  (
    n1979,
    n1794,
    n1806,
    n1834,
    n1835
  );


  xor
  g1892
  (
    n1914,
    n1870,
    n1795,
    n1790,
    n1828
  );


  nand
  g1893
  (
    n1912,
    n1839,
    n1887,
    n1874,
    n1869
  );


  and
  g1894
  (
    n1902,
    n1875,
    n1871,
    n1888,
    n1868
  );


  nor
  g1895
  (
    n1959,
    n1806,
    n1799,
    n1830,
    n1807
  );


  and
  g1896
  (
    n1958,
    n1799,
    n1813,
    n1802,
    n1812
  );


  and
  g1897
  (
    n1917,
    n1878,
    n1843,
    n1795,
    n1891
  );


  nor
  g1898
  (
    n1900,
    n1834,
    n1880,
    n1786,
    n1785
  );


  xnor
  g1899
  (
    n1923,
    n1783,
    n1832,
    n1867,
    n1785
  );


  nand
  g1900
  (
    n1938,
    n1897,
    n1818,
    n1829,
    n1804
  );


  nor
  g1901
  (
    n1960,
    n1823,
    n1792,
    n1825,
    n1826
  );


  nand
  g1902
  (
    n1968,
    n1887,
    n1878,
    n1833,
    n1786
  );


  and
  g1903
  (
    n1974,
    n1818,
    n1837,
    n1826
  );


  nor
  g1904
  (
    n1919,
    n1832,
    n1824,
    n1805,
    n1823
  );


  and
  g1905
  (
    n1951,
    n1881,
    n1867,
    n1869,
    n1797
  );


  or
  g1906
  (
    n1905,
    n1890,
    n1801,
    n1865,
    n1887
  );


  xor
  g1907
  (
    n1936,
    n1832,
    n1810,
    n1788,
    n1805
  );


  or
  g1908
  (
    n1944,
    n1823,
    n1892,
    n1796,
    n1800
  );


  and
  g1909
  (
    n1915,
    n1868,
    n1876,
    n1798,
    n1817
  );


  and
  g1910
  (
    n1921,
    n1819,
    n1796,
    n1870,
    n1808
  );


  nor
  g1911
  (
    n1920,
    n1824,
    n1891,
    n1894,
    n1789
  );


  or
  g1912
  (
    n1927,
    n1793,
    n1810,
    n1879,
    n1803
  );


  xnor
  g1913
  (
    n1948,
    n1877,
    n1784,
    n1809,
    n1838
  );


  xor
  g1914
  (
    n1908,
    n1839,
    n1819,
    n1838,
    n1814
  );


  nand
  g1915
  (
    n1977,
    n1813,
    n1835,
    n1820,
    n1799
  );


  nand
  g1916
  (
    n1911,
    n1815,
    n1879,
    n1831,
    n1790
  );


  xor
  g1917
  (
    n1975,
    n1897,
    n1895,
    n1836,
    n1822
  );


  nor
  g1918
  (
    n1981,
    n1889,
    n1788,
    n1817,
    n1864
  );


  and
  g1919
  (
    n1955,
    n1784,
    n1825,
    n1787,
    n1873
  );


  and
  g1920
  (
    n1956,
    n1803,
    n1784,
    n1819,
    n1829
  );


  xor
  g1921
  (
    n1980,
    n1864,
    n1797,
    n1842,
    n1791
  );


  xnor
  g1922
  (
    n1929,
    n1868,
    n1874,
    n1841,
    n1798
  );


  xor
  g1923
  (
    n1945,
    n1787,
    n1877,
    n1813,
    n1788
  );


  nor
  g1924
  (
    n1934,
    n1806,
    n1834,
    n1787,
    n1842
  );


  and
  g1925
  (
    n1898,
    n1891,
    n1839,
    n1803,
    n1889
  );


  or
  g1926
  (
    n1939,
    n1829,
    n1830,
    n1804,
    n1833
  );


  nand
  g1927
  (
    KeyWire_0_32,
    n1885,
    n1800,
    n1806,
    n1865
  );


  and
  g1928
  (
    n1918,
    n1824,
    n1873,
    n1878,
    n1884
  );


  or
  g1929
  (
    n1928,
    n1809,
    n1841,
    n1811,
    n1808
  );


  nor
  g1930
  (
    n1967,
    n1822,
    n1812,
    n1875,
    n1788
  );


  xnor
  g1931
  (
    n1910,
    n1816,
    n1876,
    n1838,
    n1877
  );


  and
  g1932
  (
    n1904,
    n1811,
    n1820,
    n1824,
    n1803
  );


  xor
  g1933
  (
    n1943,
    n1818,
    n1804,
    n1793,
    n1826
  );


  and
  g1934
  (
    n1961,
    n1791,
    n1791,
    n1886,
    n1828
  );


  and
  g1935
  (
    n1930,
    n1885,
    n1810,
    n1805,
    n1840
  );


  nor
  g1936
  (
    n1962,
    n1833,
    n1836,
    n1866,
    n1890
  );


  or
  g1937
  (
    n1952,
    n1886,
    n1817,
    n1827,
    n1867
  );


  nor
  g1938
  (
    n1901,
    n1886,
    n1798,
    n1839,
    n1876
  );


  nor
  g1939
  (
    n1899,
    n1799,
    n1896,
    n1814,
    n1809
  );


  nor
  g1940
  (
    n1982,
    n1884,
    n1794,
    n1801
  );


  and
  g1941
  (
    n1909,
    n1796,
    n1880,
    n1794,
    n1816
  );


  xor
  g1942
  (
    n1935,
    n1893,
    n1827,
    n1842,
    n1787
  );


  nand
  g1943
  (
    n1947,
    n1814,
    n1880,
    n1816,
    n1802
  );


  nor
  g1944
  (
    KeyWire_0_20,
    n1801,
    n1786,
    n1835,
    n1815
  );


  nor
  g1945
  (
    n1937,
    n1797,
    n1872,
    n1885,
    n1836
  );


  xnor
  g1946
  (
    n1913,
    n1821,
    n1785,
    n1783,
    n1896
  );


  or
  g1947
  (
    n1906,
    n1833,
    n1866,
    n1869,
    n1798
  );


  xor
  g1948
  (
    n1965,
    n1813,
    n1796,
    n1790,
    n1811
  );


  nand
  g1949
  (
    n1941,
    n1816,
    n1871,
    n1872,
    n1894
  );


  nand
  g1950
  (
    n1954,
    n1802,
    n1820,
    n1812,
    n1823
  );


  xor
  g1951
  (
    n2009,
    n1855,
    n1975,
    n1980,
    n1929
  );


  and
  g1952
  (
    n2012,
    n1910,
    n1899,
    n1906,
    n1974
  );


  or
  g1953
  (
    n2000,
    n1848,
    n1959,
    n1845,
    n1843
  );


  nand
  g1954
  (
    n1997,
    n1907,
    n1855,
    n1845,
    n1909
  );


  xnor
  g1955
  (
    n1986,
    n1914,
    n1956,
    n1931,
    n1852
  );


  and
  g1956
  (
    n1988,
    n1947,
    n1951,
    n1926,
    n1848
  );


  or
  g1957
  (
    n1993,
    n1912,
    n1977,
    n1844,
    n1845
  );


  and
  g1958
  (
    n2016,
    n1928,
    n1983,
    n1854,
    n1976
  );


  or
  g1959
  (
    n2013,
    n1979,
    n1940,
    n1946,
    n1962
  );


  xor
  g1960
  (
    n1985,
    n1904,
    n1972,
    n1856,
    n1849
  );


  or
  g1961
  (
    n1999,
    n1924,
    n1856,
    n1852,
    n1971
  );


  nand
  g1962
  (
    n2010,
    n1844,
    n1943,
    n1941,
    n1965
  );


  nand
  g1963
  (
    n1992,
    n1853,
    n1853,
    n1923,
    n1844
  );


  nand
  g1964
  (
    n1996,
    n1913,
    n1954,
    n1967,
    n1955
  );


  xor
  g1965
  (
    n2014,
    n1966,
    n1905,
    n1953,
    n1957
  );


  nor
  g1966
  (
    n2008,
    n1902,
    n1937,
    n1968,
    n1961
  );


  xor
  g1967
  (
    n1984,
    n1920,
    n1949,
    n1981,
    n1930
  );


  nor
  g1968
  (
    n1994,
    n1845,
    n1936,
    n1848,
    n1973
  );


  xnor
  g1969
  (
    n2015,
    n1846,
    n1852,
    n1850
  );


  nor
  g1970
  (
    n1995,
    n1908,
    n1935,
    n1850,
    n1969
  );


  or
  g1971
  (
    n1991,
    n1958,
    n1942,
    n1944,
    n1849
  );


  and
  g1972
  (
    n2018,
    n1847,
    n1933,
    n1854,
    n1932
  );


  nor
  g1973
  (
    n1987,
    n1851,
    n1900,
    n1848,
    n1854
  );


  and
  g1974
  (
    n1998,
    n1939,
    n1960,
    n1851,
    n1847
  );


  nand
  g1975
  (
    n2011,
    n1855,
    n1844,
    n1950,
    n1854
  );


  xnor
  g1976
  (
    n2004,
    n1847,
    n1927,
    n1970,
    n1901
  );


  xnor
  g1977
  (
    n2003,
    n1853,
    n1843,
    n1852,
    n1851
  );


  xnor
  g1978
  (
    n2005,
    n1855,
    n1934,
    n1963,
    n1851
  );


  and
  g1979
  (
    n1990,
    n1849,
    n1938,
    n1916,
    n1915
  );


  or
  g1980
  (
    n2002,
    n1919,
    n1948,
    n1898,
    n1846
  );


  xor
  g1981
  (
    n2007,
    n1846,
    n1846,
    n1925,
    n1917
  );


  nand
  g1982
  (
    n2017,
    n1921,
    n1850,
    n1978,
    n1964
  );


  xor
  g1983
  (
    n1989,
    n1982,
    n1952,
    n1903,
    n1922
  );


  xor
  g1984
  (
    n2006,
    n1847,
    n1918,
    n1945,
    n1853
  );


  and
  g1985
  (
    n2001,
    n32,
    n1849,
    n1911,
    n1856
  );


  xnor
  g1986
  (
    n2030,
    n1991,
    n1986,
    n2005,
    n2003
  );


  xor
  g1987
  (
    n2028,
    n1995,
    n2010,
    n1859,
    n1984
  );


  xor
  g1988
  (
    n2020,
    n1861,
    n2000,
    n1856,
    n1858
  );


  nand
  g1989
  (
    n2027,
    n1861,
    n1987,
    n2002,
    n1985
  );


  or
  g1990
  (
    n2023,
    n2014,
    n2013,
    n1857,
    n1861
  );


  xor
  g1991
  (
    n2022,
    n2016,
    n2004,
    n1988,
    n2009
  );


  xnor
  g1992
  (
    n2021,
    n1859,
    n1859,
    n1992,
    n1857
  );


  xnor
  g1993
  (
    n2024,
    n1996,
    n1858,
    n1860
  );


  nor
  g1994
  (
    n2029,
    n1858,
    n1860,
    n1994,
    n2015
  );


  and
  g1995
  (
    n2032,
    n1990,
    n2012,
    n2001,
    n2018
  );


  or
  g1996
  (
    n2031,
    n1858,
    n2008,
    n1999,
    n1998
  );


  xor
  g1997
  (
    n2025,
    n1989,
    n1993,
    n2006,
    n1860
  );


  nor
  g1998
  (
    n2019,
    n1859,
    n1997,
    n1861,
    n2011
  );


  xnor
  g1999
  (
    n2026,
    n2007,
    n1857,
    n2017
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1106,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1253,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n424,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1602,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n285,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1275,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1462,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1664,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1609,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1304,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n239,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n91,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n126,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1041,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1895,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n194,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n1539,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n170,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n1033,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n1074,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1933,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n616,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n999,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1809,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n972,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1331,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n491,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1649,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n907,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1621,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n538,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1249,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n1946,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n40,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n1157,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n602,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n1261,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n1137,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n1579,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n1694,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n1298,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n1704,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n1487,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n1775,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n241,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n919,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n1563,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n563,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1440,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n1696,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n697,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n222,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n672,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n1301,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n1464,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n476,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n404,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n1823,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n1416,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n811,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n1118,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n1607,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n315,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n1795,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


