

module Stat_3000_302
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2790,
  n2796,
  n2802,
  n2800,
  n2801,
  n2797,
  n2795,
  n2805,
  n2881,
  n2882,
  n2889,
  n2893,
  n2892,
  n2888,
  n2883,
  n2890,
  n2880,
  n2885,
  n2969,
  n2961,
  n2966,
  n2968,
  n2959,
  n2967,
  n2970,
  n2962,
  n2964,
  n2960,
  n3030,
  n3031,
  n3032,
  n3029,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n2790;
  output n2796;
  output n2802;
  output n2800;
  output n2801;
  output n2797;
  output n2795;
  output n2805;
  output n2881;
  output n2882;
  output n2889;
  output n2893;
  output n2892;
  output n2888;
  output n2883;
  output n2890;
  output n2880;
  output n2885;
  output n2969;
  output n2961;
  output n2966;
  output n2968;
  output n2959;
  output n2967;
  output n2970;
  output n2962;
  output n2964;
  output n2960;
  output n3030;
  output n3031;
  output n3032;
  output n3029;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2798;
  wire n2799;
  wire n2803;
  wire n2804;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2884;
  wire n2886;
  wire n2887;
  wire n2891;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2963;
  wire n2965;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n157,
    n20
  );


  buf
  g1
  (
    n66,
    n9
  );


  buf
  g2
  (
    n62,
    n12
  );


  buf
  g3
  (
    n104,
    n28
  );


  not
  g4
  (
    n94,
    n1
  );


  buf
  g5
  (
    n106,
    n31
  );


  buf
  g6
  (
    n124,
    n8
  );


  buf
  g7
  (
    n117,
    n19
  );


  not
  g8
  (
    KeyWire_0_18,
    n22
  );


  not
  g9
  (
    n129,
    n21
  );


  not
  g10
  (
    n153,
    n11
  );


  buf
  g11
  (
    n155,
    n10
  );


  not
  g12
  (
    n37,
    n11
  );


  buf
  g13
  (
    n47,
    n14
  );


  buf
  g14
  (
    n123,
    n25
  );


  buf
  g15
  (
    n128,
    n23
  );


  not
  g16
  (
    n93,
    n5
  );


  buf
  g17
  (
    n73,
    n6
  );


  not
  g18
  (
    n34,
    n32
  );


  buf
  g19
  (
    n126,
    n22
  );


  not
  g20
  (
    n150,
    n5
  );


  buf
  g21
  (
    n109,
    n8
  );


  buf
  g22
  (
    n36,
    n13
  );


  buf
  g23
  (
    n46,
    n2
  );


  not
  g24
  (
    n127,
    n6
  );


  not
  g25
  (
    n156,
    n24
  );


  not
  g26
  (
    KeyWire_0_42,
    n20
  );


  not
  g27
  (
    n39,
    n13
  );


  buf
  g28
  (
    n121,
    n6
  );


  not
  g29
  (
    n143,
    n2
  );


  not
  g30
  (
    n85,
    n3
  );


  not
  g31
  (
    n101,
    n26
  );


  buf
  g32
  (
    n60,
    n9
  );


  buf
  g33
  (
    n74,
    n21
  );


  not
  g34
  (
    n59,
    n6
  );


  buf
  g35
  (
    n145,
    n25
  );


  buf
  g36
  (
    n45,
    n4
  );


  not
  g37
  (
    n67,
    n23
  );


  not
  g38
  (
    n154,
    n27
  );


  buf
  g39
  (
    n42,
    n3
  );


  buf
  g40
  (
    n54,
    n28
  );


  buf
  g41
  (
    n105,
    n8
  );


  buf
  g42
  (
    n71,
    n14
  );


  not
  g43
  (
    n148,
    n10
  );


  not
  g44
  (
    n115,
    n24
  );


  buf
  g45
  (
    n75,
    n22
  );


  buf
  g46
  (
    n112,
    n22
  );


  buf
  g47
  (
    n140,
    n30
  );


  buf
  g48
  (
    n65,
    n7
  );


  not
  g49
  (
    n111,
    n30
  );


  buf
  g50
  (
    n134,
    n19
  );


  not
  g51
  (
    n103,
    n23
  );


  not
  g52
  (
    n41,
    n24
  );


  not
  g53
  (
    n88,
    n1
  );


  buf
  g54
  (
    n53,
    n4
  );


  buf
  g55
  (
    n159,
    n16
  );


  buf
  g56
  (
    n110,
    n7
  );


  not
  g57
  (
    n97,
    n32
  );


  not
  g58
  (
    n95,
    n21
  );


  buf
  g59
  (
    n113,
    n4
  );


  not
  g60
  (
    n78,
    n26
  );


  buf
  g61
  (
    n70,
    n14
  );


  buf
  g62
  (
    n108,
    n15
  );


  not
  g63
  (
    n56,
    n12
  );


  not
  g64
  (
    n142,
    n10
  );


  not
  g65
  (
    n63,
    n32
  );


  buf
  g66
  (
    n116,
    n29
  );


  buf
  g67
  (
    n141,
    n27
  );


  not
  g68
  (
    n118,
    n31
  );


  buf
  g69
  (
    n61,
    n1
  );


  buf
  g70
  (
    n87,
    n9
  );


  not
  g71
  (
    n83,
    n27
  );


  not
  g72
  (
    n79,
    n18
  );


  not
  g73
  (
    n81,
    n16
  );


  not
  g74
  (
    n135,
    n4
  );


  not
  g75
  (
    n38,
    n21
  );


  not
  g76
  (
    n160,
    n25
  );


  not
  g77
  (
    n114,
    n3
  );


  not
  g78
  (
    n144,
    n14
  );


  buf
  g79
  (
    n90,
    n18
  );


  not
  g80
  (
    n152,
    n12
  );


  not
  g81
  (
    n69,
    n30
  );


  not
  g82
  (
    n80,
    n9
  );


  not
  g83
  (
    n33,
    n23
  );


  buf
  g84
  (
    n48,
    n17
  );


  not
  g85
  (
    n136,
    n1
  );


  not
  g86
  (
    n58,
    n11
  );


  not
  g87
  (
    n131,
    n15
  );


  not
  g88
  (
    n130,
    n29
  );


  not
  g89
  (
    n158,
    n30
  );


  not
  g90
  (
    n44,
    n29
  );


  not
  g91
  (
    n137,
    n28
  );


  not
  g92
  (
    n100,
    n24
  );


  not
  g93
  (
    n50,
    n25
  );


  not
  g94
  (
    n149,
    n13
  );


  not
  g95
  (
    n119,
    n18
  );


  not
  g96
  (
    n133,
    n19
  );


  buf
  g97
  (
    n107,
    n26
  );


  not
  g98
  (
    n138,
    n8
  );


  not
  g99
  (
    n35,
    n11
  );


  not
  g100
  (
    n151,
    n10
  );


  buf
  g101
  (
    n55,
    n13
  );


  buf
  g102
  (
    KeyWire_0_25,
    n29
  );


  not
  g103
  (
    n64,
    n26
  );


  not
  g104
  (
    n86,
    n7
  );


  not
  g105
  (
    n92,
    n16
  );


  buf
  g106
  (
    n139,
    n5
  );


  buf
  g107
  (
    n89,
    n20
  );


  buf
  g108
  (
    n40,
    n19
  );


  buf
  g109
  (
    n77,
    n16
  );


  not
  g110
  (
    n68,
    n28
  );


  not
  g111
  (
    n120,
    n12
  );


  not
  g112
  (
    n57,
    n31
  );


  buf
  g113
  (
    n102,
    n18
  );


  not
  g114
  (
    n84,
    n3
  );


  buf
  g115
  (
    n98,
    n31
  );


  not
  g116
  (
    n91,
    n15
  );


  buf
  g117
  (
    n96,
    n32
  );


  not
  g118
  (
    n125,
    n15
  );


  not
  g119
  (
    n147,
    n2
  );


  not
  g120
  (
    n43,
    n20
  );


  not
  g121
  (
    n99,
    n17
  );


  buf
  g122
  (
    n76,
    n17
  );


  not
  g123
  (
    n52,
    n27
  );


  buf
  g124
  (
    n51,
    n2
  );


  buf
  g125
  (
    n122,
    n17
  );


  buf
  g126
  (
    n146,
    n5
  );


  buf
  g127
  (
    n132,
    n7
  );


  not
  g128
  (
    n475,
    n140
  );


  buf
  g129
  (
    n317,
    n98
  );


  not
  g130
  (
    n326,
    n92
  );


  not
  g131
  (
    n559,
    n47
  );


  buf
  g132
  (
    n602,
    n80
  );


  not
  g133
  (
    n456,
    n86
  );


  buf
  g134
  (
    n356,
    n44
  );


  buf
  g135
  (
    n569,
    n140
  );


  buf
  g136
  (
    n222,
    n150
  );


  not
  g137
  (
    n395,
    n48
  );


  buf
  g138
  (
    n409,
    n117
  );


  not
  g139
  (
    n198,
    n156
  );


  buf
  g140
  (
    n443,
    n82
  );


  not
  g141
  (
    n309,
    n105
  );


  buf
  g142
  (
    n273,
    n136
  );


  not
  g143
  (
    n499,
    n123
  );


  buf
  g144
  (
    n177,
    n157
  );


  buf
  g145
  (
    n289,
    n34
  );


  not
  g146
  (
    n388,
    n35
  );


  buf
  g147
  (
    n663,
    n78
  );


  buf
  g148
  (
    n563,
    n78
  );


  not
  g149
  (
    n374,
    n79
  );


  buf
  g150
  (
    KeyWire_0_37,
    n144
  );


  buf
  g151
  (
    n653,
    n72
  );


  buf
  g152
  (
    n301,
    n142
  );


  not
  g153
  (
    n438,
    n158
  );


  buf
  g154
  (
    n349,
    n63
  );


  not
  g155
  (
    n230,
    n68
  );


  not
  g156
  (
    n300,
    n158
  );


  buf
  g157
  (
    n302,
    n79
  );


  buf
  g158
  (
    n629,
    n157
  );


  not
  g159
  (
    n308,
    n119
  );


  not
  g160
  (
    n515,
    n149
  );


  buf
  g161
  (
    n468,
    n115
  );


  not
  g162
  (
    n633,
    n130
  );


  not
  g163
  (
    n195,
    n55
  );


  not
  g164
  (
    n321,
    n50
  );


  buf
  g165
  (
    n616,
    n107
  );


  not
  g166
  (
    n322,
    n81
  );


  not
  g167
  (
    n422,
    n151
  );


  not
  g168
  (
    n566,
    n159
  );


  not
  g169
  (
    n202,
    n50
  );


  buf
  g170
  (
    n310,
    n77
  );


  not
  g171
  (
    n491,
    n102
  );


  not
  g172
  (
    n223,
    n69
  );


  buf
  g173
  (
    n411,
    n36
  );


  not
  g174
  (
    n334,
    n68
  );


  buf
  g175
  (
    n446,
    n132
  );


  not
  g176
  (
    n557,
    n150
  );


  not
  g177
  (
    n262,
    n90
  );


  buf
  g178
  (
    n614,
    n94
  );


  buf
  g179
  (
    n472,
    n103
  );


  buf
  g180
  (
    n351,
    n87
  );


  buf
  g181
  (
    n283,
    n38
  );


  buf
  g182
  (
    n474,
    n139
  );


  not
  g183
  (
    n543,
    n89
  );


  buf
  g184
  (
    n413,
    n111
  );


  buf
  g185
  (
    n184,
    n36
  );


  buf
  g186
  (
    n550,
    n90
  );


  not
  g187
  (
    n190,
    n88
  );


  buf
  g188
  (
    n266,
    n44
  );


  not
  g189
  (
    n626,
    n63
  );


  buf
  g190
  (
    n303,
    n116
  );


  buf
  g191
  (
    KeyWire_0_19,
    n34
  );


  buf
  g192
  (
    n481,
    n33
  );


  not
  g193
  (
    n344,
    n96
  );


  buf
  g194
  (
    n380,
    n62
  );


  not
  g195
  (
    n384,
    n134
  );


  not
  g196
  (
    n178,
    n91
  );


  not
  g197
  (
    n448,
    n53
  );


  not
  g198
  (
    KeyWire_0_34,
    n49
  );


  not
  g199
  (
    n286,
    n149
  );


  buf
  g200
  (
    n618,
    n97
  );


  buf
  g201
  (
    n207,
    n153
  );


  buf
  g202
  (
    n292,
    n116
  );


  buf
  g203
  (
    n263,
    n117
  );


  buf
  g204
  (
    n587,
    n55
  );


  not
  g205
  (
    n311,
    n38
  );


  not
  g206
  (
    n607,
    n38
  );


  buf
  g207
  (
    n352,
    n119
  );


  buf
  g208
  (
    n161,
    n159
  );


  not
  g209
  (
    n488,
    n60
  );


  buf
  g210
  (
    n608,
    n51
  );


  not
  g211
  (
    n549,
    n73
  );


  buf
  g212
  (
    n221,
    n100
  );


  buf
  g213
  (
    n539,
    n85
  );


  not
  g214
  (
    n217,
    n144
  );


  buf
  g215
  (
    n586,
    n80
  );


  not
  g216
  (
    n165,
    n108
  );


  not
  g217
  (
    n164,
    n146
  );


  buf
  g218
  (
    n526,
    n148
  );


  not
  g219
  (
    n414,
    n56
  );


  buf
  g220
  (
    n167,
    n137
  );


  not
  g221
  (
    n383,
    n125
  );


  not
  g222
  (
    n619,
    n151
  );


  not
  g223
  (
    n427,
    n154
  );


  buf
  g224
  (
    n442,
    n57
  );


  not
  g225
  (
    n335,
    n122
  );


  buf
  g226
  (
    n593,
    n156
  );


  not
  g227
  (
    n632,
    n139
  );


  not
  g228
  (
    n329,
    n146
  );


  not
  g229
  (
    n592,
    n131
  );


  not
  g230
  (
    KeyWire_0_30,
    n128
  );


  buf
  g231
  (
    n243,
    n122
  );


  buf
  g232
  (
    n174,
    n34
  );


  buf
  g233
  (
    n245,
    n104
  );


  not
  g234
  (
    n522,
    n33
  );


  buf
  g235
  (
    n657,
    n117
  );


  not
  g236
  (
    n429,
    n60
  );


  not
  g237
  (
    n229,
    n131
  );


  buf
  g238
  (
    n290,
    n100
  );


  not
  g239
  (
    n623,
    n35
  );


  buf
  g240
  (
    n340,
    n50
  );


  buf
  g241
  (
    n267,
    n69
  );


  buf
  g242
  (
    n664,
    n54
  );


  buf
  g243
  (
    n306,
    n96
  );


  not
  g244
  (
    n354,
    n147
  );


  not
  g245
  (
    n285,
    n139
  );


  not
  g246
  (
    n574,
    n105
  );


  not
  g247
  (
    n502,
    n91
  );


  not
  g248
  (
    n247,
    n47
  );


  buf
  g249
  (
    n180,
    n145
  );


  buf
  g250
  (
    n313,
    n66
  );


  not
  g251
  (
    n257,
    n57
  );


  buf
  g252
  (
    n556,
    n46
  );


  not
  g253
  (
    n209,
    n145
  );


  buf
  g254
  (
    n449,
    n75
  );


  buf
  g255
  (
    n324,
    n99
  );


  buf
  g256
  (
    n318,
    n130
  );


  not
  g257
  (
    n494,
    n51
  );


  buf
  g258
  (
    n523,
    n84
  );


  buf
  g259
  (
    n601,
    n93
  );


  buf
  g260
  (
    n600,
    n126
  );


  buf
  g261
  (
    n583,
    n40
  );


  not
  g262
  (
    n469,
    n61
  );


  not
  g263
  (
    n436,
    n100
  );


  not
  g264
  (
    n297,
    n84
  );


  not
  g265
  (
    n254,
    n77
  );


  not
  g266
  (
    n407,
    n118
  );


  buf
  g267
  (
    n357,
    n103
  );


  buf
  g268
  (
    n342,
    n59
  );


  buf
  g269
  (
    n447,
    n135
  );


  buf
  g270
  (
    n296,
    n127
  );


  not
  g271
  (
    n400,
    n43
  );


  not
  g272
  (
    n611,
    n81
  );


  buf
  g273
  (
    n554,
    n48
  );


  not
  g274
  (
    n460,
    n119
  );


  not
  g275
  (
    n319,
    n37
  );


  buf
  g276
  (
    n578,
    n129
  );


  buf
  g277
  (
    n432,
    n74
  );


  buf
  g278
  (
    n215,
    n52
  );


  buf
  g279
  (
    n276,
    n114
  );


  not
  g280
  (
    n662,
    n37
  );


  buf
  g281
  (
    n227,
    n75
  );


  not
  g282
  (
    n639,
    n121
  );


  buf
  g283
  (
    n337,
    n149
  );


  not
  g284
  (
    n507,
    n80
  );


  not
  g285
  (
    n505,
    n66
  );


  not
  g286
  (
    n168,
    n126
  );


  not
  g287
  (
    n571,
    n74
  );


  buf
  g288
  (
    n471,
    n142
  );


  buf
  g289
  (
    n353,
    n71
  );


  buf
  g290
  (
    n228,
    n45
  );


  not
  g291
  (
    n396,
    n75
  );


  not
  g292
  (
    n572,
    n152
  );


  not
  g293
  (
    n212,
    n86
  );


  buf
  g294
  (
    KeyWire_0_11,
    n104
  );


  not
  g295
  (
    n581,
    n125
  );


  buf
  g296
  (
    n390,
    n63
  );


  not
  g297
  (
    n369,
    n123
  );


  buf
  g298
  (
    n163,
    n124
  );


  not
  g299
  (
    n295,
    n127
  );


  not
  g300
  (
    n504,
    n35
  );


  buf
  g301
  (
    n510,
    n81
  );


  buf
  g302
  (
    n373,
    n43
  );


  not
  g303
  (
    n252,
    n54
  );


  buf
  g304
  (
    KeyWire_0_54,
    n39
  );


  buf
  g305
  (
    n484,
    n107
  );


  buf
  g306
  (
    n642,
    n133
  );


  not
  g307
  (
    n455,
    n149
  );


  buf
  g308
  (
    n540,
    n150
  );


  not
  g309
  (
    n454,
    n66
  );


  not
  g310
  (
    n192,
    n59
  );


  not
  g311
  (
    n331,
    n102
  );


  not
  g312
  (
    n503,
    n156
  );


  buf
  g313
  (
    n500,
    n56
  );


  buf
  g314
  (
    n403,
    n122
  );


  buf
  g315
  (
    n216,
    n113
  );


  not
  g316
  (
    n486,
    n134
  );


  not
  g317
  (
    n193,
    n52
  );


  not
  g318
  (
    n511,
    n62
  );


  buf
  g319
  (
    n242,
    n144
  );


  buf
  g320
  (
    n451,
    n129
  );


  buf
  g321
  (
    n235,
    n155
  );


  buf
  g322
  (
    n624,
    n42
  );


  not
  g323
  (
    n382,
    n55
  );


  not
  g324
  (
    n220,
    n51
  );


  not
  g325
  (
    n535,
    n76
  );


  buf
  g326
  (
    n232,
    n120
  );


  not
  g327
  (
    n564,
    n157
  );


  buf
  g328
  (
    n635,
    n41
  );


  buf
  g329
  (
    n333,
    n39
  );


  not
  g330
  (
    n570,
    n90
  );


  not
  g331
  (
    n197,
    n101
  );


  buf
  g332
  (
    n291,
    n51
  );


  not
  g333
  (
    n599,
    n120
  );


  buf
  g334
  (
    n250,
    n92
  );


  buf
  g335
  (
    n363,
    n60
  );


  not
  g336
  (
    n631,
    n96
  );


  not
  g337
  (
    n325,
    n84
  );


  not
  g338
  (
    n424,
    n70
  );


  not
  g339
  (
    n490,
    n143
  );


  buf
  g340
  (
    n465,
    n76
  );


  buf
  g341
  (
    n253,
    n37
  );


  not
  g342
  (
    n375,
    n140
  );


  not
  g343
  (
    n501,
    n112
  );


  buf
  g344
  (
    n498,
    n141
  );


  buf
  g345
  (
    n181,
    n135
  );


  not
  g346
  (
    n487,
    n129
  );


  buf
  g347
  (
    n204,
    n87
  );


  not
  g348
  (
    n213,
    n56
  );


  not
  g349
  (
    n269,
    n49
  );


  buf
  g350
  (
    n385,
    n61
  );


  buf
  g351
  (
    n647,
    n66
  );


  buf
  g352
  (
    n594,
    n73
  );


  not
  g353
  (
    n561,
    n36
  );


  buf
  g354
  (
    n196,
    n35
  );


  buf
  g355
  (
    n457,
    n125
  );


  not
  g356
  (
    n582,
    n146
  );


  not
  g357
  (
    n421,
    n111
  );


  not
  g358
  (
    n378,
    n81
  );


  buf
  g359
  (
    n450,
    n115
  );


  buf
  g360
  (
    n381,
    n74
  );


  not
  g361
  (
    n398,
    n64
  );


  not
  g362
  (
    n265,
    n151
  );


  buf
  g363
  (
    n558,
    n56
  );


  buf
  g364
  (
    n187,
    n34
  );


  not
  g365
  (
    n555,
    n128
  );


  buf
  g366
  (
    KeyWire_0_4,
    n62
  );


  buf
  g367
  (
    n173,
    n152
  );


  buf
  g368
  (
    n434,
    n83
  );


  not
  g369
  (
    n660,
    n39
  );


  not
  g370
  (
    n650,
    n143
  );


  not
  g371
  (
    KeyWire_0_35,
    n111
  );


  not
  g372
  (
    n237,
    n147
  );


  not
  g373
  (
    n358,
    n63
  );


  buf
  g374
  (
    n408,
    n78
  );


  not
  g375
  (
    n651,
    n158
  );


  buf
  g376
  (
    n590,
    n53
  );


  buf
  g377
  (
    n275,
    n133
  );


  buf
  g378
  (
    n546,
    n153
  );


  buf
  g379
  (
    n169,
    n154
  );


  buf
  g380
  (
    n392,
    n52
  );


  not
  g381
  (
    n645,
    n95
  );


  not
  g382
  (
    n580,
    n77
  );


  buf
  g383
  (
    n444,
    n114
  );


  buf
  g384
  (
    n270,
    n116
  );


  buf
  g385
  (
    KeyWire_0_29,
    n126
  );


  buf
  g386
  (
    n506,
    n126
  );


  buf
  g387
  (
    n667,
    n38
  );


  not
  g388
  (
    n332,
    n95
  );


  not
  g389
  (
    n654,
    n90
  );


  not
  g390
  (
    n406,
    n154
  );


  not
  g391
  (
    n576,
    n148
  );


  buf
  g392
  (
    n347,
    n110
  );


  not
  g393
  (
    n338,
    n62
  );


  not
  g394
  (
    n244,
    n154
  );


  buf
  g395
  (
    n512,
    n106
  );


  not
  g396
  (
    n365,
    n84
  );


  buf
  g397
  (
    n366,
    n65
  );


  not
  g398
  (
    n359,
    n141
  );


  buf
  g399
  (
    n462,
    n74
  );


  buf
  g400
  (
    n541,
    n54
  );


  buf
  g401
  (
    n516,
    n139
  );


  not
  g402
  (
    n404,
    n64
  );


  buf
  g403
  (
    n588,
    n124
  );


  not
  g404
  (
    KeyWire_0_7,
    n52
  );


  buf
  g405
  (
    n477,
    n99
  );


  not
  g406
  (
    n622,
    n45
  );


  not
  g407
  (
    n547,
    n99
  );


  buf
  g408
  (
    n649,
    n46
  );


  not
  g409
  (
    n470,
    n42
  );


  not
  g410
  (
    n278,
    n44
  );


  not
  g411
  (
    n458,
    n120
  );


  buf
  g412
  (
    n264,
    n135
  );


  not
  g413
  (
    n316,
    n93
  );


  buf
  g414
  (
    n360,
    n118
  );


  buf
  g415
  (
    n194,
    n33
  );


  buf
  g416
  (
    n534,
    n82
  );


  not
  g417
  (
    n415,
    n101
  );


  buf
  g418
  (
    n479,
    n113
  );


  buf
  g419
  (
    n508,
    n97
  );


  buf
  g420
  (
    n418,
    n76
  );


  not
  g421
  (
    n552,
    n46
  );


  not
  g422
  (
    n659,
    n77
  );


  buf
  g423
  (
    n636,
    n87
  );


  not
  g424
  (
    n568,
    n123
  );


  not
  g425
  (
    KeyWire_0_55,
    n85
  );


  not
  g426
  (
    n251,
    n101
  );


  not
  g427
  (
    n287,
    n40
  );


  buf
  g428
  (
    KeyWire_0_1,
    n156
  );


  buf
  g429
  (
    n225,
    n48
  );


  buf
  g430
  (
    n162,
    n136
  );


  buf
  g431
  (
    n182,
    n33
  );


  buf
  g432
  (
    n485,
    n41
  );


  buf
  g433
  (
    n394,
    n151
  );


  buf
  g434
  (
    n280,
    n102
  );


  not
  g435
  (
    n648,
    n97
  );


  buf
  g436
  (
    n387,
    n89
  );


  buf
  g437
  (
    n417,
    n109
  );


  not
  g438
  (
    n282,
    n58
  );


  not
  g439
  (
    n525,
    n94
  );


  buf
  g440
  (
    n589,
    n104
  );


  not
  g441
  (
    n298,
    n142
  );


  not
  g442
  (
    n489,
    n54
  );


  not
  g443
  (
    n612,
    n153
  );


  buf
  g444
  (
    n307,
    n108
  );


  buf
  g445
  (
    n565,
    n72
  );


  not
  g446
  (
    n620,
    n110
  );


  buf
  g447
  (
    n249,
    n58
  );


  not
  g448
  (
    n189,
    n109
  );


  not
  g449
  (
    n439,
    n98
  );


  not
  g450
  (
    n405,
    n121
  );


  buf
  g451
  (
    n440,
    n148
  );


  not
  g452
  (
    n323,
    n67
  );


  buf
  g453
  (
    n538,
    n45
  );


  buf
  g454
  (
    n493,
    n134
  );


  buf
  g455
  (
    n379,
    n116
  );


  not
  g456
  (
    n463,
    n107
  );


  not
  g457
  (
    n258,
    n155
  );


  buf
  g458
  (
    n628,
    n152
  );


  buf
  g459
  (
    n402,
    n40
  );


  not
  g460
  (
    n656,
    n98
  );


  buf
  g461
  (
    n312,
    n110
  );


  not
  g462
  (
    n236,
    n60
  );


  not
  g463
  (
    n625,
    n43
  );


  buf
  g464
  (
    n513,
    n67
  );


  buf
  g465
  (
    n345,
    n150
  );


  buf
  g466
  (
    n452,
    n106
  );


  buf
  g467
  (
    n336,
    n107
  );


  buf
  g468
  (
    n288,
    n58
  );


  not
  g469
  (
    n652,
    n41
  );


  not
  g470
  (
    n531,
    n83
  );


  not
  g471
  (
    n638,
    n122
  );


  not
  g472
  (
    n661,
    n100
  );


  not
  g473
  (
    n524,
    n79
  );


  buf
  g474
  (
    n529,
    n75
  );


  buf
  g475
  (
    n179,
    n155
  );


  not
  g476
  (
    n208,
    n47
  );


  buf
  g477
  (
    n497,
    n121
  );


  buf
  g478
  (
    n637,
    n145
  );


  not
  g479
  (
    n170,
    n141
  );


  not
  g480
  (
    n372,
    n37
  );


  not
  g481
  (
    n246,
    n137
  );


  buf
  g482
  (
    n431,
    n53
  );


  buf
  g483
  (
    n364,
    n115
  );


  buf
  g484
  (
    n277,
    n97
  );


  buf
  g485
  (
    n314,
    n137
  );


  buf
  g486
  (
    n260,
    n147
  );


  not
  g487
  (
    n476,
    n71
  );


  buf
  g488
  (
    n166,
    n98
  );


  not
  g489
  (
    n259,
    n124
  );


  not
  g490
  (
    n606,
    n71
  );


  not
  g491
  (
    KeyWire_0_12,
    n118
  );


  not
  g492
  (
    n527,
    n102
  );


  buf
  g493
  (
    n185,
    n69
  );


  not
  g494
  (
    n370,
    n121
  );


  buf
  g495
  (
    n261,
    n108
  );


  not
  g496
  (
    n294,
    n114
  );


  buf
  g497
  (
    n416,
    n91
  );


  not
  g498
  (
    n544,
    n68
  );


  buf
  g499
  (
    n241,
    n128
  );


  buf
  g500
  (
    n367,
    n112
  );


  buf
  g501
  (
    n517,
    n40
  );


  not
  g502
  (
    n591,
    n41
  );


  not
  g503
  (
    n453,
    n57
  );


  buf
  g504
  (
    n536,
    n138
  );


  not
  g505
  (
    n200,
    n36
  );


  not
  g506
  (
    n410,
    n83
  );


  not
  g507
  (
    n519,
    n132
  );


  not
  g508
  (
    n551,
    n147
  );


  not
  g509
  (
    n634,
    n112
  );


  buf
  g510
  (
    n186,
    n133
  );


  not
  g511
  (
    n478,
    n153
  );


  not
  g512
  (
    n603,
    n124
  );


  buf
  g513
  (
    n579,
    n155
  );


  buf
  g514
  (
    n483,
    n68
  );


  buf
  g515
  (
    n665,
    n143
  );


  buf
  g516
  (
    n655,
    n119
  );


  not
  g517
  (
    n274,
    n64
  );


  not
  g518
  (
    n562,
    n146
  );


  not
  g519
  (
    n239,
    n42
  );


  buf
  g520
  (
    n376,
    n120
  );


  buf
  g521
  (
    n435,
    n132
  );


  not
  g522
  (
    KeyWire_0_10,
    n115
  );


  buf
  g523
  (
    n426,
    n86
  );


  not
  g524
  (
    n214,
    n49
  );


  not
  g525
  (
    n205,
    n96
  );


  not
  g526
  (
    n545,
    n103
  );


  not
  g527
  (
    n238,
    n94
  );


  buf
  g528
  (
    n459,
    n152
  );


  buf
  g529
  (
    n521,
    n138
  );


  not
  g530
  (
    n553,
    n82
  );


  not
  g531
  (
    n610,
    n132
  );


  not
  g532
  (
    n350,
    n69
  );


  buf
  g533
  (
    n495,
    n88
  );


  buf
  g534
  (
    n482,
    n58
  );


  not
  g535
  (
    n256,
    n65
  );


  buf
  g536
  (
    n339,
    n123
  );


  not
  g537
  (
    n533,
    n127
  );


  not
  g538
  (
    n377,
    n125
  );


  not
  g539
  (
    n397,
    n136
  );


  not
  g540
  (
    n305,
    n85
  );


  not
  g541
  (
    n548,
    n157
  );


  buf
  g542
  (
    n666,
    n65
  );


  buf
  g543
  (
    n218,
    n88
  );


  not
  g544
  (
    n330,
    n135
  );


  buf
  g545
  (
    n419,
    n87
  );


  not
  g546
  (
    n598,
    n137
  );


  not
  g547
  (
    n412,
    n111
  );


  not
  g548
  (
    n437,
    n43
  );


  not
  g549
  (
    n284,
    n59
  );


  buf
  g550
  (
    n423,
    n109
  );


  not
  g551
  (
    n248,
    n65
  );


  not
  g552
  (
    n240,
    n134
  );


  not
  g553
  (
    n341,
    n83
  );


  not
  g554
  (
    n210,
    n95
  );


  not
  g555
  (
    n467,
    n128
  );


  buf
  g556
  (
    n268,
    n46
  );


  not
  g557
  (
    n368,
    n129
  );


  not
  g558
  (
    n389,
    n57
  );


  buf
  g559
  (
    n615,
    n94
  );


  not
  g560
  (
    n644,
    n92
  );


  buf
  g561
  (
    n643,
    n88
  );


  not
  g562
  (
    n641,
    n113
  );


  not
  g563
  (
    n279,
    n45
  );


  buf
  g564
  (
    n371,
    n89
  );


  not
  g565
  (
    n272,
    n59
  );


  not
  g566
  (
    n613,
    n67
  );


  buf
  g567
  (
    n595,
    n61
  );


  buf
  g568
  (
    n201,
    n71
  );


  buf
  g569
  (
    n188,
    n78
  );


  buf
  g570
  (
    n393,
    n99
  );


  buf
  g571
  (
    n355,
    n53
  );


  buf
  g572
  (
    n518,
    n113
  );


  buf
  g573
  (
    n542,
    n80
  );


  not
  g574
  (
    n597,
    n145
  );


  buf
  g575
  (
    n348,
    n73
  );


  buf
  g576
  (
    n464,
    n105
  );


  not
  g577
  (
    n532,
    n159
  );


  not
  g578
  (
    n585,
    n91
  );


  not
  g579
  (
    n171,
    n70
  );


  buf
  g580
  (
    n428,
    n49
  );


  buf
  g581
  (
    n425,
    n127
  );


  buf
  g582
  (
    n441,
    n47
  );


  buf
  g583
  (
    n627,
    n79
  );


  buf
  g584
  (
    n528,
    n118
  );


  buf
  g585
  (
    n520,
    n109
  );


  not
  g586
  (
    n445,
    n142
  );


  buf
  g587
  (
    n433,
    n130
  );


  buf
  g588
  (
    n183,
    n140
  );


  buf
  g589
  (
    n420,
    n143
  );


  not
  g590
  (
    n509,
    n82
  );


  not
  g591
  (
    n343,
    n108
  );


  buf
  g592
  (
    n386,
    n136
  );


  not
  g593
  (
    n658,
    n93
  );


  not
  g594
  (
    n492,
    n103
  );


  buf
  g595
  (
    n255,
    n130
  );


  not
  g596
  (
    n401,
    n44
  );


  buf
  g597
  (
    n567,
    n104
  );


  not
  g598
  (
    n320,
    n70
  );


  buf
  g599
  (
    n233,
    n106
  );


  buf
  g600
  (
    n577,
    n92
  );


  not
  g601
  (
    n461,
    n67
  );


  buf
  g602
  (
    n496,
    n76
  );


  not
  g603
  (
    n199,
    n117
  );


  buf
  g604
  (
    n646,
    n105
  );


  buf
  g605
  (
    n473,
    n85
  );


  not
  g606
  (
    n224,
    n70
  );


  buf
  g607
  (
    n299,
    n138
  );


  not
  g608
  (
    n514,
    n48
  );


  buf
  g609
  (
    n176,
    n133
  );


  not
  g610
  (
    n621,
    n148
  );


  not
  g611
  (
    n219,
    n72
  );


  not
  g612
  (
    n530,
    n112
  );


  not
  g613
  (
    n596,
    n64
  );


  buf
  g614
  (
    n281,
    n158
  );


  not
  g615
  (
    n206,
    n93
  );


  buf
  g616
  (
    n346,
    n131
  );


  buf
  g617
  (
    n191,
    n141
  );


  not
  g618
  (
    n315,
    n131
  );


  not
  g619
  (
    n211,
    n144
  );


  buf
  g620
  (
    n327,
    n95
  );


  buf
  g621
  (
    n480,
    n86
  );


  buf
  g622
  (
    n466,
    n101
  );


  buf
  g623
  (
    KeyWire_0_46,
    n114
  );


  buf
  g624
  (
    n391,
    n55
  );


  buf
  g625
  (
    n537,
    n39
  );


  buf
  g626
  (
    n605,
    n110
  );


  buf
  g627
  (
    n293,
    n106
  );


  not
  g628
  (
    n573,
    n89
  );


  not
  g629
  (
    n226,
    n138
  );


  buf
  g630
  (
    n584,
    n61
  );


  buf
  g631
  (
    n430,
    n73
  );


  buf
  g632
  (
    n640,
    n42
  );


  not
  g633
  (
    n630,
    n50
  );


  buf
  g634
  (
    n617,
    n72
  );


  buf
  g635
  (
    n1166,
    n287
  );


  buf
  g636
  (
    n1123,
    n584
  );


  buf
  g637
  (
    n672,
    n162
  );


  not
  g638
  (
    n1412,
    n276
  );


  buf
  g639
  (
    n1540,
    n243
  );


  buf
  g640
  (
    n1325,
    n461
  );


  buf
  g641
  (
    n1193,
    n556
  );


  buf
  g642
  (
    n1405,
    n186
  );


  not
  g643
  (
    n2039,
    n483
  );


  buf
  g644
  (
    n940,
    n298
  );


  not
  g645
  (
    n681,
    n512
  );


  not
  g646
  (
    n1900,
    n343
  );


  not
  g647
  (
    n2048,
    n248
  );


  buf
  g648
  (
    n1105,
    n442
  );


  not
  g649
  (
    n2045,
    n362
  );


  buf
  g650
  (
    n1919,
    n396
  );


  buf
  g651
  (
    n1554,
    n320
  );


  not
  g652
  (
    n1593,
    n256
  );


  not
  g653
  (
    n2052,
    n290
  );


  buf
  g654
  (
    n827,
    n481
  );


  buf
  g655
  (
    n1794,
    n311
  );


  not
  g656
  (
    n1298,
    n571
  );


  buf
  g657
  (
    n1397,
    n318
  );


  not
  g658
  (
    n1760,
    n229
  );


  not
  g659
  (
    n1312,
    n214
  );


  not
  g660
  (
    n1659,
    n370
  );


  buf
  g661
  (
    n1102,
    n454
  );


  buf
  g662
  (
    n1385,
    n534
  );


  not
  g663
  (
    n1493,
    n415
  );


  buf
  g664
  (
    n890,
    n580
  );


  buf
  g665
  (
    n1229,
    n538
  );


  not
  g666
  (
    n1783,
    n274
  );


  buf
  g667
  (
    n745,
    n358
  );


  buf
  g668
  (
    n1471,
    n257
  );


  buf
  g669
  (
    n1004,
    n194
  );


  not
  g670
  (
    n1637,
    n424
  );


  buf
  g671
  (
    n1628,
    n381
  );


  buf
  g672
  (
    n1578,
    n422
  );


  buf
  g673
  (
    n671,
    n509
  );


  not
  g674
  (
    n1551,
    n517
  );


  not
  g675
  (
    n1662,
    n610
  );


  not
  g676
  (
    n1445,
    n591
  );


  not
  g677
  (
    n1145,
    n656
  );


  buf
  g678
  (
    n1805,
    n527
  );


  buf
  g679
  (
    n2040,
    n399
  );


  not
  g680
  (
    n1894,
    n386
  );


  buf
  g681
  (
    n686,
    n535
  );


  buf
  g682
  (
    n1721,
    n463
  );


  not
  g683
  (
    n712,
    n620
  );


  not
  g684
  (
    n1311,
    n248
  );


  buf
  g685
  (
    n2005,
    n340
  );


  buf
  g686
  (
    n1120,
    n326
  );


  not
  g687
  (
    n1726,
    n423
  );


  not
  g688
  (
    n1083,
    n604
  );


  not
  g689
  (
    n791,
    n238
  );


  not
  g690
  (
    n1428,
    n595
  );


  buf
  g691
  (
    n888,
    n305
  );


  not
  g692
  (
    n785,
    n401
  );


  buf
  g693
  (
    n1916,
    n437
  );


  buf
  g694
  (
    n1613,
    n612
  );


  not
  g695
  (
    n1347,
    n572
  );


  not
  g696
  (
    n1778,
    n302
  );


  not
  g697
  (
    n1513,
    n545
  );


  not
  g698
  (
    n1737,
    n322
  );


  not
  g699
  (
    n1108,
    n513
  );


  not
  g700
  (
    n1795,
    n218
  );


  buf
  g701
  (
    n1252,
    n618
  );


  buf
  g702
  (
    n1764,
    n658
  );


  buf
  g703
  (
    n1885,
    n427
  );


  buf
  g704
  (
    n2056,
    n410
  );


  buf
  g705
  (
    n1463,
    n538
  );


  not
  g706
  (
    n1130,
    n310
  );


  not
  g707
  (
    n1107,
    n261
  );


  buf
  g708
  (
    n1742,
    n499
  );


  not
  g709
  (
    n1801,
    n193
  );


  buf
  g710
  (
    n994,
    n223
  );


  buf
  g711
  (
    n1183,
    n246
  );


  buf
  g712
  (
    n874,
    n181
  );


  buf
  g713
  (
    n1433,
    n383
  );


  buf
  g714
  (
    n1806,
    n217
  );


  buf
  g715
  (
    n1909,
    n240
  );


  buf
  g716
  (
    n1887,
    n367
  );


  buf
  g717
  (
    n1202,
    n349
  );


  buf
  g718
  (
    n919,
    n261
  );


  not
  g719
  (
    n1976,
    n633
  );


  buf
  g720
  (
    n1310,
    n246
  );


  buf
  g721
  (
    n1355,
    n328
  );


  buf
  g722
  (
    n2008,
    n272
  );


  buf
  g723
  (
    n1218,
    n315
  );


  not
  g724
  (
    n2023,
    n181
  );


  buf
  g725
  (
    n868,
    n547
  );


  buf
  g726
  (
    n884,
    n266
  );


  not
  g727
  (
    n1625,
    n194
  );


  not
  g728
  (
    n1803,
    n546
  );


  buf
  g729
  (
    n959,
    n536
  );


  buf
  g730
  (
    n1063,
    n501
  );


  not
  g731
  (
    n1978,
    n654
  );


  buf
  g732
  (
    n1251,
    n641
  );


  not
  g733
  (
    n1039,
    n629
  );


  not
  g734
  (
    n2053,
    n436
  );


  buf
  g735
  (
    n1907,
    n579
  );


  buf
  g736
  (
    KeyWire_0_39,
    n536
  );


  not
  g737
  (
    n1373,
    n476
  );


  buf
  g738
  (
    n1830,
    n510
  );


  buf
  g739
  (
    n1963,
    n180
  );


  buf
  g740
  (
    n1423,
    n180
  );


  buf
  g741
  (
    n1623,
    n505
  );


  buf
  g742
  (
    n1016,
    n514
  );


  buf
  g743
  (
    n1117,
    n232
  );


  not
  g744
  (
    n1652,
    n379
  );


  not
  g745
  (
    n1159,
    n581
  );


  buf
  g746
  (
    n1380,
    n205
  );


  buf
  g747
  (
    n1605,
    n550
  );


  not
  g748
  (
    n1324,
    n525
  );


  buf
  g749
  (
    n1537,
    n616
  );


  not
  g750
  (
    n1781,
    n558
  );


  not
  g751
  (
    n1481,
    n599
  );


  buf
  g752
  (
    n1786,
    n262
  );


  not
  g753
  (
    n693,
    n539
  );


  not
  g754
  (
    n1636,
    n533
  );


  not
  g755
  (
    n1555,
    n273
  );


  buf
  g756
  (
    n825,
    n420
  );


  not
  g757
  (
    n931,
    n434
  );


  buf
  g758
  (
    n1644,
    n210
  );


  not
  g759
  (
    n1695,
    n244
  );


  not
  g760
  (
    n687,
    n255
  );


  not
  g761
  (
    n1379,
    n628
  );


  not
  g762
  (
    n947,
    n252
  );


  not
  g763
  (
    KeyWire_0_3,
    n629
  );


  not
  g764
  (
    n2060,
    n305
  );


  not
  g765
  (
    n1844,
    n625
  );


  not
  g766
  (
    n1530,
    n161
  );


  buf
  g767
  (
    n1138,
    n296
  );


  not
  g768
  (
    n720,
    n580
  );


  not
  g769
  (
    n1059,
    n347
  );


  not
  g770
  (
    n877,
    n446
  );


  not
  g771
  (
    n1182,
    n486
  );


  not
  g772
  (
    n1404,
    n569
  );


  not
  g773
  (
    n751,
    n492
  );


  buf
  g774
  (
    KeyWire_0_20,
    n171
  );


  buf
  g775
  (
    n1687,
    n520
  );


  buf
  g776
  (
    n723,
    n421
  );


  not
  g777
  (
    n1585,
    n561
  );


  buf
  g778
  (
    n1727,
    n313
  );


  buf
  g779
  (
    n1848,
    n489
  );


  buf
  g780
  (
    n1686,
    n577
  );


  buf
  g781
  (
    n1874,
    n347
  );


  not
  g782
  (
    n1579,
    n310
  );


  buf
  g783
  (
    n1257,
    n200
  );


  buf
  g784
  (
    n944,
    n491
  );


  buf
  g785
  (
    n698,
    n607
  );


  buf
  g786
  (
    n1349,
    n549
  );


  not
  g787
  (
    n1739,
    n610
  );


  not
  g788
  (
    n1612,
    n389
  );


  buf
  g789
  (
    n1892,
    n229
  );


  not
  g790
  (
    n908,
    n297
  );


  not
  g791
  (
    n1583,
    n462
  );


  buf
  g792
  (
    n1003,
    n458
  );


  not
  g793
  (
    n1790,
    n273
  );


  not
  g794
  (
    n1465,
    n645
  );


  not
  g795
  (
    n1072,
    n402
  );


  not
  g796
  (
    n807,
    n402
  );


  not
  g797
  (
    n1871,
    n635
  );


  buf
  g798
  (
    n1890,
    n585
  );


  not
  g799
  (
    n984,
    n507
  );


  buf
  g800
  (
    n1993,
    n574
  );


  not
  g801
  (
    n1563,
    n642
  );


  not
  g802
  (
    n1034,
    n562
  );


  buf
  g803
  (
    n673,
    n581
  );


  buf
  g804
  (
    n1482,
    n513
  );


  not
  g805
  (
    n1996,
    n233
  );


  not
  g806
  (
    n1852,
    n649
  );


  not
  g807
  (
    n796,
    n274
  );


  buf
  g808
  (
    n1119,
    n224
  );


  buf
  g809
  (
    n1046,
    n529
  );


  buf
  g810
  (
    KeyWire_0_63,
    n344
  );


  buf
  g811
  (
    n1490,
    n381
  );


  buf
  g812
  (
    n1525,
    n348
  );


  not
  g813
  (
    n2000,
    n652
  );


  buf
  g814
  (
    n1424,
    n191
  );


  buf
  g815
  (
    n1167,
    n569
  );


  buf
  g816
  (
    n2050,
    n592
  );


  buf
  g817
  (
    n1330,
    n384
  );


  buf
  g818
  (
    n852,
    n612
  );


  not
  g819
  (
    n1562,
    n212
  );


  not
  g820
  (
    n1384,
    n237
  );


  buf
  g821
  (
    n1126,
    n438
  );


  buf
  g822
  (
    n1337,
    n566
  );


  not
  g823
  (
    n1431,
    n357
  );


  not
  g824
  (
    n806,
    n654
  );


  buf
  g825
  (
    n1222,
    n299
  );


  not
  g826
  (
    n1589,
    n624
  );


  not
  g827
  (
    n1366,
    n453
  );


  not
  g828
  (
    n2062,
    n617
  );


  buf
  g829
  (
    n2064,
    n550
  );


  not
  g830
  (
    n1580,
    n531
  );


  not
  g831
  (
    n1041,
    n554
  );


  not
  g832
  (
    n702,
    n236
  );


  not
  g833
  (
    n1260,
    n341
  );


  buf
  g834
  (
    n1084,
    n200
  );


  buf
  g835
  (
    n808,
    n287
  );


  not
  g836
  (
    n830,
    n295
  );


  not
  g837
  (
    n1219,
    n592
  );


  not
  g838
  (
    n1817,
    n594
  );


  buf
  g839
  (
    n1044,
    n405
  );


  not
  g840
  (
    n1376,
    n293
  );


  buf
  g841
  (
    n1671,
    n429
  );


  buf
  g842
  (
    n1870,
    n496
  );


  buf
  g843
  (
    n1581,
    n518
  );


  buf
  g844
  (
    n1655,
    n377
  );


  buf
  g845
  (
    n1591,
    n232
  );


  not
  g846
  (
    n1574,
    n188
  );


  not
  g847
  (
    n1825,
    n491
  );


  buf
  g848
  (
    n1439,
    n242
  );


  buf
  g849
  (
    n2047,
    n173
  );


  not
  g850
  (
    n1944,
    n227
  );


  not
  g851
  (
    n1058,
    n431
  );


  buf
  g852
  (
    n1715,
    n362
  );


  buf
  g853
  (
    n1104,
    n212
  );


  not
  g854
  (
    n1435,
    n229
  );


  not
  g855
  (
    n1019,
    n498
  );


  not
  g856
  (
    n933,
    n394
  );


  buf
  g857
  (
    n1519,
    n532
  );


  buf
  g858
  (
    n1277,
    n597
  );


  not
  g859
  (
    n1055,
    n419
  );


  buf
  g860
  (
    n1970,
    n254
  );


  not
  g861
  (
    n861,
    n426
  );


  not
  g862
  (
    n1352,
    n588
  );


  buf
  g863
  (
    n1827,
    n244
  );


  not
  g864
  (
    n1565,
    n224
  );


  buf
  g865
  (
    n1576,
    n485
  );


  not
  g866
  (
    n1881,
    n573
  );


  not
  g867
  (
    n2049,
    n314
  );


  buf
  g868
  (
    n1535,
    n653
  );


  not
  g869
  (
    n1416,
    n620
  );


  buf
  g870
  (
    n1955,
    n194
  );


  not
  g871
  (
    n1680,
    n324
  );


  not
  g872
  (
    n1784,
    n560
  );


  buf
  g873
  (
    n855,
    n326
  );


  buf
  g874
  (
    n1747,
    n444
  );


  buf
  g875
  (
    n1789,
    n427
  );


  buf
  g876
  (
    n1953,
    n581
  );


  buf
  g877
  (
    n1816,
    n303
  );


  not
  g878
  (
    n1168,
    n308
  );


  buf
  g879
  (
    n951,
    n463
  );


  buf
  g880
  (
    n1334,
    n363
  );


  not
  g881
  (
    n1032,
    n608
  );


  not
  g882
  (
    n1908,
    n164
  );


  buf
  g883
  (
    n1914,
    n211
  );


  buf
  g884
  (
    n1195,
    n223
  );


  not
  g885
  (
    n977,
    n460
  );


  buf
  g886
  (
    n1876,
    n267
  );


  buf
  g887
  (
    n1823,
    n303
  );


  buf
  g888
  (
    KeyWire_0_6,
    n256
  );


  not
  g889
  (
    n1300,
    n553
  );


  buf
  g890
  (
    n1474,
    n457
  );


  not
  g891
  (
    n1399,
    n571
  );


  not
  g892
  (
    n1141,
    n352
  );


  not
  g893
  (
    n1160,
    n566
  );


  not
  g894
  (
    n911,
    n425
  );


  not
  g895
  (
    n927,
    n624
  );


  not
  g896
  (
    n882,
    n553
  );


  buf
  g897
  (
    n1668,
    n543
  );


  not
  g898
  (
    n1429,
    n234
  );


  buf
  g899
  (
    n1223,
    n162
  );


  not
  g900
  (
    n930,
    n492
  );


  not
  g901
  (
    n773,
    n204
  );


  buf
  g902
  (
    n1889,
    n269
  );


  buf
  g903
  (
    n1089,
    n306
  );


  not
  g904
  (
    n1146,
    n495
  );


  buf
  g905
  (
    n753,
    n428
  );


  not
  g906
  (
    n771,
    n179
  );


  buf
  g907
  (
    n1045,
    n530
  );


  not
  g908
  (
    n840,
    n541
  );


  not
  g909
  (
    n1199,
    n247
  );


  not
  g910
  (
    n2055,
    n341
  );


  buf
  g911
  (
    n1246,
    n572
  );


  not
  g912
  (
    n1539,
    n619
  );


  buf
  g913
  (
    n1922,
    n396
  );


  not
  g914
  (
    KeyWire_0_0,
    n600
  );


  buf
  g915
  (
    n777,
    n302
  );


  not
  g916
  (
    n1279,
    n653
  );


  not
  g917
  (
    n1174,
    n206
  );


  not
  g918
  (
    n815,
    n646
  );


  buf
  g919
  (
    n1931,
    n293
  );


  buf
  g920
  (
    n1499,
    n431
  );


  buf
  g921
  (
    n1171,
    n600
  );


  buf
  g922
  (
    n838,
    n402
  );


  buf
  g923
  (
    n1175,
    n311
  );


  not
  g924
  (
    n737,
    n648
  );


  not
  g925
  (
    n1484,
    n558
  );


  buf
  g926
  (
    n1736,
    n249
  );


  buf
  g927
  (
    n797,
    n379
  );


  buf
  g928
  (
    n859,
    n265
  );


  buf
  g929
  (
    n725,
    n215
  );


  buf
  g930
  (
    n2016,
    n236
  );


  buf
  g931
  (
    n1047,
    n242
  );


  buf
  g932
  (
    n1440,
    n202
  );


  buf
  g933
  (
    n1078,
    n225
  );


  buf
  g934
  (
    n701,
    n476
  );


  not
  g935
  (
    n1014,
    n365
  );


  buf
  g936
  (
    n1618,
    n358
  );


  not
  g937
  (
    n1271,
    n561
  );


  not
  g938
  (
    n750,
    n528
  );


  not
  g939
  (
    n1708,
    n318
  );


  buf
  g940
  (
    n722,
    n254
  );


  not
  g941
  (
    n689,
    n475
  );


  buf
  g942
  (
    n2034,
    n472
  );


  not
  g943
  (
    n1609,
    n342
  );


  not
  g944
  (
    n1648,
    n585
  );


  not
  g945
  (
    n1491,
    n261
  );


  not
  g946
  (
    n1319,
    n517
  );


  not
  g947
  (
    n821,
    n560
  );


  buf
  g948
  (
    n1828,
    n601
  );


  buf
  g949
  (
    n1883,
    n334
  );


  buf
  g950
  (
    n858,
    n584
  );


  not
  g951
  (
    KeyWire_0_38,
    n580
  );


  not
  g952
  (
    n1149,
    n494
  );


  not
  g953
  (
    n1582,
    n593
  );


  not
  g954
  (
    n1520,
    n163
  );


  not
  g955
  (
    KeyWire_0_57,
    n605
  );


  not
  g956
  (
    n1851,
    n448
  );


  not
  g957
  (
    n1443,
    n175
  );


  buf
  g958
  (
    n894,
    n214
  );


  buf
  g959
  (
    n814,
    n609
  );


  buf
  g960
  (
    n670,
    n486
  );


  not
  g961
  (
    n1163,
    n174
  );


  not
  g962
  (
    n820,
    n241
  );


  buf
  g963
  (
    n1457,
    n265
  );


  buf
  g964
  (
    n1284,
    n228
  );


  buf
  g965
  (
    n1452,
    n238
  );


  not
  g966
  (
    n1239,
    n263
  );


  buf
  g967
  (
    n849,
    n483
  );


  buf
  g968
  (
    n709,
    n569
  );


  buf
  g969
  (
    n870,
    n282
  );


  not
  g970
  (
    n1450,
    n532
  );


  buf
  g971
  (
    n1361,
    n317
  );


  not
  g972
  (
    n2011,
    n332
  );


  buf
  g973
  (
    n1940,
    n631
  );


  buf
  g974
  (
    n1928,
    n401
  );


  not
  g975
  (
    n1545,
    n427
  );


  buf
  g976
  (
    n1626,
    n374
  );


  not
  g977
  (
    n1902,
    n186
  );


  not
  g978
  (
    n1321,
    n582
  );


  buf
  g979
  (
    n1873,
    n176
  );


  not
  g980
  (
    n1897,
    n367
  );


  buf
  g981
  (
    n983,
    n295
  );


  not
  g982
  (
    n1552,
    n559
  );


  not
  g983
  (
    n1392,
    n485
  );


  not
  g984
  (
    n776,
    n643
  );


  buf
  g985
  (
    n1432,
    n656
  );


  not
  g986
  (
    n1531,
    n431
  );


  not
  g987
  (
    n679,
    n479
  );


  not
  g988
  (
    n1469,
    n549
  );


  not
  g989
  (
    n762,
    n639
  );


  not
  g990
  (
    n740,
    n200
  );


  not
  g991
  (
    n1676,
    n559
  );


  not
  g992
  (
    n1086,
    n309
  );


  not
  g993
  (
    n924,
    n329
  );


  not
  g994
  (
    n1864,
    n392
  );


  not
  g995
  (
    n1462,
    n575
  );


  not
  g996
  (
    n1548,
    n308
  );


  not
  g997
  (
    n1233,
    n645
  );


  not
  g998
  (
    n1225,
    n273
  );


  buf
  g999
  (
    n1473,
    n166
  );


  buf
  g1000
  (
    n829,
    n567
  );


  not
  g1001
  (
    n789,
    n552
  );


  not
  g1002
  (
    n975,
    n657
  );


  not
  g1003
  (
    n1918,
    n543
  );


  buf
  g1004
  (
    n1254,
    n630
  );


  not
  g1005
  (
    n1365,
    n363
  );


  buf
  g1006
  (
    n2041,
    n458
  );


  not
  g1007
  (
    n1112,
    n477
  );


  not
  g1008
  (
    n1913,
    n364
  );


  not
  g1009
  (
    n986,
    n223
  );


  not
  g1010
  (
    n1453,
    n464
  );


  buf
  g1011
  (
    n1950,
    n226
  );


  buf
  g1012
  (
    n764,
    n631
  );


  buf
  g1013
  (
    n889,
    n532
  );


  not
  g1014
  (
    n2018,
    n507
  );


  buf
  g1015
  (
    n993,
    n506
  );


  buf
  g1016
  (
    n1504,
    n559
  );


  not
  g1017
  (
    n1994,
    n326
  );


  buf
  g1018
  (
    n1189,
    n318
  );


  buf
  g1019
  (
    n1678,
    n412
  );


  not
  g1020
  (
    n1688,
    n166
  );


  not
  g1021
  (
    n1466,
    n187
  );


  buf
  g1022
  (
    n863,
    n473
  );


  not
  g1023
  (
    n998,
    n457
  );


  buf
  g1024
  (
    n1326,
    n311
  );


  buf
  g1025
  (
    n792,
    n578
  );


  buf
  g1026
  (
    n989,
    n202
  );


  buf
  g1027
  (
    n891,
    n626
  );


  buf
  g1028
  (
    n1304,
    n604
  );


  not
  g1029
  (
    n1230,
    n389
  );


  buf
  g1030
  (
    n1467,
    n422
  );


  not
  g1031
  (
    n968,
    n399
  );


  not
  g1032
  (
    n923,
    n296
  );


  buf
  g1033
  (
    n1584,
    n573
  );


  not
  g1034
  (
    n1372,
    n508
  );


  not
  g1035
  (
    n842,
    n559
  );


  not
  g1036
  (
    n860,
    n576
  );


  buf
  g1037
  (
    n1653,
    n425
  );


  buf
  g1038
  (
    n990,
    n424
  );


  not
  g1039
  (
    n1840,
    n584
  );


  buf
  g1040
  (
    n822,
    n467
  );


  not
  g1041
  (
    n783,
    n511
  );


  not
  g1042
  (
    n1698,
    n316
  );


  buf
  g1043
  (
    n1705,
    n221
  );


  not
  g1044
  (
    n1062,
    n516
  );


  buf
  g1045
  (
    n1723,
    n314
  );


  buf
  g1046
  (
    n1756,
    n617
  );


  buf
  g1047
  (
    n1176,
    n497
  );


  not
  g1048
  (
    n1620,
    n387
  );


  buf
  g1049
  (
    n1483,
    n400
  );


  not
  g1050
  (
    n1656,
    n390
  );


  not
  g1051
  (
    n1394,
    n602
  );


  not
  g1052
  (
    n744,
    n230
  );


  buf
  g1053
  (
    n1422,
    n259
  );


  buf
  g1054
  (
    n1588,
    n442
  );


  not
  g1055
  (
    n2044,
    n324
  );


  buf
  g1056
  (
    n1192,
    n657
  );


  not
  g1057
  (
    n1170,
    n454
  );


  buf
  g1058
  (
    n1538,
    n575
  );


  not
  g1059
  (
    n1947,
    n215
  );


  buf
  g1060
  (
    n1038,
    n333
  );


  buf
  g1061
  (
    KeyWire_0_48,
    n615
  );


  not
  g1062
  (
    n1140,
    n590
  );


  buf
  g1063
  (
    n904,
    n522
  );


  not
  g1064
  (
    n969,
    n475
  );


  buf
  g1065
  (
    n1703,
    n369
  );


  buf
  g1066
  (
    n1964,
    n216
  );


  not
  g1067
  (
    KeyWire_0_14,
    n505
  );


  not
  g1068
  (
    n950,
    n573
  );


  buf
  g1069
  (
    n1081,
    n285
  );


  buf
  g1070
  (
    n1920,
    n555
  );


  not
  g1071
  (
    n1670,
    n447
  );


  not
  g1072
  (
    n2022,
    n620
  );


  buf
  g1073
  (
    n1846,
    n306
  );


  not
  g1074
  (
    n850,
    n634
  );


  not
  g1075
  (
    n1200,
    n477
  );


  not
  g1076
  (
    n1426,
    n220
  );


  not
  g1077
  (
    n1501,
    n484
  );


  buf
  g1078
  (
    n1037,
    n356
  );


  not
  g1079
  (
    n748,
    n611
  );


  buf
  g1080
  (
    n1353,
    n177
  );


  buf
  g1081
  (
    n1370,
    n319
  );


  not
  g1082
  (
    n1549,
    n310
  );


  not
  g1083
  (
    KeyWire_0_22,
    n526
  );


  buf
  g1084
  (
    n811,
    n191
  );


  buf
  g1085
  (
    n1363,
    n564
  );


  buf
  g1086
  (
    n2033,
    n462
  );


  buf
  g1087
  (
    n768,
    n573
  );


  buf
  g1088
  (
    n1697,
    n257
  );


  buf
  g1089
  (
    n2043,
    n582
  );


  buf
  g1090
  (
    n668,
    n544
  );


  not
  g1091
  (
    n1657,
    n633
  );


  buf
  g1092
  (
    n1543,
    n184
  );


  buf
  g1093
  (
    n1728,
    n491
  );


  not
  g1094
  (
    n1398,
    n520
  );


  buf
  g1095
  (
    n1268,
    n551
  );


  not
  g1096
  (
    n2029,
    n242
  );


  buf
  g1097
  (
    n938,
    n605
  );


  buf
  g1098
  (
    n1459,
    n430
  );


  not
  g1099
  (
    n1401,
    n218
  );


  not
  g1100
  (
    n1293,
    n161
  );


  buf
  g1101
  (
    n1956,
    n578
  );


  buf
  g1102
  (
    n1295,
    n631
  );


  buf
  g1103
  (
    n1489,
    n348
  );


  not
  g1104
  (
    n1027,
    n172
  );


  buf
  g1105
  (
    n1270,
    n656
  );


  not
  g1106
  (
    n1345,
    n165
  );


  not
  g1107
  (
    n1028,
    n416
  );


  buf
  g1108
  (
    n1194,
    n332
  );


  buf
  g1109
  (
    n1523,
    n363
  );


  not
  g1110
  (
    n1796,
    n520
  );


  buf
  g1111
  (
    n1810,
    n410
  );


  buf
  g1112
  (
    n2004,
    n315
  );


  not
  g1113
  (
    n1356,
    n340
  );


  not
  g1114
  (
    n1734,
    n641
  );


  buf
  g1115
  (
    n1822,
    n555
  );


  buf
  g1116
  (
    n1346,
    n425
  );


  not
  g1117
  (
    n758,
    n373
  );


  not
  g1118
  (
    n1294,
    n586
  );


  not
  g1119
  (
    n1461,
    n276
  );


  buf
  g1120
  (
    n1224,
    n654
  );


  buf
  g1121
  (
    n1629,
    n425
  );


  not
  g1122
  (
    n1559,
    n613
  );


  buf
  g1123
  (
    n1673,
    n231
  );


  not
  g1124
  (
    n1834,
    n528
  );


  buf
  g1125
  (
    n833,
    n351
  );


  not
  g1126
  (
    n1097,
    n439
  );


  buf
  g1127
  (
    n1843,
    n359
  );


  not
  g1128
  (
    n960,
    n394
  );


  not
  g1129
  (
    n738,
    n608
  );


  buf
  g1130
  (
    n921,
    n354
  );


  not
  g1131
  (
    n1702,
    n644
  );


  not
  g1132
  (
    n1558,
    n507
  );


  buf
  g1133
  (
    n1709,
    n515
  );


  buf
  g1134
  (
    n1568,
    n385
  );


  buf
  g1135
  (
    n1616,
    n616
  );


  buf
  g1136
  (
    n1318,
    n258
  );


  not
  g1137
  (
    n1930,
    n458
  );


  not
  g1138
  (
    n2002,
    n167
  );


  not
  g1139
  (
    n2017,
    n643
  );


  not
  g1140
  (
    n1905,
    n562
  );


  buf
  g1141
  (
    n717,
    n545
  );


  buf
  g1142
  (
    n1941,
    n278
  );


  not
  g1143
  (
    n976,
    n393
  );


  buf
  g1144
  (
    n1173,
    n539
  );


  buf
  g1145
  (
    n1237,
    n424
  );


  buf
  g1146
  (
    n731,
    n465
  );


  not
  g1147
  (
    n1516,
    n587
  );


  not
  g1148
  (
    n932,
    n343
  );


  buf
  g1149
  (
    n1155,
    n503
  );


  buf
  g1150
  (
    n1820,
    n480
  );


  buf
  g1151
  (
    n824,
    n623
  );


  buf
  g1152
  (
    n1065,
    n611
  );


  buf
  g1153
  (
    n1243,
    n441
  );


  not
  g1154
  (
    n1975,
    n165
  );


  buf
  g1155
  (
    n961,
    n285
  );


  not
  g1156
  (
    n1071,
    n300
  );


  not
  g1157
  (
    n1446,
    n426
  );


  buf
  g1158
  (
    n1910,
    n624
  );


  not
  g1159
  (
    n684,
    n541
  );


  not
  g1160
  (
    n2026,
    n330
  );


  not
  g1161
  (
    n1035,
    n266
  );


  not
  g1162
  (
    n1600,
    n270
  );


  not
  g1163
  (
    n1402,
    n262
  );


  not
  g1164
  (
    n752,
    n445
  );


  buf
  g1165
  (
    n866,
    n185
  );


  buf
  g1166
  (
    n1275,
    n288
  );


  buf
  g1167
  (
    n1377,
    n251
  );


  buf
  g1168
  (
    n2037,
    n631
  );


  buf
  g1169
  (
    n907,
    n449
  );


  not
  g1170
  (
    n728,
    n463
  );


  buf
  g1171
  (
    n1599,
    n531
  );


  not
  g1172
  (
    n1536,
    n488
  );


  not
  g1173
  (
    KeyWire_0_8,
    n211
  );


  buf
  g1174
  (
    n1925,
    n653
  );


  buf
  g1175
  (
    n913,
    n225
  );


  not
  g1176
  (
    n1660,
    n328
  );


  not
  g1177
  (
    n971,
    n516
  );


  buf
  g1178
  (
    n1814,
    n288
  );


  buf
  g1179
  (
    n1464,
    n557
  );


  buf
  g1180
  (
    n1946,
    n283
  );


  not
  g1181
  (
    n688,
    n622
  );


  buf
  g1182
  (
    n945,
    n397
  );


  buf
  g1183
  (
    n920,
    n382
  );


  not
  g1184
  (
    n1100,
    n375
  );


  buf
  g1185
  (
    n1966,
    n297
  );


  buf
  g1186
  (
    n1651,
    n502
  );


  not
  g1187
  (
    n1507,
    n314
  );


  buf
  g1188
  (
    n1498,
    n211
  );


  buf
  g1189
  (
    n1235,
    n504
  );


  not
  g1190
  (
    n1276,
    n321
  );


  not
  g1191
  (
    n1896,
    n552
  );


  not
  g1192
  (
    n1681,
    n178
  );


  not
  g1193
  (
    n1116,
    n634
  );


  not
  g1194
  (
    n848,
    n320
  );


  buf
  g1195
  (
    n881,
    n456
  );


  not
  g1196
  (
    n793,
    n515
  );


  buf
  g1197
  (
    n1407,
    n216
  );


  buf
  g1198
  (
    n1357,
    n429
  );


  buf
  g1199
  (
    n1350,
    n629
  );


  buf
  g1200
  (
    n1258,
    n534
  );


  not
  g1201
  (
    n1241,
    n286
  );


  buf
  g1202
  (
    n1860,
    n231
  );


  buf
  g1203
  (
    n1775,
    n293
  );


  not
  g1204
  (
    n818,
    n231
  );


  not
  g1205
  (
    n1906,
    n587
  );


  buf
  g1206
  (
    n1307,
    n398
  );


  not
  g1207
  (
    n1152,
    n524
  );


  not
  g1208
  (
    n2067,
    n527
  );


  buf
  g1209
  (
    n1001,
    n506
  );


  not
  g1210
  (
    n1060,
    n626
  );


  buf
  g1211
  (
    n1634,
    n317
  );


  not
  g1212
  (
    n1135,
    n225
  );


  buf
  g1213
  (
    n1043,
    n246
  );


  not
  g1214
  (
    n1190,
    n369
  );


  not
  g1215
  (
    n1121,
    n611
  );


  not
  g1216
  (
    n1073,
    n615
  );


  buf
  g1217
  (
    n928,
    n400
  );


  buf
  g1218
  (
    n1767,
    n357
  );


  buf
  g1219
  (
    n1777,
    n497
  );


  buf
  g1220
  (
    n1017,
    n603
  );


  not
  g1221
  (
    n1389,
    n279
  );


  not
  g1222
  (
    n1912,
    n180
  );


  not
  g1223
  (
    n1212,
    n221
  );


  not
  g1224
  (
    n917,
    n327
  );


  buf
  g1225
  (
    n1632,
    n567
  );


  not
  g1226
  (
    n1962,
    n593
  );


  not
  g1227
  (
    n1948,
    n254
  );


  buf
  g1228
  (
    n1454,
    n192
  );


  not
  g1229
  (
    n979,
    n595
  );


  buf
  g1230
  (
    n1147,
    n245
  );


  buf
  g1231
  (
    n1408,
    n490
  );


  buf
  g1232
  (
    n2066,
    n331
  );


  not
  g1233
  (
    n756,
    n640
  );


  buf
  g1234
  (
    n1406,
    n437
  );


  buf
  g1235
  (
    n1051,
    n583
  );


  buf
  g1236
  (
    n1798,
    n335
  );


  not
  g1237
  (
    n1952,
    n229
  );


  not
  g1238
  (
    n1561,
    n638
  );


  not
  g1239
  (
    KeyWire_0_28,
    n636
  );


  not
  g1240
  (
    n909,
    n287
  );


  buf
  g1241
  (
    n1185,
    n596
  );


  not
  g1242
  (
    n1633,
    n543
  );


  not
  g1243
  (
    n1641,
    n535
  );


  not
  g1244
  (
    n1023,
    n437
  );


  not
  g1245
  (
    n1460,
    n288
  );


  buf
  g1246
  (
    n1746,
    n474
  );


  not
  g1247
  (
    n1476,
    n170
  );


  not
  g1248
  (
    n1811,
    n364
  );


  buf
  g1249
  (
    n696,
    n602
  );


  buf
  g1250
  (
    n1765,
    n621
  );


  buf
  g1251
  (
    n1831,
    n561
  );


  not
  g1252
  (
    n1569,
    n491
  );


  buf
  g1253
  (
    n1979,
    n512
  );


  not
  g1254
  (
    n779,
    n398
  );


  not
  g1255
  (
    n835,
    n167
  );


  buf
  g1256
  (
    n1521,
    n500
  );


  not
  g1257
  (
    n1750,
    n568
  );


  not
  g1258
  (
    n1977,
    n384
  );


  not
  g1259
  (
    n1244,
    n249
  );


  buf
  g1260
  (
    n1511,
    n470
  );


  buf
  g1261
  (
    n1541,
    n421
  );


  buf
  g1262
  (
    n1631,
    n198
  );


  not
  g1263
  (
    n1101,
    n644
  );


  buf
  g1264
  (
    n1942,
    n266
  );


  buf
  g1265
  (
    n1221,
    n263
  );


  not
  g1266
  (
    n1344,
    n207
  );


  not
  g1267
  (
    n966,
    n355
  );


  not
  g1268
  (
    n1730,
    n278
  );


  not
  g1269
  (
    n1154,
    n470
  );


  buf
  g1270
  (
    n845,
    n432
  );


  not
  g1271
  (
    n804,
    n194
  );


  buf
  g1272
  (
    n1619,
    n358
  );


  buf
  g1273
  (
    n805,
    n290
  );


  not
  g1274
  (
    n957,
    n172
  );


  buf
  g1275
  (
    n1502,
    n635
  );


  not
  g1276
  (
    n1510,
    n365
  );


  not
  g1277
  (
    n2003,
    n344
  );


  not
  g1278
  (
    n1187,
    n197
  );


  buf
  g1279
  (
    n1603,
    n393
  );


  not
  g1280
  (
    n1699,
    n473
  );


  not
  g1281
  (
    n1639,
    n615
  );


  not
  g1282
  (
    n1413,
    n391
  );


  buf
  g1283
  (
    n1720,
    n361
  );


  not
  g1284
  (
    n1437,
    n558
  );


  buf
  g1285
  (
    n1191,
    n515
  );


  not
  g1286
  (
    n1472,
    n383
  );


  buf
  g1287
  (
    n2012,
    n423
  );


  not
  g1288
  (
    n1951,
    n483
  );


  buf
  g1289
  (
    n1165,
    n356
  );


  buf
  g1290
  (
    n1694,
    n409
  );


  buf
  g1291
  (
    n1068,
    n640
  );


  not
  g1292
  (
    n1049,
    n367
  );


  not
  g1293
  (
    n1506,
    n338
  );


  buf
  g1294
  (
    n1761,
    n222
  );


  buf
  g1295
  (
    n1779,
    n536
  );


  not
  g1296
  (
    n1480,
    n266
  );


  buf
  g1297
  (
    n1438,
    n528
  );


  not
  g1298
  (
    n1759,
    n350
  );


  not
  g1299
  (
    n1571,
    n274
  );


  not
  g1300
  (
    n1306,
    n171
  );


  not
  g1301
  (
    n1999,
    n178
  );


  not
  g1302
  (
    n1248,
    n304
  );


  not
  g1303
  (
    KeyWire_0_60,
    n464
  );


  buf
  g1304
  (
    n1867,
    n445
  );


  buf
  g1305
  (
    n1283,
    n219
  );


  buf
  g1306
  (
    n826,
    n544
  );


  not
  g1307
  (
    n1934,
    n304
  );


  buf
  g1308
  (
    n1855,
    n468
  );


  buf
  g1309
  (
    n1606,
    n397
  );


  buf
  g1310
  (
    KeyWire_0_47,
    n513
  );


  not
  g1311
  (
    n1391,
    n302
  );


  not
  g1312
  (
    n1247,
    n184
  );


  not
  g1313
  (
    n1316,
    n464
  );


  not
  g1314
  (
    n1837,
    n333
  );


  buf
  g1315
  (
    n1974,
    n213
  );


  not
  g1316
  (
    n1309,
    n465
  );


  buf
  g1317
  (
    n1522,
    n519
  );


  not
  g1318
  (
    n1085,
    n381
  );


  buf
  g1319
  (
    n1362,
    n544
  );


  not
  g1320
  (
    n1297,
    n565
  );


  buf
  g1321
  (
    n1780,
    n385
  );


  buf
  g1322
  (
    n1114,
    n366
  );


  buf
  g1323
  (
    n1933,
    n417
  );


  not
  g1324
  (
    n1103,
    n284
  );


  buf
  g1325
  (
    n1025,
    n414
  );


  buf
  g1326
  (
    n942,
    n564
  );


  not
  g1327
  (
    n1213,
    n583
  );


  buf
  g1328
  (
    n1259,
    n285
  );


  buf
  g1329
  (
    n1351,
    n277
  );


  buf
  g1330
  (
    n1087,
    n235
  );


  not
  g1331
  (
    n1968,
    n355
  );


  buf
  g1332
  (
    n857,
    n406
  );


  buf
  g1333
  (
    n1797,
    n588
  );


  not
  g1334
  (
    n885,
    n366
  );


  buf
  g1335
  (
    n1770,
    n365
  );


  buf
  g1336
  (
    n1745,
    n368
  );


  buf
  g1337
  (
    n1577,
    n356
  );


  buf
  g1338
  (
    n1106,
    n426
  );


  not
  g1339
  (
    n1718,
    n416
  );


  not
  g1340
  (
    n1587,
    n438
  );


  not
  g1341
  (
    n1341,
    n478
  );


  not
  g1342
  (
    n1133,
    n650
  );


  buf
  g1343
  (
    KeyWire_0_17,
    n455
  );


  buf
  g1344
  (
    n915,
    n612
  );


  buf
  g1345
  (
    n1169,
    n628
  );


  buf
  g1346
  (
    n1762,
    n240
  );


  not
  g1347
  (
    n1512,
    n336
  );


  buf
  g1348
  (
    n946,
    n209
  );


  not
  g1349
  (
    n982,
    n193
  );


  not
  g1350
  (
    n705,
    n448
  );


  not
  g1351
  (
    n733,
    n405
  );


  buf
  g1352
  (
    KeyWire_0_51,
    n403
  );


  buf
  g1353
  (
    n1148,
    n303
  );


  buf
  g1354
  (
    n1725,
    n330
  );


  buf
  g1355
  (
    n1809,
    n529
  );


  not
  g1356
  (
    n1232,
    n503
  );


  buf
  g1357
  (
    n1348,
    n250
  );


  buf
  g1358
  (
    n1204,
    n360
  );


  not
  g1359
  (
    n1020,
    n606
  );


  not
  g1360
  (
    n1669,
    n567
  );


  not
  g1361
  (
    n1371,
    n466
  );


  buf
  g1362
  (
    n900,
    n595
  );


  buf
  g1363
  (
    n1597,
    n441
  );


  not
  g1364
  (
    n1701,
    n219
  );


  not
  g1365
  (
    n1006,
    n189
  );


  not
  g1366
  (
    n1804,
    n171
  );


  not
  g1367
  (
    n1961,
    n575
  );


  buf
  g1368
  (
    n1691,
    n599
  );


  buf
  g1369
  (
    n967,
    n518
  );


  buf
  g1370
  (
    n1273,
    n442
  );


  not
  g1371
  (
    n1184,
    n447
  );


  buf
  g1372
  (
    n669,
    n509
  );


  not
  g1373
  (
    n1649,
    n632
  );


  buf
  g1374
  (
    n1732,
    n230
  );


  buf
  g1375
  (
    n949,
    n549
  );


  buf
  g1376
  (
    n1518,
    n319
  );


  not
  g1377
  (
    n1289,
    n606
  );


  buf
  g1378
  (
    n1090,
    n312
  );


  not
  g1379
  (
    n1033,
    n275
  );


  not
  g1380
  (
    n743,
    n215
  );


  buf
  g1381
  (
    n721,
    n444
  );


  not
  g1382
  (
    n1080,
    n343
  );


  buf
  g1383
  (
    n1282,
    n256
  );


  buf
  g1384
  (
    n1939,
    n375
  );


  not
  g1385
  (
    n1079,
    n484
  );


  buf
  g1386
  (
    n1208,
    n355
  );


  buf
  g1387
  (
    n1553,
    n281
  );


  buf
  g1388
  (
    n988,
    n447
  );


  not
  g1389
  (
    n736,
    n163
  );


  not
  g1390
  (
    n922,
    n174
  );


  buf
  g1391
  (
    n1665,
    n195
  );


  not
  g1392
  (
    n1711,
    n376
  );


  not
  g1393
  (
    n2059,
    n645
  );


  buf
  g1394
  (
    n1666,
    n333
  );


  not
  g1395
  (
    n1381,
    n434
  );


  buf
  g1396
  (
    n2031,
    n299
  );


  not
  g1397
  (
    n934,
    n339
  );


  buf
  g1398
  (
    n875,
    n617
  );


  buf
  g1399
  (
    n1841,
    n623
  );


  buf
  g1400
  (
    n1360,
    n249
  );


  buf
  g1401
  (
    n1982,
    n444
  );


  not
  g1402
  (
    n1927,
    n544
  );


  not
  g1403
  (
    n1327,
    n164
  );


  buf
  g1404
  (
    n937,
    n547
  );


  not
  g1405
  (
    n1706,
    n208
  );


  not
  g1406
  (
    n970,
    n372
  );


  not
  g1407
  (
    n1752,
    n387
  );


  buf
  g1408
  (
    n1744,
    n488
  );


  buf
  g1409
  (
    n1415,
    n393
  );


  buf
  g1410
  (
    n1899,
    n286
  );


  not
  g1411
  (
    n1216,
    n197
  );


  not
  g1412
  (
    n1542,
    n519
  );


  not
  g1413
  (
    n1624,
    n633
  );


  not
  g1414
  (
    n1729,
    n435
  );


  not
  g1415
  (
    n716,
    n245
  );


  not
  g1416
  (
    n853,
    n650
  );


  buf
  g1417
  (
    n1800,
    n400
  );


  buf
  g1418
  (
    n1076,
    n173
  );


  buf
  g1419
  (
    n1122,
    n492
  );


  not
  g1420
  (
    n1859,
    n207
  );


  not
  g1421
  (
    n1007,
    n558
  );


  not
  g1422
  (
    n1040,
    n169
  );


  not
  g1423
  (
    n772,
    n454
  );


  not
  g1424
  (
    n1128,
    n264
  );


  not
  g1425
  (
    n1642,
    n362
  );


  not
  g1426
  (
    n1924,
    n296
  );


  buf
  g1427
  (
    n1375,
    n439
  );


  not
  g1428
  (
    n1393,
    n340
  );


  buf
  g1429
  (
    n892,
    n330
  );


  not
  g1430
  (
    n962,
    n597
  );


  not
  g1431
  (
    n1061,
    n321
  );


  buf
  g1432
  (
    KeyWire_0_61,
    n459
  );


  not
  g1433
  (
    n2010,
    n598
  );


  buf
  g1434
  (
    n1264,
    n350
  );


  buf
  g1435
  (
    n1139,
    n432
  );


  buf
  g1436
  (
    n1557,
    n236
  );


  buf
  g1437
  (
    n1923,
    n352
  );


  buf
  g1438
  (
    n1515,
    n616
  );


  buf
  g1439
  (
    n1904,
    n210
  );


  buf
  g1440
  (
    n871,
    n237
  );


  buf
  g1441
  (
    n2021,
    n637
  );


  not
  g1442
  (
    n864,
    n211
  );


  not
  g1443
  (
    n695,
    n384
  );


  not
  g1444
  (
    n1320,
    n387
  );


  buf
  g1445
  (
    n948,
    n250
  );


  not
  g1446
  (
    n1712,
    n500
  );


  not
  g1447
  (
    n800,
    n334
  );


  not
  g1448
  (
    n1514,
    n652
  );


  buf
  g1449
  (
    n1486,
    n407
  );


  not
  g1450
  (
    n828,
    n235
  );


  not
  g1451
  (
    n678,
    n396
  );


  not
  g1452
  (
    n851,
    n327
  );


  not
  g1453
  (
    n1836,
    n411
  );


  not
  g1454
  (
    n1125,
    n242
  );


  not
  g1455
  (
    n1833,
    n415
  );


  not
  g1456
  (
    n1787,
    n469
  );


  buf
  g1457
  (
    n1799,
    n533
  );


  not
  g1458
  (
    n1877,
    n468
  );


  buf
  g1459
  (
    n1477,
    n506
  );


  buf
  g1460
  (
    n926,
    n244
  );


  not
  g1461
  (
    n742,
    n204
  );


  not
  g1462
  (
    n1026,
    n640
  );


  buf
  g1463
  (
    n799,
    n353
  );


  buf
  g1464
  (
    n1313,
    n648
  );


  buf
  g1465
  (
    n2006,
    n226
  );


  buf
  g1466
  (
    n1274,
    n456
  );


  not
  g1467
  (
    n1095,
    n627
  );


  buf
  g1468
  (
    n1808,
    n216
  );


  buf
  g1469
  (
    n1985,
    n352
  );


  buf
  g1470
  (
    n1567,
    n436
  );


  not
  g1471
  (
    n846,
    n651
  );


  buf
  g1472
  (
    n1710,
    n406
  );


  buf
  g1473
  (
    n1733,
    n501
  );


  buf
  g1474
  (
    n954,
    n375
  );


  buf
  g1475
  (
    n2007,
    n436
  );


  not
  g1476
  (
    n1015,
    n217
  );


  buf
  g1477
  (
    n813,
    n353
  );


  buf
  g1478
  (
    n1005,
    n537
  );


  not
  g1479
  (
    n1544,
    n213
  );


  buf
  g1480
  (
    n1987,
    n340
  );


  not
  g1481
  (
    n1829,
    n619
  );


  not
  g1482
  (
    n1434,
    n230
  );


  not
  g1483
  (
    n1792,
    n349
  );


  not
  g1484
  (
    n862,
    n283
  );


  not
  g1485
  (
    n1788,
    n292
  );


  buf
  g1486
  (
    n1611,
    n529
  );


  not
  g1487
  (
    n1658,
    n537
  );


  not
  g1488
  (
    n1615,
    n399
  );


  buf
  g1489
  (
    n1505,
    n502
  );


  not
  g1490
  (
    n1031,
    n183
  );


  not
  g1491
  (
    n719,
    n359
  );


  not
  g1492
  (
    n1418,
    n263
  );


  buf
  g1493
  (
    n1302,
    n635
  );


  buf
  g1494
  (
    n1868,
    n431
  );


  buf
  g1495
  (
    n910,
    n168
  );


  not
  g1496
  (
    n1442,
    n651
  );


  buf
  g1497
  (
    n1812,
    n224
  );


  not
  g1498
  (
    n1242,
    n473
  );


  not
  g1499
  (
    n749,
    n450
  );


  buf
  g1500
  (
    n1054,
    n548
  );


  not
  g1501
  (
    n1990,
    n390
  );


  not
  g1502
  (
    n1495,
    n270
  );


  buf
  g1503
  (
    n1802,
    n651
  );


  not
  g1504
  (
    n974,
    n472
  );


  not
  g1505
  (
    n1714,
    n429
  );


  not
  g1506
  (
    n876,
    n368
  );


  buf
  g1507
  (
    n916,
    n462
  );


  buf
  g1508
  (
    n1592,
    n386
  );


  buf
  g1509
  (
    n1610,
    n182
  );


  not
  g1510
  (
    n1675,
    n220
  );


  not
  g1511
  (
    n823,
    n195
  );


  not
  g1512
  (
    n1724,
    n501
  );


  buf
  g1513
  (
    n760,
    n218
  );


  buf
  g1514
  (
    KeyWire_0_24,
    n196
  );


  not
  g1515
  (
    n784,
    n550
  );


  not
  g1516
  (
    n1134,
    n224
  );


  buf
  g1517
  (
    n1991,
    n164
  );


  buf
  g1518
  (
    n1269,
    n201
  );


  buf
  g1519
  (
    n981,
    n542
  );


  buf
  g1520
  (
    n918,
    n205
  );


  not
  g1521
  (
    n1253,
    n497
  );


  not
  g1522
  (
    n1957,
    n436
  );


  buf
  g1523
  (
    n953,
    n227
  );


  not
  g1524
  (
    n2015,
    n525
  );


  buf
  g1525
  (
    n786,
    n627
  );


  buf
  g1526
  (
    n1292,
    n325
  );


  not
  g1527
  (
    n2036,
    n210
  );


  buf
  g1528
  (
    n1959,
    n652
  );


  not
  g1529
  (
    n839,
    n555
  );


  not
  g1530
  (
    n726,
    n607
  );


  buf
  g1531
  (
    n1880,
    n269
  );


  not
  g1532
  (
    n1343,
    n172
  );


  not
  g1533
  (
    n1425,
    n551
  );


  not
  g1534
  (
    n1564,
    n475
  );


  buf
  g1535
  (
    n878,
    n322
  );


  not
  g1536
  (
    n1332,
    n167
  );


  buf
  g1537
  (
    n1479,
    n401
  );


  buf
  g1538
  (
    n1700,
    n646
  );


  not
  g1539
  (
    n1854,
    n493
  );


  not
  g1540
  (
    n2065,
    n479
  );


  not
  g1541
  (
    n985,
    n271
  );


  not
  g1542
  (
    n1875,
    n271
  );


  buf
  g1543
  (
    n996,
    n337
  );


  buf
  g1544
  (
    n1333,
    n543
  );


  not
  g1545
  (
    n1064,
    n443
  );


  not
  g1546
  (
    n1436,
    n188
  );


  not
  g1547
  (
    n1771,
    n331
  );


  buf
  g1548
  (
    n1291,
    n253
  );


  buf
  g1549
  (
    n1323,
    n527
  );


  buf
  g1550
  (
    n1932,
    n195
  );


  buf
  g1551
  (
    n1835,
    n621
  );


  buf
  g1552
  (
    n1111,
    n411
  );


  buf
  g1553
  (
    n2013,
    n299
  );


  buf
  g1554
  (
    n856,
    n502
  );


  not
  g1555
  (
    n1207,
    n533
  );


  buf
  g1556
  (
    n697,
    n450
  );


  buf
  g1557
  (
    n2019,
    n196
  );


  not
  g1558
  (
    n1858,
    n510
  );


  not
  g1559
  (
    n1328,
    n530
  );


  buf
  g1560
  (
    n914,
    n411
  );


  not
  g1561
  (
    n1672,
    n418
  );


  buf
  g1562
  (
    n832,
    n324
  );


  buf
  g1563
  (
    n755,
    n473
  );


  not
  g1564
  (
    n958,
    n489
  );


  not
  g1565
  (
    n1400,
    n193
  );


  buf
  g1566
  (
    n2025,
    n272
  );


  buf
  g1567
  (
    n1757,
    n237
  );


  not
  g1568
  (
    n1679,
    n433
  );


  not
  g1569
  (
    n1878,
    n542
  );


  not
  g1570
  (
    n1917,
    n321
  );


  not
  g1571
  (
    n1621,
    n433
  );


  not
  g1572
  (
    n754,
    n234
  );


  not
  g1573
  (
    n1824,
    n459
  );


  buf
  g1574
  (
    n1082,
    n556
  );


  not
  g1575
  (
    n2038,
    n422
  );


  buf
  g1576
  (
    n912,
    n252
  );


  buf
  g1577
  (
    n1958,
    n315
  );


  not
  g1578
  (
    n680,
    n243
  );


  not
  g1579
  (
    n817,
    n475
  );


  not
  g1580
  (
    n1647,
    n442
  );


  buf
  g1581
  (
    n1598,
    n600
  );


  not
  g1582
  (
    n1118,
    n504
  );


  buf
  g1583
  (
    n905,
    n580
  );


  not
  g1584
  (
    n746,
    n506
  );


  buf
  g1585
  (
    n1556,
    n438
  );


  not
  g1586
  (
    n1901,
    n332
  );


  buf
  g1587
  (
    n1077,
    n258
  );


  not
  g1588
  (
    n1444,
    n280
  );


  buf
  g1589
  (
    n1217,
    n327
  );


  buf
  g1590
  (
    n1198,
    n472
  );


  buf
  g1591
  (
    n795,
    n486
  );


  buf
  g1592
  (
    n1879,
    n282
  );


  buf
  g1593
  (
    n1500,
    n398
  );


  buf
  g1594
  (
    n1967,
    n323
  );


  not
  g1595
  (
    n1000,
    n176
  );


  not
  g1596
  (
    n1127,
    n654
  );


  buf
  g1597
  (
    n1865,
    n407
  );


  buf
  g1598
  (
    n1201,
    n551
  );


  buf
  g1599
  (
    n1509,
    n169
  );


  buf
  g1600
  (
    n1524,
    n450
  );


  buf
  g1601
  (
    KeyWire_0_33,
    n275
  );


  buf
  g1602
  (
    n1265,
    n259
  );


  buf
  g1603
  (
    n1382,
    n361
  );


  buf
  g1604
  (
    KeyWire_0_36,
    n279
  );


  buf
  g1605
  (
    n1211,
    n208
  );


  buf
  g1606
  (
    n1288,
    n649
  );


  buf
  g1607
  (
    n1278,
    n298
  );


  not
  g1608
  (
    n1308,
    n535
  );


  buf
  g1609
  (
    n1374,
    n248
  );


  buf
  g1610
  (
    n1898,
    n319
  );


  buf
  g1611
  (
    n995,
    n596
  );


  buf
  g1612
  (
    KeyWire_0_56,
    n219
  );


  not
  g1613
  (
    KeyWire_0_27,
    n250
  );


  not
  g1614
  (
    n1663,
    n238
  );


  buf
  g1615
  (
    n865,
    n598
  );


  not
  g1616
  (
    n1018,
    n161
  );


  buf
  g1617
  (
    n1630,
    n212
  );


  buf
  g1618
  (
    n1150,
    n233
  );


  buf
  g1619
  (
    n1884,
    n170
  );


  buf
  g1620
  (
    n1042,
    n275
  );


  not
  g1621
  (
    n1617,
    n238
  );


  buf
  g1622
  (
    n1098,
    n208
  );


  not
  g1623
  (
    n1387,
    n162
  );


  buf
  g1624
  (
    n1013,
    n168
  );


  not
  g1625
  (
    n1738,
    n565
  );


  buf
  g1626
  (
    n1915,
    n330
  );


  not
  g1627
  (
    n707,
    n563
  );


  buf
  g1628
  (
    n1021,
    n440
  );


  not
  g1629
  (
    n699,
    n233
  );


  not
  g1630
  (
    n1067,
    n279
  );


  not
  g1631
  (
    n2042,
    n213
  );


  buf
  g1632
  (
    n2058,
    n362
  );


  not
  g1633
  (
    n1682,
    n456
  );


  buf
  g1634
  (
    n1713,
    n557
  );


  not
  g1635
  (
    n1684,
    n613
  );


  not
  g1636
  (
    n902,
    n635
  );


  buf
  g1637
  (
    n1335,
    n307
  );


  buf
  g1638
  (
    n1943,
    n488
  );


  not
  g1639
  (
    n1793,
    n368
  );


  buf
  g1640
  (
    n781,
    n181
  );


  buf
  g1641
  (
    n1847,
    n177
  );


  buf
  g1642
  (
    n1249,
    n523
  );


  buf
  g1643
  (
    n1088,
    n335
  );


  buf
  g1644
  (
    n1158,
    n360
  );


  not
  g1645
  (
    n1743,
    n283
  );


  not
  g1646
  (
    n1980,
    n453
  );


  not
  g1647
  (
    n1969,
    n305
  );


  not
  g1648
  (
    n1162,
    n493
  );


  not
  g1649
  (
    n1299,
    n239
  );


  not
  g1650
  (
    n1819,
    n453
  );


  buf
  g1651
  (
    n735,
    n240
  );


  not
  g1652
  (
    n1863,
    n267
  );


  not
  g1653
  (
    n1573,
    n292
  );


  not
  g1654
  (
    n1638,
    n505
  );


  buf
  g1655
  (
    n1151,
    n486
  );


  buf
  g1656
  (
    n1430,
    n590
  );


  not
  g1657
  (
    n803,
    n199
  );


  buf
  g1658
  (
    n1607,
    n314
  );


  buf
  g1659
  (
    n1441,
    n625
  );


  buf
  g1660
  (
    n1998,
    n448
  );


  buf
  g1661
  (
    KeyWire_0_9,
    n313
  );


  buf
  g1662
  (
    n1813,
    n462
  );


  not
  g1663
  (
    n1547,
    n524
  );


  not
  g1664
  (
    n1857,
    n577
  );


  buf
  g1665
  (
    n674,
    n370
  );


  buf
  g1666
  (
    n1255,
    n298
  );


  buf
  g1667
  (
    n1240,
    n619
  );


  buf
  g1668
  (
    n1231,
    n289
  );


  buf
  g1669
  (
    n2063,
    n418
  );


  buf
  g1670
  (
    n1096,
    n517
  );


  not
  g1671
  (
    n1215,
    n400
  );


  buf
  g1672
  (
    n778,
    n604
  );


  not
  g1673
  (
    n1590,
    n540
  );


  buf
  g1674
  (
    n1785,
    n269
  );


  buf
  g1675
  (
    n2051,
    n655
  );


  not
  g1676
  (
    n1396,
    n386
  );


  buf
  g1677
  (
    n1110,
    n258
  );


  not
  g1678
  (
    n1142,
    n227
  );


  not
  g1679
  (
    n1109,
    n512
  );


  not
  g1680
  (
    n1056,
    n260
  );


  not
  g1681
  (
    n1093,
    n346
  );


  not
  g1682
  (
    n1414,
    n591
  );


  buf
  g1683
  (
    n973,
    n285
  );


  buf
  g1684
  (
    n1604,
    n438
  );


  not
  g1685
  (
    n1053,
    n539
  );


  buf
  g1686
  (
    n1526,
    n452
  );


  not
  g1687
  (
    n690,
    n307
  );


  buf
  g1688
  (
    n1754,
    n516
  );


  buf
  g1689
  (
    n1903,
    n554
  );


  buf
  g1690
  (
    n1314,
    n554
  );


  not
  g1691
  (
    n1369,
    n639
  );


  buf
  g1692
  (
    n1997,
    n295
  );


  not
  g1693
  (
    n1988,
    n280
  );


  not
  g1694
  (
    n1973,
    n504
  );


  buf
  g1695
  (
    n1758,
    n622
  );


  not
  g1696
  (
    n1226,
    n471
  );


  not
  g1697
  (
    n1685,
    n403
  );


  buf
  g1698
  (
    n1862,
    n326
  );


  buf
  g1699
  (
    n887,
    n627
  );


  buf
  g1700
  (
    n837,
    n342
  );


  not
  g1701
  (
    n770,
    n253
  );


  not
  g1702
  (
    n935,
    n322
  );


  not
  g1703
  (
    n1872,
    n215
  );


  not
  g1704
  (
    n1532,
    n603
  );


  buf
  g1705
  (
    n1303,
    n613
  );


  buf
  g1706
  (
    n1689,
    n518
  );


  not
  g1707
  (
    n1074,
    n259
  );


  buf
  g1708
  (
    n1748,
    n418
  );


  not
  g1709
  (
    KeyWire_0_15,
    n264
  );


  buf
  g1710
  (
    n1161,
    n564
  );


  not
  g1711
  (
    n1266,
    n567
  );


  buf
  g1712
  (
    n809,
    n546
  );


  not
  g1713
  (
    n1256,
    n389
  );


  buf
  g1714
  (
    n1417,
    n251
  );


  buf
  g1715
  (
    n1322,
    n655
  );


  not
  g1716
  (
    n1853,
    n477
  );


  not
  g1717
  (
    n1972,
    n354
  );


  not
  g1718
  (
    n1342,
    n541
  );


  buf
  g1719
  (
    n1181,
    n168
  );


  not
  g1720
  (
    n1113,
    n572
  );


  buf
  g1721
  (
    n816,
    n465
  );


  buf
  g1722
  (
    n1650,
    n397
  );


  buf
  g1723
  (
    n1981,
    n255
  );


  not
  g1724
  (
    n1069,
    n278
  );


  buf
  g1725
  (
    n1011,
    n255
  );


  not
  g1726
  (
    n1132,
    n585
  );


  not
  g1727
  (
    n734,
    n280
  );


  buf
  g1728
  (
    n1227,
    n616
  );


  buf
  g1729
  (
    n1497,
    n312
  );


  not
  g1730
  (
    n1368,
    n411
  );


  buf
  g1731
  (
    n739,
    n498
  );


  not
  g1732
  (
    n676,
    n534
  );


  buf
  g1733
  (
    n1528,
    n300
  );


  not
  g1734
  (
    n1586,
    n528
  );


  buf
  g1735
  (
    n1722,
    n531
  );


  not
  g1736
  (
    KeyWire_0_40,
    n560
  );


  buf
  g1737
  (
    n1992,
    n618
  );


  buf
  g1738
  (
    n1177,
    n274
  );


  buf
  g1739
  (
    n682,
    n633
  );


  buf
  g1740
  (
    n1179,
    n382
  );


  not
  g1741
  (
    n1066,
    n655
  );


  not
  g1742
  (
    n1458,
    n494
  );


  not
  g1743
  (
    n897,
    n590
  );


  buf
  g1744
  (
    n2028,
    n532
  );


  buf
  g1745
  (
    n1949,
    n566
  );


  not
  g1746
  (
    n1338,
    n217
  );


  not
  g1747
  (
    n1960,
    n574
  );


  buf
  g1748
  (
    n1210,
    n260
  );


  buf
  g1749
  (
    n1180,
    n435
  );


  buf
  g1750
  (
    n1895,
    n523
  );


  buf
  g1751
  (
    n1156,
    n525
  );


  not
  g1752
  (
    n1409,
    n571
  );


  not
  g1753
  (
    n1468,
    n467
  );


  not
  g1754
  (
    n1807,
    n522
  );


  not
  g1755
  (
    n1419,
    n198
  );


  not
  g1756
  (
    n741,
    n287
  );


  not
  g1757
  (
    n1839,
    n460
  );


  buf
  g1758
  (
    n757,
    n245
  );


  not
  g1759
  (
    n1774,
    n521
  );


  not
  g1760
  (
    n1643,
    n278
  );


  buf
  g1761
  (
    n1317,
    n415
  );


  not
  g1762
  (
    n1024,
    n495
  );


  buf
  g1763
  (
    n1172,
    n353
  );


  buf
  g1764
  (
    n879,
    n440
  );


  buf
  g1765
  (
    n1367,
    n396
  );


  not
  g1766
  (
    n1386,
    n338
  );


  buf
  g1767
  (
    n1888,
    n261
  );


  buf
  g1768
  (
    n1832,
    n421
  );


  not
  g1769
  (
    n1470,
    n308
  );


  not
  g1770
  (
    n1842,
    n189
  );


  buf
  g1771
  (
    n1821,
    n170
  );


  buf
  g1772
  (
    n1124,
    n449
  );


  buf
  g1773
  (
    n761,
    n592
  );


  not
  g1774
  (
    n1594,
    n325
  );


  buf
  g1775
  (
    n1735,
    n395
  );


  buf
  g1776
  (
    n1075,
    n177
  );


  buf
  g1777
  (
    n1517,
    n547
  );


  buf
  g1778
  (
    n991,
    n607
  );


  not
  g1779
  (
    n1503,
    n343
  );


  buf
  g1780
  (
    n780,
    n455
  );


  buf
  g1781
  (
    n955,
    n605
  );


  not
  g1782
  (
    n886,
    n495
  );


  not
  g1783
  (
    KeyWire_0_49,
    n482
  );


  buf
  g1784
  (
    n963,
    n433
  );


  buf
  g1785
  (
    n972,
    n523
  );


  not
  g1786
  (
    n1575,
    n460
  );


  not
  g1787
  (
    n1717,
    n269
  );


  buf
  g1788
  (
    n765,
    n361
  );


  buf
  g1789
  (
    n1696,
    n345
  );


  not
  g1790
  (
    n1234,
    n342
  );


  buf
  g1791
  (
    n802,
    n357
  );


  not
  g1792
  (
    n2027,
    n268
  );


  buf
  g1793
  (
    n1410,
    n333
  );


  not
  g1794
  (
    n729,
    n301
  );


  buf
  g1795
  (
    n965,
    n632
  );


  buf
  g1796
  (
    n1716,
    n383
  );


  not
  g1797
  (
    n1921,
    n455
  );


  buf
  g1798
  (
    n896,
    n584
  );


  buf
  g1799
  (
    n801,
    n196
  );


  not
  g1800
  (
    n1882,
    n464
  );


  buf
  g1801
  (
    n787,
    n534
  );


  not
  g1802
  (
    n1527,
    n372
  );


  not
  g1803
  (
    n939,
    n552
  );


  buf
  g1804
  (
    n1704,
    n637
  );


  not
  g1805
  (
    n1094,
    n192
  );


  buf
  g1806
  (
    n831,
    n347
  );


  not
  g1807
  (
    n1228,
    n366
  );


  not
  g1808
  (
    n2024,
    n286
  );


  buf
  g1809
  (
    n1560,
    n570
  );


  not
  g1810
  (
    n2009,
    n521
  );


  not
  g1811
  (
    n1983,
    n192
  );


  buf
  g1812
  (
    n941,
    n591
  );


  not
  g1813
  (
    n854,
    n337
  );


  not
  g1814
  (
    n1776,
    n252
  );


  buf
  g1815
  (
    n1719,
    n443
  );


  buf
  g1816
  (
    n1845,
    n163
  );


  not
  g1817
  (
    n763,
    n163
  );


  not
  g1818
  (
    n1455,
    n179
  );


  not
  g1819
  (
    n1203,
    n311
  );


  buf
  g1820
  (
    KeyWire_0_32,
    n230
  );


  buf
  g1821
  (
    n2046,
    n363
  );


  not
  g1822
  (
    n2001,
    n498
  );


  not
  g1823
  (
    n1340,
    n247
  );


  not
  g1824
  (
    n790,
    n175
  );


  buf
  g1825
  (
    n1280,
    n253
  );


  not
  g1826
  (
    n1755,
    n391
  );


  buf
  g1827
  (
    n1099,
    n524
  );


  not
  g1828
  (
    n1236,
    n329
  );


  not
  g1829
  (
    n1209,
    n470
  );


  not
  g1830
  (
    n1421,
    n412
  );


  buf
  g1831
  (
    n895,
    n611
  );


  not
  g1832
  (
    n1768,
    n621
  );


  buf
  g1833
  (
    n1137,
    n429
  );


  buf
  g1834
  (
    n901,
    n181
  );


  buf
  g1835
  (
    n1635,
    n565
  );


  buf
  g1836
  (
    n747,
    n414
  );


  not
  g1837
  (
    n980,
    n325
  );


  not
  g1838
  (
    n1627,
    n576
  );


  xnor
  g1839
  (
    n1766,
    n222,
    n169,
    n509,
    n617
  );


  nand
  g1840
  (
    n710,
    n279,
    n538,
    n174,
    n537
  );


  nor
  g1841
  (
    n683,
    n471,
    n190,
    n355,
    n385
  );


  or
  g1842
  (
    n1290,
    n613,
    n459,
    n320,
    n489
  );


  xnor
  g1843
  (
    n1420,
    n568,
    n282,
    n376,
    n561
  );


  xor
  g1844
  (
    n1664,
    n323,
    n634,
    n446,
    n169
  );


  nand
  g1845
  (
    n685,
    n319,
    n295,
    n538,
    n289
  );


  or
  g1846
  (
    n714,
    n243,
    n657,
    n199,
    n405
  );


  nand
  g1847
  (
    n898,
    n299,
    n420,
    n336,
    n587
  );


  xnor
  g1848
  (
    n1390,
    n350,
    n480,
    n380
  );


  nor
  g1849
  (
    n1971,
    n371,
    n289,
    n251,
    n267
  );


  xnor
  g1850
  (
    n992,
    n345,
    n531,
    n167,
    n496
  );


  nand
  g1851
  (
    n1815,
    n174,
    n388,
    n198,
    n231
  );


  or
  g1852
  (
    n834,
    n186,
    n214,
    n308,
    n618
  );


  xnor
  g1853
  (
    n1595,
    n329,
    n389,
    n284,
    n545
  );


  xnor
  g1854
  (
    n1926,
    n371,
    n643,
    n594,
    n328
  );


  xnor
  g1855
  (
    n704,
    n420,
    n556,
    n510,
    n178
  );


  xnor
  g1856
  (
    n956,
    n378,
    n393,
    n625,
    n471
  );


  xnor
  g1857
  (
    n2068,
    n571,
    n410,
    n641,
    n240
  );


  or
  g1858
  (
    n1645,
    n344,
    n619,
    n280,
    n508
  );


  or
  g1859
  (
    n1614,
    n598,
    n245,
    n221,
    n307
  );


  nor
  g1860
  (
    n2020,
    n293,
    n487,
    n331
  );


  nor
  g1861
  (
    n1529,
    n337,
    n200,
    n297,
    n452
  );


  nor
  g1862
  (
    n1427,
    n185,
    n402,
    n599,
    n591
  );


  xor
  g1863
  (
    n1378,
    n496,
    n281,
    n179,
    n216
  );


  nand
  g1864
  (
    n1206,
    n647,
    n369,
    n653,
    n416
  );


  xnor
  g1865
  (
    n711,
    n576,
    n595,
    n605,
    n408
  );


  xor
  g1866
  (
    n1456,
    n331,
    n570,
    n614,
    n563
  );


  nor
  g1867
  (
    n1214,
    n586,
    n179,
    n599,
    n639
  );


  nand
  g1868
  (
    n964,
    n632,
    n469,
    n629,
    n414
  );


  xor
  g1869
  (
    n1331,
    n644,
    n397,
    n594,
    n263
  );


  nand
  g1870
  (
    n1449,
    n316,
    n478,
    n449,
    n262
  );


  xnor
  g1871
  (
    n1447,
    n625,
    n575,
    n637,
    n332
  );


  xnor
  g1872
  (
    n929,
    n239,
    n368,
    n447,
    n203
  );


  nand
  g1873
  (
    n978,
    n267,
    n341,
    n540,
    n186
  );


  nand
  g1874
  (
    n1263,
    n346,
    n377,
    n583,
    n398
  );


  or
  g1875
  (
    n675,
    n208,
    n301,
    n382,
    n632
  );


  or
  g1876
  (
    n732,
    n199,
    n434,
    n284,
    n255
  );


  xor
  g1877
  (
    n843,
    n649,
    n376,
    n374,
    n281
  );


  xor
  g1878
  (
    n1286,
    n419,
    n346,
    n498,
    n503
  );


  xnor
  g1879
  (
    n943,
    n526,
    n191,
    n265,
    n451
  );


  xor
  g1880
  (
    n1305,
    n239,
    n312,
    n597,
    n515
  );


  nor
  g1881
  (
    n1281,
    n297,
    n161,
    n446,
    n421
  );


  and
  g1882
  (
    n788,
    n203,
    n166,
    n195,
    n638
  );


  nand
  g1883
  (
    n1205,
    n564,
    n526,
    n461,
    n489
  );


  nand
  g1884
  (
    n715,
    n213,
    n334,
    n339,
    n206
  );


  nor
  g1885
  (
    n1050,
    n227,
    n388,
    n373,
    n383
  );


  and
  g1886
  (
    n713,
    n548,
    n493,
    n349,
    n226
  );


  nand
  g1887
  (
    n1475,
    n658,
    n360,
    n335,
    n568
  );


  nand
  g1888
  (
    n1856,
    n395,
    n657,
    n514,
    n300
  );


  nor
  g1889
  (
    n1601,
    n271,
    n523,
    n600,
    n474
  );


  xor
  g1890
  (
    n769,
    n305,
    n187,
    n655,
    n469
  );


  and
  g1891
  (
    n1861,
    n187,
    n450,
    n417,
    n220
  );


  or
  g1892
  (
    n718,
    n387,
    n443,
    n413,
    n509
  );


  and
  g1893
  (
    n1935,
    n410,
    n173,
    n457,
    n589
  );


  or
  g1894
  (
    n1534,
    n366,
    n206,
    n406,
    n223
  );


  nand
  g1895
  (
    n1995,
    n458,
    n568,
    n334,
    n417
  );


  xor
  g1896
  (
    n1674,
    n404,
    n183,
    n508,
    n185
  );


  nor
  g1897
  (
    n1984,
    n586,
    n563,
    n508,
    n492
  );


  or
  g1898
  (
    n1570,
    n176,
    n602,
    n437,
    n537
  );


  nand
  g1899
  (
    n1272,
    n623,
    n505,
    n294,
    n296
  );


  and
  g1900
  (
    n1359,
    n236,
    n560,
    n277,
    n247
  );


  and
  g1901
  (
    n836,
    n265,
    n405,
    n290,
    n277
  );


  xor
  g1902
  (
    n1763,
    n306,
    n272,
    n499,
    n336
  );


  and
  g1903
  (
    n1741,
    n407,
    n435,
    n539,
    n504
  );


  nor
  g1904
  (
    n2054,
    n351,
    n656,
    n607,
    n291
  );


  xnor
  g1905
  (
    n880,
    n235,
    n424,
    n203,
    n640
  );


  xnor
  g1906
  (
    n1364,
    n309,
    n379,
    n418,
    n165
  );


  nand
  g1907
  (
    n1339,
    n521,
    n466,
    n350,
    n510
  );


  nand
  g1908
  (
    n1057,
    n345,
    n289,
    n428,
    n275
  );


  xor
  g1909
  (
    n819,
    n378,
    n190,
    n551,
    n566
  );


  nand
  g1910
  (
    n1354,
    n354,
    n630,
    n391,
    n338
  );


  nor
  g1911
  (
    n899,
    n268,
    n371,
    n612,
    n204
  );


  xnor
  g1912
  (
    n2032,
    n524,
    n288,
    n501,
    n449
  );


  xor
  g1913
  (
    n1048,
    n557,
    n638,
    n344,
    n328
  );


  or
  g1914
  (
    n774,
    n461,
    n248,
    n453,
    n614
  );


  xor
  g1915
  (
    n841,
    n301,
    n384,
    n430,
    n380
  );


  and
  g1916
  (
    n1261,
    n481,
    n217,
    n412,
    n484
  );


  or
  g1917
  (
    n844,
    n542,
    n260,
    n210,
    n220
  );


  xor
  g1918
  (
    n1052,
    n205,
    n456,
    n250,
    n546
  );


  nor
  g1919
  (
    n1153,
    n415,
    n351,
    n433,
    n628
  );


  nand
  g1920
  (
    n1036,
    n202,
    n188,
    n488,
    n379
  );


  nand
  g1921
  (
    n1478,
    n448,
    n563,
    n403,
    n603
  );


  nor
  g1922
  (
    n1315,
    n409,
    n312,
    n317,
    n609
  );


  or
  g1923
  (
    n798,
    n500,
    n175,
    n651,
    n406
  );


  xnor
  g1924
  (
    n1002,
    n394,
    n642,
    n191,
    n258
  );


  and
  g1925
  (
    n782,
    n360,
    n553,
    n316,
    n252
  );


  or
  g1926
  (
    n1220,
    n241,
    n408,
    n359,
    n601
  );


  nand
  g1927
  (
    n1989,
    n596,
    n184,
    n183,
    n557
  );


  nand
  g1928
  (
    n1188,
    n374,
    n359,
    n313,
    n636
  );


  or
  g1929
  (
    n677,
    n540,
    n392,
    n602,
    n536
  );


  nor
  g1930
  (
    n952,
    n268,
    n173,
    n511,
    n371
  );


  xor
  g1931
  (
    n2035,
    n386,
    n171,
    n556,
    n446
  );


  xor
  g1932
  (
    n847,
    n601,
    n232,
    n307,
    n414
  );


  nor
  g1933
  (
    n1654,
    n370,
    n452,
    n209,
    n272
  );


  or
  g1934
  (
    n1769,
    n336,
    n219,
    n205,
    n188
  );


  and
  g1935
  (
    n1965,
    n589,
    n306,
    n337,
    n562
  );


  nand
  g1936
  (
    n1296,
    n614,
    n234,
    n445,
    n292
  );


  or
  g1937
  (
    n1029,
    n378,
    n316,
    n428,
    n548
  );


  or
  g1938
  (
    n1818,
    n608,
    n369,
    n646,
    n282
  );


  and
  g1939
  (
    n1937,
    n190,
    n481,
    n212,
    n457
  );


  nor
  g1940
  (
    n810,
    n466,
    n338,
    n187,
    n259
  );


  and
  g1941
  (
    n1329,
    n180,
    n365,
    n335,
    n375
  );


  nor
  g1942
  (
    n1012,
    n467,
    n650,
    n380,
    n474
  );


  xor
  g1943
  (
    n1115,
    n166,
    n264,
    n646,
    n270
  );


  xor
  g1944
  (
    n1485,
    n658,
    n540,
    n321,
    n579
  );


  and
  g1945
  (
    n794,
    n601,
    n641,
    n618,
    n373
  );


  xnor
  g1946
  (
    n1186,
    n320,
    n317,
    n478,
    n358
  );


  xor
  g1947
  (
    n759,
    n470,
    n182,
    n325,
    n522
  );


  or
  g1948
  (
    n1740,
    n399,
    n376,
    n459,
    n241
  );


  or
  g1949
  (
    n1091,
    n535,
    n409,
    n327,
    n451
  );


  or
  g1950
  (
    n1403,
    n395,
    n298,
    n356,
    n652
  );


  xnor
  g1951
  (
    n1197,
    n650,
    n419,
    n226,
    n581
  );


  xor
  g1952
  (
    n775,
    n533,
    n372,
    n626,
    n444
  );


  xnor
  g1953
  (
    KeyWire_0_41,
    n494,
    n465,
    n482,
    n377
  );


  xnor
  g1954
  (
    n1494,
    n207,
    n590,
    n228,
    n586
  );


  xor
  g1955
  (
    n1009,
    n589,
    n606,
    n246,
    n594
  );


  nor
  g1956
  (
    n1411,
    n391,
    n577,
    n209,
    n521
  );


  xnor
  g1957
  (
    n1826,
    n430,
    n439,
    n372,
    n175
  );


  xor
  g1958
  (
    n1030,
    n323,
    n574,
    n482,
    n256
  );


  nand
  g1959
  (
    n1136,
    n349,
    n392,
    n503,
    n583
  );


  xor
  g1960
  (
    n1849,
    n388,
    n460,
    n461,
    n413
  );


  xor
  g1961
  (
    n1677,
    n648,
    n313,
    n514,
    n499
  );


  xor
  g1962
  (
    n1661,
    n339,
    n409,
    n630,
    n207
  );


  xnor
  g1963
  (
    n1533,
    n494,
    n445,
    n520,
    n184
  );


  nor
  g1964
  (
    n2057,
    n647,
    n345,
    n493,
    n517
  );


  or
  g1965
  (
    n1693,
    n468,
    n370,
    n628,
    n214
  );


  xnor
  g1966
  (
    n724,
    n598,
    n183,
    n232,
    n434
  );


  nand
  g1967
  (
    n1749,
    n373,
    n162,
    n264,
    n392
  );


  nor
  g1968
  (
    n873,
    n522,
    n218,
    n609,
    n185
  );


  nand
  g1969
  (
    n1850,
    n233,
    n352,
    n647,
    n485
  );


  xor
  g1970
  (
    n1267,
    n525,
    n323,
    n606,
    n251
  );


  xnor
  g1971
  (
    n1022,
    n198,
    n500,
    n610,
    n647
  );


  and
  g1972
  (
    n1395,
    n479,
    n364,
    n203,
    n511
  );


  or
  g1973
  (
    n1388,
    n550,
    n626,
    n578,
    n620
  );


  xnor
  g1974
  (
    n767,
    n197,
    n562,
    n639,
    n182
  );


  and
  g1975
  (
    n1753,
    n380,
    n570,
    n592,
    n439
  );


  and
  g1976
  (
    n1508,
    n454,
    n511,
    n367,
    n209
  );


  xnor
  g1977
  (
    n893,
    n644,
    n519,
    n490,
    n572
  );


  and
  g1978
  (
    n1143,
    n268,
    n168,
    n206,
    n593
  );


  or
  g1979
  (
    n1690,
    n649,
    n570,
    n423,
    n518
  );


  and
  g1980
  (
    n1070,
    n480,
    n419,
    n603,
    n426
  );


  and
  g1981
  (
    n1751,
    n530,
    n329,
    n374,
    n197
  );


  xnor
  g1982
  (
    n812,
    n294,
    n622,
    n423,
    n273
  );


  nand
  g1983
  (
    n2030,
    n432,
    n413,
    n364,
    n290
  );


  and
  g1984
  (
    n1245,
    n253,
    n642,
    n526,
    n502
  );


  or
  g1985
  (
    n1157,
    n512,
    n348,
    n164,
    n478
  );


  nand
  g1986
  (
    n694,
    n441,
    n585,
    n609,
    n499
  );


  xnor
  g1987
  (
    n1891,
    n577,
    n318,
    n582,
    n467
  );


  nand
  g1988
  (
    n703,
    n582,
    n301,
    n390,
    n294
  );


  nor
  g1989
  (
    n1773,
    n357,
    n490,
    n257,
    n172
  );


  or
  g1990
  (
    n1488,
    n634,
    n541,
    n202,
    n286
  );


  and
  g1991
  (
    n730,
    n291,
    n597,
    n468,
    n627
  );


  nor
  g1992
  (
    n1496,
    n596,
    n382,
    n302,
    n579
  );


  nand
  g1993
  (
    n997,
    n354,
    n346,
    n474,
    n270
  );


  nor
  g1994
  (
    n1911,
    n189,
    n552,
    n271,
    n624
  );


  and
  g1995
  (
    n1646,
    n471,
    n529,
    n249,
    n469
  );


  or
  g1996
  (
    n1546,
    n303,
    n427,
    n441,
    n643
  );


  and
  g1997
  (
    n1550,
    n622,
    n574,
    n381,
    n472
  );


  xnor
  g1998
  (
    n727,
    n385,
    n484,
    n339,
    n555
  );


  nand
  g1999
  (
    n1144,
    n404,
    n404,
    n322,
    n241
  );


  xor
  g2000
  (
    n1986,
    n190,
    n576,
    n452,
    n324
  );


  nand
  g2001
  (
    n766,
    n604,
    n403,
    n377,
    n440
  );


  nand
  g2002
  (
    n706,
    n228,
    n412,
    n260,
    n610
  );


  or
  g2003
  (
    n1358,
    n201,
    n482,
    n615,
    n292
  );


  xor
  g2004
  (
    n692,
    n530,
    n170,
    n636,
    n476
  );


  and
  g2005
  (
    n1869,
    n353,
    n281,
    n637,
    n588
  );


  nand
  g2006
  (
    n1448,
    n507,
    n276,
    n204,
    n378
  );


  xor
  g2007
  (
    n999,
    n262,
    n497,
    n623,
    n196
  );


  nor
  g2008
  (
    n1667,
    n291,
    n182,
    n479,
    n408
  );


  and
  g2009
  (
    n1492,
    n277,
    n636,
    n451,
    n284
  );


  nand
  g2010
  (
    n2061,
    n432,
    n304,
    n589,
    n416
  );


  or
  g2011
  (
    n708,
    n315,
    n239,
    n404,
    n451
  );


  xnor
  g2012
  (
    n1596,
    n192,
    n257,
    n309,
    n422
  );


  nor
  g2013
  (
    n903,
    n658,
    n565,
    n351,
    n487
  );


  xnor
  g2014
  (
    n1938,
    n648,
    n413,
    n614,
    n481
  );


  and
  g2015
  (
    n1287,
    n417,
    n516,
    n553,
    n390
  );


  xor
  g2016
  (
    n1487,
    n477,
    n178,
    n495,
    n435
  );


  xnor
  g2017
  (
    n1945,
    n201,
    n455,
    n225,
    n542
  );


  xor
  g2018
  (
    n700,
    n304,
    n283,
    n496,
    n548
  );


  xnor
  g2019
  (
    n1791,
    n645,
    n630,
    n578,
    n554
  );


  and
  g2020
  (
    n872,
    n420,
    n545,
    n428,
    n443
  );


  xor
  g2021
  (
    n1608,
    n587,
    n513,
    n244,
    n342
  );


  xor
  g2022
  (
    n1451,
    n237,
    n638,
    n519,
    n176
  );


  or
  g2023
  (
    n1683,
    n608,
    n388,
    n247,
    n347
  );


  xnor
  g2024
  (
    n1383,
    n487,
    n569,
    n642,
    n309
  );


  xnor
  g2025
  (
    n1731,
    n341,
    n463,
    n440,
    n588
  );


  nor
  g2026
  (
    n1164,
    n201,
    n243,
    n476,
    n254
  );


  xnor
  g2027
  (
    n691,
    n235,
    n222,
    n579,
    n234
  );


  xnor
  g2028
  (
    n1692,
    n549,
    n621,
    n527,
    n361
  );


  nor
  g2029
  (
    n1929,
    n593,
    n514,
    n483,
    n276
  );


  xnor
  g2030
  (
    n1092,
    n466,
    n348,
    n547,
    n407
  );


  and
  g2031
  (
    n1954,
    n193,
    n294,
    n490,
    n221
  );


  xnor
  g2032
  (
    n883,
    n408,
    n199,
    n401,
    n300
  );


  and
  g2033
  (
    n925,
    n394,
    n291,
    n189,
    n485
  );


  or
  g2034
  (
    n1936,
    n310,
    n177,
    n228,
    n165
  );


  xnor
  g2035
  (
    n1129,
    n430,
    n395,
    n222,
    n546
  );


  and
  g2036
  (
    n2091,
    n1053,
    n1710,
    n1627,
    n1158
  );


  nand
  g2037
  (
    n2310,
    n714,
    n2008,
    n1893,
    n1816
  );


  xnor
  g2038
  (
    n2228,
    n1771,
    n1906,
    n1687,
    n765
  );


  xor
  g2039
  (
    n2226,
    n2027,
    n1909,
    n1154,
    n1836
  );


  or
  g2040
  (
    n2267,
    n1117,
    n781,
    n1438,
    n724
  );


  xnor
  g2041
  (
    n2083,
    n681,
    n732,
    n741,
    n1880
  );


  xnor
  g2042
  (
    n2215,
    n758,
    n2044,
    n708,
    n1014
  );


  xor
  g2043
  (
    n2407,
    n1400,
    n1731,
    n1573,
    n1297
  );


  nand
  g2044
  (
    n2271,
    n1510,
    n1564,
    n1931,
    n1020
  );


  xor
  g2045
  (
    n2232,
    n1613,
    n1256,
    n1363,
    n951
  );


  or
  g2046
  (
    n2438,
    n862,
    n1244,
    n2042,
    n2048
  );


  nand
  g2047
  (
    n2393,
    n1775,
    n1268,
    n1646,
    n1553
  );


  xor
  g2048
  (
    n2390,
    n1022,
    n1887,
    n1427,
    n1676
  );


  xnor
  g2049
  (
    n2391,
    n1692,
    n1389,
    n1420,
    n2005
  );


  and
  g2050
  (
    n2224,
    n1583,
    n1640,
    n1941,
    n763
  );


  xnor
  g2051
  (
    n2192,
    n746,
    n1795,
    n824,
    n1575
  );


  or
  g2052
  (
    n2243,
    n1959,
    n1747,
    n1950,
    n1760
  );


  nand
  g2053
  (
    n2106,
    n960,
    n1821,
    n1405,
    n1937
  );


  or
  g2054
  (
    n2355,
    n1052,
    n1361,
    n1184,
    n1074
  );


  xnor
  g2055
  (
    n2331,
    n1064,
    n1622,
    n1375,
    n1313
  );


  nand
  g2056
  (
    n2311,
    n1292,
    n1658,
    n1720,
    n1900
  );


  or
  g2057
  (
    n2346,
    n1426,
    n1418,
    n697,
    n1848
  );


  nor
  g2058
  (
    n2216,
    n1249,
    n786,
    n1849,
    n1248
  );


  nand
  g2059
  (
    n2095,
    n1855,
    n721,
    n1350,
    n784
  );


  xor
  g2060
  (
    n2400,
    n1076,
    n1278,
    n1940,
    n1041
  );


  xor
  g2061
  (
    n2342,
    n1987,
    n1414,
    n986,
    n2045
  );


  or
  g2062
  (
    n2160,
    n1057,
    n1072,
    n1499,
    n992
  );


  xnor
  g2063
  (
    n2459,
    n2051,
    n1441,
    n1119,
    n1230
  );


  nand
  g2064
  (
    n2155,
    n1634,
    n1923,
    n710,
    n974
  );


  and
  g2065
  (
    n2466,
    n880,
    n1274,
    n1419,
    n670
  );


  xnor
  g2066
  (
    n2456,
    n1630,
    n692,
    n1183,
    n1545
  );


  or
  g2067
  (
    n2314,
    n962,
    n1942,
    n2014,
    n1029
  );


  or
  g2068
  (
    n2248,
    n949,
    n1560,
    n854,
    n1989
  );


  xnor
  g2069
  (
    n2103,
    n1311,
    n1901,
    n1973,
    n1533
  );


  nand
  g2070
  (
    n2209,
    n2030,
    n1580,
    n2001,
    n720
  );


  nand
  g2071
  (
    n2108,
    n827,
    n1101,
    n899,
    n1936
  );


  xor
  g2072
  (
    n2387,
    n916,
    n1245,
    n2012,
    n1595
  );


  xor
  g2073
  (
    n2269,
    n1145,
    n2014,
    n874,
    n912
  );


  nor
  g2074
  (
    n2385,
    n752,
    n797,
    n1772,
    n1150
  );


  nand
  g2075
  (
    n2265,
    n1899,
    n1066,
    n1301,
    n1099
  );


  nand
  g2076
  (
    n2225,
    n1915,
    n1370,
    n1661,
    n926
  );


  or
  g2077
  (
    n2462,
    n1601,
    n1380,
    n1196,
    n2029
  );


  nor
  g2078
  (
    n2341,
    n861,
    n1035,
    n1168,
    n975
  );


  nand
  g2079
  (
    n2098,
    n1970,
    n1240,
    n2027,
    n2013
  );


  nand
  g2080
  (
    n2211,
    n1246,
    n1558,
    n1843,
    n1779
  );


  and
  g2081
  (
    n2425,
    n1492,
    n896,
    n1343,
    n1740
  );


  xnor
  g2082
  (
    n2277,
    n990,
    n863,
    n1901,
    n836
  );


  nand
  g2083
  (
    n2383,
    n911,
    n1004,
    n1176,
    n1265
  );


  xor
  g2084
  (
    n2227,
    n2009,
    n1452,
    n1938,
    n1999
  );


  nand
  g2085
  (
    n2244,
    n1454,
    n950,
    n887,
    n1486
  );


  and
  g2086
  (
    n2329,
    n1349,
    n1237,
    n748,
    n979
  );


  xor
  g2087
  (
    n2093,
    n1156,
    n1220,
    n1762,
    n1068
  );


  xnor
  g2088
  (
    n2444,
    n671,
    n1432,
    n849,
    n908
  );


  and
  g2089
  (
    n2455,
    n2050,
    n2025,
    n1104,
    n1989
  );


  xnor
  g2090
  (
    n2181,
    n703,
    n1137,
    n2050,
    n1830
  );


  xor
  g2091
  (
    n2251,
    n917,
    n1143,
    n1670,
    n1723
  );


  xor
  g2092
  (
    n2102,
    n779,
    n726,
    n1907,
    n1012
  );


  or
  g2093
  (
    n2401,
    n1289,
    n789,
    n2048,
    n1587
  );


  or
  g2094
  (
    n2430,
    n1636,
    n2033,
    n1952,
    n1386
  );


  or
  g2095
  (
    n2259,
    n1439,
    n1243,
    n1996,
    n914
  );


  xor
  g2096
  (
    n2193,
    n1195,
    n1565,
    n1933,
    n1146
  );


  and
  g2097
  (
    n2379,
    n715,
    n775,
    n1743,
    n774
  );


  nor
  g2098
  (
    n2365,
    n1136,
    n869,
    n1153,
    n2018
  );


  or
  g2099
  (
    n2448,
    n1546,
    n755,
    n873,
    n1062
  );


  nor
  g2100
  (
    n2240,
    n1908,
    n1189,
    n1059,
    n941
  );


  or
  g2101
  (
    n2075,
    n1091,
    n1257,
    n1352,
    n1685
  );


  or
  g2102
  (
    n2332,
    n1186,
    n1190,
    n1912,
    n761
  );


  xnor
  g2103
  (
    n2368,
    n2012,
    n2033,
    n1011,
    n1511
  );


  xor
  g2104
  (
    n2195,
    n988,
    n1907,
    n696,
    n1071
  );


  and
  g2105
  (
    n2377,
    n1532,
    n1535,
    n1684,
    n1472
  );


  or
  g2106
  (
    n2394,
    n1986,
    n1130,
    n865,
    n1395
  );


  xor
  g2107
  (
    n2419,
    n1173,
    n1031,
    n1234,
    n1015
  );


  nor
  g2108
  (
    n2289,
    n963,
    n1916,
    n1883,
    n1488
  );


  nand
  g2109
  (
    n2389,
    n1138,
    n1980,
    n707,
    n1247
  );


  nor
  g2110
  (
    n2237,
    n812,
    n1475,
    n1403,
    n2040
  );


  or
  g2111
  (
    n2122,
    n1120,
    n1042,
    n1991,
    n1251
  );


  or
  g2112
  (
    n2307,
    n2044,
    n747,
    n1148,
    n1463
  );


  nand
  g2113
  (
    n2437,
    n754,
    n2028,
    n1934,
    n1235
  );


  xnor
  g2114
  (
    n2435,
    n1898,
    n2028,
    n1121,
    n1703
  );


  xnor
  g2115
  (
    n2364,
    n791,
    n1134,
    n923,
    n1100
  );


  xnor
  g2116
  (
    n2114,
    n1797,
    n943,
    n2052,
    n1948
  );


  nand
  g2117
  (
    n2361,
    n1967,
    n1700,
    n1067,
    n940
  );


  or
  g2118
  (
    n2337,
    n691,
    n1815,
    n2040,
    n1938
  );


  or
  g2119
  (
    n2070,
    n1114,
    n1886,
    n1953,
    n2023
  );


  xor
  g2120
  (
    n2413,
    n1678,
    n872,
    n944,
    n1621
  );


  or
  g2121
  (
    n2135,
    n1216,
    n1372,
    n901,
    n1947
  );


  xnor
  g2122
  (
    n2109,
    n1976,
    n1913,
    n1956,
    n1506
  );


  nor
  g2123
  (
    n2079,
    n694,
    n1734,
    n1645,
    n1603
  );


  nand
  g2124
  (
    n2351,
    n1733,
    n1429,
    n1314,
    n1893
  );


  nor
  g2125
  (
    n2352,
    n1949,
    n1548,
    n1562,
    n686
  );


  nor
  g2126
  (
    n2399,
    n1526,
    n1659,
    n2046,
    n1933
  );


  nand
  g2127
  (
    n2176,
    n2007,
    n1838,
    n2035,
    n1958
  );


  or
  g2128
  (
    n2324,
    n1727,
    n1782,
    n1063,
    n1077
  );


  and
  g2129
  (
    n2316,
    n728,
    n1943,
    n1271,
    n2031
  );


  or
  g2130
  (
    n2194,
    n970,
    n825,
    n738,
    n1778
  );


  nor
  g2131
  (
    n2107,
    n1468,
    n1479,
    n1152,
    n712
  );


  or
  g2132
  (
    n2128,
    n679,
    n1625,
    n1721,
    n1903
  );


  xor
  g2133
  (
    n2417,
    n1503,
    n1597,
    n1112,
    n1382
  );


  nor
  g2134
  (
    n2221,
    n2025,
    n668,
    n1612,
    n1928
  );


  xnor
  g2135
  (
    n2201,
    n782,
    n1858,
    n1803,
    n1316
  );


  xor
  g2136
  (
    n2085,
    n1366,
    n1222,
    n1997,
    n1284
  );


  or
  g2137
  (
    n2447,
    n1940,
    n1713,
    n1518,
    n1302
  );


  nor
  g2138
  (
    n2446,
    n1914,
    n2046,
    n793,
    n1941
  );


  nand
  g2139
  (
    n2319,
    n1976,
    n1990,
    n1281,
    n1748
  );


  xor
  g2140
  (
    n2443,
    n1096,
    n846,
    n972,
    n1217
  );


  xor
  g2141
  (
    n2129,
    n1856,
    n1219,
    n722,
    n1936
  );


  nor
  g2142
  (
    n2283,
    n1416,
    n819,
    n994,
    n1959
  );


  nand
  g2143
  (
    n2092,
    n876,
    n977,
    n953,
    n1770
  );


  xnor
  g2144
  (
    n2273,
    n2027,
    n1730,
    n1385,
    n1951
  );


  nand
  g2145
  (
    n2077,
    n1852,
    n1774,
    n829,
    n830
  );


  nor
  g2146
  (
    n2469,
    n834,
    n1862,
    n2045,
    n2050
  );


  or
  g2147
  (
    KeyWire_0_31,
    n999,
    n1007,
    n1097,
    n1339
  );


  and
  g2148
  (
    n2349,
    n2026,
    n919,
    n2049,
    n1755
  );


  xor
  g2149
  (
    n2428,
    n1436,
    n2052,
    n706,
    n1377
  );


  and
  g2150
  (
    n2223,
    n1962,
    n809,
    n935,
    n1214
  );


  nand
  g2151
  (
    n2431,
    n1846,
    n687,
    n2011,
    n1899
  );


  nor
  g2152
  (
    n2285,
    n1529,
    n1181,
    n1309,
    n1261
  );


  nand
  g2153
  (
    n2140,
    n895,
    n1501,
    n2029,
    n1924
  );


  or
  g2154
  (
    n2260,
    n1332,
    n1598,
    n682,
    n1460
  );


  xnor
  g2155
  (
    n2247,
    n930,
    n1824,
    n1983,
    n1177
  );


  xnor
  g2156
  (
    n2143,
    n1844,
    n1790,
    n1667,
    n2033
  );


  nand
  g2157
  (
    n2465,
    n1725,
    n948,
    n1258,
    n983
  );


  nand
  g2158
  (
    KeyWire_0_59,
    n1135,
    n2026,
    n676,
    n1996
  );


  xor
  g2159
  (
    n2111,
    n1393,
    n1210,
    n801,
    n844
  );


  or
  g2160
  (
    n2410,
    n1079,
    n1030,
    n1085,
    n1863
  );


  nand
  g2161
  (
    n2336,
    n1997,
    n877,
    n1293,
    n1507
  );


  xnor
  g2162
  (
    n2278,
    n1956,
    n1726,
    n1351,
    n1491
  );


  xnor
  g2163
  (
    n2212,
    n1974,
    n1555,
    n1891,
    n2024
  );


  xnor
  g2164
  (
    n2188,
    n1756,
    n1524,
    n1592,
    n1691
  );


  and
  g2165
  (
    n2069,
    n1909,
    n1178,
    n702,
    n1635
  );


  xor
  g2166
  (
    n2113,
    n1149,
    n1614,
    n1127,
    n2019
  );


  nor
  g2167
  (
    n2152,
    n813,
    n2040,
    n1780,
    n1025
  );


  xor
  g2168
  (
    n2149,
    n1364,
    n1045,
    n1910,
    n1428
  );


  xnor
  g2169
  (
    n2270,
    n1967,
    n1896,
    n1514,
    n1897
  );


  xor
  g2170
  (
    n2142,
    n1861,
    n1371,
    n1800,
    n1576
  );


  xor
  g2171
  (
    n2262,
    n770,
    n1594,
    n1490,
    n1906
  );


  xor
  g2172
  (
    n2461,
    n1801,
    n778,
    n2041,
    n1473
  );


  xor
  g2173
  (
    n2214,
    n1509,
    n1056,
    n1988,
    n2000
  );


  and
  g2174
  (
    n2133,
    n1758,
    n1991,
    n1399,
    n1001
  );


  and
  g2175
  (
    n2239,
    n760,
    n2034,
    n1252,
    n965
  );


  nand
  g2176
  (
    n2139,
    n1903,
    n1865,
    n785,
    n1295
  );


  nand
  g2177
  (
    n2220,
    n2020,
    n841,
    n1920,
    n1878
  );


  nand
  g2178
  (
    n2238,
    n2011,
    n2016,
    n1530,
    n1369
  );


  nand
  g2179
  (
    n2235,
    n1859,
    n1890,
    n1980,
    n1390
  );


  or
  g2180
  (
    n2445,
    n1904,
    n759,
    n1043,
    n832
  );


  and
  g2181
  (
    n2320,
    n1746,
    n1051,
    n1572,
    n1707
  );


  xor
  g2182
  (
    n2422,
    n934,
    n1945,
    n2038,
    n2006
  );


  nor
  g2183
  (
    n2156,
    n2029,
    n716,
    n1718,
    n1192
  );


  nand
  g2184
  (
    n2296,
    n2041,
    n1679,
    n1935,
    n1487
  );


  nor
  g2185
  (
    n2080,
    n1182,
    n807,
    n1242,
    n902
  );


  xnor
  g2186
  (
    n2326,
    n1812,
    n1408,
    n2037,
    n1513
  );


  and
  g2187
  (
    n2101,
    n1430,
    n1638,
    n1525,
    n1674
  );


  nand
  g2188
  (
    n2124,
    n1753,
    n685,
    n1517,
    n2010
  );


  nand
  g2189
  (
    n2163,
    n1927,
    n1307,
    n976,
    n1541
  );


  nand
  g2190
  (
    n2170,
    n1698,
    n1159,
    n2043,
    n1966
  );


  or
  g2191
  (
    n2317,
    n1550,
    n987,
    n1781,
    n1722
  );


  nand
  g2192
  (
    n2177,
    n1892,
    n1742,
    n892,
    n1116
  );


  or
  g2193
  (
    n2414,
    n1706,
    n1449,
    n680,
    n1964
  );


  xnor
  g2194
  (
    n2118,
    n733,
    n1276,
    n1662,
    n1126
  );


  xor
  g2195
  (
    n2275,
    n1516,
    n795,
    n1600,
    n878
  );


  nor
  g2196
  (
    n2268,
    n742,
    n1992,
    n1105,
    n1643
  );


  xnor
  g2197
  (
    n2348,
    n1425,
    n1884,
    n1785,
    n851
  );


  xor
  g2198
  (
    n2460,
    n1663,
    n1038,
    n1003,
    n2017
  );


  xor
  g2199
  (
    n2301,
    n1017,
    n1373,
    n1140,
    n1329
  );


  or
  g2200
  (
    n2427,
    n699,
    n1037,
    n858,
    n1123
  );


  xor
  g2201
  (
    n2290,
    n2044,
    n1660,
    n1765,
    n1098
  );


  and
  g2202
  (
    n2436,
    n1632,
    n1671,
    n1819,
    n1777
  );


  or
  g2203
  (
    n2322,
    n1609,
    n2044,
    n1599,
    n2036
  );


  xor
  g2204
  (
    n2345,
    n1853,
    n1170,
    n2031,
    n1995
  );


  and
  g2205
  (
    n2468,
    n1552,
    n1736,
    n1000,
    n1484
  );


  nand
  g2206
  (
    n2249,
    n890,
    n727,
    n2022,
    n1900
  );


  xnor
  g2207
  (
    n2137,
    n993,
    n1639,
    n1021,
    n1954
  );


  nand
  g2208
  (
    n2409,
    n1789,
    n1424,
    n956,
    n1090
  );


  nand
  g2209
  (
    n2408,
    n1335,
    n980,
    n2030,
    n1683
  );


  xor
  g2210
  (
    n2339,
    n698,
    n1433,
    n1238,
    n1624
  );


  xnor
  g2211
  (
    n2297,
    n1241,
    n2036,
    n1589,
    n1916
  );


  nand
  g2212
  (
    n2246,
    n800,
    n689,
    n1194,
    n1571
  );


  and
  g2213
  (
    n2340,
    n1212,
    n1935,
    n1291,
    n1867
  );


  and
  g2214
  (
    n2199,
    n898,
    n1554,
    n1005,
    n2036
  );


  xor
  g2215
  (
    n2125,
    n1344,
    n2035,
    n1929,
    n2021
  );


  nor
  g2216
  (
    n2374,
    n1682,
    n1203,
    n2037,
    n804
  );


  xnor
  g2217
  (
    n2190,
    n852,
    n1327,
    n1939,
    n1157
  );


  nand
  g2218
  (
    n2241,
    n1055,
    n1569,
    n1811,
    n1719
  );


  nand
  g2219
  (
    n2454,
    n773,
    n964,
    n1282,
    n1397
  );


  or
  g2220
  (
    n2250,
    n1891,
    n1505,
    n1283,
    n1118
  );


  or
  g2221
  (
    n2266,
    n1087,
    n1111,
    n1966,
    n1911
  );


  xnor
  g2222
  (
    n2218,
    n1574,
    n1286,
    n2034,
    n1922
  );


  and
  g2223
  (
    KeyWire_0_5,
    n822,
    n1255,
    n1358,
    n2029
  );


  and
  g2224
  (
    n2323,
    n1465,
    n1467,
    n1163,
    n913
  );


  nor
  g2225
  (
    n2150,
    n831,
    n1680,
    n739,
    n850
  );


  xor
  g2226
  (
    n2168,
    n1102,
    n672,
    n1481,
    n2043
  );


  xor
  g2227
  (
    n2229,
    n1926,
    n2013,
    n2042,
    n1677
  );


  and
  g2228
  (
    n2406,
    n1808,
    n1885,
    n1969,
    n1191
  );


  nand
  g2229
  (
    n2360,
    n1175,
    n1981,
    n875,
    n1462
  );


  or
  g2230
  (
    n2432,
    n1890,
    n1131,
    n835,
    n1898
  );


  or
  g2231
  (
    n2180,
    n802,
    n1006,
    n1421,
    n1620
  );


  xnor
  g2232
  (
    n2115,
    n1187,
    n796,
    n1934,
    n1260
  );


  xnor
  g2233
  (
    n2376,
    n1489,
    n2038,
    n1809,
    n1791
  );


  nand
  g2234
  (
    n2302,
    n837,
    n1201,
    n1711,
    n870
  );


  nor
  g2235
  (
    n2242,
    n1990,
    n1398,
    n1315,
    n1995
  );


  xor
  g2236
  (
    n2325,
    n855,
    n718,
    n1902,
    n1226
  );


  xor
  g2237
  (
    n2164,
    n1764,
    n1331,
    n764,
    n968
  );


  nor
  g2238
  (
    n2334,
    n1984,
    n1943,
    n1768,
    n1732
  );


  xnor
  g2239
  (
    n2146,
    n2039,
    n1290,
    n1457,
    n1032
  );


  xnor
  g2240
  (
    n2126,
    n932,
    n1961,
    n1147,
    n1054
  );


  nand
  g2241
  (
    n2198,
    n725,
    n1911,
    n1083,
    n833
  );


  nor
  g2242
  (
    n2076,
    n1978,
    n1827,
    n1879,
    n1568
  );


  or
  g2243
  (
    n2230,
    n723,
    n1641,
    n1270,
    n1229
  );


  xor
  g2244
  (
    n2415,
    n2047,
    n1690,
    n1729,
    n1832
  );


  xnor
  g2245
  (
    n2169,
    n1310,
    n1211,
    n1374,
    n997
  );


  xnor
  g2246
  (
    n2100,
    n1160,
    n1889,
    n2041,
    n995
  );


  xnor
  g2247
  (
    n2309,
    n1963,
    n1476,
    n1413,
    n1813
  );


  nor
  g2248
  (
    n2353,
    n1233,
    n1478,
    n1642,
    n1082
  );


  and
  g2249
  (
    n2219,
    n2005,
    n1932,
    n1666,
    n1818
  );


  and
  g2250
  (
    n2356,
    n961,
    n1267,
    n1977,
    n1434
  );


  nand
  g2251
  (
    n2452,
    n1735,
    n1987,
    n1287,
    n751
  );


  xnor
  g2252
  (
    n2127,
    n1950,
    n1502,
    n1317,
    n1320
  );


  nor
  g2253
  (
    n2234,
    n1665,
    n2046,
    n1303,
    n1285
  );


  and
  g2254
  (
    n2094,
    n1988,
    n847,
    n954,
    n1953
  );


  xnor
  g2255
  (
    n2412,
    n1851,
    n1180,
    n2019,
    n1799
  );


  nand
  g2256
  (
    n2305,
    n669,
    n1608,
    n927,
    n2026
  );


  xnor
  g2257
  (
    n2151,
    n1443,
    n1961,
    n709,
    n1681
  );


  nand
  g2258
  (
    n2450,
    n1912,
    n1955,
    n1048,
    n701
  );


  xor
  g2259
  (
    n2371,
    n1461,
    n1929,
    n1368,
    n1845
  );


  xor
  g2260
  (
    n2279,
    n1384,
    n2007,
    n1129,
    n1688
  );


  nor
  g2261
  (
    n2350,
    n1829,
    n1132,
    n1590,
    n1537
  );


  xnor
  g2262
  (
    n2207,
    n1557,
    n1993,
    n1823,
    n1124
  );


  or
  g2263
  (
    n2449,
    n1155,
    n947,
    n2047,
    n1767
  );


  xor
  g2264
  (
    n2358,
    n820,
    n1346,
    n1367,
    n1868
  );


  and
  g2265
  (
    n2172,
    n966,
    n1944,
    n1992,
    n1239
  );


  or
  g2266
  (
    n2402,
    n1080,
    n777,
    n1355,
    n1628
  );


  xor
  g2267
  (
    n2105,
    n1084,
    n1889,
    n1095,
    n1539
  );


  nand
  g2268
  (
    n2304,
    n1984,
    n1401,
    n1169,
    n1167
  );


  or
  g2269
  (
    n2404,
    n1294,
    n1915,
    n1543,
    n1515
  );


  nand
  g2270
  (
    n2295,
    n2034,
    n1820,
    n996,
    n2024
  );


  nand
  g2271
  (
    n2173,
    n1894,
    n1593,
    n1979,
    n1275
  );


  nand
  g2272
  (
    n2179,
    n1975,
    n1133,
    n1874,
    n1334
  );


  nand
  g2273
  (
    n2470,
    n1205,
    n1918,
    n1411,
    n1070
  );


  or
  g2274
  (
    n2202,
    n1847,
    n881,
    n1221,
    n1657
  );


  xnor
  g2275
  (
    n2148,
    n1971,
    n1567,
    n1209,
    n1277
  );


  xnor
  g2276
  (
    n2084,
    n1027,
    n1174,
    n1607,
    n675
  );


  and
  g2277
  (
    n2116,
    n907,
    n1814,
    n1741,
    n1834
  );


  or
  g2278
  (
    n2191,
    n1376,
    n1921,
    n1796,
    n1456
  );


  xnor
  g2279
  (
    n2375,
    n2031,
    n1977,
    n1435,
    n1648
  );


  xor
  g2280
  (
    n2388,
    n1236,
    n1142,
    n792,
    n1857
  );


  xor
  g2281
  (
    n2363,
    n1952,
    n1047,
    n745,
    n1325
  );


  xnor
  g2282
  (
    n2381,
    n1647,
    n1365,
    n1833,
    n1404
  );


  xor
  g2283
  (
    n2395,
    n1300,
    n859,
    n1321,
    n1534
  );


  or
  g2284
  (
    n2457,
    n978,
    n891,
    n1549,
    n937
  );


  or
  g2285
  (
    n2421,
    n2043,
    n1306,
    n1757,
    n922
  );


  nand
  g2286
  (
    n2318,
    n772,
    n729,
    n1616,
    n1944
  );


  nand
  g2287
  (
    n2369,
    n816,
    n1787,
    n1615,
    n673
  );


  nand
  g2288
  (
    n2261,
    n1918,
    n1709,
    n936,
    n1651
  );


  xnor
  g2289
  (
    n2138,
    n735,
    n814,
    n828,
    n883
  );


  xnor
  g2290
  (
    n2208,
    n1474,
    n2049,
    n1470,
    n1694
  );


  and
  g2291
  (
    n2380,
    n1431,
    n1206,
    n1994,
    n1026
  );


  xnor
  g2292
  (
    n2217,
    n1391,
    n1407,
    n1860,
    n1280
  );


  nand
  g2293
  (
    n2231,
    n767,
    n1570,
    n798,
    n1122
  );


  xnor
  g2294
  (
    n2464,
    n787,
    n1039,
    n1109,
    n1299
  );


  nor
  g2295
  (
    n2293,
    n1802,
    n1793,
    n1551,
    n920
  );


  nand
  g2296
  (
    n2099,
    n1652,
    n1686,
    n1822,
    n2048
  );


  nor
  g2297
  (
    n2372,
    n1324,
    n1360,
    n2017,
    n1982
  );


  and
  g2298
  (
    n2132,
    n1716,
    n711,
    n734,
    n2030
  );


  xor
  g2299
  (
    n2121,
    n998,
    n1250,
    n815,
    n1523
  );


  nand
  g2300
  (
    n2258,
    n2031,
    n1873,
    n918,
    n1092
  );


  nor
  g2301
  (
    n2144,
    n731,
    n783,
    n1617,
    n674
  );


  or
  g2302
  (
    n2123,
    n1304,
    n973,
    n1078,
    n1342
  );


  and
  g2303
  (
    n2392,
    n1538,
    n719,
    n704,
    n1008
  );


  nand
  g2304
  (
    n2233,
    n1605,
    n766,
    n1745,
    n1269
  );


  xnor
  g2305
  (
    n2157,
    n1065,
    n1455,
    n2003,
    n1223
  );


  xor
  g2306
  (
    n2073,
    n1654,
    n1761,
    n1922,
    n871
  );


  xnor
  g2307
  (
    n2222,
    n1296,
    n688,
    n1669,
    n1009
  );


  nor
  g2308
  (
    n2291,
    n1914,
    n1752,
    n1942,
    n946
  );


  nor
  g2309
  (
    n2359,
    n1094,
    n1672,
    n2048,
    n1081
  );


  xnor
  g2310
  (
    n2338,
    n1161,
    n1125,
    n1347,
    n1699
  );


  and
  g2311
  (
    n2166,
    n2035,
    n1999,
    n1536,
    n1960
  );


  and
  g2312
  (
    n2178,
    n1266,
    n1697,
    n821,
    n1939
  );


  nor
  g2313
  (
    n2255,
    n2033,
    n1872,
    n1751,
    n1406
  );


  nor
  g2314
  (
    KeyWire_0_21,
    n1655,
    n1337,
    n839,
    n1958
  );


  and
  g2315
  (
    n2347,
    n1817,
    n1262,
    n1895,
    n1379
  );


  and
  g2316
  (
    n2458,
    n969,
    n842,
    n1409,
    n2042
  );


  xnor
  g2317
  (
    n2335,
    n1892,
    n1749,
    n1932,
    n1586
  );


  nor
  g2318
  (
    n2086,
    n1402,
    n1588,
    n1604,
    n2015
  );


  and
  g2319
  (
    n2434,
    n1920,
    n1086,
    n904,
    n955
  );


  xor
  g2320
  (
    n2288,
    n1807,
    n1493,
    n894,
    n1519
  );


  xor
  g2321
  (
    n2090,
    n1224,
    n1036,
    n1910,
    n2052
  );


  nand
  g2322
  (
    n2354,
    n1930,
    n2024,
    n1704,
    n1088
  );


  or
  g2323
  (
    n2321,
    n845,
    n958,
    n1925,
    n1263
  );


  and
  g2324
  (
    n2313,
    n1982,
    n2026,
    n1965,
    n1396
  );


  and
  g2325
  (
    n2333,
    n1656,
    n1483,
    n1970,
    n1423
  );


  xnor
  g2326
  (
    n2096,
    n1596,
    n1016,
    n1715,
    n749
  );


  or
  g2327
  (
    n2467,
    n1695,
    n1540,
    n1913,
    n931
  );


  or
  g2328
  (
    n2205,
    n1166,
    n1919,
    n939,
    n1957
  );


  xor
  g2329
  (
    n2071,
    n1610,
    n1326,
    n1972,
    n1387
  );


  xor
  g2330
  (
    n2120,
    n1259,
    n1179,
    n808,
    n985
  );


  xnor
  g2331
  (
    n2183,
    n1305,
    n1839,
    n1113,
    n730
  );


  nand
  g2332
  (
    n2104,
    n1144,
    n1664,
    n915,
    n1579
  );


  and
  g2333
  (
    n2300,
    n1049,
    n1061,
    n1050,
    n924
  );


  and
  g2334
  (
    n2184,
    n1653,
    n1837,
    n933,
    n1228
  );


  nand
  g2335
  (
    n2154,
    n1835,
    n1650,
    n1924,
    n1308
  );


  nor
  g2336
  (
    n2161,
    n1875,
    n1921,
    n2039,
    n1446
  );


  xnor
  g2337
  (
    n2286,
    n1496,
    n1328,
    n1805,
    n1378
  );


  xnor
  g2338
  (
    n2440,
    n2008,
    n1784,
    n1069,
    n929
  );


  nand
  g2339
  (
    n2136,
    n868,
    n984,
    n1482,
    n743
  );


  xnor
  g2340
  (
    n2423,
    n2010,
    n1556,
    n753,
    n1415
  );


  or
  g2341
  (
    n2263,
    n1962,
    n780,
    n2028,
    n1357
  );


  nor
  g2342
  (
    n2362,
    n1383,
    n2022,
    n695,
    n1831
  );


  xor
  g2343
  (
    n2429,
    n1544,
    n1728,
    n736,
    n1520
  );


  xor
  g2344
  (
    n2287,
    n1629,
    n1948,
    n1040,
    n1759
  );


  xnor
  g2345
  (
    n2097,
    n1232,
    n2025,
    n2027,
    n1675
  );


  xor
  g2346
  (
    n2405,
    n942,
    n1881,
    n2038,
    n1497
  );


  nor
  g2347
  (
    n2370,
    n1869,
    n1495,
    n897,
    n799
  );


  or
  g2348
  (
    n2367,
    n1188,
    n1561,
    n971,
    n2051
  );


  nor
  g2349
  (
    n2072,
    n879,
    n2018,
    n1323,
    n1786
  );


  nor
  g2350
  (
    n2378,
    n1107,
    n2032,
    n1696,
    n1340
  );


  or
  g2351
  (
    n2254,
    n823,
    n737,
    n2009,
    n1458
  );


  nor
  g2352
  (
    n2245,
    n882,
    n991,
    n2049,
    n1923
  );


  or
  g2353
  (
    n2312,
    n740,
    n938,
    n1231,
    n1888
  );


  or
  g2354
  (
    n2130,
    n2037,
    n1139,
    n1611,
    n817
  );


  nand
  g2355
  (
    n2403,
    n1422,
    n1559,
    n1960,
    n893
  );


  xor
  g2356
  (
    n2386,
    n1410,
    n1288,
    n1864,
    n1500
  );


  or
  g2357
  (
    n2252,
    n1312,
    n1945,
    n1673,
    n1521
  );


  xnor
  g2358
  (
    n2330,
    n1273,
    n713,
    n2025,
    n1850
  );


  xnor
  g2359
  (
    n2110,
    n1018,
    n2032,
    n2000,
    n1448
  );


  and
  g2360
  (
    n2282,
    n803,
    n909,
    n769,
    n1471
  );


  xnor
  g2361
  (
    n2089,
    n757,
    n1917,
    n1566,
    n1794
  );


  nor
  g2362
  (
    n2411,
    n2023,
    n2035,
    n1902,
    n1577
  );


  or
  g2363
  (
    n2112,
    n957,
    n925,
    n1766,
    n1033
  );


  xnor
  g2364
  (
    n2074,
    n886,
    n1019,
    n2036,
    n810
  );


  and
  g2365
  (
    n2366,
    n1165,
    n1034,
    n776,
    n1108
  );


  xnor
  g2366
  (
    n2420,
    n1024,
    n1998,
    n1951,
    n1060
  );


  and
  g2367
  (
    n2439,
    n788,
    n1527,
    n1798,
    n1585
  );


  and
  g2368
  (
    n2442,
    n1985,
    n2001,
    n867,
    n1637
  );


  nand
  g2369
  (
    n2210,
    n1973,
    n2052,
    n1563,
    n853
  );


  and
  g2370
  (
    n2141,
    n921,
    n1013,
    n1969,
    n1788
  );


  xor
  g2371
  (
    n2078,
    n1469,
    n818,
    n1689,
    n1141
  );


  nor
  g2372
  (
    n2162,
    n1870,
    n1046,
    n1512,
    n1986
  );


  nor
  g2373
  (
    n2451,
    n848,
    n1618,
    n744,
    n888
  );


  nand
  g2374
  (
    n2159,
    n1957,
    n1348,
    n1894,
    n1714
  );


  xor
  g2375
  (
    n2357,
    n678,
    n2037,
    n1581,
    n1508
  );


  and
  g2376
  (
    n2174,
    n1164,
    n1578,
    n1606,
    n1336
  );


  nor
  g2377
  (
    n2294,
    n1264,
    n1840,
    n1965,
    n1925
  );


  xnor
  g2378
  (
    n2253,
    n1480,
    n1955,
    n2002,
    n1171
  );


  xnor
  g2379
  (
    n2281,
    n1322,
    n2004,
    n1073,
    n1947
  );


  or
  g2380
  (
    n2264,
    n1876,
    n1994,
    n1946,
    n900
  );


  and
  g2381
  (
    n2196,
    n1623,
    n2041,
    n1466,
    n690
  );


  and
  g2382
  (
    n2426,
    n1253,
    n1737,
    n2051,
    n1353
  );


  nor
  g2383
  (
    n2206,
    n1450,
    n1693,
    n1412,
    n1895
  );


  nor
  g2384
  (
    n2441,
    n750,
    n1531,
    n982,
    n1750
  );


  or
  g2385
  (
    KeyWire_0_13,
    n1773,
    n1272,
    n1075,
    n1225
  );


  nand
  g2386
  (
    n2398,
    n2040,
    n1877,
    n1002,
    n1954
  );


  and
  g2387
  (
    n2424,
    n1631,
    n1602,
    n1668,
    n2006
  );


  or
  g2388
  (
    n2081,
    n1198,
    n1172,
    n1792,
    n1093
  );


  xnor
  g2389
  (
    n2306,
    n952,
    n2045,
    n2034,
    n885
  );


  and
  g2390
  (
    n2396,
    n2039,
    n1345,
    n1985,
    n1447
  );


  xor
  g2391
  (
    n2200,
    n889,
    n1633,
    n1841,
    n2047
  );


  xnor
  g2392
  (
    n2131,
    n1908,
    n1227,
    n1044,
    n838
  );


  or
  g2393
  (
    n2274,
    n884,
    n1362,
    n1359,
    n1341
  );


  xor
  g2394
  (
    n2257,
    n1804,
    n805,
    n1417,
    n1769
  );


  nor
  g2395
  (
    n2167,
    n1381,
    n2004,
    n1993,
    n1584
  );


  nor
  g2396
  (
    n2256,
    n1494,
    n1333,
    n1542,
    n1724
  );


  xor
  g2397
  (
    n2182,
    n1477,
    n811,
    n1972,
    n2003
  );


  nor
  g2398
  (
    n2189,
    n1701,
    n1998,
    n1254,
    n928
  );


  and
  g2399
  (
    KeyWire_0_62,
    n2024,
    n1930,
    n1825,
    n1451
  );


  xor
  g2400
  (
    n2213,
    n1437,
    n1905,
    n1783,
    n1866
  );


  nand
  g2401
  (
    n2373,
    n2015,
    n1547,
    n1937,
    n1582
  );


  or
  g2402
  (
    n2308,
    n1979,
    n1522,
    n1193,
    n1388
  );


  nand
  g2403
  (
    n2171,
    n1649,
    n1028,
    n762,
    n1103
  );


  xnor
  g2404
  (
    n2315,
    n1927,
    n2030,
    n717,
    n945
  );


  nand
  g2405
  (
    n2134,
    n1440,
    n1854,
    n1394,
    n1963
  );


  and
  g2406
  (
    n2298,
    n1591,
    n1744,
    n1442,
    n1356
  );


  and
  g2407
  (
    n2175,
    n1888,
    n1626,
    n1202,
    n790
  );


  nand
  g2408
  (
    n2082,
    n1464,
    n1968,
    n856,
    n2051
  );


  nor
  g2409
  (
    n2327,
    n2021,
    n1200,
    n1971,
    n1197
  );


  nand
  g2410
  (
    n2088,
    n1485,
    n700,
    n1826,
    n1702
  );


  and
  g2411
  (
    n2197,
    n2046,
    n1810,
    n1498,
    n959
  );


  nand
  g2412
  (
    n2280,
    n1983,
    n1754,
    n2039,
    n826
  );


  and
  g2413
  (
    n2276,
    n1199,
    n2032,
    n1207,
    n1705
  );


  nor
  g2414
  (
    n2165,
    n1964,
    n794,
    n1338,
    n1712
  );


  nand
  g2415
  (
    n2147,
    n1981,
    n2028,
    n1904,
    n705
  );


  xor
  g2416
  (
    n2185,
    n2002,
    n1776,
    n1208,
    n1978
  );


  nor
  g2417
  (
    n2236,
    n1318,
    n1354,
    n1444,
    n693
  );


  nor
  g2418
  (
    n2453,
    n1330,
    n768,
    n2042,
    n1928
  );


  nand
  g2419
  (
    n2119,
    n860,
    n1763,
    n1453,
    n1023
  );


  or
  g2420
  (
    n2204,
    n1151,
    n1828,
    n1946,
    n1896
  );


  nand
  g2421
  (
    n2087,
    n1806,
    n903,
    n1298,
    n1905
  );


  and
  g2422
  (
    n2292,
    n1319,
    n1897,
    n806,
    n1213
  );


  and
  g2423
  (
    n2384,
    n1010,
    n1162,
    n677,
    n1528
  );


  and
  g2424
  (
    n2145,
    n2049,
    n2047,
    n1739,
    n1504
  );


  nand
  g2425
  (
    n2303,
    n857,
    n683,
    n1644,
    n2032
  );


  and
  g2426
  (
    n2284,
    n1185,
    n2020,
    n1058,
    n1392
  );


  nor
  g2427
  (
    n2416,
    n1128,
    n1215,
    n1842,
    n771
  );


  xor
  g2428
  (
    n2397,
    n1931,
    n1882,
    n905,
    n2016
  );


  nand
  g2429
  (
    n2186,
    n1445,
    n843,
    n1619,
    n906
  );


  and
  g2430
  (
    n2433,
    n981,
    n1917,
    n1115,
    n1106
  );


  nand
  g2431
  (
    n2418,
    n1871,
    n1110,
    n1717,
    n1974
  );


  or
  g2432
  (
    n2328,
    n840,
    n2038,
    n1926,
    n1089
  );


  xor
  g2433
  (
    n2343,
    n1968,
    n866,
    n684,
    n2045
  );


  xor
  g2434
  (
    n2463,
    n1919,
    n1708,
    n2050,
    n1975
  );


  xor
  g2435
  (
    n2158,
    n989,
    n910,
    n2043,
    n756
  );


  xnor
  g2436
  (
    n2344,
    n1738,
    n1949,
    n1279,
    n967
  );


  or
  g2437
  (
    KeyWire_0_58,
    n864,
    n1204,
    n1218,
    n1459
  );


  buf
  g2438
  (
    n2487,
    n2074
  );


  not
  g2439
  (
    n2479,
    n2098
  );


  not
  g2440
  (
    n2471,
    n2091
  );


  buf
  g2441
  (
    n2484,
    n2077
  );


  or
  g2442
  (
    n2472,
    n2072,
    n2082
  );


  and
  g2443
  (
    n2475,
    n2076,
    n2080
  );


  xnor
  g2444
  (
    n2481,
    n2097,
    n2087
  );


  nor
  g2445
  (
    n2476,
    n2096,
    n2085
  );


  or
  g2446
  (
    n2473,
    n2069,
    n2079
  );


  nand
  g2447
  (
    n2485,
    n2094,
    n2073
  );


  nor
  g2448
  (
    n2480,
    n2090,
    n2092
  );


  xor
  g2449
  (
    n2474,
    n2081,
    n2075
  );


  nor
  g2450
  (
    n2483,
    n2086,
    n2084
  );


  xnor
  g2451
  (
    n2486,
    n2088,
    n2089
  );


  and
  g2452
  (
    KeyWire_0_53,
    n2095,
    n2071
  );


  nor
  g2453
  (
    n2482,
    n2070,
    n2078
  );


  xnor
  g2454
  (
    n2477,
    n2083,
    n2093
  );


  nor
  g2455
  (
    n2501,
    n2057,
    n2061,
    n2055,
    n2058
  );


  and
  g2456
  (
    n2505,
    n2059,
    n2055,
    n2471,
    n2061
  );


  xor
  g2457
  (
    n2495,
    n2062,
    n2059,
    n2053,
    n2063
  );


  and
  g2458
  (
    n2500,
    n2483,
    n2061,
    n2064,
    n2053
  );


  nor
  g2459
  (
    n2493,
    n2060,
    n2057,
    n2485,
    n2472
  );


  xor
  g2460
  (
    n2497,
    n2480,
    n2061,
    n2057,
    n2060
  );


  or
  g2461
  (
    n2502,
    n2054,
    n2053,
    n2056,
    n2055
  );


  and
  g2462
  (
    n2496,
    n2099,
    n2063,
    n2487,
    n2475
  );


  xor
  g2463
  (
    n2492,
    n2064,
    n2055,
    n2060,
    n2059
  );


  xor
  g2464
  (
    n2498,
    n2100,
    n2058,
    n2059,
    n2481
  );


  xor
  g2465
  (
    n2503,
    n2060,
    n2058,
    n2482,
    n2053
  );


  nand
  g2466
  (
    n2491,
    n2056,
    n2054,
    n2477,
    n2103
  );


  or
  g2467
  (
    n2489,
    n2478,
    n2487,
    n2479,
    n2062
  );


  nor
  g2468
  (
    n2490,
    n2473,
    n2062,
    n2054
  );


  nor
  g2469
  (
    n2499,
    n2063,
    n2104,
    n2064,
    n2062
  );


  xor
  g2470
  (
    n2488,
    n2057,
    n2484,
    n2056,
    n2474
  );


  xor
  g2471
  (
    n2494,
    n2486,
    n2063,
    n2101,
    n2058
  );


  xor
  g2472
  (
    n2504,
    n2056,
    n2476,
    n2064,
    n2102
  );


  buf
  g2473
  (
    n2511,
    n2494
  );


  buf
  g2474
  (
    n2508,
    n2105
  );


  nor
  g2475
  (
    n2507,
    n2110,
    n2114
  );


  nand
  g2476
  (
    n2512,
    n2488,
    n2116,
    n2117,
    n2492
  );


  xor
  g2477
  (
    n2509,
    n2491,
    n2108,
    n2113,
    n2493
  );


  or
  g2478
  (
    KeyWire_0_43,
    n2111,
    n2489,
    n2107,
    n2112
  );


  nor
  g2479
  (
    n2510,
    n2490,
    n2106,
    n2109,
    n2115
  );


  buf
  g2480
  (
    n2536,
    n2509
  );


  buf
  g2481
  (
    n2533,
    n2507
  );


  nand
  g2482
  (
    n2527,
    n2506,
    n2177
  );


  nor
  g2483
  (
    n2519,
    n2173,
    n2172,
    n2508,
    n2510
  );


  xnor
  g2484
  (
    n2530,
    n2162,
    n2511,
    n2158
  );


  nand
  g2485
  (
    n2523,
    n2128,
    n2130,
    n2123,
    n2150
  );


  or
  g2486
  (
    n2514,
    n2512,
    n2155,
    n2119,
    n2139
  );


  and
  g2487
  (
    n2532,
    n2185,
    n2159,
    n2171,
    n2136
  );


  and
  g2488
  (
    n2522,
    n2129,
    n2175,
    n2153,
    n2131
  );


  or
  g2489
  (
    n2528,
    n2127,
    n2509,
    n2168,
    n2142
  );


  xor
  g2490
  (
    n2526,
    n2187,
    n2149,
    n2512
  );


  xor
  g2491
  (
    n2529,
    n2147,
    n2508,
    n2132,
    n2176
  );


  xor
  g2492
  (
    n2538,
    n2164,
    n2161,
    n2124,
    n2507
  );


  xnor
  g2493
  (
    n2513,
    n2508,
    n2506,
    n2126,
    n2509
  );


  and
  g2494
  (
    n2524,
    n2156,
    n2140,
    n2174,
    n2180
  );


  nor
  g2495
  (
    n2534,
    n2510,
    n2507,
    n2133,
    n2182
  );


  xnor
  g2496
  (
    n2531,
    n2163,
    n2178,
    n2146,
    n2179
  );


  or
  g2497
  (
    n2521,
    n2511,
    n2170,
    n2186,
    n2120
  );


  nand
  g2498
  (
    n2515,
    n2181,
    n2167,
    n2144,
    n2135
  );


  nand
  g2499
  (
    n2537,
    n2151,
    n2169,
    n2125,
    n2118
  );


  nand
  g2500
  (
    n2535,
    n2152,
    n2507,
    n2511,
    n2184
  );


  nor
  g2501
  (
    n2517,
    n2134,
    n2121,
    n2137,
    n2183
  );


  xnor
  g2502
  (
    n2518,
    n2510,
    n2143,
    n2122,
    n2509
  );


  nor
  g2503
  (
    n2520,
    n2160,
    n2166,
    n2510,
    n2141
  );


  xnor
  g2504
  (
    n2525,
    n2154,
    n2148,
    n2157,
    n2145
  );


  nor
  g2505
  (
    n2516,
    n2138,
    n2165,
    n2512,
    n2508
  );


  not
  g2506
  (
    n2616,
    n2535
  );


  not
  g2507
  (
    n2582,
    n2531
  );


  buf
  g2508
  (
    n2545,
    n2522
  );


  not
  g2509
  (
    n2540,
    n2524
  );


  not
  g2510
  (
    n2585,
    n2522
  );


  buf
  g2511
  (
    n2548,
    n2521
  );


  not
  g2512
  (
    n2639,
    n2528
  );


  buf
  g2513
  (
    n2575,
    n2521
  );


  buf
  g2514
  (
    n2561,
    n2513
  );


  buf
  g2515
  (
    n2592,
    n2532
  );


  not
  g2516
  (
    n2635,
    n2515
  );


  buf
  g2517
  (
    n2539,
    n2534
  );


  not
  g2518
  (
    n2601,
    n660
  );


  not
  g2519
  (
    n2543,
    n2532
  );


  not
  g2520
  (
    n2593,
    n2520
  );


  not
  g2521
  (
    n2572,
    n2524
  );


  buf
  g2522
  (
    n2594,
    n662
  );


  buf
  g2523
  (
    n2620,
    n2518
  );


  not
  g2524
  (
    n2636,
    n2519
  );


  not
  g2525
  (
    n2608,
    n2521
  );


  not
  g2526
  (
    n2596,
    n2537
  );


  buf
  g2527
  (
    n2640,
    n2516
  );


  not
  g2528
  (
    n2588,
    n2527
  );


  buf
  g2529
  (
    n2604,
    n2536
  );


  buf
  g2530
  (
    n2621,
    n2496
  );


  buf
  g2531
  (
    n2549,
    n2532
  );


  buf
  g2532
  (
    n2562,
    n2516
  );


  not
  g2533
  (
    n2544,
    n2516
  );


  buf
  g2534
  (
    n2547,
    n659
  );


  buf
  g2535
  (
    n2614,
    n2537
  );


  not
  g2536
  (
    n2618,
    n2527
  );


  not
  g2537
  (
    KeyWire_0_52,
    n2525
  );


  buf
  g2538
  (
    n2587,
    n2518
  );


  not
  g2539
  (
    n2598,
    n2190
  );


  buf
  g2540
  (
    n2558,
    n2528
  );


  buf
  g2541
  (
    n2581,
    n2523
  );


  not
  g2542
  (
    n2609,
    n2525
  );


  not
  g2543
  (
    n2624,
    n2188
  );


  not
  g2544
  (
    n2566,
    n2529
  );


  not
  g2545
  (
    n2641,
    n2526
  );


  not
  g2546
  (
    n2637,
    n2515
  );


  buf
  g2547
  (
    n2571,
    n2522
  );


  buf
  g2548
  (
    n2597,
    n2519
  );


  not
  g2549
  (
    n2600,
    n661
  );


  not
  g2550
  (
    n2578,
    n2536
  );


  not
  g2551
  (
    n2634,
    n2535
  );


  buf
  g2552
  (
    n2573,
    n2514
  );


  buf
  g2553
  (
    n2615,
    n2531
  );


  not
  g2554
  (
    n2611,
    n2530
  );


  buf
  g2555
  (
    n2579,
    n2530
  );


  not
  g2556
  (
    n2546,
    n2520
  );


  buf
  g2557
  (
    n2550,
    n659
  );


  not
  g2558
  (
    n2542,
    n2526
  );


  not
  g2559
  (
    n2628,
    n2519
  );


  not
  g2560
  (
    n2602,
    n2514
  );


  not
  g2561
  (
    n2569,
    n2530
  );


  not
  g2562
  (
    n2580,
    n2531
  );


  not
  g2563
  (
    n2556,
    n2533
  );


  buf
  g2564
  (
    n2619,
    n2538
  );


  not
  g2565
  (
    n2627,
    n2533
  );


  not
  g2566
  (
    n2570,
    n660
  );


  not
  g2567
  (
    n2589,
    n2525
  );


  not
  g2568
  (
    n2554,
    n2516
  );


  buf
  g2569
  (
    n2563,
    n661
  );


  not
  g2570
  (
    n2590,
    n2513
  );


  not
  g2571
  (
    n2625,
    n2531
  );


  buf
  g2572
  (
    n2613,
    n2527
  );


  not
  g2573
  (
    n2583,
    n2513
  );


  not
  g2574
  (
    n2632,
    n2524
  );


  buf
  g2575
  (
    n2567,
    n2533
  );


  not
  g2576
  (
    n2552,
    n2514
  );


  not
  g2577
  (
    n2586,
    n2525
  );


  not
  g2578
  (
    n2577,
    n2528
  );


  buf
  g2579
  (
    n2617,
    n2536
  );


  not
  g2580
  (
    n2638,
    n2523
  );


  buf
  g2581
  (
    n2629,
    n2520
  );


  buf
  g2582
  (
    n2607,
    n2517
  );


  buf
  g2583
  (
    n2605,
    n2524
  );


  not
  g2584
  (
    n2553,
    n2520
  );


  buf
  g2585
  (
    n2630,
    n2538
  );


  buf
  g2586
  (
    n2557,
    n2518
  );


  not
  g2587
  (
    n2568,
    n2515
  );


  not
  g2588
  (
    n2574,
    n2536
  );


  buf
  g2589
  (
    n2584,
    n661
  );


  not
  g2590
  (
    n2560,
    n659
  );


  buf
  g2591
  (
    n2633,
    n2528
  );


  not
  g2592
  (
    n2622,
    n2499
  );


  not
  g2593
  (
    n2595,
    n2518
  );


  not
  g2594
  (
    n2606,
    n2534
  );


  not
  g2595
  (
    n2591,
    n2537
  );


  not
  g2596
  (
    n2551,
    n2497
  );


  buf
  g2597
  (
    n2559,
    n660
  );


  buf
  g2598
  (
    n2564,
    n2527
  );


  buf
  g2599
  (
    n2623,
    n2534
  );


  not
  g2600
  (
    n2642,
    n2532
  );


  buf
  g2601
  (
    n2555,
    n2523
  );


  not
  g2602
  (
    n2603,
    n661
  );


  xnor
  g2603
  (
    n2565,
    n2495,
    n2513,
    n2535,
    n2526
  );


  nor
  g2604
  (
    n2541,
    n2529,
    n2515,
    n2534,
    n660
  );


  nor
  g2605
  (
    n2610,
    n2535,
    n2538,
    n2533,
    n2529
  );


  and
  g2606
  (
    n2626,
    n2189,
    n2517,
    n2529,
    n2523
  );


  nor
  g2607
  (
    n2612,
    n2522,
    n2517,
    n2519,
    n2526
  );


  or
  g2608
  (
    n2599,
    n2537,
    n2517,
    n2514,
    n659
  );


  xor
  g2609
  (
    n2631,
    n2530,
    n2538,
    n2498,
    n2521
  );


  buf
  g2610
  (
    n2644,
    n2546
  );


  buf
  g2611
  (
    n2655,
    n2539
  );


  buf
  g2612
  (
    n2660,
    n2503
  );


  not
  g2613
  (
    n2662,
    n2502
  );


  nand
  g2614
  (
    n2647,
    n2196,
    n2546
  );


  xnor
  g2615
  (
    n2648,
    n2544,
    n2503
  );


  or
  g2616
  (
    n2658,
    n2542,
    n2539
  );


  nand
  g2617
  (
    n2657,
    n2547,
    n2548
  );


  or
  g2618
  (
    n2656,
    n2544,
    n2541
  );


  xor
  g2619
  (
    n2661,
    n2191,
    n2502
  );


  and
  g2620
  (
    n2646,
    n2540,
    n2192
  );


  nand
  g2621
  (
    n2653,
    n2547,
    n2501
  );


  xnor
  g2622
  (
    n2645,
    n2500,
    n2543
  );


  nor
  g2623
  (
    n2643,
    n2543,
    n2505
  );


  and
  g2624
  (
    n2650,
    n2548,
    n2504
  );


  xor
  g2625
  (
    KeyWire_0_26,
    n2194,
    n2545
  );


  and
  g2626
  (
    n2652,
    n2505,
    n2195
  );


  nor
  g2627
  (
    KeyWire_0_50,
    n2504,
    n2545
  );


  xnor
  g2628
  (
    n2649,
    n2542,
    n2541
  );


  or
  g2629
  (
    n2651,
    n2540,
    n2193
  );


  buf
  g2630
  (
    n2676,
    n2643
  );


  not
  g2631
  (
    n2663,
    n2650
  );


  not
  g2632
  (
    n2673,
    n2644
  );


  buf
  g2633
  (
    n2665,
    n2654
  );


  buf
  g2634
  (
    n2671,
    n2657
  );


  not
  g2635
  (
    n2672,
    n2651
  );


  not
  g2636
  (
    n2674,
    n2646
  );


  not
  g2637
  (
    n2667,
    n2645
  );


  not
  g2638
  (
    n2668,
    n2649
  );


  not
  g2639
  (
    n2678,
    n2652
  );


  buf
  g2640
  (
    n2675,
    n2658
  );


  buf
  g2641
  (
    n2666,
    n2648
  );


  buf
  g2642
  (
    n2670,
    n2653
  );


  not
  g2643
  (
    n2669,
    n2647
  );


  not
  g2644
  (
    n2677,
    n2655
  );


  buf
  g2645
  (
    n2664,
    n2656
  );


  and
  g2646
  (
    n2679,
    n2566,
    n2553,
    n2197,
    n2589
  );


  or
  g2647
  (
    n2688,
    n2668,
    n2556,
    n2198,
    n2664
  );


  or
  g2648
  (
    n2708,
    n2592,
    n2568,
    n2558,
    n2564
  );


  and
  g2649
  (
    n2701,
    n2604,
    n2669,
    n2602,
    n2567
  );


  nor
  g2650
  (
    n2690,
    n2562,
    n2663,
    n2549,
    n2585
  );


  xor
  g2651
  (
    n2721,
    n2675,
    n2599,
    n2605,
    n2596
  );


  nor
  g2652
  (
    n2713,
    n2593,
    n2602,
    n2576,
    n2561
  );


  nand
  g2653
  (
    n2685,
    n2669,
    n2563,
    n2663,
    n2667
  );


  and
  g2654
  (
    n2703,
    n2670,
    n2566,
    n2671,
    n2587
  );


  xnor
  g2655
  (
    n2689,
    n2578,
    n2598,
    n2665,
    n2563
  );


  and
  g2656
  (
    n2710,
    n2665,
    n2577,
    n2586,
    n2591
  );


  xor
  g2657
  (
    n2730,
    n2575,
    n2554,
    n2594,
    n2669
  );


  xor
  g2658
  (
    n2682,
    n2591,
    n2572,
    n2560,
    n2675
  );


  or
  g2659
  (
    n2694,
    n2603,
    n2674,
    n2672,
    n2552
  );


  and
  g2660
  (
    n2686,
    n2606,
    n2664,
    n2581,
    n2573
  );


  xnor
  g2661
  (
    n2704,
    n2555,
    n2665,
    n2603,
    n2553
  );


  xor
  g2662
  (
    n2715,
    n2666,
    n2597,
    n2570,
    n2601
  );


  nand
  g2663
  (
    n2684,
    n2666,
    n2598,
    n2557,
    n2600
  );


  or
  g2664
  (
    n2705,
    n2674,
    n2560,
    n2592,
    n2671
  );


  and
  g2665
  (
    n2706,
    n2586,
    n2577,
    n2589,
    n2598
  );


  nor
  g2666
  (
    n2725,
    n2606,
    n2557,
    n2671,
    n2601
  );


  or
  g2667
  (
    n2712,
    n2674,
    n2670,
    n2673,
    n2667
  );


  xnor
  g2668
  (
    n2724,
    n2590,
    n2580,
    n2569,
    n2203
  );


  nand
  g2669
  (
    n2709,
    n2600,
    n2584,
    n2663,
    n2552
  );


  and
  g2670
  (
    n2680,
    n2674,
    n2595,
    n2673,
    n2580
  );


  xor
  g2671
  (
    n2728,
    n2596,
    n2585,
    n2582,
    n2565
  );


  nor
  g2672
  (
    n2700,
    n2572,
    n2605,
    n2670,
    n2672
  );


  nor
  g2673
  (
    n2702,
    n2604,
    n2665,
    n2201,
    n2667
  );


  xnor
  g2674
  (
    n2714,
    n2595,
    n2202,
    n2550,
    n2574
  );


  xor
  g2675
  (
    n2719,
    n2604,
    n2663,
    n2596,
    n2602
  );


  and
  g2676
  (
    n2697,
    n2559,
    n2594,
    n2588,
    n2554
  );


  xor
  g2677
  (
    n2681,
    n2568,
    n2675,
    n2605,
    n2583
  );


  xor
  g2678
  (
    n2723,
    n2668,
    n2550,
    n2673,
    n2561
  );


  and
  g2679
  (
    n2726,
    n2606,
    n2668,
    n2596,
    n2205
  );


  and
  g2680
  (
    n2711,
    n2583,
    n2559,
    n2666,
    n2575
  );


  and
  g2681
  (
    n2727,
    n2594,
    n2551,
    n2565,
    n2571
  );


  xor
  g2682
  (
    n2699,
    n2206,
    n2562,
    n2582,
    n2558
  );


  or
  g2683
  (
    n2695,
    n2664,
    n2594,
    n2579,
    n2567
  );


  nor
  g2684
  (
    n2683,
    n2601,
    n2564,
    n2555,
    n2599
  );


  xnor
  g2685
  (
    n2720,
    n2570,
    n2581,
    n2601,
    n2590
  );


  xor
  g2686
  (
    n2692,
    n2603,
    n2593,
    n2606
  );


  xor
  g2687
  (
    n2716,
    n2600,
    n2668,
    n2593,
    n2671
  );


  xor
  g2688
  (
    n2691,
    n2600,
    n2669,
    n2673,
    n2672
  );


  or
  g2689
  (
    n2698,
    n2597,
    n2207,
    n2670,
    n2602
  );


  xnor
  g2690
  (
    n2696,
    n2549,
    n2604,
    n2599,
    n2598
  );


  xnor
  g2691
  (
    n2722,
    n2576,
    n2595,
    n2551,
    n2584
  );


  nor
  g2692
  (
    n2718,
    n2587,
    n2556,
    n2599,
    n2603
  );


  nor
  g2693
  (
    n2717,
    n2574,
    n2605,
    n2672,
    n2578
  );


  or
  g2694
  (
    n2729,
    n2597,
    n2204,
    n2595,
    n2208
  );


  xnor
  g2695
  (
    n2687,
    n2666,
    n2200,
    n2569,
    n2664
  );


  xor
  g2696
  (
    n2707,
    n2579,
    n2199,
    n2573,
    n2667
  );


  xor
  g2697
  (
    n2693,
    n2588,
    n2571,
    n2675,
    n2597
  );


  or
  g2698
  (
    n2758,
    n2626,
    n2628,
    n2622,
    n2619
  );


  or
  g2699
  (
    n2773,
    n2616,
    n2636,
    n2721,
    n2705
  );


  xnor
  g2700
  (
    n2766,
    n2699,
    n2621,
    n2224,
    n2640
  );


  or
  g2701
  (
    n2779,
    n2679,
    n2730,
    n2622,
    n2617
  );


  xor
  g2702
  (
    n2749,
    n2689,
    n2684,
    n2726,
    n2640
  );


  and
  g2703
  (
    n2739,
    n2718,
    n2630,
    n2625,
    n2680
  );


  xor
  g2704
  (
    n2753,
    n2632,
    n2704,
    n2696,
    n2694
  );


  and
  g2705
  (
    n2761,
    n2724,
    n2661,
    n2213,
    n2710
  );


  nor
  g2706
  (
    n2751,
    n2631,
    n2717,
    n2635,
    n2609
  );


  nor
  g2707
  (
    n2744,
    n2702,
    n2728,
    n2613,
    n2703
  );


  xor
  g2708
  (
    n2765,
    n2700,
    n2637,
    n2628,
    n2682
  );


  nand
  g2709
  (
    n2757,
    n2720,
    n2688,
    n2714,
    n2618
  );


  nand
  g2710
  (
    n2778,
    n2218,
    n2611,
    n2636,
    n2708
  );


  xor
  g2711
  (
    n2740,
    n2640,
    n2612,
    n2615,
    n2620
  );


  xor
  g2712
  (
    n2769,
    n2613,
    n2633,
    n2627,
    n2614
  );


  xnor
  g2713
  (
    n2776,
    n2638,
    n2221,
    n2685,
    n2626
  );


  and
  g2714
  (
    n2762,
    n2729,
    n2623,
    n2719,
    n2707
  );


  xor
  g2715
  (
    n2748,
    n2616,
    n2615,
    n2636,
    n2706
  );


  xnor
  g2716
  (
    n2756,
    n2608,
    n2691,
    n2614,
    n2615
  );


  and
  g2717
  (
    n2736,
    n2690,
    n2722,
    n2609,
    n2623
  );


  xor
  g2718
  (
    n2767,
    n2622,
    n2634,
    n2614,
    n2716
  );


  xor
  g2719
  (
    n2770,
    n2629,
    n2624,
    n2610
  );


  nor
  g2720
  (
    n2764,
    n2635,
    n2659,
    n2618,
    n2632
  );


  xnor
  g2721
  (
    n2741,
    n2637,
    n2215,
    n2621,
    n2611
  );


  xnor
  g2722
  (
    n2782,
    n2609,
    n2612,
    n2607,
    n2619
  );


  nor
  g2723
  (
    n2781,
    n2629,
    n2609,
    n2695,
    n2608
  );


  xor
  g2724
  (
    n2760,
    n2662,
    n2610,
    n2634,
    n2620
  );


  nand
  g2725
  (
    n2752,
    n2628,
    n2686,
    n2219,
    n2216
  );


  and
  g2726
  (
    n2745,
    n2217,
    n2627,
    n2607,
    n2626
  );


  nand
  g2727
  (
    n2777,
    n2608,
    n2621,
    n2626,
    n2616
  );


  nand
  g2728
  (
    n2774,
    n2222,
    n2615,
    n2698,
    n2210
  );


  or
  g2729
  (
    n2755,
    n2693,
    n2638,
    n2683,
    n2620
  );


  and
  g2730
  (
    n2759,
    n2629,
    n2636,
    n2712,
    n2623
  );


  and
  g2731
  (
    n2731,
    n2624,
    n2607,
    n2621,
    n2692
  );


  or
  g2732
  (
    n2754,
    n2612,
    n2633,
    n2723,
    n2613
  );


  xor
  g2733
  (
    n2737,
    n2638,
    n2607,
    n2614,
    n2637
  );


  xor
  g2734
  (
    n2768,
    n2211,
    n2610,
    n2611,
    n2629
  );


  and
  g2735
  (
    n2775,
    n2639,
    n2634,
    n2617,
    n2640
  );


  or
  g2736
  (
    n2742,
    n2613,
    n2209,
    n2632,
    n2610
  );


  xor
  g2737
  (
    n2733,
    n2625,
    n2624,
    n2681,
    n2715
  );


  or
  g2738
  (
    n2746,
    n2639,
    n2616,
    n2617,
    n2611
  );


  nand
  g2739
  (
    n2734,
    n2214,
    n2638,
    n2637,
    n2625
  );


  nor
  g2740
  (
    n2747,
    n2633,
    n2625,
    n2639,
    n2619
  );


  or
  g2741
  (
    n2743,
    n2701,
    n2631,
    n2623,
    n2630
  );


  xnor
  g2742
  (
    n2732,
    n2632,
    n2634,
    n2608,
    n2633
  );


  xor
  g2743
  (
    n2771,
    n2618,
    n2631,
    n2630,
    n2628
  );


  nand
  g2744
  (
    n2750,
    n2631,
    n2630,
    n2639,
    n2617
  );


  nor
  g2745
  (
    n2772,
    n2612,
    n2709,
    n2727,
    n2619
  );


  and
  g2746
  (
    n2738,
    n2220,
    n2725,
    n2622,
    n2223
  );


  nand
  g2747
  (
    n2763,
    n2713,
    n2635,
    n2627,
    n2618
  );


  xor
  g2748
  (
    n2780,
    n2711,
    n2627,
    n2212,
    n2620
  );


  and
  g2749
  (
    n2735,
    n2687,
    n2635,
    n2660,
    n2697
  );


  not
  g2750
  (
    n2789,
    n2733
  );


  buf
  g2751
  (
    n2784,
    n2731
  );


  buf
  g2752
  (
    n2787,
    n2731
  );


  not
  g2753
  (
    n2786,
    n2734
  );


  not
  g2754
  (
    n2788,
    n2733
  );


  not
  g2755
  (
    n2785,
    n2225
  );


  buf
  g2756
  (
    n2783,
    n2732
  );


  and
  g2757
  (
    n2792,
    n2788,
    n2786,
    n2783,
    n2787
  );


  nor
  g2758
  (
    n2799,
    n2249,
    n2238,
    n2786
  );


  nor
  g2759
  (
    n2793,
    n2246,
    n2230,
    n2789,
    n2229
  );


  or
  g2760
  (
    n2794,
    n2785,
    n2784,
    n2231,
    n2227
  );


  xor
  g2761
  (
    n2798,
    n2783,
    n2783,
    n2785,
    n2784
  );


  xnor
  g2762
  (
    n2796,
    n2234,
    n2789,
    n2787
  );


  nor
  g2763
  (
    n2804,
    n2784,
    n2678,
    n2785
  );


  or
  g2764
  (
    n2791,
    n2243,
    n2676,
    n2245,
    n2786
  );


  xor
  g2765
  (
    n2803,
    n2248,
    n2250,
    n2233,
    n2788
  );


  nor
  g2766
  (
    n2797,
    n2226,
    n2783,
    n2785,
    n2677
  );


  xnor
  g2767
  (
    n2800,
    n2677,
    n2247,
    n2676,
    n2239
  );


  nor
  g2768
  (
    n2801,
    n2232,
    n2677,
    n2244,
    n2242
  );


  xnor
  g2769
  (
    n2795,
    n2676,
    n2240,
    n2241,
    n2228
  );


  or
  g2770
  (
    n2790,
    n2235,
    n2237,
    n2678,
    n2788
  );


  xnor
  g2771
  (
    n2805,
    n2678,
    n2784,
    n2677,
    n2788
  );


  and
  g2772
  (
    n2802,
    n2236,
    n2676,
    n2787,
    n2789
  );


  and
  g2773
  (
    n2809,
    n2260,
    n2253,
    n2803,
    n2805
  );


  nor
  g2774
  (
    n2810,
    n2737,
    n2259,
    n2735,
    n2252
  );


  and
  g2775
  (
    n2806,
    n2254,
    n2736,
    n2258,
    n2735
  );


  nor
  g2776
  (
    n2812,
    n2255,
    n2801,
    n2737,
    n2256
  );


  xor
  g2777
  (
    n2811,
    n2262,
    n2798,
    n2734,
    n2736
  );


  or
  g2778
  (
    n2807,
    n2802,
    n2266,
    n2799,
    n2800
  );


  nor
  g2779
  (
    n2813,
    n2267,
    n2251,
    n2257,
    n2804
  );


  nand
  g2780
  (
    n2808,
    n2265,
    n2263,
    n2264,
    n2261
  );


  xor
  g2781
  (
    n2820,
    n2808,
    n2750,
    n2811,
    n2758
  );


  or
  g2782
  (
    n2824,
    n2808,
    n2806,
    n2770,
    n2274
  );


  xor
  g2783
  (
    n2815,
    n2743,
    n2762,
    n2761
  );


  nor
  g2784
  (
    n2828,
    n2781,
    n2743,
    n2752,
    n2751
  );


  and
  g2785
  (
    n2832,
    n2813,
    n2773,
    n2753,
    n2755
  );


  nor
  g2786
  (
    n2835,
    n2769,
    n2276,
    n2763,
    n2776
  );


  and
  g2787
  (
    n2842,
    n2746,
    n2745,
    n2754,
    n2772
  );


  or
  g2788
  (
    n2823,
    n2809,
    n2764,
    n2738,
    n2756
  );


  nand
  g2789
  (
    n2841,
    n2760,
    n2808,
    n2809,
    n2780
  );


  nor
  g2790
  (
    n2843,
    n2754,
    n2748,
    n2272,
    n2757
  );


  nor
  g2791
  (
    n2822,
    n2780,
    n2773,
    n2807,
    n2755
  );


  or
  g2792
  (
    n2821,
    n2769,
    n2759,
    n2812,
    n2771
  );


  xor
  g2793
  (
    n2827,
    n2747,
    n2739,
    n2809,
    n2751
  );


  xor
  g2794
  (
    n2834,
    n2812,
    n2760,
    n2749,
    n2741
  );


  nand
  g2795
  (
    n2829,
    n2756,
    n2745,
    n2270,
    n2810
  );


  or
  g2796
  (
    n2845,
    n2766,
    n2752,
    n2777,
    n2763
  );


  nand
  g2797
  (
    n2825,
    n2268,
    n2740,
    n2807,
    n2774
  );


  xor
  g2798
  (
    n2819,
    n2765,
    n2269,
    n2759,
    n2774
  );


  nor
  g2799
  (
    n2837,
    n2810,
    n2271,
    n2806
  );


  and
  g2800
  (
    n2838,
    n2750,
    n2765,
    n2771,
    n2761
  );


  nor
  g2801
  (
    n2836,
    n2753,
    n2767,
    n2740,
    n2810
  );


  xnor
  g2802
  (
    n2833,
    n2808,
    n2778,
    n2275,
    n2809
  );


  xor
  g2803
  (
    n2826,
    n2775,
    n2273,
    n2744,
    n2768
  );


  and
  g2804
  (
    n2831,
    n2757,
    n2746,
    n2813
  );


  xnor
  g2805
  (
    n2830,
    n2813,
    n2811,
    n2739,
    n2747
  );


  nor
  g2806
  (
    n2814,
    n2811,
    n2778,
    n2810,
    n2779
  );


  nand
  g2807
  (
    KeyWire_0_45,
    n2807,
    n2806,
    n2811,
    n2779
  );


  xor
  g2808
  (
    n2816,
    n2768,
    n2812,
    n2770
  );


  or
  g2809
  (
    n2844,
    n2807,
    n2766,
    n2775,
    n2776
  );


  and
  g2810
  (
    KeyWire_0_23,
    n2742,
    n2749,
    n2777,
    n2767
  );


  nand
  g2811
  (
    n2818,
    n2764,
    n2772,
    n2738,
    n2744
  );


  and
  g2812
  (
    n2840,
    n2758,
    n2741,
    n2742,
    n2748
  );


  not
  g2813
  (
    n2867,
    n2815
  );


  not
  g2814
  (
    n2847,
    n2825
  );


  not
  g2815
  (
    n2874,
    n2829
  );


  not
  g2816
  (
    n2848,
    n2822
  );


  not
  g2817
  (
    n2861,
    n2826
  );


  buf
  g2818
  (
    n2864,
    n2827
  );


  buf
  g2819
  (
    n2872,
    n2818
  );


  not
  g2820
  (
    n2865,
    n2816
  );


  not
  g2821
  (
    n2855,
    n2821
  );


  buf
  g2822
  (
    n2851,
    n2822
  );


  buf
  g2823
  (
    n2870,
    n2824
  );


  buf
  g2824
  (
    n2873,
    n2826
  );


  buf
  g2825
  (
    n2857,
    n2818
  );


  buf
  g2826
  (
    n2877,
    n2829
  );


  not
  g2827
  (
    n2850,
    n2828
  );


  buf
  g2828
  (
    n2852,
    n2827
  );


  buf
  g2829
  (
    n2869,
    n2825
  );


  buf
  g2830
  (
    n2854,
    n2824
  );


  buf
  g2831
  (
    n2863,
    n2789
  );


  not
  g2832
  (
    n2875,
    n2820
  );


  not
  g2833
  (
    n2860,
    n2815
  );


  buf
  g2834
  (
    n2856,
    n2830
  );


  buf
  g2835
  (
    n2859,
    n2821
  );


  buf
  g2836
  (
    n2853,
    n2814
  );


  buf
  g2837
  (
    n2868,
    n2820
  );


  not
  g2838
  (
    n2876,
    n2814
  );


  buf
  g2839
  (
    n2878,
    n2830
  );


  not
  g2840
  (
    n2871,
    n2823
  );


  buf
  g2841
  (
    n2866,
    n2819
  );


  not
  g2842
  (
    n2858,
    n2823
  );


  not
  g2843
  (
    n2849,
    n2817
  );


  buf
  g2844
  (
    n2862,
    n2817
  );


  xor
  g2845
  (
    n2846,
    n2816,
    n2277
  );


  and
  g2846
  (
    n2879,
    n2828,
    n2819
  );


  nand
  g2847
  (
    n2883,
    n664,
    n666
  );


  nand
  g2848
  (
    n2894,
    n2847,
    n2846,
    n662,
    n2864
  );


  xnor
  g2849
  (
    n2885,
    n2855,
    n2851,
    n667,
    n2875
  );


  or
  g2850
  (
    n2880,
    n667,
    n2852,
    n663,
    n665
  );


  or
  g2851
  (
    n2887,
    n2869,
    n665,
    n2866,
    n2849
  );


  xor
  g2852
  (
    n2884,
    n2854,
    n663,
    n662,
    n664
  );


  xor
  g2853
  (
    n2881,
    n664,
    n2873,
    n2858,
    n667
  );


  and
  g2854
  (
    n2886,
    n2865,
    n2874,
    n2856,
    n663
  );


  nor
  g2855
  (
    n2891,
    n2850,
    n666,
    n2867,
    n2862
  );


  nor
  g2856
  (
    n2890,
    n2872,
    n2278,
    n2860,
    n2868
  );


  or
  g2857
  (
    n2882,
    n664,
    n663,
    n2861,
    n2832
  );


  xnor
  g2858
  (
    n2888,
    n662,
    n666,
    n2859
  );


  or
  g2859
  (
    n2893,
    n2870,
    n665,
    n667,
    n2857
  );


  xnor
  g2860
  (
    n2889,
    n2831,
    n2832,
    n665,
    n2853
  );


  xor
  g2861
  (
    n2892,
    n2871,
    n2848,
    n2863,
    n2831
  );


  nand
  g2862
  (
    n2896,
    n2890,
    n2839,
    n2833,
    n2834
  );


  nor
  g2863
  (
    n2899,
    n2893,
    n2836,
    n2892,
    n2839
  );


  xor
  g2864
  (
    n2897,
    n2836,
    n2833,
    n2834,
    n2835
  );


  or
  g2865
  (
    n2895,
    n2840,
    n2837,
    n2838
  );


  nand
  g2866
  (
    n2898,
    n2835,
    n2837,
    n2891,
    n2894
  );


  xor
  g2867
  (
    n2912,
    n2329,
    n2895,
    n2294,
    n2297
  );


  nand
  g2868
  (
    n2909,
    n2899,
    n2898,
    n2321,
    n2841
  );


  xor
  g2869
  (
    n2908,
    n2896,
    n2842,
    n2322,
    n2326
  );


  xnor
  g2870
  (
    n2910,
    n2304,
    n2316,
    n2330,
    n2290
  );


  nand
  g2871
  (
    n2916,
    n2898,
    n2840,
    n2314,
    n2301
  );


  or
  g2872
  (
    n2906,
    n2897,
    n2302,
    n2289,
    n2312
  );


  xor
  g2873
  (
    n2917,
    n2298,
    n2279,
    n2318,
    n2323
  );


  or
  g2874
  (
    n2919,
    n2306,
    n2899,
    n2315,
    n2305
  );


  xor
  g2875
  (
    n2913,
    n2281,
    n2328,
    n2309,
    n2895
  );


  or
  g2876
  (
    n2907,
    n2283,
    n2319,
    n2300,
    n2286
  );


  nor
  g2877
  (
    n2914,
    n2282,
    n2299,
    n2296,
    n2325
  );


  xnor
  g2878
  (
    n2903,
    n2303,
    n2293,
    n2897,
    n2334
  );


  nand
  g2879
  (
    n2900,
    n2896,
    n2331,
    n2841,
    n2899
  );


  xnor
  g2880
  (
    n2918,
    n2327,
    n2311,
    n2295,
    n2333
  );


  nand
  g2881
  (
    n2905,
    n2320,
    n2895,
    n2307,
    n2288
  );


  xor
  g2882
  (
    n2915,
    n2899,
    n2285,
    n2313,
    n2280
  );


  nand
  g2883
  (
    n2904,
    n2332,
    n2291,
    n2324,
    n2898
  );


  nand
  g2884
  (
    n2901,
    n2898,
    n2284,
    n2308,
    n2310
  );


  nand
  g2885
  (
    n2911,
    n2896,
    n2287,
    n2292,
    n2895
  );


  xor
  g2886
  (
    n2902,
    n2317,
    n2897,
    n2896
  );


  buf
  g2887
  (
    n2921,
    n2900
  );


  not
  g2888
  (
    n2923,
    n2877
  );


  not
  g2889
  (
    n2922,
    n2876
  );


  nand
  g2890
  (
    n2924,
    n2335,
    n2902,
    n2879
  );


  xnor
  g2891
  (
    n2920,
    n2878,
    n2901,
    n2902
  );


  nor
  g2892
  (
    n2941,
    n2642,
    n2338,
    n2068
  );


  or
  g2893
  (
    n2940,
    n2342,
    n2920,
    n2068
  );


  xor
  g2894
  (
    n2937,
    n160,
    n2845,
    n2920
  );


  or
  g2895
  (
    n2925,
    n2341,
    n2921,
    n2920
  );


  xor
  g2896
  (
    n2935,
    n160,
    n2068,
    n2067
  );


  xor
  g2897
  (
    n2943,
    n2921,
    n2922,
    n2066
  );


  or
  g2898
  (
    n2932,
    n2339,
    n2781,
    n2344
  );


  or
  g2899
  (
    n2928,
    n2922,
    n2845,
    n2782
  );


  xnor
  g2900
  (
    n2942,
    n2782,
    n2067,
    n2642,
    n2340
  );


  nor
  g2901
  (
    n2939,
    n2641,
    n2641,
    n2922,
    n2343
  );


  and
  g2902
  (
    n2944,
    n2922,
    n2781,
    n2065,
    n2921
  );


  and
  g2903
  (
    n2930,
    n160,
    n2066,
    n2920
  );


  nand
  g2904
  (
    n2929,
    n159,
    n2923,
    n160,
    n2066
  );


  and
  g2905
  (
    n2931,
    n2924,
    n2924,
    n2781,
    n2782
  );


  xnor
  g2906
  (
    n2936,
    n2336,
    n2844,
    n2923
  );


  xnor
  g2907
  (
    n2933,
    n2068,
    n2843,
    n2065
  );


  xnor
  g2908
  (
    n2934,
    n2924,
    n2842,
    n2641,
    n2923
  );


  nor
  g2909
  (
    n2926,
    n2065,
    n2921,
    n2843,
    n2924
  );


  nor
  g2910
  (
    n2927,
    n2641,
    n2844,
    n2067,
    n2782
  );


  xor
  g2911
  (
    n2938,
    n2067,
    n2337,
    n2642
  );


  buf
  g2912
  (
    n2948,
    n2935
  );


  buf
  g2913
  (
    n2952,
    n2930
  );


  not
  g2914
  (
    n2954,
    n2932
  );


  buf
  g2915
  (
    n2950,
    n2936
  );


  not
  g2916
  (
    n2947,
    n2931
  );


  not
  g2917
  (
    n2953,
    n2927
  );


  and
  g2918
  (
    n2946,
    n2935,
    n2929
  );


  nand
  g2919
  (
    n2958,
    n2930,
    n2934,
    n2925
  );


  xor
  g2920
  (
    n2957,
    n2932,
    n2931,
    n2928,
    n2929
  );


  nor
  g2921
  (
    n2951,
    n2933,
    n2936,
    n2931,
    n2932
  );


  and
  g2922
  (
    n2949,
    n2931,
    n2933,
    n2934
  );


  or
  g2923
  (
    n2945,
    n2933,
    n2926
  );


  xnor
  g2924
  (
    n2956,
    n2932,
    n2935,
    n2925
  );


  or
  g2925
  (
    n2955,
    n2928,
    n2936,
    n2927
  );


  and
  g2926
  (
    n2961,
    n2909,
    n2913,
    n2903,
    n2919
  );


  xnor
  g2927
  (
    n2963,
    n2904,
    n2945,
    n2905,
    n2907
  );


  xor
  g2928
  (
    n2959,
    n2914,
    n2904,
    n2937,
    n2918
  );


  xnor
  g2929
  (
    n2970,
    n2948,
    n2918,
    n2946,
    n2917
  );


  or
  g2930
  (
    n2966,
    n2954,
    n2911,
    n2956,
    n2919
  );


  nor
  g2931
  (
    n2968,
    n2909,
    n2905,
    n2908
  );


  xor
  g2932
  (
    n2960,
    n2916,
    n2953,
    n2906,
    n2911
  );


  nand
  g2933
  (
    n2965,
    n2913,
    n2951,
    n2910,
    n2952
  );


  and
  g2934
  (
    n2969,
    n2903,
    n2912,
    n2937,
    n2949
  );


  xor
  g2935
  (
    n2967,
    n2950,
    n2947,
    n2912,
    n2907
  );


  and
  g2936
  (
    n2962,
    n2910,
    n2915,
    n2916,
    n2955
  );


  xor
  g2937
  (
    n2964,
    n2914,
    n2915,
    n2906,
    n2917
  );


  xnor
  g2938
  (
    n2972,
    n2969,
    n2938,
    n2937
  );


  or
  g2939
  (
    n2971,
    n2937,
    n2970,
    n2938
  );


  or
  g2940
  (
    n2979,
    n2971,
    n2941,
    n2939
  );


  and
  g2941
  (
    n2977,
    n2972,
    n2939,
    n2942,
    n2971
  );


  nand
  g2942
  (
    n2975,
    n2944,
    n2971,
    n2972,
    n2940
  );


  nor
  g2943
  (
    n2973,
    n2939,
    n2942,
    n2944
  );


  and
  g2944
  (
    n2974,
    n2972,
    n2940,
    n2941,
    n2942
  );


  or
  g2945
  (
    n2976,
    n2972,
    n2939,
    n2943
  );


  and
  g2946
  (
    n2978,
    n2941,
    n2944,
    n2942,
    n2940
  );


  or
  g2947
  (
    n2980,
    n2971,
    n2940,
    n2943
  );


  xnor
  g2948
  (
    KeyWire_0_16,
    n2978,
    n2977,
    n2425,
    n2390
  );


  xnor
  g2949
  (
    n2997,
    n2975,
    n2973,
    n2957,
    n2958
  );


  and
  g2950
  (
    n3008,
    n2980,
    n2363,
    n2979,
    n2391
  );


  xor
  g2951
  (
    n2999,
    n2351,
    n2977,
    n2411,
    n2976
  );


  xnor
  g2952
  (
    n3011,
    n2423,
    n2422,
    n2980,
    n2978
  );


  nor
  g2953
  (
    n2982,
    n2413,
    n2379,
    n2438,
    n2360
  );


  or
  g2954
  (
    n3001,
    n2358,
    n2979,
    n2435,
    n2978
  );


  nand
  g2955
  (
    n2989,
    n2402,
    n2398,
    n2359,
    n2389
  );


  nor
  g2956
  (
    n2984,
    n2978,
    n2419,
    n2433,
    n2349
  );


  or
  g2957
  (
    n3003,
    n2406,
    n2980,
    n2421
  );


  nand
  g2958
  (
    n3000,
    n2353,
    n2408,
    n2405,
    n2977
  );


  nor
  g2959
  (
    n3004,
    n2975,
    n2373,
    n2394,
    n2385
  );


  xnor
  g2960
  (
    KeyWire_0_44,
    n2375,
    n2361,
    n2410,
    n2377
  );


  xnor
  g2961
  (
    n2993,
    n2381,
    n2365,
    n2437,
    n2973
  );


  nor
  g2962
  (
    n3009,
    n2370,
    n2362,
    n2357,
    n2369
  );


  nand
  g2963
  (
    n2992,
    n2388,
    n2974,
    n2367,
    n2348
  );


  nand
  g2964
  (
    n2985,
    n2436,
    n2975,
    n2417,
    n2976
  );


  nor
  g2965
  (
    n2996,
    n2430,
    n2976,
    n2974,
    n2354
  );


  or
  g2966
  (
    n2991,
    n2364,
    n2979,
    n2401,
    n2352
  );


  nor
  g2967
  (
    n3005,
    n2345,
    n2384,
    n2979,
    n2431
  );


  nor
  g2968
  (
    n2988,
    n2386,
    n2371,
    n2397,
    n2409
  );


  xor
  g2969
  (
    n3010,
    n2355,
    n2974,
    n2382,
    n2374
  );


  xnor
  g2970
  (
    n3007,
    n2347,
    n2387,
    n2372,
    n2350
  );


  and
  g2971
  (
    n2983,
    n2396,
    n2976,
    n2393,
    n2429
  );


  nor
  g2972
  (
    n2994,
    n2412,
    n2376,
    n2399,
    n2415
  );


  nand
  g2973
  (
    n3006,
    n2427,
    n2346,
    n2426,
    n2974
  );


  or
  g2974
  (
    n2998,
    n2395,
    n2356,
    n2977,
    n2424
  );


  and
  g2975
  (
    n3002,
    n2432,
    n2973,
    n2380,
    n2392
  );


  nor
  g2976
  (
    n2990,
    n2975,
    n2407,
    n2428,
    n2416
  );


  or
  g2977
  (
    n2986,
    n2368,
    n2973,
    n2434,
    n2400
  );


  nor
  g2978
  (
    n2995,
    n2420,
    n2418,
    n2383,
    n2366
  );


  xor
  g2979
  (
    n2987,
    n2378,
    n2403,
    n2414,
    n2404
  );


  xnor
  g2980
  (
    n3022,
    n2449,
    n2987,
    n2981,
    n2470
  );


  nand
  g2981
  (
    n3023,
    n2986,
    n2445,
    n2992,
    n2467
  );


  or
  g2982
  (
    n3015,
    n3005,
    n2455,
    n2458,
    n2452
  );


  nor
  g2983
  (
    n3026,
    n2453,
    n3004,
    n2469,
    n3010
  );


  nand
  g2984
  (
    n3013,
    n2998,
    n2444,
    n2991,
    n2446
  );


  nor
  g2985
  (
    n3020,
    n3002,
    n2448,
    n3003,
    n2440
  );


  xor
  g2986
  (
    n3019,
    n2464,
    n2463,
    n3009,
    n2442
  );


  or
  g2987
  (
    n3028,
    n2995,
    n2460,
    n2441,
    n2450
  );


  nor
  g2988
  (
    KeyWire_0_2,
    n2468,
    n2451,
    n2999,
    n3012
  );


  nor
  g2989
  (
    n3024,
    n3001,
    n3006,
    n2990,
    n2456
  );


  xor
  g2990
  (
    n3016,
    n2462,
    n2454,
    n2985,
    n2996
  );


  nor
  g2991
  (
    n3027,
    n2457,
    n2439,
    n2994,
    n2466
  );


  or
  g2992
  (
    n3025,
    n2993,
    n2461,
    n3011,
    n2989
  );


  or
  g2993
  (
    n3018,
    n3000,
    n2982,
    n2459,
    n2997
  );


  nor
  g2994
  (
    n3017,
    n3007,
    n2447,
    n2983,
    n2443
  );


  nor
  g2995
  (
    n3014,
    n2988,
    n2984,
    n3008,
    n2465
  );


  nand
  g2996
  (
    n3030,
    n3019,
    n3027,
    n3013,
    n3023
  );


  xor
  g2997
  (
    n3031,
    n3026,
    n3014,
    n3016,
    n3020
  );


  or
  g2998
  (
    n3032,
    n3017,
    n3015,
    n3021,
    n3022
  );


  xnor
  g2999
  (
    n3029,
    n3025,
    n3018,
    n3028,
    n3024
  );


  xor
  KeyGate_0_0
  (
    n1196,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n399,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n3021,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1602,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n203,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n2153,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1238,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n362,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1893,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1285,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n271,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n328,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n604,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n2382,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1178,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n2014,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n3012,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1866,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n49,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n234,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1336,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n2187,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1250,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n2817,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n867,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n82,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n2659,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1131,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n906,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n560,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n609,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n2203,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n1622,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n987,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n172,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n231,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n1566,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n575,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n1772,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n1886,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n1262,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n1782,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n72,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n2506,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n2981,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n2839,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n304,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n1838,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n1640,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n936,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n2654,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n1301,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n2576,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n2478,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n361,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n175,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n1010,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n869,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n2272,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n2299,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n1008,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n1707,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n2117,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n1572,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

