

module Stat_489_535
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n508,
  n492,
  n495,
  n490,
  n489,
  n496,
  n510,
  n507,
  n503,
  n491,
  n504,
  n514,
  n497,
  n505,
  n513,
  n494,
  n506,
  n500,
  n502,
  n512,
  n487,
  n509,
  n499,
  n498,
  n488,
  n501,
  n493,
  n511,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;
  output n508;output n492;output n495;output n490;output n489;output n496;output n510;output n507;output n503;output n491;output n504;output n514;output n497;output n505;output n513;output n494;output n506;output n500;output n502;output n512;output n487;output n509;output n499;output n498;output n488;output n501;output n493;output n511;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n97,
    n23
  );


  buf
  g1
  (
    n101,
    n5
  );


  not
  g2
  (
    n50,
    n18
  );


  buf
  g3
  (
    n72,
    n5
  );


  buf
  g4
  (
    n26,
    n6
  );


  not
  g5
  (
    n34,
    n24
  );


  not
  g6
  (
    n64,
    n25
  );


  buf
  g7
  (
    n122,
    n14
  );


  not
  g8
  (
    n56,
    n9
  );


  not
  g9
  (
    n27,
    n23
  );


  not
  g10
  (
    n109,
    n16
  );


  buf
  g11
  (
    n114,
    n3
  );


  not
  g12
  (
    n108,
    n5
  );


  buf
  g13
  (
    n118,
    n16
  );


  buf
  g14
  (
    n115,
    n1
  );


  not
  g15
  (
    n43,
    n12
  );


  buf
  g16
  (
    n52,
    n10
  );


  not
  g17
  (
    n57,
    n22
  );


  not
  g18
  (
    n41,
    n14
  );


  not
  g19
  (
    n91,
    n14
  );


  buf
  g20
  (
    n71,
    n7
  );


  buf
  g21
  (
    n48,
    n9
  );


  not
  g22
  (
    n106,
    n8
  );


  not
  g23
  (
    n86,
    n25
  );


  buf
  g24
  (
    n38,
    n21
  );


  not
  g25
  (
    n53,
    n22
  );


  buf
  g26
  (
    n47,
    n5
  );


  not
  g27
  (
    n110,
    n1
  );


  not
  g28
  (
    n42,
    n17
  );


  buf
  g29
  (
    n55,
    n8
  );


  not
  g30
  (
    n84,
    n16
  );


  not
  g31
  (
    n94,
    n11
  );


  not
  g32
  (
    n98,
    n16
  );


  not
  g33
  (
    n61,
    n15
  );


  not
  g34
  (
    n36,
    n14
  );


  buf
  g35
  (
    n113,
    n18
  );


  not
  g36
  (
    n74,
    n23
  );


  buf
  g37
  (
    n104,
    n20
  );


  buf
  g38
  (
    n121,
    n7
  );


  not
  g39
  (
    n85,
    n23
  );


  not
  g40
  (
    n105,
    n13
  );


  buf
  g41
  (
    n81,
    n21
  );


  not
  g42
  (
    n66,
    n10
  );


  buf
  g43
  (
    n83,
    n4
  );


  not
  g44
  (
    n70,
    n10
  );


  buf
  g45
  (
    n30,
    n19
  );


  buf
  g46
  (
    n111,
    n7
  );


  buf
  g47
  (
    n68,
    n2
  );


  buf
  g48
  (
    n73,
    n3
  );


  not
  g49
  (
    n90,
    n11
  );


  buf
  g50
  (
    n67,
    n24
  );


  buf
  g51
  (
    n93,
    n6
  );


  not
  g52
  (
    n82,
    n11
  );


  buf
  g53
  (
    n87,
    n21
  );


  not
  g54
  (
    n77,
    n1
  );


  not
  g55
  (
    n120,
    n15
  );


  buf
  g56
  (
    n116,
    n9
  );


  not
  g57
  (
    n100,
    n4
  );


  buf
  g58
  (
    n46,
    n7
  );


  not
  g59
  (
    n95,
    n17
  );


  not
  g60
  (
    n33,
    n18
  );


  buf
  g61
  (
    n69,
    n19
  );


  not
  g62
  (
    n60,
    n24
  );


  buf
  g63
  (
    n79,
    n17
  );


  buf
  g64
  (
    n99,
    n13
  );


  buf
  g65
  (
    n102,
    n2
  );


  buf
  g66
  (
    n89,
    n19
  );


  not
  g67
  (
    n37,
    n13
  );


  buf
  g68
  (
    n80,
    n25
  );


  not
  g69
  (
    n39,
    n9
  );


  not
  g70
  (
    n123,
    n17
  );


  not
  g71
  (
    n112,
    n12
  );


  buf
  g72
  (
    n92,
    n1
  );


  buf
  g73
  (
    n32,
    n12
  );


  not
  g74
  (
    n35,
    n22
  );


  not
  g75
  (
    n45,
    n21
  );


  buf
  g76
  (
    n62,
    n3
  );


  buf
  g77
  (
    n125,
    n4
  );


  not
  g78
  (
    n31,
    n10
  );


  not
  g79
  (
    n78,
    n15
  );


  buf
  g80
  (
    n51,
    n8
  );


  buf
  g81
  (
    n65,
    n8
  );


  buf
  g82
  (
    n75,
    n12
  );


  not
  g83
  (
    n103,
    n25
  );


  not
  g84
  (
    n44,
    n18
  );


  buf
  g85
  (
    n96,
    n22
  );


  buf
  g86
  (
    n58,
    n2
  );


  buf
  g87
  (
    n54,
    n20
  );


  buf
  g88
  (
    n76,
    n15
  );


  not
  g89
  (
    n119,
    n4
  );


  not
  g90
  (
    n29,
    n24
  );


  buf
  g91
  (
    n59,
    n6
  );


  buf
  g92
  (
    n107,
    n3
  );


  not
  g93
  (
    n117,
    n6
  );


  not
  g94
  (
    n40,
    n19
  );


  buf
  g95
  (
    n88,
    n13
  );


  not
  g96
  (
    n49,
    n20
  );


  not
  g97
  (
    n28,
    n20
  );


  not
  g98
  (
    n124,
    n11
  );


  buf
  g99
  (
    n63,
    n2
  );


  not
  g100
  (
    n216,
    n96
  );


  buf
  g101
  (
    n179,
    n95
  );


  buf
  g102
  (
    n270,
    n55
  );


  buf
  g103
  (
    n231,
    n35
  );


  not
  g104
  (
    n274,
    n33
  );


  not
  g105
  (
    n271,
    n105
  );


  not
  g106
  (
    n193,
    n101
  );


  not
  g107
  (
    n161,
    n110
  );


  not
  g108
  (
    n261,
    n52
  );


  not
  g109
  (
    n176,
    n70
  );


  not
  g110
  (
    n206,
    n84
  );


  not
  g111
  (
    n165,
    n76
  );


  buf
  g112
  (
    n152,
    n70
  );


  not
  g113
  (
    n217,
    n83
  );


  not
  g114
  (
    n214,
    n118
  );


  buf
  g115
  (
    n177,
    n48
  );


  not
  g116
  (
    n245,
    n108
  );


  buf
  g117
  (
    n221,
    n89
  );


  not
  g118
  (
    n131,
    n60
  );


  not
  g119
  (
    n138,
    n38
  );


  not
  g120
  (
    n196,
    n117
  );


  not
  g121
  (
    n141,
    n123
  );


  not
  g122
  (
    n126,
    n77
  );


  buf
  g123
  (
    n247,
    n46
  );


  buf
  g124
  (
    n254,
    n112
  );


  not
  g125
  (
    n209,
    n88
  );


  not
  g126
  (
    n192,
    n56
  );


  not
  g127
  (
    n160,
    n117
  );


  not
  g128
  (
    n218,
    n110
  );


  not
  g129
  (
    n267,
    n35
  );


  not
  g130
  (
    n148,
    n107
  );


  buf
  g131
  (
    n255,
    n87
  );


  not
  g132
  (
    n275,
    n113
  );


  not
  g133
  (
    n129,
    n74
  );


  not
  g134
  (
    n128,
    n85
  );


  buf
  g135
  (
    n248,
    n44
  );


  not
  g136
  (
    n240,
    n37
  );


  buf
  g137
  (
    n151,
    n85
  );


  not
  g138
  (
    n185,
    n61
  );


  not
  g139
  (
    n205,
    n55
  );


  not
  g140
  (
    n225,
    n52
  );


  buf
  g141
  (
    n158,
    n80
  );


  not
  g142
  (
    n145,
    n104
  );


  buf
  g143
  (
    n210,
    n67
  );


  buf
  g144
  (
    n224,
    n63
  );


  buf
  g145
  (
    n219,
    n32
  );


  buf
  g146
  (
    n264,
    n59
  );


  not
  g147
  (
    n149,
    n122
  );


  buf
  g148
  (
    n234,
    n116
  );


  buf
  g149
  (
    n189,
    n32
  );


  not
  g150
  (
    n220,
    n73
  );


  not
  g151
  (
    n213,
    n56
  );


  buf
  g152
  (
    n178,
    n42
  );


  not
  g153
  (
    n139,
    n105
  );


  not
  g154
  (
    n134,
    n51
  );


  not
  g155
  (
    n146,
    n86
  );


  not
  g156
  (
    n142,
    n41
  );


  not
  g157
  (
    n182,
    n125
  );


  buf
  g158
  (
    n239,
    n91
  );


  buf
  g159
  (
    n170,
    n81
  );


  not
  g160
  (
    n262,
    n110
  );


  buf
  g161
  (
    n135,
    n93
  );


  buf
  g162
  (
    n243,
    n110
  );


  not
  g163
  (
    n187,
    n28
  );


  not
  g164
  (
    n195,
    n26
  );


  buf
  g165
  (
    n164,
    n108
  );


  not
  g166
  (
    n207,
    n36
  );


  buf
  g167
  (
    n252,
    n39
  );


  buf
  g168
  (
    n166,
    n68
  );


  buf
  g169
  (
    n222,
    n43
  );


  not
  g170
  (
    n269,
    n89
  );


  buf
  g171
  (
    n258,
    n46
  );


  not
  g172
  (
    n265,
    n119
  );


  buf
  g173
  (
    n150,
    n34
  );


  or
  g174
  (
    n147,
    n40,
    n92
  );


  xor
  g175
  (
    n136,
    n89,
    n66,
    n75,
    n79
  );


  nand
  g176
  (
    n184,
    n72,
    n39,
    n103,
    n107
  );


  xnor
  g177
  (
    n276,
    n120,
    n27,
    n111,
    n81
  );


  nor
  g178
  (
    n186,
    n107,
    n34,
    n105,
    n59
  );


  nand
  g179
  (
    n257,
    n45,
    n115,
    n114
  );


  or
  g180
  (
    n169,
    n119,
    n106,
    n72,
    n79
  );


  nor
  g181
  (
    n223,
    n29,
    n64,
    n99,
    n82
  );


  nand
  g182
  (
    n143,
    n75,
    n80,
    n96,
    n91
  );


  nor
  g183
  (
    n175,
    n81,
    n120,
    n79,
    n68
  );


  and
  g184
  (
    n227,
    n54,
    n58,
    n86
  );


  nand
  g185
  (
    n171,
    n55,
    n53,
    n85,
    n107
  );


  or
  g186
  (
    n235,
    n73,
    n97,
    n72,
    n76
  );


  nor
  g187
  (
    n236,
    n102,
    n36,
    n120,
    n123
  );


  and
  g188
  (
    n191,
    n50,
    n43,
    n62,
    n123
  );


  or
  g189
  (
    n260,
    n44,
    n121,
    n94
  );


  xor
  g190
  (
    n279,
    n121,
    n112,
    n60,
    n45
  );


  or
  g191
  (
    n215,
    n37,
    n40,
    n82,
    n115
  );


  xor
  g192
  (
    n268,
    n65,
    n50,
    n58,
    n69
  );


  nor
  g193
  (
    n263,
    n90,
    n78,
    n29,
    n42
  );


  and
  g194
  (
    n278,
    n102,
    n36,
    n90,
    n58
  );


  xor
  g195
  (
    n156,
    n31,
    n115,
    n108,
    n104
  );


  nor
  g196
  (
    n157,
    n47,
    n56,
    n101,
    n27
  );


  xnor
  g197
  (
    n155,
    n95,
    n93,
    n77,
    n79
  );


  nor
  g198
  (
    n201,
    n76,
    n116,
    n92,
    n49
  );


  and
  g199
  (
    n249,
    n42,
    n74,
    n90,
    n61
  );


  or
  g200
  (
    n242,
    n43,
    n38,
    n90,
    n67
  );


  xnor
  g201
  (
    n266,
    n94,
    n73,
    n37,
    n33
  );


  nor
  g202
  (
    n253,
    n91,
    n68,
    n71
  );


  xor
  g203
  (
    n277,
    n84,
    n66,
    n34,
    n116
  );


  xor
  g204
  (
    n163,
    n65,
    n109,
    n42,
    n27
  );


  nor
  g205
  (
    n204,
    n74,
    n113,
    n88
  );


  or
  g206
  (
    n140,
    n30,
    n69,
    n63,
    n53
  );


  and
  g207
  (
    n256,
    n99,
    n59,
    n26,
    n30
  );


  and
  g208
  (
    n172,
    n57,
    n31,
    n30,
    n41
  );


  xnor
  g209
  (
    n228,
    n32,
    n118,
    n49,
    n63
  );


  xor
  g210
  (
    n246,
    n104,
    n43,
    n116,
    n118
  );


  nor
  g211
  (
    n190,
    n106,
    n121,
    n113,
    n69
  );


  or
  g212
  (
    n280,
    n38,
    n71,
    n95,
    n45
  );


  and
  g213
  (
    n168,
    n64,
    n86,
    n87,
    n111
  );


  nand
  g214
  (
    n198,
    n66,
    n124,
    n54
  );


  nand
  g215
  (
    n244,
    n91,
    n75,
    n103,
    n84
  );


  and
  g216
  (
    n183,
    n72,
    n33,
    n63,
    n39
  );


  nand
  g217
  (
    n154,
    n106,
    n92,
    n27,
    n67
  );


  nor
  g218
  (
    n188,
    n64,
    n31,
    n36,
    n98
  );


  and
  g219
  (
    n208,
    n125,
    n96,
    n109,
    n102
  );


  or
  g220
  (
    n232,
    n122,
    n44,
    n124,
    n81
  );


  or
  g221
  (
    n167,
    n46,
    n64,
    n55,
    n103
  );


  and
  g222
  (
    n281,
    n97,
    n124,
    n111,
    n35
  );


  xnor
  g223
  (
    n137,
    n103,
    n97,
    n83,
    n123
  );


  nor
  g224
  (
    n229,
    n28,
    n84,
    n113,
    n93
  );


  xor
  g225
  (
    n199,
    n80,
    n61,
    n106,
    n82
  );


  and
  g226
  (
    n194,
    n71,
    n65,
    n49,
    n96
  );


  or
  g227
  (
    n238,
    n117,
    n109,
    n29,
    n87
  );


  or
  g228
  (
    n251,
    n83,
    n50,
    n45,
    n112
  );


  nor
  g229
  (
    n202,
    n62,
    n100,
    n52,
    n56
  );


  and
  g230
  (
    n174,
    n39,
    n49,
    n51,
    n114
  );


  xor
  g231
  (
    n162,
    n61,
    n98,
    n48,
    n99
  );


  xnor
  g232
  (
    n153,
    n46,
    n75,
    n37,
    n58
  );


  and
  g233
  (
    n159,
    n26,
    n111,
    n100,
    n119
  );


  nand
  g234
  (
    n200,
    n53,
    n94,
    n80,
    n104
  );


  nand
  g235
  (
    n226,
    n101,
    n92,
    n89,
    n88
  );


  or
  g236
  (
    n211,
    n119,
    n29,
    n66,
    n76
  );


  nor
  g237
  (
    n132,
    n53,
    n48,
    n41,
    n95
  );


  nand
  g238
  (
    n130,
    n51,
    n109,
    n65,
    n54
  );


  nor
  g239
  (
    n241,
    n69,
    n121,
    n100,
    n40
  );


  xnor
  g240
  (
    n197,
    n47,
    n78,
    n73,
    n122
  );


  xor
  g241
  (
    n230,
    n41,
    n101,
    n32,
    n99
  );


  xor
  g242
  (
    n237,
    n112,
    n74,
    n78,
    n54
  );


  or
  g243
  (
    n203,
    n105,
    n59,
    n57,
    n50
  );


  xor
  g244
  (
    n180,
    n62,
    n57,
    n51,
    n47
  );


  and
  g245
  (
    n259,
    n125,
    n70,
    n48,
    n114
  );


  or
  g246
  (
    n144,
    n82,
    n52,
    n60,
    n26
  );


  xor
  g247
  (
    n133,
    n62,
    n30,
    n118,
    n77
  );


  or
  g248
  (
    n250,
    n93,
    n108,
    n57,
    n71
  );


  xnor
  g249
  (
    n127,
    n100,
    n120,
    n78,
    n44
  );


  nand
  g250
  (
    n212,
    n38,
    n125,
    n85,
    n98
  );


  xor
  g251
  (
    n233,
    n33,
    n47,
    n28,
    n60
  );


  nor
  g252
  (
    n173,
    n28,
    n114,
    n83,
    n31
  );


  or
  g253
  (
    n273,
    n70,
    n97,
    n98,
    n67
  );


  xnor
  g254
  (
    n181,
    n40,
    n35,
    n122,
    n102
  );


  xnor
  g255
  (
    n272,
    n87,
    n34,
    n77,
    n117
  );


  xor
  g256
  (
    n302,
    n225,
    n218,
    n223,
    n193
  );


  xor
  g257
  (
    n339,
    n225,
    n195,
    n263,
    n234
  );


  nand
  g258
  (
    n304,
    n134,
    n232,
    n171,
    n268
  );


  nor
  g259
  (
    n287,
    n202,
    n242,
    n277,
    n214
  );


  and
  g260
  (
    n394,
    n149,
    n191,
    n241,
    n180
  );


  nand
  g261
  (
    n321,
    n249,
    n201,
    n190,
    n257
  );


  or
  g262
  (
    n355,
    n137,
    n273,
    n138,
    n200
  );


  nor
  g263
  (
    n309,
    n141,
    n152,
    n210,
    n130
  );


  nor
  g264
  (
    n317,
    n231,
    n247,
    n260,
    n137
  );


  xor
  g265
  (
    n341,
    n216,
    n200,
    n146,
    n128
  );


  and
  g266
  (
    n353,
    n159,
    n208,
    n199,
    n217
  );


  xor
  g267
  (
    n319,
    n195,
    n163,
    n206,
    n147
  );


  and
  g268
  (
    n306,
    n224,
    n180,
    n176,
    n202
  );


  nand
  g269
  (
    n376,
    n155,
    n145,
    n218,
    n167
  );


  xnor
  g270
  (
    n395,
    n182,
    n264,
    n192,
    n189
  );


  or
  g271
  (
    n298,
    n221,
    n191,
    n151,
    n132
  );


  and
  g272
  (
    n369,
    n185,
    n197,
    n141,
    n260
  );


  xnor
  g273
  (
    n359,
    n272,
    n272,
    n266,
    n274
  );


  or
  g274
  (
    n337,
    n267,
    n211,
    n243,
    n227
  );


  and
  g275
  (
    n311,
    n152,
    n272,
    n133,
    n233
  );


  xnor
  g276
  (
    n357,
    n247,
    n223,
    n204,
    n203
  );


  nand
  g277
  (
    n354,
    n247,
    n127,
    n212,
    n246
  );


  or
  g278
  (
    n385,
    n214,
    n267,
    n183,
    n129
  );


  nand
  g279
  (
    n324,
    n270,
    n264,
    n278,
    n251
  );


  nor
  g280
  (
    n331,
    n207,
    n213,
    n221,
    n181
  );


  xnor
  g281
  (
    n282,
    n193,
    n275,
    n248,
    n234
  );


  or
  g282
  (
    n293,
    n147,
    n168,
    n252,
    n251
  );


  xnor
  g283
  (
    n351,
    n280,
    n160,
    n281,
    n153
  );


  or
  g284
  (
    n368,
    n178,
    n194,
    n269,
    n163
  );


  nand
  g285
  (
    n398,
    n148,
    n252,
    n245,
    n166
  );


  nor
  g286
  (
    n328,
    n270,
    n280,
    n164,
    n224
  );


  and
  g287
  (
    n325,
    n217,
    n249,
    n171,
    n144
  );


  and
  g288
  (
    n338,
    n207,
    n240,
    n187,
    n204
  );


  nand
  g289
  (
    n315,
    n181,
    n144,
    n174
  );


  and
  g290
  (
    n292,
    n239,
    n235,
    n156,
    n212
  );


  xor
  g291
  (
    n374,
    n196,
    n228,
    n256,
    n229
  );


  xor
  g292
  (
    n362,
    n134,
    n254,
    n220,
    n135
  );


  or
  g293
  (
    n314,
    n153,
    n258,
    n273,
    n178
  );


  nand
  g294
  (
    n387,
    n251,
    n195,
    n157,
    n196
  );


  or
  g295
  (
    n379,
    n261,
    n145,
    n126,
    n191
  );


  or
  g296
  (
    n386,
    n198,
    n273,
    n241,
    n259
  );


  xnor
  g297
  (
    n361,
    n225,
    n245,
    n184,
    n222
  );


  nor
  g298
  (
    n390,
    n266,
    n205,
    n176,
    n206
  );


  nor
  g299
  (
    n378,
    n183,
    n236,
    n259,
    n127
  );


  or
  g300
  (
    n344,
    n211,
    n169,
    n255,
    n192
  );


  or
  g301
  (
    n373,
    n208,
    n226,
    n209,
    n231
  );


  nand
  g302
  (
    n388,
    n140,
    n150,
    n215,
    n174
  );


  xor
  g303
  (
    n358,
    n232,
    n190,
    n131,
    n235
  );


  or
  g304
  (
    n397,
    n175,
    n230,
    n244,
    n243
  );


  and
  g305
  (
    n366,
    n223,
    n153,
    n128,
    n269
  );


  nand
  g306
  (
    n389,
    n170,
    n276,
    n147,
    n186
  );


  xnor
  g307
  (
    n323,
    n219,
    n168,
    n265,
    n154
  );


  and
  g308
  (
    n380,
    n215,
    n254,
    n207,
    n182
  );


  xor
  g309
  (
    n286,
    n133,
    n239,
    n138,
    n271
  );


  and
  g310
  (
    n305,
    n186,
    n242,
    n209,
    n263
  );


  or
  g311
  (
    n329,
    n268,
    n237,
    n244,
    n136
  );


  xor
  g312
  (
    n384,
    n260,
    n188,
    n184,
    n136
  );


  xor
  g313
  (
    n318,
    n162,
    n219,
    n186,
    n210
  );


  xnor
  g314
  (
    n303,
    n198,
    n175,
    n154,
    n248
  );


  or
  g315
  (
    n375,
    n131,
    n242,
    n279,
    n248
  );


  or
  g316
  (
    n365,
    n255,
    n267,
    n228,
    n128
  );


  xor
  g317
  (
    n347,
    n213,
    n150,
    n250,
    n240
  );


  or
  g318
  (
    n313,
    n257,
    n148,
    n280,
    n182
  );


  nand
  g319
  (
    n392,
    n271,
    n196,
    n215,
    n243
  );


  xnor
  g320
  (
    n335,
    n236,
    n154,
    n270,
    n277
  );


  and
  g321
  (
    n290,
    n268,
    n190,
    n137,
    n161
  );


  or
  g322
  (
    n330,
    n226,
    n150,
    n224,
    n261
  );


  xnor
  g323
  (
    n346,
    n180,
    n158,
    n178,
    n262
  );


  nor
  g324
  (
    n336,
    n149,
    n146,
    n173,
    n221
  );


  nand
  g325
  (
    n312,
    n141,
    n275,
    n143,
    n250
  );


  xor
  g326
  (
    n334,
    n220,
    n140,
    n160
  );


  nand
  g327
  (
    n370,
    n143,
    n238,
    n135,
    n198
  );


  and
  g328
  (
    n352,
    n155,
    n220,
    n240,
    n156
  );


  xnor
  g329
  (
    n364,
    n194,
    n271,
    n161,
    n266
  );


  xnor
  g330
  (
    n371,
    n170,
    n226,
    n232,
    n158
  );


  xnor
  g331
  (
    n297,
    n135,
    n250,
    n246,
    n278
  );


  or
  g332
  (
    n342,
    n230,
    n143,
    n237,
    n199
  );


  or
  g333
  (
    n345,
    n236,
    n152,
    n222,
    n206
  );


  and
  g334
  (
    n301,
    n203,
    n192,
    n157,
    n262
  );


  and
  g335
  (
    n288,
    n252,
    n139,
    n176,
    n126
  );


  xor
  g336
  (
    n377,
    n214,
    n163,
    n173,
    n167
  );


  or
  g337
  (
    n285,
    n205,
    n274,
    n139,
    n197
  );


  xnor
  g338
  (
    n340,
    n185,
    n205,
    n222,
    n166
  );


  or
  g339
  (
    n350,
    n256,
    n245,
    n149,
    n162
  );


  nor
  g340
  (
    n291,
    n218,
    n132,
    n217,
    n276
  );


  nand
  g341
  (
    n294,
    n263,
    n172,
    n193,
    n230
  );


  nor
  g342
  (
    n327,
    n227,
    n256,
    n177,
    n139
  );


  nand
  g343
  (
    n299,
    n175,
    n281,
    n253,
    n187
  );


  nand
  g344
  (
    n381,
    n258,
    n168,
    n189,
    n201
  );


  xor
  g345
  (
    n382,
    n167,
    n177,
    n127,
    n274
  );


  or
  g346
  (
    n393,
    n254,
    n171,
    n203,
    n130
  );


  nor
  g347
  (
    n296,
    n194,
    n211,
    n181,
    n136
  );


  xnor
  g348
  (
    n316,
    n142,
    n265,
    n155,
    n239
  );


  xnor
  g349
  (
    n308,
    n161,
    n156,
    n204,
    n238
  );


  or
  g350
  (
    n372,
    n201,
    n159,
    n129,
    n188
  );


  or
  g351
  (
    n343,
    n158,
    n189,
    n265,
    n133
  );


  xnor
  g352
  (
    n307,
    n162,
    n159,
    n157,
    n142
  );


  and
  g353
  (
    n295,
    n183,
    n275,
    n202,
    n253
  );


  or
  g354
  (
    n356,
    n172,
    n278,
    n165,
    n216
  );


  and
  g355
  (
    n349,
    n165,
    n179,
    n258,
    n187
  );


  xnor
  g356
  (
    n360,
    n255,
    n238,
    n169,
    n166
  );


  xnor
  g357
  (
    n363,
    n235,
    n142,
    n148,
    n228
  );


  xnor
  g358
  (
    n348,
    n269,
    n213,
    n209,
    n165
  );


  nand
  g359
  (
    n310,
    n237,
    n179,
    n249,
    n129
  );


  xor
  g360
  (
    n367,
    n216,
    n177,
    n231,
    n200
  );


  nand
  g361
  (
    n322,
    n145,
    n261,
    n281,
    n151
  );


  nand
  g362
  (
    n320,
    n208,
    n229,
    n227,
    n132
  );


  nor
  g363
  (
    n383,
    n229,
    n257,
    n199,
    n233
  );


  xor
  g364
  (
    n326,
    n219,
    n131,
    n184,
    n264
  );


  nor
  g365
  (
    n333,
    n277,
    n144,
    n210,
    n276
  );


  xor
  g366
  (
    n391,
    n130,
    n164,
    n279
  );


  nor
  g367
  (
    n396,
    n138,
    n185,
    n188,
    n126
  );


  or
  g368
  (
    n283,
    n212,
    n197,
    n262,
    n279
  );


  nand
  g369
  (
    n332,
    n172,
    n169,
    n134,
    n259
  );


  xor
  g370
  (
    n300,
    n170,
    n246,
    n151,
    n173
  );


  xor
  g371
  (
    n289,
    n241,
    n179,
    n233,
    n234
  );


  or
  g372
  (
    n284,
    n253,
    n146,
    n244,
    n160
  );


  nand
  g373
  (
    n481,
    n321,
    n285,
    n334
  );


  xnor
  g374
  (
    n408,
    n284,
    n321,
    n319,
    n308
  );


  xor
  g375
  (
    n474,
    n346,
    n331,
    n313,
    n339
  );


  nand
  g376
  (
    n456,
    n298,
    n325,
    n347,
    n394
  );


  xnor
  g377
  (
    n440,
    n380,
    n390,
    n326,
    n369
  );


  nand
  g378
  (
    n430,
    n342,
    n292,
    n318,
    n355
  );


  nor
  g379
  (
    n421,
    n378,
    n283,
    n381,
    n302
  );


  nor
  g380
  (
    n425,
    n320,
    n296,
    n338,
    n367
  );


  xnor
  g381
  (
    n470,
    n285,
    n337,
    n321,
    n318
  );


  nand
  g382
  (
    n410,
    n377,
    n391,
    n390,
    n358
  );


  xnor
  g383
  (
    n426,
    n380,
    n372,
    n362,
    n359
  );


  nor
  g384
  (
    n455,
    n355,
    n301,
    n309,
    n371
  );


  or
  g385
  (
    n483,
    n388,
    n290,
    n356
  );


  xor
  g386
  (
    n448,
    n373,
    n350,
    n340,
    n284
  );


  xor
  g387
  (
    n431,
    n341,
    n304,
    n300,
    n297
  );


  xor
  g388
  (
    n459,
    n305,
    n390,
    n336,
    n386
  );


  and
  g389
  (
    n458,
    n339,
    n305,
    n288,
    n333
  );


  xor
  g390
  (
    n469,
    n320,
    n375,
    n326,
    n312
  );


  and
  g391
  (
    n486,
    n357,
    n353,
    n324,
    n336
  );


  or
  g392
  (
    n419,
    n389,
    n396,
    n316,
    n294
  );


  xor
  g393
  (
    n452,
    n354,
    n353,
    n387,
    n314
  );


  or
  g394
  (
    n471,
    n341,
    n318,
    n369,
    n328
  );


  nor
  g395
  (
    n417,
    n303,
    n385,
    n351,
    n341
  );


  nor
  g396
  (
    n438,
    n357,
    n391,
    n377,
    n375
  );


  nor
  g397
  (
    n476,
    n290,
    n395,
    n315,
    n286
  );


  xnor
  g398
  (
    n433,
    n383,
    n364,
    n308,
    n327
  );


  nand
  g399
  (
    n467,
    n345,
    n307,
    n343,
    n309
  );


  xor
  g400
  (
    n473,
    n346,
    n365,
    n301,
    n293
  );


  or
  g401
  (
    n453,
    n362,
    n353,
    n380,
    n287
  );


  nor
  g402
  (
    n401,
    n330,
    n322,
    n389,
    n357
  );


  nand
  g403
  (
    n485,
    n397,
    n387,
    n322,
    n367
  );


  nand
  g404
  (
    n449,
    n366,
    n368,
    n337,
    n398
  );


  and
  g405
  (
    n444,
    n355,
    n310,
    n338,
    n361
  );


  and
  g406
  (
    n437,
    n289,
    n311,
    n327,
    n329
  );


  xor
  g407
  (
    n478,
    n289,
    n317,
    n284,
    n331
  );


  xor
  g408
  (
    n484,
    n359,
    n291,
    n311,
    n345
  );


  nor
  g409
  (
    n416,
    n366,
    n381,
    n297,
    n388
  );


  and
  g410
  (
    n427,
    n373,
    n336,
    n326,
    n364
  );


  xor
  g411
  (
    n441,
    n294,
    n371,
    n332,
    n282
  );


  xor
  g412
  (
    n446,
    n356,
    n316,
    n317,
    n361
  );


  or
  g413
  (
    n461,
    n297,
    n286,
    n396,
    n314
  );


  xnor
  g414
  (
    n429,
    n305,
    n323,
    n364,
    n375
  );


  xor
  g415
  (
    n418,
    n367,
    n382,
    n343,
    n360
  );


  nor
  g416
  (
    n402,
    n379,
    n330,
    n293,
    n352
  );


  xor
  g417
  (
    n423,
    n313,
    n295,
    n389,
    n370
  );


  xor
  g418
  (
    n405,
    n312,
    n383,
    n319,
    n330
  );


  nand
  g419
  (
    n466,
    n302,
    n323,
    n392,
    n344
  );


  and
  g420
  (
    n413,
    n395,
    n288,
    n370,
    n302
  );


  nor
  g421
  (
    n443,
    n317,
    n334,
    n290,
    n379
  );


  and
  g422
  (
    n435,
    n361,
    n299,
    n301,
    n386
  );


  xor
  g423
  (
    n428,
    n324,
    n393,
    n391,
    n329
  );


  xnor
  g424
  (
    n482,
    n300,
    n352,
    n371,
    n363
  );


  or
  g425
  (
    n454,
    n315,
    n288,
    n351,
    n291
  );


  nand
  g426
  (
    n460,
    n366,
    n299,
    n370,
    n289
  );


  or
  g427
  (
    n415,
    n328,
    n306,
    n325,
    n374
  );


  and
  g428
  (
    n462,
    n300,
    n381,
    n382,
    n398
  );


  xnor
  g429
  (
    n479,
    n303,
    n287,
    n340,
    n360
  );


  or
  g430
  (
    n465,
    n333,
    n349,
    n395,
    n348
  );


  nor
  g431
  (
    n414,
    n382,
    n360,
    n379,
    n283
  );


  xor
  g432
  (
    n457,
    n350,
    n335,
    n323,
    n307
  );


  or
  g433
  (
    n472,
    n348,
    n308,
    n294,
    n368
  );


  nand
  g434
  (
    n403,
    n376,
    n311,
    n334,
    n392
  );


  and
  g435
  (
    n439,
    n393,
    n307,
    n358,
    n304
  );


  or
  g436
  (
    n409,
    n397,
    n335,
    n372,
    n342
  );


  and
  g437
  (
    n468,
    n369,
    n329,
    n298,
    n363
  );


  or
  g438
  (
    n436,
    n358,
    n292,
    n385,
    n392
  );


  and
  g439
  (
    n407,
    n328,
    n310,
    n332,
    n384
  );


  xnor
  g440
  (
    n480,
    n298,
    n387,
    n348,
    n286
  );


  nor
  g441
  (
    n399,
    n396,
    n349,
    n344,
    n338
  );


  nand
  g442
  (
    n442,
    n349,
    n374,
    n344,
    n324
  );


  xor
  g443
  (
    n450,
    n282,
    n345,
    n394,
    n359
  );


  xnor
  g444
  (
    n424,
    n350,
    n388,
    n304,
    n282
  );


  nor
  g445
  (
    n412,
    n339,
    n327,
    n312,
    n386
  );


  nand
  g446
  (
    n463,
    n303,
    n362,
    n296,
    n306
  );


  nand
  g447
  (
    n406,
    n397,
    n306,
    n347,
    n376
  );


  and
  g448
  (
    n422,
    n295,
    n378,
    n374,
    n335
  );


  and
  g449
  (
    n451,
    n291,
    n384,
    n365,
    n296
  );


  and
  g450
  (
    n447,
    n313,
    n310,
    n346,
    n368
  );


  nand
  g451
  (
    n432,
    n337,
    n332,
    n285,
    n342
  );


  nor
  g452
  (
    n464,
    n365,
    n299,
    n322,
    n340
  );


  or
  g453
  (
    n420,
    n354,
    n287,
    n319,
    n295
  );


  xor
  g454
  (
    n411,
    n343,
    n376,
    n385,
    n325
  );


  or
  g455
  (
    n475,
    n363,
    n315,
    n331,
    n384
  );


  nand
  g456
  (
    n400,
    n373,
    n292,
    n394,
    n383
  );


  nor
  g457
  (
    n434,
    n283,
    n293,
    n377,
    n351
  );


  or
  g458
  (
    n477,
    n378,
    n393,
    n372,
    n354
  );


  nor
  g459
  (
    n404,
    n398,
    n314,
    n333,
    n347
  );


  or
  g460
  (
    n445,
    n316,
    n320,
    n309,
    n352
  );


  nor
  g461
  (
    n491,
    n463,
    n486,
    n423,
    n411
  );


  or
  g462
  (
    n501,
    n431,
    n449,
    n459,
    n479
  );


  and
  g463
  (
    n496,
    n403,
    n414,
    n461,
    n484
  );


  xnor
  g464
  (
    n487,
    n478,
    n466,
    n400,
    n470
  );


  and
  g465
  (
    n506,
    n438,
    n432,
    n480,
    n421
  );


  xor
  g466
  (
    n489,
    n402,
    n478,
    n442,
    n457
  );


  nor
  g467
  (
    n502,
    n462,
    n418,
    n467,
    n477
  );


  xnor
  g468
  (
    n505,
    n410,
    n477,
    n460,
    n441
  );


  or
  g469
  (
    n493,
    n482,
    n426,
    n472,
    n476
  );


  nor
  g470
  (
    n503,
    n446,
    n448,
    n399,
    n429
  );


  xnor
  g471
  (
    AntiSAT_key_wire,
    n474,
    n475,
    n416,
    n479
  );


  and
  g472
  (
    n492,
    n486,
    n484,
    n405,
    n427
  );


  nor
  g473
  (
    n512,
    n435,
    n455,
    n422,
    n482
  );


  xor
  g474
  (
    n509,
    n485,
    n482,
    n430,
    n480
  );


  or
  g475
  (
    n511,
    n475,
    n484,
    n409,
    n445
  );


  nor
  g476
  (
    n513,
    n420,
    n417,
    n454,
    n406
  );


  and
  g477
  (
    n497,
    n465,
    n437,
    n483,
    n478
  );


  or
  g478
  (
    n490,
    n443,
    n433,
    n444,
    n412
  );


  xor
  g479
  (
    n498,
    n428,
    n456,
    n481,
    n485
  );


  xnor
  g480
  (
    n507,
    n479,
    n477,
    n476,
    n481
  );


  or
  g481
  (
    n494,
    n483,
    n483,
    n485,
    n439
  );


  nor
  g482
  (
    n500,
    n458,
    n404,
    n469,
    n481
  );


  xnor
  g483
  (
    n499,
    n425,
    n450,
    n436,
    n447
  );


  xor
  g484
  (
    n488,
    n468,
    n419,
    n434,
    n415
  );


  and
  g485
  (
    n495,
    n473,
    n424,
    n413,
    n464
  );


  nor
  g486
  (
    n504,
    n486,
    n401,
    n476,
    n407
  );


  and
  g487
  (
    n508,
    n471,
    n440,
    n451,
    n452
  );


  nor
  g488
  (
    n514,
    n475,
    n408,
    n453,
    n480
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_25
  (
    gbar_input_0_0,
    keyIn_0_25,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_1,
    keyIn_0_26,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_2,
    keyIn_0_27,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_3,
    keyIn_0_28,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_4,
    keyIn_0_29,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_5,
    keyIn_0_30,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_6,
    keyIn_0_31,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_7,
    keyIn_0_32,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_8,
    keyIn_0_33,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_9,
    keyIn_0_34,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_10,
    keyIn_0_35,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_11,
    keyIn_0_36,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_12,
    keyIn_0_37,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_13,
    keyIn_0_38,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_14,
    keyIn_0_39,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_15,
    keyIn_0_40,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_16,
    keyIn_0_41,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_17,
    keyIn_0_42,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_18,
    keyIn_0_43,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_19,
    keyIn_0_44,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_20,
    keyIn_0_45,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_21,
    keyIn_0_46,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_22,
    keyIn_0_47,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_23,
    keyIn_0_48,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_24,
    keyIn_0_49,
    n25
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n510,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

