

module Stat_821_382
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n571,
  n767,
  n766,
  n764,
  n760,
  n765,
  n770,
  n762,
  n768,
  n771,
  n759,
  n758,
  n796,
  n798,
  n803,
  n802,
  n811,
  n815,
  n828,
  n832,
  n833,
  n839,
  n840,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;
  output n571;output n767;output n766;output n764;output n760;output n765;output n770;output n762;output n768;output n771;output n759;output n758;output n796;output n798;output n803;output n802;output n811;output n815;output n828;output n832;output n833;output n839;output n840;
  wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n761;wire n763;wire n769;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n797;wire n799;wire n800;wire n801;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n812;wire n813;wire n814;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n829;wire n830;wire n831;wire n834;wire n835;wire n836;wire n837;wire n838;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n32,
    n7
  );


  buf
  g1
  (
    n89,
    n9
  );


  buf
  g2
  (
    n64,
    n18
  );


  buf
  g3
  (
    n42,
    n6
  );


  not
  g4
  (
    n54,
    n6
  );


  buf
  g5
  (
    n90,
    n15
  );


  buf
  g6
  (
    n22,
    n19
  );


  buf
  g7
  (
    n67,
    n19
  );


  buf
  g8
  (
    n36,
    n17
  );


  not
  g9
  (
    n71,
    n3
  );


  buf
  g10
  (
    n33,
    n12
  );


  not
  g11
  (
    n52,
    n2
  );


  buf
  g12
  (
    n44,
    n10
  );


  buf
  g13
  (
    n28,
    n19
  );


  buf
  g14
  (
    n20,
    n16
  );


  buf
  g15
  (
    n46,
    n18
  );


  not
  g16
  (
    n94,
    n8
  );


  buf
  g17
  (
    n25,
    n17
  );


  not
  g18
  (
    n24,
    n8
  );


  buf
  g19
  (
    n91,
    n13
  );


  buf
  g20
  (
    n70,
    n6
  );


  not
  g21
  (
    n57,
    n16
  );


  not
  g22
  (
    n84,
    n12
  );


  not
  g23
  (
    n85,
    n10
  );


  buf
  g24
  (
    n48,
    n1
  );


  buf
  g25
  (
    n88,
    n14
  );


  buf
  g26
  (
    n50,
    n2
  );


  buf
  g27
  (
    n75,
    n13
  );


  buf
  g28
  (
    n30,
    n7
  );


  not
  g29
  (
    n79,
    n2
  );


  not
  g30
  (
    n56,
    n18
  );


  buf
  g31
  (
    n77,
    n14
  );


  not
  g32
  (
    n87,
    n4
  );


  not
  g33
  (
    n51,
    n5
  );


  not
  g34
  (
    n39,
    n14
  );


  not
  g35
  (
    n45,
    n8
  );


  not
  g36
  (
    n23,
    n9
  );


  buf
  g37
  (
    n72,
    n18
  );


  not
  g38
  (
    n93,
    n6
  );


  buf
  g39
  (
    n73,
    n14
  );


  not
  g40
  (
    n78,
    n12
  );


  buf
  g41
  (
    n60,
    n15
  );


  buf
  g42
  (
    n41,
    n4
  );


  not
  g43
  (
    n61,
    n8
  );


  not
  g44
  (
    n63,
    n17
  );


  buf
  g45
  (
    n95,
    n2
  );


  not
  g46
  (
    n81,
    n4
  );


  not
  g47
  (
    n34,
    n11
  );


  buf
  g48
  (
    n38,
    n5
  );


  not
  g49
  (
    n40,
    n3
  );


  not
  g50
  (
    n59,
    n13
  );


  buf
  g51
  (
    n69,
    n16
  );


  buf
  g52
  (
    n35,
    n9
  );


  buf
  g53
  (
    n27,
    n3
  );


  not
  g54
  (
    n68,
    n5
  );


  not
  g55
  (
    n76,
    n4
  );


  not
  g56
  (
    n49,
    n17
  );


  not
  g57
  (
    n47,
    n11
  );


  buf
  g58
  (
    n58,
    n15
  );


  not
  g59
  (
    n37,
    n7
  );


  not
  g60
  (
    n83,
    n11
  );


  buf
  g61
  (
    n82,
    n15
  );


  not
  g62
  (
    n21,
    n7
  );


  not
  g63
  (
    n86,
    n10
  );


  buf
  g64
  (
    n74,
    n1
  );


  not
  g65
  (
    n65,
    n12
  );


  not
  g66
  (
    n29,
    n1
  );


  buf
  g67
  (
    n43,
    n13
  );


  buf
  g68
  (
    n55,
    n3
  );


  not
  g69
  (
    n66,
    n11
  );


  not
  g70
  (
    n53,
    n10
  );


  not
  g71
  (
    n31,
    n19
  );


  buf
  g72
  (
    n80,
    n1
  );


  not
  g73
  (
    n62,
    n9
  );


  buf
  g74
  (
    n26,
    n16
  );


  not
  g75
  (
    n92,
    n5
  );


  buf
  g76
  (
    n339,
    n73
  );


  buf
  g77
  (
    n137,
    n23
  );


  not
  g78
  (
    n219,
    n26
  );


  buf
  g79
  (
    n112,
    n20
  );


  buf
  g80
  (
    n125,
    n53
  );


  buf
  g81
  (
    n244,
    n70
  );


  not
  g82
  (
    n308,
    n69
  );


  not
  g83
  (
    n202,
    n24
  );


  not
  g84
  (
    n126,
    n70
  );


  buf
  g85
  (
    n325,
    n59
  );


  buf
  g86
  (
    n225,
    n37
  );


  not
  g87
  (
    n314,
    n71
  );


  not
  g88
  (
    n114,
    n81
  );


  not
  g89
  (
    n343,
    n59
  );


  buf
  g90
  (
    n212,
    n85
  );


  not
  g91
  (
    n352,
    n71
  );


  buf
  g92
  (
    n159,
    n22
  );


  buf
  g93
  (
    n139,
    n21
  );


  buf
  g94
  (
    n122,
    n41
  );


  buf
  g95
  (
    n100,
    n23
  );


  buf
  g96
  (
    n330,
    n42
  );


  buf
  g97
  (
    n111,
    n21
  );


  buf
  g98
  (
    n163,
    n58
  );


  buf
  g99
  (
    n151,
    n28
  );


  not
  g100
  (
    n260,
    n90
  );


  not
  g101
  (
    n318,
    n47
  );


  buf
  g102
  (
    n108,
    n88
  );


  not
  g103
  (
    n104,
    n82
  );


  buf
  g104
  (
    n121,
    n48
  );


  buf
  g105
  (
    n147,
    n84
  );


  not
  g106
  (
    n350,
    n89
  );


  not
  g107
  (
    n313,
    n25
  );


  not
  g108
  (
    n205,
    n22
  );


  buf
  g109
  (
    n256,
    n37
  );


  buf
  g110
  (
    n110,
    n88
  );


  buf
  g111
  (
    n236,
    n46
  );


  not
  g112
  (
    n182,
    n48
  );


  buf
  g113
  (
    n134,
    n49
  );


  buf
  g114
  (
    n243,
    n67
  );


  not
  g115
  (
    n266,
    n67
  );


  not
  g116
  (
    n380,
    n68
  );


  not
  g117
  (
    n262,
    n55
  );


  buf
  g118
  (
    n378,
    n61
  );


  buf
  g119
  (
    n310,
    n38
  );


  buf
  g120
  (
    n162,
    n77
  );


  buf
  g121
  (
    n117,
    n36
  );


  buf
  g122
  (
    n297,
    n87
  );


  not
  g123
  (
    n257,
    n43
  );


  not
  g124
  (
    n322,
    n31
  );


  not
  g125
  (
    n274,
    n60
  );


  buf
  g126
  (
    n319,
    n55
  );


  buf
  g127
  (
    n148,
    n54
  );


  buf
  g128
  (
    n311,
    n76
  );


  buf
  g129
  (
    n307,
    n74
  );


  buf
  g130
  (
    n127,
    n45
  );


  not
  g131
  (
    n279,
    n34
  );


  not
  g132
  (
    n269,
    n58
  );


  buf
  g133
  (
    n255,
    n39
  );


  not
  g134
  (
    n119,
    n36
  );


  buf
  g135
  (
    n200,
    n24
  );


  not
  g136
  (
    n348,
    n43
  );


  not
  g137
  (
    n193,
    n69
  );


  buf
  g138
  (
    n99,
    n67
  );


  buf
  g139
  (
    n216,
    n41
  );


  buf
  g140
  (
    n240,
    n36
  );


  not
  g141
  (
    n101,
    n38
  );


  not
  g142
  (
    n364,
    n30
  );


  not
  g143
  (
    n359,
    n47
  );


  buf
  g144
  (
    n340,
    n25
  );


  not
  g145
  (
    n323,
    n42
  );


  buf
  g146
  (
    n238,
    n39
  );


  buf
  g147
  (
    n250,
    n50
  );


  not
  g148
  (
    n172,
    n33
  );


  buf
  g149
  (
    n227,
    n22
  );


  buf
  g150
  (
    n189,
    n29
  );


  not
  g151
  (
    n371,
    n87
  );


  not
  g152
  (
    n267,
    n70
  );


  buf
  g153
  (
    n366,
    n76
  );


  buf
  g154
  (
    n261,
    n31
  );


  not
  g155
  (
    n303,
    n70
  );


  not
  g156
  (
    n105,
    n64
  );


  not
  g157
  (
    n334,
    n66
  );


  buf
  g158
  (
    n210,
    n51
  );


  not
  g159
  (
    n248,
    n80
  );


  buf
  g160
  (
    n146,
    n40
  );


  not
  g161
  (
    n342,
    n74
  );


  buf
  g162
  (
    n284,
    n34
  );


  not
  g163
  (
    n177,
    n56
  );


  not
  g164
  (
    n170,
    n80
  );


  buf
  g165
  (
    n191,
    n45
  );


  not
  g166
  (
    n158,
    n68
  );


  not
  g167
  (
    n188,
    n46
  );


  not
  g168
  (
    n229,
    n82
  );


  buf
  g169
  (
    n135,
    n82
  );


  not
  g170
  (
    n226,
    n24
  );


  buf
  g171
  (
    n301,
    n86
  );


  buf
  g172
  (
    n192,
    n34
  );


  buf
  g173
  (
    n120,
    n49
  );


  buf
  g174
  (
    n207,
    n30
  );


  buf
  g175
  (
    n259,
    n60
  );


  buf
  g176
  (
    n183,
    n66
  );


  not
  g177
  (
    n263,
    n60
  );


  buf
  g178
  (
    n252,
    n40
  );


  buf
  g179
  (
    n335,
    n22
  );


  buf
  g180
  (
    n357,
    n50
  );


  buf
  g181
  (
    n295,
    n43
  );


  buf
  g182
  (
    n345,
    n35
  );


  not
  g183
  (
    n132,
    n85
  );


  buf
  g184
  (
    n312,
    n51
  );


  buf
  g185
  (
    n361,
    n40
  );


  buf
  g186
  (
    n228,
    n55
  );


  not
  g187
  (
    n247,
    n52
  );


  buf
  g188
  (
    n285,
    n85
  );


  not
  g189
  (
    n201,
    n31
  );


  buf
  g190
  (
    n116,
    n49
  );


  buf
  g191
  (
    n195,
    n75
  );


  buf
  g192
  (
    n281,
    n59
  );


  not
  g193
  (
    n254,
    n86
  );


  not
  g194
  (
    n271,
    n24
  );


  buf
  g195
  (
    n234,
    n32
  );


  not
  g196
  (
    n346,
    n63
  );


  buf
  g197
  (
    n175,
    n75
  );


  not
  g198
  (
    n242,
    n35
  );


  buf
  g199
  (
    n180,
    n46
  );


  not
  g200
  (
    n272,
    n44
  );


  buf
  g201
  (
    n290,
    n84
  );


  buf
  g202
  (
    n324,
    n30
  );


  not
  g203
  (
    n153,
    n45
  );


  not
  g204
  (
    n160,
    n54
  );


  not
  g205
  (
    n249,
    n88
  );


  buf
  g206
  (
    n245,
    n35
  );


  buf
  g207
  (
    n214,
    n63
  );


  not
  g208
  (
    n265,
    n50
  );


  buf
  g209
  (
    n376,
    n28
  );


  not
  g210
  (
    n333,
    n74
  );


  not
  g211
  (
    n296,
    n32
  );


  not
  g212
  (
    n231,
    n77
  );


  buf
  g213
  (
    n369,
    n56
  );


  not
  g214
  (
    n109,
    n46
  );


  not
  g215
  (
    n161,
    n62
  );


  not
  g216
  (
    n143,
    n52
  );


  not
  g217
  (
    n288,
    n89
  );


  not
  g218
  (
    n302,
    n53
  );


  not
  g219
  (
    n351,
    n28
  );


  buf
  g220
  (
    n298,
    n45
  );


  not
  g221
  (
    n115,
    n79
  );


  not
  g222
  (
    n239,
    n66
  );


  not
  g223
  (
    n128,
    n90
  );


  not
  g224
  (
    n203,
    n47
  );


  buf
  g225
  (
    n331,
    n91
  );


  buf
  g226
  (
    n184,
    n81
  );


  not
  g227
  (
    n332,
    n78
  );


  buf
  g228
  (
    n190,
    n86
  );


  buf
  g229
  (
    n368,
    n61
  );


  buf
  g230
  (
    n118,
    n65
  );


  buf
  g231
  (
    n168,
    n57
  );


  buf
  g232
  (
    n291,
    n82
  );


  not
  g233
  (
    n321,
    n71
  );


  not
  g234
  (
    n251,
    n65
  );


  buf
  g235
  (
    n338,
    n21
  );


  buf
  g236
  (
    n198,
    n47
  );


  not
  g237
  (
    n140,
    n39
  );


  not
  g238
  (
    n370,
    n44
  );


  buf
  g239
  (
    n286,
    n77
  );


  not
  g240
  (
    n181,
    n87
  );


  not
  g241
  (
    n154,
    n31
  );


  buf
  g242
  (
    n336,
    n56
  );


  buf
  g243
  (
    n379,
    n57
  );


  buf
  g244
  (
    n164,
    n77
  );


  not
  g245
  (
    n123,
    n43
  );


  buf
  g246
  (
    n316,
    n20
  );


  not
  g247
  (
    n133,
    n40
  );


  buf
  g248
  (
    n169,
    n33
  );


  not
  g249
  (
    n152,
    n72
  );


  buf
  g250
  (
    n98,
    n54
  );


  buf
  g251
  (
    n355,
    n71
  );


  buf
  g252
  (
    n241,
    n74
  );


  not
  g253
  (
    n328,
    n61
  );


  not
  g254
  (
    n171,
    n62
  );


  not
  g255
  (
    n194,
    n37
  );


  buf
  g256
  (
    n309,
    n80
  );


  buf
  g257
  (
    n124,
    n38
  );


  buf
  g258
  (
    n329,
    n64
  );


  not
  g259
  (
    n280,
    n84
  );


  not
  g260
  (
    n317,
    n67
  );


  not
  g261
  (
    n287,
    n61
  );


  buf
  g262
  (
    n213,
    n59
  );


  not
  g263
  (
    n220,
    n73
  );


  not
  g264
  (
    n344,
    n20
  );


  not
  g265
  (
    n306,
    n51
  );


  not
  g266
  (
    n327,
    n83
  );


  not
  g267
  (
    n206,
    n23
  );


  not
  g268
  (
    n320,
    n76
  );


  not
  g269
  (
    n142,
    n87
  );


  not
  g270
  (
    n246,
    n27
  );


  not
  g271
  (
    n103,
    n69
  );


  buf
  g272
  (
    n315,
    n33
  );


  not
  g273
  (
    n136,
    n34
  );


  not
  g274
  (
    n326,
    n73
  );


  buf
  g275
  (
    n337,
    n79
  );


  buf
  g276
  (
    n106,
    n91
  );


  buf
  g277
  (
    n282,
    n42
  );


  buf
  g278
  (
    n157,
    n29
  );


  buf
  g279
  (
    n372,
    n80
  );


  buf
  g280
  (
    n176,
    n26
  );


  not
  g281
  (
    n173,
    n29
  );


  buf
  g282
  (
    n349,
    n83
  );


  not
  g283
  (
    n197,
    n32
  );


  not
  g284
  (
    n299,
    n66
  );


  not
  g285
  (
    n382,
    n78
  );


  buf
  g286
  (
    n276,
    n72
  );


  not
  g287
  (
    n373,
    n36
  );


  buf
  g288
  (
    n365,
    n64
  );


  not
  g289
  (
    n300,
    n72
  );


  buf
  g290
  (
    n293,
    n65
  );


  not
  g291
  (
    n253,
    n78
  );


  not
  g292
  (
    n199,
    n42
  );


  buf
  g293
  (
    n196,
    n25
  );


  not
  g294
  (
    n289,
    n54
  );


  not
  g295
  (
    n150,
    n32
  );


  buf
  g296
  (
    n341,
    n75
  );


  not
  g297
  (
    n165,
    n53
  );


  not
  g298
  (
    n167,
    n64
  );


  buf
  g299
  (
    n264,
    n89
  );


  not
  g300
  (
    n149,
    n78
  );


  not
  g301
  (
    n278,
    n23
  );


  buf
  g302
  (
    n97,
    n65
  );


  not
  g303
  (
    n374,
    n53
  );


  buf
  g304
  (
    n347,
    n63
  );


  buf
  g305
  (
    n131,
    n84
  );


  not
  g306
  (
    n353,
    n85
  );


  buf
  g307
  (
    n178,
    n56
  );


  buf
  g308
  (
    n96,
    n30
  );


  buf
  g309
  (
    n179,
    n72
  );


  not
  g310
  (
    n218,
    n29
  );


  not
  g311
  (
    n215,
    n27
  );


  buf
  g312
  (
    n367,
    n86
  );


  not
  g313
  (
    n208,
    n39
  );


  buf
  g314
  (
    n305,
    n91
  );


  not
  g315
  (
    n277,
    n81
  );


  buf
  g316
  (
    n155,
    n58
  );


  buf
  g317
  (
    n356,
    n41
  );


  not
  g318
  (
    n230,
    n52
  );


  buf
  g319
  (
    n360,
    n35
  );


  not
  g320
  (
    n221,
    n62
  );


  buf
  g321
  (
    n224,
    n27
  );


  not
  g322
  (
    n283,
    n89
  );


  not
  g323
  (
    n145,
    n58
  );


  buf
  g324
  (
    n294,
    n37
  );


  not
  g325
  (
    n102,
    n26
  );


  not
  g326
  (
    n363,
    n73
  );


  not
  g327
  (
    n268,
    n48
  );


  not
  g328
  (
    n237,
    n68
  );


  buf
  g329
  (
    n107,
    n21
  );


  not
  g330
  (
    n113,
    n51
  );


  buf
  g331
  (
    n375,
    n88
  );


  buf
  g332
  (
    n235,
    n79
  );


  buf
  g333
  (
    n304,
    n26
  );


  not
  g334
  (
    n174,
    n83
  );


  not
  g335
  (
    n129,
    n68
  );


  buf
  g336
  (
    n233,
    n33
  );


  buf
  g337
  (
    n258,
    n38
  );


  not
  g338
  (
    n377,
    n62
  );


  buf
  g339
  (
    n187,
    n57
  );


  buf
  g340
  (
    n186,
    n57
  );


  not
  g341
  (
    n144,
    n63
  );


  buf
  g342
  (
    n381,
    n79
  );


  buf
  g343
  (
    n138,
    n69
  );


  buf
  g344
  (
    n292,
    n90
  );


  buf
  g345
  (
    n275,
    n44
  );


  not
  g346
  (
    n362,
    n60
  );


  buf
  g347
  (
    n217,
    n81
  );


  not
  g348
  (
    n141,
    n76
  );


  buf
  g349
  (
    n211,
    n25
  );


  not
  g350
  (
    n166,
    n55
  );


  not
  g351
  (
    n354,
    n50
  );


  buf
  g352
  (
    n222,
    n20
  );


  buf
  g353
  (
    n358,
    n83
  );


  not
  g354
  (
    n130,
    n41
  );


  not
  g355
  (
    n204,
    n28
  );


  not
  g356
  (
    n273,
    n52
  );


  not
  g357
  (
    n232,
    n27
  );


  not
  g358
  (
    n209,
    n90
  );


  buf
  g359
  (
    n223,
    n75
  );


  buf
  g360
  (
    n185,
    n48
  );


  buf
  g361
  (
    n270,
    n49
  );


  buf
  g362
  (
    n156,
    n44
  );


  buf
  g363
  (
    n493,
    n134
  );


  buf
  g364
  (
    n496,
    n101
  );


  buf
  g365
  (
    n428,
    n107
  );


  not
  g366
  (
    n384,
    n208
  );


  buf
  g367
  (
    n441,
    n129
  );


  not
  g368
  (
    n474,
    n123
  );


  not
  g369
  (
    n407,
    n138
  );


  buf
  g370
  (
    n383,
    n111
  );


  not
  g371
  (
    n410,
    n113
  );


  buf
  g372
  (
    n417,
    n136
  );


  not
  g373
  (
    n397,
    n195
  );


  not
  g374
  (
    n477,
    n178
  );


  buf
  g375
  (
    n473,
    n110
  );


  not
  g376
  (
    n448,
    n96
  );


  not
  g377
  (
    n423,
    n179
  );


  buf
  g378
  (
    n475,
    n186
  );


  not
  g379
  (
    n454,
    n166
  );


  buf
  g380
  (
    n486,
    n102
  );


  buf
  g381
  (
    n433,
    n106
  );


  not
  g382
  (
    n459,
    n148
  );


  buf
  g383
  (
    n395,
    n172
  );


  not
  g384
  (
    n430,
    n205
  );


  not
  g385
  (
    n385,
    n156
  );


  buf
  g386
  (
    n472,
    n190
  );


  not
  g387
  (
    n398,
    n127
  );


  not
  g388
  (
    n427,
    n118
  );


  not
  g389
  (
    n403,
    n109
  );


  buf
  g390
  (
    n438,
    n206
  );


  not
  g391
  (
    n451,
    n202
  );


  not
  g392
  (
    n396,
    n177
  );


  not
  g393
  (
    n445,
    n146
  );


  buf
  g394
  (
    n484,
    n188
  );


  buf
  g395
  (
    n447,
    n126
  );


  buf
  g396
  (
    n411,
    n97
  );


  buf
  g397
  (
    n388,
    n122
  );


  not
  g398
  (
    n401,
    n204
  );


  buf
  g399
  (
    n429,
    n100
  );


  buf
  g400
  (
    n476,
    n198
  );


  not
  g401
  (
    n482,
    n183
  );


  buf
  g402
  (
    n439,
    n163
  );


  not
  g403
  (
    n400,
    n170
  );


  buf
  g404
  (
    n444,
    n191
  );


  buf
  g405
  (
    n487,
    n207
  );


  buf
  g406
  (
    n413,
    n193
  );


  buf
  g407
  (
    n479,
    n135
  );


  not
  g408
  (
    n471,
    n174
  );


  not
  g409
  (
    n489,
    n209
  );


  buf
  g410
  (
    n440,
    n168
  );


  not
  g411
  (
    n488,
    n104
  );


  buf
  g412
  (
    n421,
    n200
  );


  buf
  g413
  (
    n463,
    n171
  );


  buf
  g414
  (
    n446,
    n120
  );


  not
  g415
  (
    n394,
    n133
  );


  buf
  g416
  (
    n412,
    n162
  );


  not
  g417
  (
    n453,
    n128
  );


  buf
  g418
  (
    n452,
    n151
  );


  not
  g419
  (
    n460,
    n119
  );


  buf
  g420
  (
    n478,
    n192
  );


  not
  g421
  (
    n455,
    n203
  );


  not
  g422
  (
    n422,
    n189
  );


  not
  g423
  (
    n409,
    n181
  );


  not
  g424
  (
    n464,
    n141
  );


  buf
  g425
  (
    n490,
    n167
  );


  not
  g426
  (
    n443,
    n132
  );


  buf
  g427
  (
    n420,
    n196
  );


  buf
  g428
  (
    n461,
    n152
  );


  not
  g429
  (
    n434,
    n153
  );


  not
  g430
  (
    n470,
    n98
  );


  not
  g431
  (
    n457,
    n160
  );


  not
  g432
  (
    n492,
    n155
  );


  buf
  g433
  (
    n469,
    n164
  );


  buf
  g434
  (
    n418,
    n149
  );


  buf
  g435
  (
    n467,
    n161
  );


  not
  g436
  (
    n416,
    n142
  );


  not
  g437
  (
    n495,
    n115
  );


  buf
  g438
  (
    n392,
    n103
  );


  buf
  g439
  (
    n432,
    n150
  );


  buf
  g440
  (
    n419,
    n199
  );


  buf
  g441
  (
    n481,
    n185
  );


  not
  g442
  (
    n437,
    n180
  );


  not
  g443
  (
    n480,
    n112
  );


  not
  g444
  (
    n415,
    n182
  );


  buf
  g445
  (
    n431,
    n157
  );


  buf
  g446
  (
    n390,
    n154
  );


  not
  g447
  (
    n386,
    n173
  );


  buf
  g448
  (
    n425,
    n99
  );


  not
  g449
  (
    n414,
    n158
  );


  buf
  g450
  (
    n435,
    n175
  );


  not
  g451
  (
    n442,
    n130
  );


  not
  g452
  (
    n402,
    n184
  );


  buf
  g453
  (
    n462,
    n147
  );


  buf
  g454
  (
    n391,
    n131
  );


  buf
  g455
  (
    n456,
    n187
  );


  buf
  g456
  (
    n408,
    n121
  );


  buf
  g457
  (
    n436,
    n159
  );


  buf
  g458
  (
    n491,
    n108
  );


  not
  g459
  (
    n387,
    n124
  );


  not
  g460
  (
    n494,
    n145
  );


  not
  g461
  (
    n449,
    n117
  );


  buf
  g462
  (
    n458,
    n143
  );


  buf
  g463
  (
    n405,
    n144
  );


  not
  g464
  (
    n404,
    n125
  );


  not
  g465
  (
    n483,
    n169
  );


  buf
  g466
  (
    n468,
    n197
  );


  buf
  g467
  (
    n465,
    n137
  );


  buf
  g468
  (
    n399,
    n114
  );


  buf
  g469
  (
    n424,
    n140
  );


  buf
  g470
  (
    n393,
    n116
  );


  buf
  g471
  (
    n450,
    n201
  );


  buf
  g472
  (
    n426,
    n105
  );


  not
  g473
  (
    n466,
    n194
  );


  buf
  g474
  (
    n406,
    n165
  );


  not
  g475
  (
    n485,
    n176
  );


  buf
  g476
  (
    n389,
    n139
  );


  or
  g477
  (
    n501,
    n423,
    n417,
    n386,
    n416
  );


  nand
  g478
  (
    n518,
    n413,
    n387,
    n391,
    n403
  );


  xor
  g479
  (
    n508,
    n420,
    n385,
    n425,
    n394
  );


  and
  g480
  (
    n510,
    n422,
    n397,
    n393,
    n390
  );


  nand
  g481
  (
    n511,
    n408,
    n419,
    n389,
    n406
  );


  nand
  g482
  (
    n507,
    n399,
    n415,
    n422,
    n384
  );


  xnor
  g483
  (
    n500,
    n412,
    n397,
    n387,
    n392
  );


  xor
  g484
  (
    n515,
    n386,
    n405,
    n425,
    n407
  );


  nand
  g485
  (
    n505,
    n409,
    n409,
    n408,
    n388
  );


  nand
  g486
  (
    n498,
    n418,
    n398,
    n399,
    n407
  );


  nor
  g487
  (
    n509,
    n394,
    n412,
    n393,
    n402
  );


  and
  g488
  (
    n506,
    n417,
    n426,
    n398,
    n411
  );


  or
  g489
  (
    n503,
    n388,
    n413,
    n400
  );


  xnor
  g490
  (
    n497,
    n384,
    n396,
    n427,
    n410
  );


  or
  g491
  (
    n517,
    n396,
    n406,
    n418,
    n421
  );


  xnor
  g492
  (
    n513,
    n395,
    n421,
    n416,
    n426
  );


  or
  g493
  (
    n499,
    n404,
    n385,
    n420,
    n403
  );


  xnor
  g494
  (
    n502,
    n390,
    n424,
    n404,
    n401
  );


  or
  g495
  (
    n516,
    n391,
    n419,
    n415,
    n423
  );


  nor
  g496
  (
    n512,
    n410,
    n401,
    n383,
    n392
  );


  nand
  g497
  (
    n504,
    n389,
    n402,
    n414,
    n405
  );


  nand
  g498
  (
    n514,
    n395,
    n411,
    n414,
    n424
  );


  buf
  g499
  (
    n522,
    n499
  );


  buf
  g500
  (
    n528,
    n504
  );


  not
  g501
  (
    n523,
    n502
  );


  not
  g502
  (
    n521,
    n507
  );


  buf
  g503
  (
    n520,
    n500
  );


  not
  g504
  (
    n519,
    n498
  );


  not
  g505
  (
    n527,
    n501
  );


  not
  g506
  (
    n525,
    n506
  );


  buf
  g507
  (
    n524,
    n503
  );


  xor
  g508
  (
    n526,
    n505,
    n497
  );


  not
  g509
  (
    n537,
    n524
  );


  buf
  g510
  (
    n531,
    n520
  );


  buf
  g511
  (
    n533,
    n521
  );


  buf
  g512
  (
    n536,
    n523
  );


  not
  g513
  (
    n532,
    n525
  );


  not
  g514
  (
    n529,
    n522
  );


  buf
  g515
  (
    n535,
    n519
  );


  buf
  g516
  (
    n534,
    n527
  );


  not
  g517
  (
    n530,
    n526
  );


  not
  g518
  (
    n542,
    n214
  );


  buf
  g519
  (
    n546,
    n533
  );


  xnor
  g520
  (
    n539,
    n229,
    n530,
    n213,
    n242
  );


  xnor
  g521
  (
    n550,
    n235,
    n210,
    n530,
    n220
  );


  and
  g522
  (
    n548,
    n225,
    n238,
    n221,
    n533
  );


  xor
  g523
  (
    n544,
    n234,
    n532,
    n228
  );


  xnor
  g524
  (
    n540,
    n240,
    n239,
    n534,
    n212
  );


  xnor
  g525
  (
    n547,
    n223,
    n232,
    n237,
    n533
  );


  nand
  g526
  (
    n538,
    n211,
    n224,
    n215,
    n533
  );


  or
  g527
  (
    n545,
    n230,
    n529,
    n218,
    n227
  );


  or
  g528
  (
    n549,
    n241,
    n219,
    n531,
    n217
  );


  or
  g529
  (
    n541,
    n236,
    n216,
    n226,
    n531
  );


  nor
  g530
  (
    n543,
    n222,
    n534,
    n233,
    n231
  );


  nand
  g531
  (
    n562,
    n445,
    n538,
    n543,
    n430
  );


  nand
  g532
  (
    n554,
    n244,
    n445,
    n539,
    n439
  );


  nand
  g533
  (
    n560,
    n541,
    n443,
    n540,
    n428
  );


  xor
  g534
  (
    n557,
    n544,
    n443,
    n542,
    n245
  );


  or
  g535
  (
    n558,
    n444,
    n541,
    n441,
    n538
  );


  nor
  g536
  (
    n552,
    n543,
    n431,
    n247,
    n539
  );


  nor
  g537
  (
    n551,
    n429,
    n540,
    n440,
    n434
  );


  xor
  g538
  (
    n559,
    n435,
    n436,
    n440,
    n446
  );


  or
  g539
  (
    n555,
    n433,
    n442,
    n432,
    n542
  );


  or
  g540
  (
    n561,
    n544,
    n437,
    n246,
    n248
  );


  and
  g541
  (
    n564,
    n434,
    n442,
    n545,
    n437
  );


  xor
  g542
  (
    n563,
    n441,
    n430,
    n428,
    n433
  );


  and
  g543
  (
    n565,
    n439,
    n429,
    n243,
    n427
  );


  nor
  g544
  (
    n553,
    n436,
    n431,
    n432,
    n435
  );


  nand
  g545
  (
    n556,
    n446,
    n438,
    n444
  );


  xnor
  g546
  (
    n569,
    n563,
    n565,
    n553,
    n253
  );


  nand
  g547
  (
    n581,
    n551,
    n272,
    n258,
    n289
  );


  xor
  g548
  (
    n577,
    n264,
    n259,
    n260,
    n292
  );


  nor
  g549
  (
    n566,
    n254,
    n564,
    n558,
    n559
  );


  xor
  g550
  (
    n575,
    n556,
    n280,
    n285,
    n279
  );


  nor
  g551
  (
    n576,
    n283,
    n273,
    n261,
    n278
  );


  xor
  g552
  (
    n580,
    n267,
    n266,
    n296,
    n557
  );


  xor
  g553
  (
    n579,
    n269,
    n562,
    n277,
    n560
  );


  nor
  g554
  (
    n578,
    n270,
    n286,
    n565,
    n555
  );


  nand
  g555
  (
    n567,
    n295,
    n282,
    n256,
    n255
  );


  or
  g556
  (
    n574,
    n291,
    n249,
    n271,
    n288
  );


  and
  g557
  (
    n570,
    n268,
    n275,
    n265,
    n294
  );


  xor
  g558
  (
    n572,
    n257,
    n561,
    n284,
    n274
  );


  xor
  g559
  (
    n571,
    n552,
    n251,
    n262,
    n293
  );


  nor
  g560
  (
    n573,
    n554,
    n290,
    n281,
    n250
  );


  or
  g561
  (
    n568,
    n252,
    n263,
    n276,
    n287
  );


  buf
  g562
  (
    n613,
    n450
  );


  buf
  g563
  (
    n619,
    n476
  );


  buf
  g564
  (
    n607,
    n473
  );


  not
  g565
  (
    n597,
    n570
  );


  not
  g566
  (
    n609,
    n573
  );


  not
  g567
  (
    n594,
    n453
  );


  buf
  g568
  (
    n588,
    n465
  );


  buf
  g569
  (
    n623,
    n576
  );


  buf
  g570
  (
    n617,
    n458
  );


  not
  g571
  (
    n601,
    n460
  );


  not
  g572
  (
    n583,
    n567
  );


  not
  g573
  (
    n602,
    n465
  );


  buf
  g574
  (
    n608,
    n572
  );


  not
  g575
  (
    n626,
    n468
  );


  not
  g576
  (
    n598,
    n451
  );


  not
  g577
  (
    n604,
    n458
  );


  xor
  g578
  (
    n621,
    n471,
    n468
  );


  nand
  g579
  (
    n620,
    n469,
    n572,
    n452,
    n463
  );


  xor
  g580
  (
    n618,
    n478,
    n472,
    n484,
    n464
  );


  nor
  g581
  (
    n589,
    n460,
    n575,
    n482,
    n566
  );


  or
  g582
  (
    n593,
    n489,
    n568,
    n455,
    n478
  );


  xnor
  g583
  (
    n603,
    n487,
    n570,
    n566,
    n568
  );


  xor
  g584
  (
    n610,
    n575,
    n574,
    n450,
    n571
  );


  xor
  g585
  (
    n615,
    n453,
    n566,
    n492,
    n569
  );


  nor
  g586
  (
    n611,
    n576,
    n467,
    n569
  );


  nand
  g587
  (
    n595,
    n470,
    n577,
    n483,
    n459
  );


  nand
  g588
  (
    n587,
    n577,
    n571,
    n463,
    n459
  );


  or
  g589
  (
    n614,
    n487,
    n448,
    n477,
    n485
  );


  nand
  g590
  (
    n605,
    n488,
    n572,
    n452,
    n569
  );


  nor
  g591
  (
    n627,
    n451,
    n569,
    n457,
    n567
  );


  xor
  g592
  (
    n592,
    n568,
    n573,
    n570,
    n477
  );


  nand
  g593
  (
    n628,
    n577,
    n462,
    n574,
    n479
  );


  or
  g594
  (
    n599,
    n456,
    n490,
    n447,
    n480
  );


  or
  g595
  (
    n586,
    n568,
    n474,
    n567,
    n489
  );


  xor
  g596
  (
    n591,
    n574,
    n461,
    n466,
    n475
  );


  nor
  g597
  (
    n590,
    n469,
    n449,
    n472,
    n576
  );


  or
  g598
  (
    n585,
    n479,
    n571,
    n481
  );


  xnor
  g599
  (
    n596,
    n490,
    n572,
    n475,
    n575
  );


  or
  g600
  (
    n582,
    n456,
    n576,
    n574,
    n491
  );


  xnor
  g601
  (
    n584,
    n470,
    n571,
    n454,
    n573
  );


  xor
  g602
  (
    n600,
    n567,
    n471,
    n491,
    n575
  );


  or
  g603
  (
    n616,
    n447,
    n455,
    n573,
    n486
  );


  nor
  g604
  (
    n612,
    n464,
    n474,
    n473,
    n482
  );


  and
  g605
  (
    n606,
    n485,
    n454,
    n476,
    n577
  );


  xnor
  g606
  (
    n622,
    n483,
    n449,
    n484,
    n570
  );


  nor
  g607
  (
    n624,
    n488,
    n462,
    n457,
    n486
  );


  or
  g608
  (
    n625,
    n448,
    n466,
    n461,
    n480
  );


  not
  g609
  (
    n630,
    n591
  );


  buf
  g610
  (
    n635,
    n584
  );


  not
  g611
  (
    n633,
    n597
  );


  not
  g612
  (
    n638,
    n583
  );


  not
  g613
  (
    n629,
    n598
  );


  buf
  g614
  (
    n637,
    n593
  );


  nor
  g615
  (
    n631,
    n589,
    n590
  );


  and
  g616
  (
    n636,
    n587,
    n596,
    n595,
    n598
  );


  xnor
  g617
  (
    n634,
    n596,
    n586,
    n592,
    n594
  );


  or
  g618
  (
    n632,
    n595,
    n588,
    n597,
    n585
  );


  buf
  g619
  (
    n642,
    n606
  );


  buf
  g620
  (
    n647,
    n606
  );


  nor
  g621
  (
    n641,
    n637,
    n610
  );


  nand
  g622
  (
    n640,
    n631,
    n630,
    n607,
    n632
  );


  xnor
  g623
  (
    n648,
    n638,
    n603,
    n599,
    n602
  );


  nor
  g624
  (
    n649,
    n492,
    n638,
    n602,
    n600
  );


  nand
  g625
  (
    n646,
    n604,
    n599,
    n600,
    n608
  );


  or
  g626
  (
    n639,
    n607,
    n601,
    n610
  );


  nor
  g627
  (
    n643,
    n603,
    n605,
    n608,
    n635
  );


  xor
  g628
  (
    n644,
    n604,
    n609,
    n605
  );


  and
  g629
  (
    n645,
    n633,
    n629,
    n634,
    n636
  );


  not
  g630
  (
    n666,
    n643
  );


  not
  g631
  (
    n670,
    n308
  );


  buf
  g632
  (
    n657,
    n322
  );


  not
  g633
  (
    n678,
    n508
  );


  not
  g634
  (
    n689,
    n642
  );


  buf
  g635
  (
    n668,
    n309
  );


  not
  g636
  (
    n677,
    n611
  );


  buf
  g637
  (
    n671,
    n648
  );


  not
  g638
  (
    n655,
    n647
  );


  not
  g639
  (
    n676,
    n641
  );


  not
  g640
  (
    n669,
    n649
  );


  not
  g641
  (
    n674,
    n648
  );


  buf
  g642
  (
    n662,
    n644
  );


  not
  g643
  (
    n651,
    n319
  );


  buf
  g644
  (
    n686,
    n327
  );


  not
  g645
  (
    n681,
    n645
  );


  buf
  g646
  (
    n656,
    n303
  );


  not
  g647
  (
    n688,
    n649
  );


  buf
  g648
  (
    n690,
    n640
  );


  not
  g649
  (
    n665,
    n644
  );


  not
  g650
  (
    n658,
    n611
  );


  buf
  g651
  (
    n683,
    n647
  );


  buf
  g652
  (
    n679,
    n616
  );


  buf
  g653
  (
    n692,
    n645
  );


  not
  g654
  (
    n652,
    n648
  );


  not
  g655
  (
    n663,
    n318
  );


  nor
  g656
  (
    n673,
    n644,
    n639
  );


  nor
  g657
  (
    n672,
    n617,
    n613,
    n534,
    n301
  );


  xnor
  g658
  (
    n661,
    n512,
    n614,
    n314,
    n642
  );


  xnor
  g659
  (
    n687,
    n649,
    n614,
    n640,
    n325
  );


  xnor
  g660
  (
    n653,
    n513,
    n643,
    n645,
    n305
  );


  nand
  g661
  (
    n680,
    n640,
    n641,
    n509,
    n647
  );


  and
  g662
  (
    n650,
    n615,
    n320,
    n317,
    n311
  );


  nand
  g663
  (
    n660,
    n315,
    n612,
    n298
  );


  nor
  g664
  (
    n691,
    n639,
    n645,
    n646,
    n321
  );


  or
  g665
  (
    n675,
    n534,
    n299,
    n313,
    n312
  );


  and
  g666
  (
    n684,
    n642,
    n646,
    n511,
    n310
  );


  xnor
  g667
  (
    n667,
    n640,
    n326,
    n641,
    n324
  );


  and
  g668
  (
    n664,
    n510,
    n297,
    n646,
    n316
  );


  nand
  g669
  (
    n685,
    n647,
    n306,
    n646,
    n323
  );


  or
  g670
  (
    n693,
    n307,
    n649,
    n643,
    n304
  );


  and
  g671
  (
    n654,
    n644,
    n615,
    n616,
    n639
  );


  nor
  g672
  (
    n659,
    n643,
    n642,
    n613,
    n641
  );


  xnor
  g673
  (
    n682,
    n300,
    n639,
    n648,
    n302
  );


  buf
  g674
  (
    n710,
    n336
  );


  buf
  g675
  (
    n728,
    n674
  );


  buf
  g676
  (
    n734,
    n680
  );


  buf
  g677
  (
    n711,
    n535
  );


  not
  g678
  (
    n736,
    n496
  );


  buf
  g679
  (
    n703,
    n659
  );


  buf
  g680
  (
    n696,
    n665
  );


  not
  g681
  (
    n733,
    n689
  );


  buf
  g682
  (
    n708,
    n670
  );


  not
  g683
  (
    n724,
    n494
  );


  buf
  g684
  (
    n741,
    n618
  );


  buf
  g685
  (
    n718,
    n536
  );


  not
  g686
  (
    n705,
    n536
  );


  not
  g687
  (
    n697,
    n658
  );


  not
  g688
  (
    n720,
    n693
  );


  not
  g689
  (
    n706,
    n681
  );


  xnor
  g690
  (
    n699,
    n656,
    n683
  );


  xnor
  g691
  (
    n716,
    n679,
    n686,
    n682,
    n662
  );


  nand
  g692
  (
    n702,
    n673,
    n545,
    n680,
    n332
  );


  nand
  g693
  (
    n719,
    n536,
    n518,
    n687,
    n671
  );


  and
  g694
  (
    n713,
    n339,
    n328,
    n653,
    n514
  );


  nor
  g695
  (
    n709,
    n537,
    n689,
    n676,
    n549
  );


  nand
  g696
  (
    n739,
    n684,
    n692,
    n579,
    n650
  );


  nor
  g697
  (
    n725,
    n677,
    n495,
    n651,
    n493
  );


  xnor
  g698
  (
    n715,
    n618,
    n338,
    n688,
    n546
  );


  xor
  g699
  (
    n722,
    n342,
    n550,
    n330,
    n678
  );


  xnor
  g700
  (
    n695,
    n578,
    n684,
    n516,
    n580
  );


  xnor
  g701
  (
    n737,
    n537,
    n621,
    n691
  );


  xnor
  g702
  (
    n738,
    n578,
    n334,
    n495,
    n654
  );


  xnor
  g703
  (
    n700,
    n675,
    n580,
    n617,
    n579
  );


  nand
  g704
  (
    n723,
    n691,
    n682,
    n528,
    n331
  );


  xor
  g705
  (
    n714,
    n579,
    n547,
    n535,
    n620
  );


  nor
  g706
  (
    n727,
    n676,
    n536,
    n664,
    n672
  );


  nor
  g707
  (
    n704,
    n335,
    n620,
    n578,
    n344
  );


  nand
  g708
  (
    n698,
    n579,
    n546,
    n687,
    n535
  );


  nand
  g709
  (
    n701,
    n580,
    n690,
    n581,
    n679
  );


  xnor
  g710
  (
    n726,
    n681,
    n581,
    n693,
    n91
  );


  xnor
  g711
  (
    n735,
    n580,
    n669,
    n667,
    n494
  );


  xnor
  g712
  (
    n717,
    n690,
    n550,
    n581,
    n677
  );


  nand
  g713
  (
    n730,
    n652,
    n329,
    n663,
    n678
  );


  nor
  g714
  (
    n740,
    n537,
    n581,
    n333,
    n340
  );


  xnor
  g715
  (
    n732,
    n661,
    n578,
    n493,
    n548
  );


  or
  g716
  (
    n712,
    n657,
    n692,
    n337,
    n686
  );


  xnor
  g717
  (
    n729,
    n619,
    n549,
    n683,
    n537
  );


  and
  g718
  (
    n694,
    n548,
    n341,
    n666,
    n517
  );


  nor
  g719
  (
    n731,
    n660,
    n515,
    n619,
    n535
  );


  or
  g720
  (
    n721,
    n343,
    n668,
    n688,
    n685
  );


  nor
  g721
  (
    n707,
    n685,
    n496,
    n547,
    n655
  );


  not
  g722
  (
    n744,
    n694
  );


  buf
  g723
  (
    n742,
    n696
  );


  xor
  g724
  (
    n743,
    n695,
    n697
  );


  or
  g725
  (
    n745,
    n744,
    n742,
    n743
  );


  not
  g726
  (
    n746,
    n745
  );


  not
  g727
  (
    n747,
    n745
  );


  not
  g728
  (
    n755,
    n746
  );


  not
  g729
  (
    n749,
    n746
  );


  not
  g730
  (
    n753,
    n747
  );


  not
  g731
  (
    n751,
    n746
  );


  buf
  g732
  (
    n748,
    n746
  );


  not
  g733
  (
    n750,
    n747
  );


  buf
  g734
  (
    n752,
    n747
  );


  not
  g735
  (
    n754,
    n747
  );


  nor
  g736
  (
    n770,
    n626,
    n703,
    n748,
    n713
  );


  or
  g737
  (
    n760,
    n729,
    n705,
    n626,
    n727
  );


  and
  g738
  (
    AntiSAT_key_wire,
    n754,
    n721,
    n753,
    n752
  );


  xnor
  g739
  (
    n758,
    n750,
    n708,
    n719,
    n753
  );


  or
  g740
  (
    n762,
    n720,
    n710,
    n716,
    n699
  );


  nand
  g741
  (
    n768,
    n623,
    n711,
    n751,
    n715
  );


  and
  g742
  (
    n771,
    n755,
    n702,
    n725,
    n751
  );


  or
  g743
  (
    n763,
    n622,
    n714,
    n754,
    n700
  );


  nand
  g744
  (
    n766,
    n712,
    n717,
    n730,
    n698
  );


  and
  g745
  (
    n767,
    n624,
    n709,
    n752,
    n724
  );


  nor
  g746
  (
    n756,
    n728,
    n750,
    n726,
    n731
  );


  nand
  g747
  (
    n761,
    n749,
    n701,
    n754,
    n723
  );


  and
  g748
  (
    n769,
    n749,
    n748,
    n718,
    n707
  );


  or
  g749
  (
    n757,
    n755,
    n623,
    n624,
    n704
  );


  xor
  g750
  (
    n759,
    n722,
    n625,
    n755,
    n706
  );


  nor
  g751
  (
    n765,
    n755,
    n622,
    n625,
    n732
  );


  not
  g752
  (
    n773,
    n767
  );


  buf
  g753
  (
    n775,
    n770
  );


  not
  g754
  (
    n776,
    n771
  );


  buf
  g755
  (
    n772,
    n345
  );


  nand
  g756
  (
    n774,
    n768,
    n769
  );


  buf
  g757
  (
    n789,
    n346
  );


  buf
  g758
  (
    n777,
    n776
  );


  not
  g759
  (
    n787,
    n93
  );


  not
  g760
  (
    n792,
    n92
  );


  buf
  g761
  (
    n793,
    n351
  );


  not
  g762
  (
    n778,
    n774
  );


  not
  g763
  (
    n784,
    n354
  );


  buf
  g764
  (
    n791,
    n93
  );


  xnor
  g765
  (
    n794,
    n773,
    n353
  );


  or
  g766
  (
    n783,
    n94,
    n734,
    n735,
    n347
  );


  or
  g767
  (
    n779,
    n348,
    n352,
    n95,
    n772
  );


  xor
  g768
  (
    n790,
    n93,
    n94,
    n92,
    n776
  );


  xor
  g769
  (
    n786,
    n94,
    n776,
    n349,
    n92
  );


  or
  g770
  (
    n788,
    n774,
    n775,
    n773
  );


  nand
  g771
  (
    n781,
    n773,
    n94,
    n772,
    n775
  );


  xor
  g772
  (
    n785,
    n93,
    n95,
    n774
  );


  nand
  g773
  (
    n782,
    n773,
    n774,
    n95,
    n775
  );


  nor
  g774
  (
    n780,
    n733,
    n350,
    n776,
    n92
  );


  not
  g775
  (
    n795,
    n778
  );


  not
  g776
  (
    n798,
    n779
  );


  buf
  g777
  (
    n797,
    n780
  );


  not
  g778
  (
    n796,
    n777
  );


  nand
  g779
  (
    n799,
    n781,
    n797,
    n798,
    n780
  );


  buf
  g780
  (
    n800,
    n799
  );


  buf
  g781
  (
    n801,
    n799
  );


  not
  g782
  (
    n803,
    n801
  );


  and
  g783
  (
    n802,
    n801,
    n800,
    n355
  );


  and
  g784
  (
    n804,
    n801,
    n357,
    n800,
    n356
  );


  nand
  g785
  (
    n805,
    n804,
    n782,
    n781
  );


  buf
  g786
  (
    n807,
    n805
  );


  not
  g787
  (
    n809,
    n784
  );


  nand
  g788
  (
    n808,
    n783,
    n358,
    n805,
    n785
  );


  nand
  g789
  (
    n806,
    n784,
    n783,
    n805
  );


  buf
  g790
  (
    n810,
    n806
  );


  not
  g791
  (
    n811,
    n806
  );


  or
  g792
  (
    n812,
    n811,
    n359
  );


  buf
  g793
  (
    n814,
    n812
  );


  buf
  g794
  (
    n813,
    n812
  );


  and
  g795
  (
    n815,
    n785,
    n786,
    n812
  );


  and
  g796
  (
    n816,
    n814,
    n787,
    n788,
    n815
  );


  nor
  g797
  (
    n817,
    n788,
    n627,
    n787,
    n786
  );


  nand
  g798
  (
    n819,
    n807,
    n807,
    n816,
    n366
  );


  and
  g799
  (
    n825,
    n361,
    n365,
    n808,
    n809
  );


  xnor
  g800
  (
    n820,
    n360,
    n809,
    n817
  );


  xor
  g801
  (
    n821,
    n370,
    n816,
    n807
  );


  xnor
  g802
  (
    n818,
    n364,
    n817,
    n368,
    n816
  );


  xnor
  g803
  (
    n823,
    n369,
    n808,
    n362,
    n809
  );


  xor
  g804
  (
    n822,
    n808,
    n808,
    n627,
    n817
  );


  xnor
  g805
  (
    n824,
    n807,
    n367,
    n363,
    n817
  );


  or
  g806
  (
    n827,
    n823,
    n825,
    n824
  );


  nand
  g807
  (
    n826,
    n822,
    n821,
    n824,
    n820
  );


  xnor
  g808
  (
    n828,
    n819,
    n371,
    n372,
    n818
  );


  xor
  g809
  (
    n830,
    n790,
    n789,
    n828
  );


  nor
  g810
  (
    n829,
    n827,
    n790,
    n791
  );


  or
  g811
  (
    n832,
    n793,
    n830,
    n738,
    n792
  );


  or
  g812
  (
    n831,
    n829,
    n793,
    n736,
    n830
  );


  nor
  g813
  (
    n833,
    n830,
    n830,
    n737,
    n792
  );


  and
  g814
  (
    n834,
    n374,
    n373,
    n628,
    n833
  );


  or
  g815
  (
    n837,
    n376,
    n375,
    n380,
    n382
  );


  nand
  g816
  (
    n836,
    n381,
    n834,
    n379,
    n377
  );


  nor
  g817
  (
    n838,
    n739,
    n740,
    n834,
    n628
  );


  xor
  g818
  (
    n835,
    n794,
    n378,
    n834
  );


  nand
  g819
  (
    n839,
    n837,
    n837,
    n838,
    n836
  );


  and
  g820
  (
    n840,
    n741,
    n835,
    n838,
    n794
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_19
  (
    gbar_input_0_0,
    keyIn_0_19,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_20
  (
    gbar_input_0_1,
    keyIn_0_20,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_21
  (
    gbar_input_0_2,
    keyIn_0_21,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_22
  (
    gbar_input_0_3,
    keyIn_0_22,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_23
  (
    gbar_input_0_4,
    keyIn_0_23,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_24
  (
    gbar_input_0_5,
    keyIn_0_24,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_25
  (
    gbar_input_0_6,
    keyIn_0_25,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_26
  (
    gbar_input_0_7,
    keyIn_0_26,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_27
  (
    gbar_input_0_8,
    keyIn_0_27,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_28
  (
    gbar_input_0_9,
    keyIn_0_28,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_10,
    keyIn_0_29,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_11,
    keyIn_0_30,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_12,
    keyIn_0_31,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_13,
    keyIn_0_32,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_14,
    keyIn_0_33,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_15,
    keyIn_0_34,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_16,
    keyIn_0_35,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_17,
    keyIn_0_36,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_18,
    keyIn_0_37,
    n19
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n764,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

