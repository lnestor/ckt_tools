

module Stat_3000_324
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2639,
  n2629,
  n2634,
  n2631,
  n2633,
  n2626,
  n2637,
  n2628,
  n2627,
  n2642,
  n2640,
  n2643,
  n2823,
  n2831,
  n2828,
  n2827,
  n2817,
  n2842,
  n2833,
  n2829,
  n2815,
  n2825,
  n3032,
  n3026,
  n3028,
  n3023,
  n3025,
  n3030,
  n3031,
  n3027,
  n3024,
  n3029,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n2639;
  output n2629;
  output n2634;
  output n2631;
  output n2633;
  output n2626;
  output n2637;
  output n2628;
  output n2627;
  output n2642;
  output n2640;
  output n2643;
  output n2823;
  output n2831;
  output n2828;
  output n2827;
  output n2817;
  output n2842;
  output n2833;
  output n2829;
  output n2815;
  output n2825;
  output n3032;
  output n3026;
  output n3028;
  output n3023;
  output n3025;
  output n3030;
  output n3031;
  output n3027;
  output n3024;
  output n3029;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2630;
  wire n2632;
  wire n2635;
  wire n2636;
  wire n2638;
  wire n2641;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2816;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2824;
  wire n2826;
  wire n2830;
  wire n2832;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    KeyWire_0_42,
    n18
  );


  buf
  g1
  (
    n154,
    n9
  );


  not
  g2
  (
    n94,
    n30
  );


  not
  g3
  (
    n144,
    n20
  );


  not
  g4
  (
    n142,
    n15
  );


  not
  g5
  (
    n63,
    n9
  );


  not
  g6
  (
    n155,
    n14
  );


  buf
  g7
  (
    n122,
    n11
  );


  buf
  g8
  (
    n124,
    n28
  );


  buf
  g9
  (
    n34,
    n17
  );


  not
  g10
  (
    n110,
    n22
  );


  buf
  g11
  (
    n151,
    n22
  );


  not
  g12
  (
    n119,
    n23
  );


  not
  g13
  (
    n57,
    n15
  );


  not
  g14
  (
    n134,
    n24
  );


  not
  g15
  (
    n59,
    n30
  );


  not
  g16
  (
    n138,
    n29
  );


  buf
  g17
  (
    n39,
    n20
  );


  not
  g18
  (
    n106,
    n12
  );


  buf
  g19
  (
    n56,
    n10
  );


  not
  g20
  (
    n81,
    n4
  );


  not
  g21
  (
    n108,
    n11
  );


  buf
  g22
  (
    n50,
    n29
  );


  buf
  g23
  (
    n36,
    n20
  );


  not
  g24
  (
    n60,
    n1
  );


  buf
  g25
  (
    n114,
    n23
  );


  buf
  g26
  (
    n121,
    n22
  );


  buf
  g27
  (
    n97,
    n12
  );


  buf
  g28
  (
    KeyWire_0_38,
    n6
  );


  not
  g29
  (
    n104,
    n24
  );


  not
  g30
  (
    n84,
    n29
  );


  not
  g31
  (
    n37,
    n30
  );


  not
  g32
  (
    n111,
    n20
  );


  buf
  g33
  (
    n147,
    n2
  );


  not
  g34
  (
    n69,
    n31
  );


  buf
  g35
  (
    n91,
    n7
  );


  not
  g36
  (
    n89,
    n9
  );


  buf
  g37
  (
    n54,
    n27
  );


  not
  g38
  (
    n82,
    n14
  );


  buf
  g39
  (
    n83,
    n26
  );


  buf
  g40
  (
    n127,
    n31
  );


  not
  g41
  (
    n80,
    n28
  );


  not
  g42
  (
    n51,
    n25
  );


  not
  g43
  (
    n139,
    n4
  );


  not
  g44
  (
    n87,
    n15
  );


  buf
  g45
  (
    n46,
    n9
  );


  not
  g46
  (
    n115,
    n3
  );


  buf
  g47
  (
    n41,
    n29
  );


  buf
  g48
  (
    n92,
    n10
  );


  buf
  g49
  (
    n49,
    n17
  );


  not
  g50
  (
    n112,
    n10
  );


  buf
  g51
  (
    n90,
    n3
  );


  not
  g52
  (
    n152,
    n1
  );


  not
  g53
  (
    n130,
    n18
  );


  not
  g54
  (
    n132,
    n11
  );


  buf
  g55
  (
    n44,
    n16
  );


  buf
  g56
  (
    n113,
    n19
  );


  not
  g57
  (
    n93,
    n2
  );


  not
  g58
  (
    n77,
    n15
  );


  buf
  g59
  (
    n71,
    n3
  );


  buf
  g60
  (
    n102,
    n31
  );


  buf
  g61
  (
    n86,
    n24
  );


  buf
  g62
  (
    n88,
    n16
  );


  buf
  g63
  (
    n73,
    n13
  );


  not
  g64
  (
    KeyWire_0_44,
    n1
  );


  not
  g65
  (
    n103,
    n14
  );


  not
  g66
  (
    n148,
    n18
  );


  buf
  g67
  (
    n85,
    n4
  );


  not
  g68
  (
    n101,
    n2
  );


  not
  g69
  (
    n143,
    n19
  );


  not
  g70
  (
    n53,
    n28
  );


  not
  g71
  (
    n72,
    n12
  );


  buf
  g72
  (
    n78,
    n6
  );


  buf
  g73
  (
    n55,
    n18
  );


  buf
  g74
  (
    n136,
    n5
  );


  not
  g75
  (
    n61,
    n23
  );


  buf
  g76
  (
    n98,
    n16
  );


  not
  g77
  (
    n141,
    n26
  );


  buf
  g78
  (
    n76,
    n5
  );


  buf
  g79
  (
    n58,
    n21
  );


  not
  g80
  (
    n62,
    n21
  );


  not
  g81
  (
    n65,
    n28
  );


  buf
  g82
  (
    n43,
    n7
  );


  not
  g83
  (
    n47,
    n17
  );


  not
  g84
  (
    n75,
    n6
  );


  buf
  g85
  (
    n107,
    n17
  );


  buf
  g86
  (
    n116,
    n13
  );


  not
  g87
  (
    n68,
    n16
  );


  not
  g88
  (
    n117,
    n2
  );


  buf
  g89
  (
    n145,
    n23
  );


  not
  g90
  (
    n33,
    n8
  );


  buf
  g91
  (
    n42,
    n5
  );


  buf
  g92
  (
    n109,
    n8
  );


  not
  g93
  (
    n153,
    n27
  );


  not
  g94
  (
    n64,
    n21
  );


  buf
  g95
  (
    n128,
    n10
  );


  not
  g96
  (
    n156,
    n27
  );


  buf
  g97
  (
    n67,
    n3
  );


  not
  g98
  (
    n66,
    n26
  );


  buf
  g99
  (
    n96,
    n25
  );


  not
  g100
  (
    n140,
    n31
  );


  not
  g101
  (
    n48,
    n25
  );


  not
  g102
  (
    n100,
    n14
  );


  buf
  g103
  (
    n118,
    n7
  );


  buf
  g104
  (
    n146,
    n19
  );


  not
  g105
  (
    n149,
    n27
  );


  buf
  g106
  (
    n150,
    n8
  );


  buf
  g107
  (
    n40,
    n11
  );


  buf
  g108
  (
    n129,
    n13
  );


  not
  g109
  (
    n38,
    n7
  );


  buf
  g110
  (
    n52,
    n25
  );


  not
  g111
  (
    n45,
    n1
  );


  not
  g112
  (
    n79,
    n6
  );


  not
  g113
  (
    n135,
    n19
  );


  not
  g114
  (
    n126,
    n26
  );


  buf
  g115
  (
    n123,
    n8
  );


  buf
  g116
  (
    n125,
    n4
  );


  not
  g117
  (
    n120,
    n21
  );


  buf
  g118
  (
    n74,
    n30
  );


  not
  g119
  (
    n105,
    n12
  );


  buf
  g120
  (
    n131,
    n22
  );


  not
  g121
  (
    n95,
    n13
  );


  not
  g122
  (
    n99,
    n5
  );


  buf
  g123
  (
    n137,
    n24
  );


  buf
  g124
  (
    n640,
    n71
  );


  buf
  g125
  (
    n223,
    n129
  );


  not
  g126
  (
    n305,
    n81
  );


  buf
  g127
  (
    n596,
    n149
  );


  not
  g128
  (
    n525,
    n105
  );


  buf
  g129
  (
    n479,
    n87
  );


  buf
  g130
  (
    n336,
    n119
  );


  not
  g131
  (
    n369,
    n96
  );


  buf
  g132
  (
    n171,
    n106
  );


  not
  g133
  (
    n163,
    n108
  );


  not
  g134
  (
    n310,
    n140
  );


  buf
  g135
  (
    n457,
    n140
  );


  not
  g136
  (
    n288,
    n99
  );


  not
  g137
  (
    n512,
    n98
  );


  buf
  g138
  (
    n562,
    n105
  );


  buf
  g139
  (
    n227,
    n119
  );


  not
  g140
  (
    n367,
    n36
  );


  buf
  g141
  (
    n545,
    n100
  );


  not
  g142
  (
    n231,
    n61
  );


  not
  g143
  (
    n488,
    n102
  );


  not
  g144
  (
    n345,
    n33
  );


  not
  g145
  (
    KeyWire_0_59,
    n83
  );


  not
  g146
  (
    n556,
    n71
  );


  not
  g147
  (
    n222,
    n80
  );


  buf
  g148
  (
    n263,
    n107
  );


  buf
  g149
  (
    n361,
    n56
  );


  buf
  g150
  (
    n358,
    n97
  );


  not
  g151
  (
    n191,
    n50
  );


  not
  g152
  (
    KeyWire_0_50,
    n79
  );


  not
  g153
  (
    n602,
    n64
  );


  buf
  g154
  (
    n604,
    n39
  );


  not
  g155
  (
    n206,
    n133
  );


  not
  g156
  (
    n301,
    n114
  );


  not
  g157
  (
    n220,
    n123
  );


  buf
  g158
  (
    n161,
    n147
  );


  not
  g159
  (
    n481,
    n108
  );


  buf
  g160
  (
    n578,
    n156
  );


  not
  g161
  (
    n572,
    n127
  );


  not
  g162
  (
    n535,
    n123
  );


  buf
  g163
  (
    n576,
    n142
  );


  not
  g164
  (
    n605,
    n69
  );


  not
  g165
  (
    n224,
    n77
  );


  buf
  g166
  (
    n182,
    n42
  );


  buf
  g167
  (
    n388,
    n92
  );


  buf
  g168
  (
    n416,
    n78
  );


  buf
  g169
  (
    n197,
    n94
  );


  not
  g170
  (
    n281,
    n134
  );


  not
  g171
  (
    n341,
    n132
  );


  not
  g172
  (
    n534,
    n57
  );


  buf
  g173
  (
    n202,
    n60
  );


  not
  g174
  (
    n378,
    n130
  );


  not
  g175
  (
    n234,
    n146
  );


  buf
  g176
  (
    n337,
    n117
  );


  not
  g177
  (
    n519,
    n90
  );


  not
  g178
  (
    n436,
    n60
  );


  buf
  g179
  (
    n507,
    n55
  );


  buf
  g180
  (
    n346,
    n81
  );


  buf
  g181
  (
    n204,
    n41
  );


  buf
  g182
  (
    n394,
    n60
  );


  not
  g183
  (
    n564,
    n124
  );


  not
  g184
  (
    n577,
    n99
  );


  buf
  g185
  (
    n628,
    n112
  );


  buf
  g186
  (
    n492,
    n110
  );


  not
  g187
  (
    n625,
    n84
  );


  not
  g188
  (
    n256,
    n137
  );


  buf
  g189
  (
    n482,
    n47
  );


  buf
  g190
  (
    n428,
    n67
  );


  not
  g191
  (
    n522,
    n149
  );


  not
  g192
  (
    n230,
    n38
  );


  not
  g193
  (
    n370,
    n114
  );


  buf
  g194
  (
    n648,
    n67
  );


  buf
  g195
  (
    n542,
    n54
  );


  buf
  g196
  (
    n299,
    n47
  );


  buf
  g197
  (
    n166,
    n115
  );


  buf
  g198
  (
    n441,
    n150
  );


  not
  g199
  (
    n473,
    n143
  );


  not
  g200
  (
    n489,
    n101
  );


  not
  g201
  (
    n459,
    n54
  );


  not
  g202
  (
    n257,
    n57
  );


  buf
  g203
  (
    n591,
    n107
  );


  not
  g204
  (
    n386,
    n51
  );


  buf
  g205
  (
    n157,
    n139
  );


  buf
  g206
  (
    n258,
    n57
  );


  not
  g207
  (
    n503,
    n35
  );


  buf
  g208
  (
    n181,
    n34
  );


  not
  g209
  (
    n550,
    n73
  );


  buf
  g210
  (
    n321,
    n138
  );


  not
  g211
  (
    n405,
    n80
  );


  buf
  g212
  (
    n438,
    n98
  );


  buf
  g213
  (
    n480,
    n143
  );


  not
  g214
  (
    n573,
    n34
  );


  not
  g215
  (
    n179,
    n141
  );


  not
  g216
  (
    n290,
    n55
  );


  buf
  g217
  (
    n174,
    n84
  );


  not
  g218
  (
    n592,
    n117
  );


  not
  g219
  (
    n353,
    n45
  );


  buf
  g220
  (
    n209,
    n44
  );


  not
  g221
  (
    n500,
    n46
  );


  buf
  g222
  (
    n348,
    n129
  );


  buf
  g223
  (
    n213,
    n155
  );


  buf
  g224
  (
    KeyWire_0_12,
    n143
  );


  not
  g225
  (
    n328,
    n72
  );


  buf
  g226
  (
    n484,
    n106
  );


  buf
  g227
  (
    n627,
    n79
  );


  not
  g228
  (
    n216,
    n145
  );


  not
  g229
  (
    n568,
    n151
  );


  not
  g230
  (
    n274,
    n127
  );


  buf
  g231
  (
    n343,
    n128
  );


  buf
  g232
  (
    n476,
    n137
  );


  buf
  g233
  (
    n311,
    n69
  );


  buf
  g234
  (
    n569,
    n127
  );


  buf
  g235
  (
    n291,
    n66
  );


  buf
  g236
  (
    n236,
    n90
  );


  not
  g237
  (
    n597,
    n111
  );


  buf
  g238
  (
    n331,
    n116
  );


  buf
  g239
  (
    n237,
    n135
  );


  not
  g240
  (
    n632,
    n53
  );


  buf
  g241
  (
    n347,
    n125
  );


  not
  g242
  (
    n211,
    n104
  );


  buf
  g243
  (
    n193,
    n66
  );


  not
  g244
  (
    n233,
    n135
  );


  not
  g245
  (
    n268,
    n132
  );


  buf
  g246
  (
    n318,
    n79
  );


  buf
  g247
  (
    n235,
    n43
  );


  buf
  g248
  (
    n371,
    n126
  );


  buf
  g249
  (
    n567,
    n93
  );


  not
  g250
  (
    n523,
    n58
  );


  buf
  g251
  (
    n521,
    n38
  );


  buf
  g252
  (
    n471,
    n129
  );


  buf
  g253
  (
    n313,
    n56
  );


  buf
  g254
  (
    n403,
    n126
  );


  not
  g255
  (
    n273,
    n128
  );


  buf
  g256
  (
    n502,
    n132
  );


  not
  g257
  (
    n376,
    n90
  );


  buf
  g258
  (
    n444,
    n67
  );


  not
  g259
  (
    n340,
    n42
  );


  not
  g260
  (
    n516,
    n65
  );


  not
  g261
  (
    n434,
    n83
  );


  buf
  g262
  (
    n410,
    n49
  );


  buf
  g263
  (
    n297,
    n152
  );


  not
  g264
  (
    n165,
    n51
  );


  buf
  g265
  (
    n284,
    n110
  );


  buf
  g266
  (
    n243,
    n124
  );


  buf
  g267
  (
    n543,
    n76
  );


  not
  g268
  (
    n399,
    n73
  );


  not
  g269
  (
    n508,
    n59
  );


  not
  g270
  (
    n391,
    n78
  );


  not
  g271
  (
    n309,
    n43
  );


  not
  g272
  (
    n635,
    n41
  );


  buf
  g273
  (
    n228,
    n36
  );


  not
  g274
  (
    n537,
    n79
  );


  not
  g275
  (
    n552,
    n53
  );


  not
  g276
  (
    n246,
    n86
  );


  buf
  g277
  (
    n218,
    n49
  );


  buf
  g278
  (
    n404,
    n58
  );


  not
  g279
  (
    n463,
    n118
  );


  not
  g280
  (
    n430,
    n112
  );


  buf
  g281
  (
    n285,
    n89
  );


  buf
  g282
  (
    n558,
    n43
  );


  buf
  g283
  (
    n506,
    n108
  );


  not
  g284
  (
    n464,
    n82
  );


  not
  g285
  (
    n520,
    n124
  );


  not
  g286
  (
    KeyWire_0_37,
    n39
  );


  not
  g287
  (
    n402,
    n62
  );


  buf
  g288
  (
    n618,
    n152
  );


  not
  g289
  (
    KeyWire_0_10,
    n136
  );


  buf
  g290
  (
    n292,
    n84
  );


  buf
  g291
  (
    n614,
    n96
  );


  not
  g292
  (
    n250,
    n104
  );


  not
  g293
  (
    n160,
    n140
  );


  buf
  g294
  (
    n574,
    n75
  );


  not
  g295
  (
    n259,
    n63
  );


  not
  g296
  (
    n276,
    n155
  );


  buf
  g297
  (
    n398,
    n147
  );


  buf
  g298
  (
    n547,
    n150
  );


  buf
  g299
  (
    n372,
    n51
  );


  not
  g300
  (
    n643,
    n154
  );


  not
  g301
  (
    n335,
    n134
  );


  not
  g302
  (
    n362,
    n71
  );


  buf
  g303
  (
    n354,
    n92
  );


  buf
  g304
  (
    n619,
    n88
  );


  buf
  g305
  (
    n269,
    n36
  );


  not
  g306
  (
    n296,
    n97
  );


  not
  g307
  (
    n580,
    n141
  );


  not
  g308
  (
    n497,
    n54
  );


  buf
  g309
  (
    n407,
    n155
  );


  buf
  g310
  (
    n515,
    n155
  );


  buf
  g311
  (
    n585,
    n72
  );


  not
  g312
  (
    n278,
    n82
  );


  buf
  g313
  (
    n423,
    n40
  );


  not
  g314
  (
    n208,
    n138
  );


  not
  g315
  (
    n418,
    n113
  );


  buf
  g316
  (
    n338,
    n89
  );


  not
  g317
  (
    n283,
    n33
  );


  buf
  g318
  (
    n559,
    n134
  );


  buf
  g319
  (
    n425,
    n77
  );


  buf
  g320
  (
    n232,
    n65
  );


  buf
  g321
  (
    n350,
    n56
  );


  buf
  g322
  (
    n650,
    n143
  );


  not
  g323
  (
    n442,
    n59
  );


  not
  g324
  (
    n526,
    n145
  );


  buf
  g325
  (
    n451,
    n136
  );


  not
  g326
  (
    n406,
    n115
  );


  not
  g327
  (
    n613,
    n85
  );


  buf
  g328
  (
    n355,
    n154
  );


  not
  g329
  (
    n393,
    n141
  );


  not
  g330
  (
    n374,
    n48
  );


  not
  g331
  (
    n189,
    n37
  );


  not
  g332
  (
    n432,
    n102
  );


  not
  g333
  (
    n470,
    n140
  );


  buf
  g334
  (
    n517,
    n141
  );


  not
  g335
  (
    n531,
    n151
  );


  not
  g336
  (
    n172,
    n51
  );


  not
  g337
  (
    n334,
    n84
  );


  not
  g338
  (
    n450,
    n82
  );


  not
  g339
  (
    n254,
    n47
  );


  buf
  g340
  (
    n575,
    n152
  );


  buf
  g341
  (
    n454,
    n78
  );


  not
  g342
  (
    n286,
    n116
  );


  buf
  g343
  (
    n443,
    n48
  );


  buf
  g344
  (
    n487,
    n108
  );


  buf
  g345
  (
    n563,
    n139
  );


  buf
  g346
  (
    n298,
    n64
  );


  not
  g347
  (
    KeyWire_0_16,
    n133
  );


  buf
  g348
  (
    n456,
    n150
  );


  buf
  g349
  (
    n581,
    n153
  );


  buf
  g350
  (
    n504,
    n53
  );


  not
  g351
  (
    n307,
    n148
  );


  buf
  g352
  (
    n415,
    n65
  );


  buf
  g353
  (
    n453,
    n85
  );


  not
  g354
  (
    KeyWire_0_43,
    n59
  );


  not
  g355
  (
    n357,
    n52
  );


  buf
  g356
  (
    n249,
    n90
  );


  buf
  g357
  (
    n413,
    n102
  );


  buf
  g358
  (
    n411,
    n95
  );


  buf
  g359
  (
    n215,
    n35
  );


  not
  g360
  (
    n637,
    n91
  );


  not
  g361
  (
    n458,
    n126
  );


  not
  g362
  (
    n158,
    n83
  );


  buf
  g363
  (
    n401,
    n98
  );


  not
  g364
  (
    n176,
    n91
  );


  buf
  g365
  (
    n483,
    n97
  );


  not
  g366
  (
    n644,
    n75
  );


  not
  g367
  (
    n198,
    n69
  );


  buf
  g368
  (
    n366,
    n76
  );


  buf
  g369
  (
    n217,
    n118
  );


  buf
  g370
  (
    n207,
    n85
  );


  buf
  g371
  (
    n266,
    n106
  );


  not
  g372
  (
    n275,
    n105
  );


  buf
  g373
  (
    n544,
    n68
  );


  not
  g374
  (
    n162,
    n156
  );


  not
  g375
  (
    n630,
    n40
  );


  not
  g376
  (
    n461,
    n133
  );


  not
  g377
  (
    n595,
    n39
  );


  not
  g378
  (
    n384,
    n87
  );


  buf
  g379
  (
    KeyWire_0_22,
    n39
  );


  not
  g380
  (
    n303,
    n144
  );


  not
  g381
  (
    n599,
    n128
  );


  not
  g382
  (
    n528,
    n61
  );


  not
  g383
  (
    n280,
    n142
  );


  not
  g384
  (
    n294,
    n151
  );


  buf
  g385
  (
    n478,
    n148
  );


  not
  g386
  (
    n560,
    n92
  );


  buf
  g387
  (
    n490,
    n35
  );


  not
  g388
  (
    n185,
    n34
  );


  not
  g389
  (
    n261,
    n117
  );


  not
  g390
  (
    n201,
    n151
  );


  not
  g391
  (
    n186,
    n115
  );


  not
  g392
  (
    n620,
    n96
  );


  not
  g393
  (
    n200,
    n116
  );


  buf
  g394
  (
    n364,
    n99
  );


  not
  g395
  (
    n329,
    n114
  );


  buf
  g396
  (
    n600,
    n60
  );


  buf
  g397
  (
    n633,
    n106
  );


  buf
  g398
  (
    n389,
    n99
  );


  buf
  g399
  (
    n326,
    n46
  );


  buf
  g400
  (
    n494,
    n119
  );


  not
  g401
  (
    n649,
    n94
  );


  not
  g402
  (
    n387,
    n38
  );


  buf
  g403
  (
    n647,
    n74
  );


  not
  g404
  (
    n565,
    n44
  );


  not
  g405
  (
    n616,
    n76
  );


  not
  g406
  (
    n606,
    n123
  );


  not
  g407
  (
    n212,
    n98
  );


  not
  g408
  (
    n629,
    n156
  );


  buf
  g409
  (
    n652,
    n116
  );


  buf
  g410
  (
    n247,
    n58
  );


  buf
  g411
  (
    n421,
    n150
  );


  buf
  g412
  (
    n486,
    n87
  );


  not
  g413
  (
    n638,
    n101
  );


  not
  g414
  (
    n412,
    n68
  );


  not
  g415
  (
    n199,
    n136
  );


  buf
  g416
  (
    n373,
    n104
  );


  not
  g417
  (
    n607,
    n118
  );


  buf
  g418
  (
    n510,
    n110
  );


  not
  g419
  (
    n539,
    n75
  );


  buf
  g420
  (
    n586,
    n146
  );


  buf
  g421
  (
    n159,
    n52
  );


  buf
  g422
  (
    n302,
    n46
  );


  not
  g423
  (
    n608,
    n129
  );


  not
  g424
  (
    n617,
    n50
  );


  buf
  g425
  (
    n594,
    n52
  );


  buf
  g426
  (
    n365,
    n68
  );


  buf
  g427
  (
    n472,
    n131
  );


  buf
  g428
  (
    n553,
    n40
  );


  buf
  g429
  (
    n448,
    n115
  );


  not
  g430
  (
    n324,
    n121
  );


  not
  g431
  (
    n501,
    n147
  );


  not
  g432
  (
    n175,
    n120
  );


  not
  g433
  (
    n610,
    n109
  );


  not
  g434
  (
    KeyWire_0_33,
    n88
  );


  buf
  g435
  (
    n327,
    n109
  );


  buf
  g436
  (
    n642,
    n88
  );


  not
  g437
  (
    n433,
    n125
  );


  buf
  g438
  (
    n351,
    n53
  );


  buf
  g439
  (
    n474,
    n144
  );


  buf
  g440
  (
    n180,
    n154
  );


  not
  g441
  (
    n452,
    n153
  );


  buf
  g442
  (
    n546,
    n94
  );


  not
  g443
  (
    n332,
    n135
  );


  buf
  g444
  (
    n214,
    n43
  );


  buf
  g445
  (
    n533,
    n131
  );


  not
  g446
  (
    n241,
    n48
  );


  not
  g447
  (
    n455,
    n118
  );


  not
  g448
  (
    n509,
    n111
  );


  buf
  g449
  (
    n349,
    n142
  );


  not
  g450
  (
    n493,
    n100
  );


  buf
  g451
  (
    n203,
    n135
  );


  not
  g452
  (
    n239,
    n130
  );


  buf
  g453
  (
    n380,
    n103
  );


  buf
  g454
  (
    n287,
    n65
  );


  not
  g455
  (
    n513,
    n86
  );


  not
  g456
  (
    n462,
    n87
  );


  buf
  g457
  (
    n333,
    n139
  );


  not
  g458
  (
    n582,
    n105
  );


  not
  g459
  (
    n272,
    n59
  );


  not
  g460
  (
    n221,
    n50
  );


  not
  g461
  (
    n551,
    n121
  );


  not
  g462
  (
    n561,
    n64
  );


  buf
  g463
  (
    n314,
    n113
  );


  not
  g464
  (
    n339,
    n63
  );


  not
  g465
  (
    n168,
    n83
  );


  not
  g466
  (
    n417,
    n95
  );


  not
  g467
  (
    n251,
    n131
  );


  not
  g468
  (
    n437,
    n42
  );


  buf
  g469
  (
    n192,
    n124
  );


  not
  g470
  (
    n465,
    n40
  );


  buf
  g471
  (
    n636,
    n55
  );


  buf
  g472
  (
    n210,
    n117
  );


  buf
  g473
  (
    n375,
    n64
  );


  not
  g474
  (
    n252,
    n107
  );


  buf
  g475
  (
    n477,
    n62
  );


  buf
  g476
  (
    n529,
    n131
  );


  buf
  g477
  (
    n612,
    n49
  );


  buf
  g478
  (
    n511,
    n67
  );


  not
  g479
  (
    n323,
    n95
  );


  buf
  g480
  (
    n316,
    n120
  );


  buf
  g481
  (
    n170,
    n152
  );


  buf
  g482
  (
    n187,
    n114
  );


  buf
  g483
  (
    n205,
    n109
  );


  not
  g484
  (
    n588,
    n86
  );


  buf
  g485
  (
    n279,
    n47
  );


  buf
  g486
  (
    n267,
    n70
  );


  buf
  g487
  (
    n485,
    n49
  );


  not
  g488
  (
    n496,
    n91
  );


  buf
  g489
  (
    n390,
    n125
  );


  buf
  g490
  (
    n536,
    n89
  );


  buf
  g491
  (
    n611,
    n100
  );


  buf
  g492
  (
    n194,
    n41
  );


  not
  g493
  (
    n368,
    n92
  );


  buf
  g494
  (
    n395,
    n52
  );


  not
  g495
  (
    n540,
    n134
  );


  not
  g496
  (
    n589,
    n58
  );


  buf
  g497
  (
    n491,
    n132
  );


  buf
  g498
  (
    n396,
    n70
  );


  buf
  g499
  (
    n169,
    n71
  );


  buf
  g500
  (
    n300,
    n56
  );


  not
  g501
  (
    n422,
    n109
  );


  buf
  g502
  (
    n248,
    n103
  );


  not
  g503
  (
    n460,
    n93
  );


  buf
  g504
  (
    n570,
    n62
  );


  not
  g505
  (
    n587,
    n113
  );


  buf
  g506
  (
    n527,
    n119
  );


  buf
  g507
  (
    n557,
    n103
  );


  buf
  g508
  (
    n356,
    n95
  );


  buf
  g509
  (
    n173,
    n80
  );


  not
  g510
  (
    n532,
    n142
  );


  not
  g511
  (
    n593,
    n153
  );


  not
  g512
  (
    n518,
    n37
  );


  not
  g513
  (
    n571,
    n145
  );


  not
  g514
  (
    n242,
    n81
  );


  buf
  g515
  (
    n315,
    n82
  );


  not
  g516
  (
    n359,
    n68
  );


  not
  g517
  (
    n549,
    n122
  );


  not
  g518
  (
    n164,
    n101
  );


  buf
  g519
  (
    n344,
    n112
  );


  buf
  g520
  (
    n603,
    n120
  );


  buf
  g521
  (
    n495,
    n73
  );


  not
  g522
  (
    n646,
    n149
  );


  not
  g523
  (
    n264,
    n148
  );


  buf
  g524
  (
    n289,
    n33
  );


  not
  g525
  (
    n190,
    n138
  );


  not
  g526
  (
    n631,
    n96
  );


  not
  g527
  (
    KeyWire_0_26,
    n81
  );


  buf
  g528
  (
    n260,
    n85
  );


  buf
  g529
  (
    n499,
    n122
  );


  buf
  g530
  (
    n626,
    n42
  );


  buf
  g531
  (
    n566,
    n110
  );


  not
  g532
  (
    n167,
    n74
  );


  not
  g533
  (
    n439,
    n111
  );


  not
  g534
  (
    n360,
    n156
  );


  buf
  g535
  (
    n178,
    n104
  );


  buf
  g536
  (
    n400,
    n88
  );


  buf
  g537
  (
    n426,
    n126
  );


  not
  g538
  (
    n196,
    n57
  );


  buf
  g539
  (
    n306,
    n107
  );


  buf
  g540
  (
    n270,
    n44
  );


  buf
  g541
  (
    n377,
    n44
  );


  not
  g542
  (
    n579,
    n34
  );


  buf
  g543
  (
    n308,
    n76
  );


  not
  g544
  (
    n609,
    n45
  );


  not
  g545
  (
    n317,
    n80
  );


  not
  g546
  (
    n583,
    n128
  );


  buf
  g547
  (
    n295,
    n46
  );


  buf
  g548
  (
    n469,
    n93
  );


  buf
  g549
  (
    n381,
    n146
  );


  buf
  g550
  (
    n431,
    n148
  );


  buf
  g551
  (
    n467,
    n89
  );


  not
  g552
  (
    n446,
    n111
  );


  not
  g553
  (
    n293,
    n145
  );


  buf
  g554
  (
    n195,
    n149
  );


  not
  g555
  (
    n621,
    n136
  );


  buf
  g556
  (
    n184,
    n33
  );


  not
  g557
  (
    n320,
    n70
  );


  buf
  g558
  (
    n304,
    n36
  );


  buf
  g559
  (
    n225,
    n93
  );


  buf
  g560
  (
    KeyWire_0_5,
    n146
  );


  buf
  g561
  (
    n409,
    n41
  );


  not
  g562
  (
    n188,
    n144
  );


  buf
  g563
  (
    n379,
    n153
  );


  buf
  g564
  (
    n639,
    n103
  );


  not
  g565
  (
    n466,
    n125
  );


  buf
  g566
  (
    n598,
    n154
  );


  buf
  g567
  (
    n330,
    n69
  );


  not
  g568
  (
    n590,
    n86
  );


  not
  g569
  (
    n414,
    n147
  );


  not
  g570
  (
    n271,
    n37
  );


  not
  g571
  (
    n641,
    n127
  );


  not
  g572
  (
    n282,
    n137
  );


  not
  g573
  (
    n245,
    n123
  );


  buf
  g574
  (
    n623,
    n97
  );


  buf
  g575
  (
    n435,
    n61
  );


  buf
  g576
  (
    n277,
    n66
  );


  not
  g577
  (
    n312,
    n77
  );


  buf
  g578
  (
    n601,
    n113
  );


  buf
  g579
  (
    n385,
    n45
  );


  buf
  g580
  (
    n427,
    n122
  );


  not
  g581
  (
    n424,
    n48
  );


  buf
  g582
  (
    n524,
    n121
  );


  not
  g583
  (
    n548,
    n63
  );


  buf
  g584
  (
    n622,
    n70
  );


  not
  g585
  (
    n408,
    n37
  );


  not
  g586
  (
    n319,
    n144
  );


  not
  g587
  (
    n651,
    n138
  );


  not
  g588
  (
    n624,
    n121
  );


  not
  g589
  (
    n352,
    n130
  );


  not
  g590
  (
    n475,
    n72
  );


  buf
  g591
  (
    n555,
    n100
  );


  not
  g592
  (
    n183,
    n38
  );


  not
  g593
  (
    n342,
    n130
  );


  not
  g594
  (
    n538,
    n91
  );


  not
  g595
  (
    n253,
    n61
  );


  not
  g596
  (
    n392,
    n35
  );


  buf
  g597
  (
    n530,
    n122
  );


  not
  g598
  (
    n440,
    n72
  );


  not
  g599
  (
    n177,
    n62
  );


  not
  g600
  (
    n449,
    n94
  );


  buf
  g601
  (
    n468,
    n133
  );


  not
  g602
  (
    n219,
    n55
  );


  buf
  g603
  (
    KeyWire_0_57,
    n73
  );


  not
  g604
  (
    n262,
    n112
  );


  buf
  g605
  (
    n382,
    n77
  );


  not
  g606
  (
    n226,
    n102
  );


  buf
  g607
  (
    n265,
    n54
  );


  not
  g608
  (
    n420,
    n50
  );


  not
  g609
  (
    n419,
    n78
  );


  buf
  g610
  (
    n229,
    n120
  );


  not
  g611
  (
    n244,
    n74
  );


  not
  g612
  (
    n615,
    n75
  );


  not
  g613
  (
    n363,
    n63
  );


  not
  g614
  (
    n584,
    n74
  );


  not
  g615
  (
    n383,
    n66
  );


  not
  g616
  (
    n505,
    n137
  );


  not
  g617
  (
    n240,
    n139
  );


  not
  g618
  (
    n238,
    n101
  );


  not
  g619
  (
    n645,
    n45
  );


  buf
  g620
  (
    n1531,
    n538
  );


  buf
  g621
  (
    n668,
    n233
  );


  buf
  g622
  (
    n1573,
    n624
  );


  not
  g623
  (
    n1592,
    n585
  );


  not
  g624
  (
    n1275,
    n269
  );


  buf
  g625
  (
    n1433,
    n286
  );


  buf
  g626
  (
    n1316,
    n372
  );


  not
  g627
  (
    n855,
    n449
  );


  not
  g628
  (
    n689,
    n264
  );


  buf
  g629
  (
    n1831,
    n435
  );


  not
  g630
  (
    n1412,
    n456
  );


  not
  g631
  (
    n746,
    n472
  );


  buf
  g632
  (
    n873,
    n400
  );


  buf
  g633
  (
    n1963,
    n307
  );


  not
  g634
  (
    n1005,
    n566
  );


  not
  g635
  (
    n1417,
    n227
  );


  not
  g636
  (
    n1273,
    n195
  );


  not
  g637
  (
    n1857,
    n323
  );


  buf
  g638
  (
    n1754,
    n380
  );


  buf
  g639
  (
    n876,
    n531
  );


  buf
  g640
  (
    n827,
    n615
  );


  buf
  g641
  (
    n676,
    n259
  );


  buf
  g642
  (
    n850,
    n394
  );


  not
  g643
  (
    n779,
    n570
  );


  not
  g644
  (
    n1509,
    n510
  );


  buf
  g645
  (
    n875,
    n264
  );


  not
  g646
  (
    n1711,
    n559
  );


  buf
  g647
  (
    n1109,
    n280
  );


  buf
  g648
  (
    n1045,
    n397
  );


  buf
  g649
  (
    n796,
    n316
  );


  not
  g650
  (
    n1585,
    n430
  );


  buf
  g651
  (
    n1123,
    n512
  );


  buf
  g652
  (
    n1448,
    n606
  );


  buf
  g653
  (
    n1097,
    n463
  );


  not
  g654
  (
    n727,
    n212
  );


  not
  g655
  (
    n1251,
    n386
  );


  not
  g656
  (
    n1313,
    n311
  );


  not
  g657
  (
    n898,
    n572
  );


  not
  g658
  (
    n1879,
    n347
  );


  not
  g659
  (
    n707,
    n381
  );


  buf
  g660
  (
    n818,
    n603
  );


  not
  g661
  (
    n1118,
    n359
  );


  buf
  g662
  (
    n1905,
    n566
  );


  buf
  g663
  (
    n1209,
    n463
  );


  buf
  g664
  (
    n891,
    n379
  );


  not
  g665
  (
    n1873,
    n494
  );


  buf
  g666
  (
    n1868,
    n528
  );


  not
  g667
  (
    n1904,
    n450
  );


  not
  g668
  (
    n1314,
    n378
  );


  not
  g669
  (
    n1012,
    n253
  );


  buf
  g670
  (
    n1895,
    n479
  );


  buf
  g671
  (
    n1815,
    n270
  );


  buf
  g672
  (
    n1874,
    n636
  );


  not
  g673
  (
    n1625,
    n237
  );


  not
  g674
  (
    n1063,
    n438
  );


  buf
  g675
  (
    n1556,
    n568
  );


  buf
  g676
  (
    n1756,
    n218
  );


  buf
  g677
  (
    n1116,
    n647
  );


  not
  g678
  (
    n1792,
    n508
  );


  not
  g679
  (
    n1630,
    n286
  );


  not
  g680
  (
    n1534,
    n470
  );


  not
  g681
  (
    n1497,
    n455
  );


  not
  g682
  (
    n1568,
    n310
  );


  buf
  g683
  (
    n993,
    n294
  );


  buf
  g684
  (
    n721,
    n218
  );


  buf
  g685
  (
    n1174,
    n602
  );


  not
  g686
  (
    n1155,
    n634
  );


  not
  g687
  (
    n1974,
    n403
  );


  buf
  g688
  (
    n1449,
    n329
  );


  buf
  g689
  (
    n777,
    n478
  );


  not
  g690
  (
    n998,
    n631
  );


  not
  g691
  (
    n1686,
    n310
  );


  buf
  g692
  (
    n1936,
    n434
  );


  not
  g693
  (
    n1616,
    n477
  );


  not
  g694
  (
    n1732,
    n628
  );


  buf
  g695
  (
    n969,
    n389
  );


  buf
  g696
  (
    n785,
    n417
  );


  buf
  g697
  (
    n1926,
    n388
  );


  buf
  g698
  (
    n683,
    n515
  );


  not
  g699
  (
    n990,
    n310
  );


  buf
  g700
  (
    n1192,
    n219
  );


  not
  g701
  (
    n1318,
    n207
  );


  not
  g702
  (
    n1539,
    n571
  );


  not
  g703
  (
    n1357,
    n160
  );


  not
  g704
  (
    n1542,
    n409
  );


  buf
  g705
  (
    n985,
    n502
  );


  buf
  g706
  (
    n695,
    n479
  );


  not
  g707
  (
    n1289,
    n402
  );


  not
  g708
  (
    n1132,
    n377
  );


  buf
  g709
  (
    n1721,
    n283
  );


  buf
  g710
  (
    n1399,
    n423
  );


  buf
  g711
  (
    n1191,
    n323
  );


  not
  g712
  (
    n1722,
    n634
  );


  buf
  g713
  (
    n817,
    n213
  );


  buf
  g714
  (
    n1353,
    n359
  );


  buf
  g715
  (
    n948,
    n369
  );


  not
  g716
  (
    n1135,
    n619
  );


  not
  g717
  (
    n1774,
    n343
  );


  not
  g718
  (
    n776,
    n171
  );


  buf
  g719
  (
    n1025,
    n274
  );


  not
  g720
  (
    n1390,
    n627
  );


  not
  g721
  (
    n1207,
    n524
  );


  buf
  g722
  (
    KeyWire_0_25,
    n642
  );


  buf
  g723
  (
    n1644,
    n496
  );


  not
  g724
  (
    n1973,
    n252
  );


  buf
  g725
  (
    n1327,
    n250
  );


  buf
  g726
  (
    n1744,
    n528
  );


  not
  g727
  (
    n1156,
    n374
  );


  buf
  g728
  (
    n1780,
    n536
  );


  not
  g729
  (
    n819,
    n551
  );


  not
  g730
  (
    n1588,
    n551
  );


  not
  g731
  (
    n872,
    n246
  );


  not
  g732
  (
    n805,
    n350
  );


  not
  g733
  (
    n987,
    n237
  );


  buf
  g734
  (
    n1258,
    n523
  );


  not
  g735
  (
    n1679,
    n638
  );


  buf
  g736
  (
    n1133,
    n356
  );


  buf
  g737
  (
    n1511,
    n458
  );


  buf
  g738
  (
    n708,
    n470
  );


  not
  g739
  (
    n1731,
    n513
  );


  buf
  g740
  (
    n976,
    n292
  );


  buf
  g741
  (
    n663,
    n614
  );


  not
  g742
  (
    n760,
    n237
  );


  not
  g743
  (
    n1799,
    n248
  );


  buf
  g744
  (
    n1001,
    n438
  );


  buf
  g745
  (
    n1030,
    n172
  );


  buf
  g746
  (
    KeyWire_0_48,
    n365
  );


  not
  g747
  (
    n1127,
    n215
  );


  not
  g748
  (
    n1858,
    n191
  );


  not
  g749
  (
    n1490,
    n581
  );


  buf
  g750
  (
    n1212,
    n211
  );


  not
  g751
  (
    n1178,
    n351
  );


  not
  g752
  (
    n1699,
    n240
  );


  not
  g753
  (
    n1690,
    n313
  );


  buf
  g754
  (
    n874,
    n396
  );


  buf
  g755
  (
    n1445,
    n323
  );


  buf
  g756
  (
    n1604,
    n290
  );


  not
  g757
  (
    n1581,
    n377
  );


  buf
  g758
  (
    n767,
    n487
  );


  not
  g759
  (
    n1682,
    n422
  );


  buf
  g760
  (
    n1834,
    n584
  );


  not
  g761
  (
    n934,
    n159
  );


  buf
  g762
  (
    n1671,
    n255
  );


  buf
  g763
  (
    n1274,
    n561
  );


  not
  g764
  (
    n1875,
    n272
  );


  buf
  g765
  (
    n705,
    n295
  );


  not
  g766
  (
    KeyWire_0_39,
    n455
  );


  not
  g767
  (
    n1771,
    n219
  );


  buf
  g768
  (
    n1820,
    n613
  );


  buf
  g769
  (
    n1003,
    n440
  );


  buf
  g770
  (
    n894,
    n521
  );


  not
  g771
  (
    n912,
    n443
  );


  not
  g772
  (
    n1597,
    n553
  );


  not
  g773
  (
    KeyWire_0_21,
    n411
  );


  buf
  g774
  (
    n1053,
    n409
  );


  not
  g775
  (
    n1341,
    n358
  );


  not
  g776
  (
    n907,
    n575
  );


  buf
  g777
  (
    n1641,
    n193
  );


  buf
  g778
  (
    n1222,
    n289
  );


  not
  g779
  (
    n1842,
    n230
  );


  buf
  g780
  (
    n1600,
    n281
  );


  buf
  g781
  (
    n1951,
    n394
  );


  buf
  g782
  (
    n1252,
    n648
  );


  buf
  g783
  (
    n871,
    n622
  );


  not
  g784
  (
    n844,
    n325
  );


  buf
  g785
  (
    KeyWire_0_61,
    n185
  );


  not
  g786
  (
    KeyWire_0_20,
    n253
  );


  not
  g787
  (
    n660,
    n562
  );


  buf
  g788
  (
    n1175,
    n580
  );


  buf
  g789
  (
    n1849,
    n291
  );


  buf
  g790
  (
    n919,
    n190
  );


  not
  g791
  (
    n1047,
    n316
  );


  not
  g792
  (
    n1478,
    n644
  );


  not
  g793
  (
    n892,
    n608
  );


  buf
  g794
  (
    n1256,
    n480
  );


  not
  g795
  (
    n1668,
    n501
  );


  not
  g796
  (
    n1878,
    n625
  );


  not
  g797
  (
    n1461,
    n465
  );


  buf
  g798
  (
    n1795,
    n424
  );


  not
  g799
  (
    n1042,
    n337
  );


  buf
  g800
  (
    n1479,
    n247
  );


  buf
  g801
  (
    n1678,
    n533
  );


  buf
  g802
  (
    n1441,
    n216
  );


  buf
  g803
  (
    n1935,
    n561
  );


  buf
  g804
  (
    n1903,
    n532
  );


  buf
  g805
  (
    n1395,
    n587
  );


  buf
  g806
  (
    n1230,
    n315
  );


  buf
  g807
  (
    n1598,
    n292
  );


  not
  g808
  (
    n1687,
    n439
  );


  not
  g809
  (
    n1570,
    n157
  );


  buf
  g810
  (
    n1655,
    n270
  );


  buf
  g811
  (
    n1176,
    n200
  );


  buf
  g812
  (
    n1893,
    n297
  );


  not
  g813
  (
    n1354,
    n321
  );


  not
  g814
  (
    n1157,
    n605
  );


  not
  g815
  (
    n975,
    n284
  );


  buf
  g816
  (
    n938,
    n320
  );


  buf
  g817
  (
    n838,
    n624
  );


  buf
  g818
  (
    n1753,
    n167
  );


  buf
  g819
  (
    n1683,
    n434
  );


  not
  g820
  (
    n718,
    n321
  );


  buf
  g821
  (
    n995,
    n265
  );


  not
  g822
  (
    n867,
    n225
  );


  not
  g823
  (
    n1602,
    n194
  );


  buf
  g824
  (
    n1205,
    n239
  );


  buf
  g825
  (
    n1526,
    n516
  );


  not
  g826
  (
    n791,
    n523
  );


  buf
  g827
  (
    n1757,
    n409
  );


  not
  g828
  (
    n1867,
    n209
  );


  buf
  g829
  (
    n1424,
    n475
  );


  not
  g830
  (
    n1697,
    n314
  );


  buf
  g831
  (
    n1688,
    n540
  );


  buf
  g832
  (
    n1606,
    n558
  );


  not
  g833
  (
    n1010,
    n206
  );


  buf
  g834
  (
    n1790,
    n364
  );


  not
  g835
  (
    n905,
    n297
  );


  not
  g836
  (
    n1802,
    n184
  );


  buf
  g837
  (
    n1218,
    n347
  );


  not
  g838
  (
    n861,
    n257
  );


  buf
  g839
  (
    n1476,
    n477
  );


  not
  g840
  (
    n1139,
    n313
  );


  not
  g841
  (
    n1324,
    n473
  );


  buf
  g842
  (
    n736,
    n546
  );


  buf
  g843
  (
    n1015,
    n177
  );


  buf
  g844
  (
    n1355,
    n610
  );


  not
  g845
  (
    n1586,
    n509
  );


  not
  g846
  (
    n1735,
    n250
  );


  buf
  g847
  (
    n1240,
    n342
  );


  not
  g848
  (
    n977,
    n208
  );


  buf
  g849
  (
    n1173,
    n347
  );


  not
  g850
  (
    n1114,
    n430
  );


  not
  g851
  (
    n1457,
    n640
  );


  not
  g852
  (
    n1826,
    n236
  );


  buf
  g853
  (
    n733,
    n163
  );


  not
  g854
  (
    n1080,
    n432
  );


  buf
  g855
  (
    n978,
    n497
  );


  not
  g856
  (
    n847,
    n244
  );


  not
  g857
  (
    n1238,
    n452
  );


  not
  g858
  (
    n1458,
    n445
  );


  not
  g859
  (
    n1729,
    n567
  );


  not
  g860
  (
    n1019,
    n226
  );


  not
  g861
  (
    n1366,
    n399
  );


  buf
  g862
  (
    n1338,
    n517
  );


  not
  g863
  (
    n1825,
    n603
  );


  not
  g864
  (
    n1898,
    n554
  );


  not
  g865
  (
    n1810,
    n508
  );


  buf
  g866
  (
    n700,
    n612
  );


  not
  g867
  (
    n780,
    n635
  );


  not
  g868
  (
    n1486,
    n247
  );


  buf
  g869
  (
    n1028,
    n475
  );


  buf
  g870
  (
    n1309,
    n442
  );


  not
  g871
  (
    n1577,
    n560
  );


  buf
  g872
  (
    n1652,
    n643
  );


  not
  g873
  (
    n1242,
    n545
  );


  not
  g874
  (
    n1545,
    n544
  );


  not
  g875
  (
    n953,
    n407
  );


  not
  g876
  (
    n1813,
    n271
  );


  not
  g877
  (
    n1818,
    n377
  );


  not
  g878
  (
    n722,
    n274
  );


  not
  g879
  (
    n1125,
    n512
  );


  not
  g880
  (
    n653,
    n398
  );


  not
  g881
  (
    n1748,
    n502
  );


  not
  g882
  (
    n1013,
    n476
  );


  not
  g883
  (
    n899,
    n499
  );


  not
  g884
  (
    n942,
    n351
  );


  buf
  g885
  (
    n1793,
    n467
  );


  not
  g886
  (
    n1980,
    n428
  );


  buf
  g887
  (
    n728,
    n485
  );


  not
  g888
  (
    n1785,
    n303
  );


  not
  g889
  (
    KeyWire_0_19,
    n617
  );


  not
  g890
  (
    n1854,
    n571
  );


  buf
  g891
  (
    n724,
    n428
  );


  buf
  g892
  (
    n1689,
    n308
  );


  not
  g893
  (
    n1337,
    n288
  );


  buf
  g894
  (
    n703,
    n172
  );


  not
  g895
  (
    n1546,
    n321
  );


  not
  g896
  (
    n792,
    n599
  );


  not
  g897
  (
    n1966,
    n173
  );


  buf
  g898
  (
    n726,
    n482
  );


  buf
  g899
  (
    n1094,
    n621
  );


  buf
  g900
  (
    n1624,
    n422
  );


  buf
  g901
  (
    n888,
    n388
  );


  not
  g902
  (
    n1208,
    n301
  );


  buf
  g903
  (
    n1405,
    n579
  );


  buf
  g904
  (
    n1612,
    n648
  );


  buf
  g905
  (
    n1103,
    n609
  );


  not
  g906
  (
    n1656,
    n207
  );


  not
  g907
  (
    KeyWire_0_62,
    n615
  );


  not
  g908
  (
    n1249,
    n537
  );


  not
  g909
  (
    n1477,
    n201
  );


  not
  g910
  (
    n1056,
    n214
  );


  buf
  g911
  (
    n936,
    n480
  );


  not
  g912
  (
    n1043,
    n416
  );


  buf
  g913
  (
    n1194,
    n259
  );


  buf
  g914
  (
    n821,
    n373
  );


  buf
  g915
  (
    n1033,
    n213
  );


  buf
  g916
  (
    n1631,
    n610
  );


  buf
  g917
  (
    n1862,
    n424
  );


  buf
  g918
  (
    n1784,
    n420
  );


  not
  g919
  (
    n1452,
    n283
  );


  buf
  g920
  (
    n1685,
    n633
  );


  not
  g921
  (
    n954,
    n217
  );


  buf
  g922
  (
    n926,
    n564
  );


  not
  g923
  (
    n834,
    n569
  );


  not
  g924
  (
    n1946,
    n224
  );


  not
  g925
  (
    n1278,
    n277
  );


  buf
  g926
  (
    n1404,
    n235
  );


  not
  g927
  (
    KeyWire_0_35,
    n369
  );


  buf
  g928
  (
    n1659,
    n237
  );


  not
  g929
  (
    n1741,
    n293
  );


  buf
  g930
  (
    n1848,
    n637
  );


  not
  g931
  (
    n967,
    n629
  );


  not
  g932
  (
    n1276,
    n546
  );


  not
  g933
  (
    n1409,
    n216
  );


  not
  g934
  (
    n1430,
    n277
  );


  not
  g935
  (
    n772,
    n306
  );


  buf
  g936
  (
    n1589,
    n486
  );


  not
  g937
  (
    n1675,
    n304
  );


  buf
  g938
  (
    n973,
    n495
  );


  buf
  g939
  (
    n1934,
    n303
  );


  buf
  g940
  (
    n880,
    n249
  );


  buf
  g941
  (
    n1937,
    n191
  );


  not
  g942
  (
    n1823,
    n453
  );


  buf
  g943
  (
    n949,
    n367
  );


  not
  g944
  (
    n1266,
    n164
  );


  not
  g945
  (
    n1809,
    n448
  );


  buf
  g946
  (
    n828,
    n507
  );


  not
  g947
  (
    n744,
    n429
  );


  buf
  g948
  (
    n751,
    n530
  );


  buf
  g949
  (
    n1185,
    n488
  );


  buf
  g950
  (
    n1093,
    n370
  );


  not
  g951
  (
    n1921,
    n192
  );


  not
  g952
  (
    n1464,
    n163
  );


  buf
  g953
  (
    n1263,
    n318
  );


  not
  g954
  (
    n1645,
    n561
  );


  buf
  g955
  (
    n1707,
    n379
  );


  not
  g956
  (
    n801,
    n644
  );


  not
  g957
  (
    n1090,
    n205
  );


  not
  g958
  (
    n1498,
    n182
  );


  not
  g959
  (
    n1106,
    n467
  );


  buf
  g960
  (
    n712,
    n354
  );


  buf
  g961
  (
    n1286,
    n604
  );


  not
  g962
  (
    n1710,
    n542
  );


  not
  g963
  (
    n1345,
    n241
  );


  buf
  g964
  (
    n1416,
    n231
  );


  not
  g965
  (
    n1669,
    n234
  );


  not
  g966
  (
    n1654,
    n428
  );


  not
  g967
  (
    n1034,
    n522
  );


  not
  g968
  (
    n740,
    n509
  );


  not
  g969
  (
    n687,
    n496
  );


  not
  g970
  (
    n1305,
    n443
  );


  not
  g971
  (
    n1911,
    n253
  );


  buf
  g972
  (
    n1277,
    n626
  );


  not
  g973
  (
    n1350,
    n426
  );


  buf
  g974
  (
    n1067,
    n308
  );


  buf
  g975
  (
    n1446,
    n459
  );


  buf
  g976
  (
    n842,
    n610
  );


  not
  g977
  (
    n1484,
    n465
  );


  not
  g978
  (
    n1703,
    n298
  );


  buf
  g979
  (
    n1952,
    n404
  );


  buf
  g980
  (
    n885,
    n512
  );


  buf
  g981
  (
    n1373,
    n330
  );


  buf
  g982
  (
    n886,
    n378
  );


  buf
  g983
  (
    n889,
    n289
  );


  buf
  g984
  (
    n1129,
    n538
  );


  not
  g985
  (
    n1643,
    n480
  );


  not
  g986
  (
    n1475,
    n386
  );


  buf
  g987
  (
    n865,
    n450
  );


  buf
  g988
  (
    n1403,
    n294
  );


  not
  g989
  (
    n1065,
    n632
  );


  not
  g990
  (
    n1510,
    n380
  );


  buf
  g991
  (
    n854,
    n586
  );


  buf
  g992
  (
    n674,
    n194
  );


  buf
  g993
  (
    n1775,
    n639
  );


  buf
  g994
  (
    n1299,
    n307
  );


  not
  g995
  (
    n1413,
    n366
  );


  buf
  g996
  (
    n901,
    n643
  );


  not
  g997
  (
    n920,
    n360
  );


  not
  g998
  (
    n1326,
    n469
  );


  buf
  g999
  (
    n909,
    n349
  );


  buf
  g1000
  (
    n1569,
    n283
  );


  buf
  g1001
  (
    n1894,
    n485
  );


  not
  g1002
  (
    n918,
    n401
  );


  not
  g1003
  (
    n1717,
    n286
  );


  buf
  g1004
  (
    n1932,
    n506
  );


  not
  g1005
  (
    n1436,
    n243
  );


  not
  g1006
  (
    n1228,
    n415
  );


  not
  g1007
  (
    n1359,
    n367
  );


  buf
  g1008
  (
    n1740,
    n382
  );


  buf
  g1009
  (
    n1215,
    n188
  );


  buf
  g1010
  (
    n1247,
    n230
  );


  not
  g1011
  (
    n666,
    n393
  );


  not
  g1012
  (
    n1673,
    n517
  );


  not
  g1013
  (
    n1899,
    n651
  );


  buf
  g1014
  (
    n1184,
    n550
  );


  buf
  g1015
  (
    n1349,
    n273
  );


  buf
  g1016
  (
    n1343,
    n582
  );


  buf
  g1017
  (
    n1949,
    n604
  );


  not
  g1018
  (
    n775,
    n260
  );


  buf
  g1019
  (
    KeyWire_0_1,
    n356
  );


  buf
  g1020
  (
    n1235,
    n411
  );


  buf
  g1021
  (
    n778,
    n624
  );


  not
  g1022
  (
    n1315,
    n322
  );


  not
  g1023
  (
    n1421,
    n210
  );


  not
  g1024
  (
    n1162,
    n505
  );


  buf
  g1025
  (
    n1102,
    n403
  );


  buf
  g1026
  (
    n896,
    n461
  );


  not
  g1027
  (
    n988,
    n288
  );


  buf
  g1028
  (
    n1776,
    n268
  );


  buf
  g1029
  (
    n939,
    n519
  );


  not
  g1030
  (
    n1027,
    n357
  );


  buf
  g1031
  (
    n1142,
    n596
  );


  not
  g1032
  (
    n1664,
    n268
  );


  not
  g1033
  (
    n1508,
    n192
  );


  buf
  g1034
  (
    n753,
    n593
  );


  buf
  g1035
  (
    n765,
    n161
  );


  buf
  g1036
  (
    n1059,
    n379
  );


  not
  g1037
  (
    n869,
    n231
  );


  not
  g1038
  (
    n750,
    n588
  );


  not
  g1039
  (
    n940,
    n552
  );


  not
  g1040
  (
    n1143,
    n434
  );


  buf
  g1041
  (
    n1302,
    n471
  );


  buf
  g1042
  (
    n1516,
    n361
  );


  not
  g1043
  (
    n678,
    n340
  );


  not
  g1044
  (
    n1112,
    n189
  );


  not
  g1045
  (
    n1041,
    n395
  );


  buf
  g1046
  (
    n1537,
    n379
  );


  not
  g1047
  (
    n1200,
    n545
  );


  not
  g1048
  (
    n1601,
    n344
  );


  buf
  g1049
  (
    n1420,
    n169
  );


  not
  g1050
  (
    n1715,
    n370
  );


  buf
  g1051
  (
    n1426,
    n375
  );


  buf
  g1052
  (
    n1367,
    n553
  );


  buf
  g1053
  (
    n686,
    n429
  );


  buf
  g1054
  (
    n853,
    n646
  );


  buf
  g1055
  (
    n1948,
    n529
  );


  buf
  g1056
  (
    n1883,
    n518
  );


  buf
  g1057
  (
    n709,
    n269
  );


  buf
  g1058
  (
    n1742,
    n353
  );


  buf
  g1059
  (
    n1877,
    n331
  );


  buf
  g1060
  (
    n1797,
    n462
  );


  not
  g1061
  (
    n1022,
    n249
  );


  not
  g1062
  (
    n1614,
    n628
  );


  buf
  g1063
  (
    n1189,
    n328
  );


  not
  g1064
  (
    n1294,
    n407
  );


  not
  g1065
  (
    n1487,
    n572
  );


  buf
  g1066
  (
    n1499,
    n254
  );


  not
  g1067
  (
    n1198,
    n336
  );


  not
  g1068
  (
    n1565,
    n244
  );


  buf
  g1069
  (
    n1626,
    n197
  );


  not
  g1070
  (
    n1765,
    n204
  );


  buf
  g1071
  (
    n1817,
    n444
  );


  buf
  g1072
  (
    n1483,
    n526
  );


  buf
  g1073
  (
    n1134,
    n264
  );


  buf
  g1074
  (
    KeyWire_0_15,
    n626
  );


  buf
  g1075
  (
    n1298,
    n481
  );


  buf
  g1076
  (
    n1725,
    n464
  );


  buf
  g1077
  (
    n1393,
    n606
  );


  buf
  g1078
  (
    n877,
    n551
  );


  not
  g1079
  (
    n719,
    n455
  );


  not
  g1080
  (
    KeyWire_0_63,
    n164
  );


  not
  g1081
  (
    n1706,
    n393
  );


  buf
  g1082
  (
    n725,
    n639
  );


  buf
  g1083
  (
    n1036,
    n565
  );


  not
  g1084
  (
    n1621,
    n464
  );


  buf
  g1085
  (
    n682,
    n470
  );


  not
  g1086
  (
    n1855,
    n165
  );


  not
  g1087
  (
    n667,
    n320
  );


  not
  g1088
  (
    n688,
    n214
  );


  buf
  g1089
  (
    n884,
    n549
  );


  buf
  g1090
  (
    n955,
    n258
  );


  buf
  g1091
  (
    n1838,
    n157
  );


  buf
  g1092
  (
    n1847,
    n563
  );


  buf
  g1093
  (
    n1213,
    n550
  );


  not
  g1094
  (
    n904,
    n391
  );


  not
  g1095
  (
    n1168,
    n467
  );


  not
  g1096
  (
    n1856,
    n279
  );


  not
  g1097
  (
    n1078,
    n163
  );


  buf
  g1098
  (
    n1957,
    n616
  );


  buf
  g1099
  (
    n1726,
    n398
  );


  not
  g1100
  (
    n1290,
    n567
  );


  buf
  g1101
  (
    n758,
    n273
  );


  not
  g1102
  (
    n1223,
    n640
  );


  buf
  g1103
  (
    n1829,
    n275
  );


  buf
  g1104
  (
    n1459,
    n557
  );


  not
  g1105
  (
    n1651,
    n288
  );


  buf
  g1106
  (
    n696,
    n383
  );


  not
  g1107
  (
    n1924,
    n289
  );


  buf
  g1108
  (
    n1300,
    n211
  );


  not
  g1109
  (
    n1061,
    n425
  );


  buf
  g1110
  (
    n1049,
    n468
  );


  buf
  g1111
  (
    n1088,
    n421
  );


  buf
  g1112
  (
    n743,
    n230
  );


  not
  g1113
  (
    n1518,
    n524
  );


  buf
  g1114
  (
    n1419,
    n165
  );


  not
  g1115
  (
    n1677,
    n381
  );


  buf
  g1116
  (
    n1559,
    n306
  );


  not
  g1117
  (
    n1255,
    n297
  );


  not
  g1118
  (
    n957,
    n183
  );


  not
  g1119
  (
    n701,
    n546
  );


  buf
  g1120
  (
    KeyWire_0_30,
    n557
  );


  not
  g1121
  (
    n866,
    n402
  );


  not
  g1122
  (
    n1591,
    n641
  );


  not
  g1123
  (
    n1469,
    n408
  );


  not
  g1124
  (
    n1226,
    n518
  );


  not
  g1125
  (
    n1066,
    n320
  );


  not
  g1126
  (
    n1613,
    n282
  );


  buf
  g1127
  (
    n1344,
    n368
  );


  buf
  g1128
  (
    n826,
    n534
  );


  not
  g1129
  (
    n1021,
    n462
  );


  buf
  g1130
  (
    n1288,
    n487
  );


  buf
  g1131
  (
    n1493,
    n450
  );


  not
  g1132
  (
    n929,
    n364
  );


  not
  g1133
  (
    n1146,
    n649
  );


  buf
  g1134
  (
    n1939,
    n224
  );


  buf
  g1135
  (
    n1901,
    n295
  );


  buf
  g1136
  (
    n1730,
    n417
  );


  buf
  g1137
  (
    n1204,
    n312
  );


  buf
  g1138
  (
    n1593,
    n593
  );


  not
  g1139
  (
    n1646,
    n560
  );


  not
  g1140
  (
    n1234,
    n631
  );


  buf
  g1141
  (
    n1976,
    n192
  );


  not
  g1142
  (
    n1772,
    n220
  );


  not
  g1143
  (
    n1060,
    n170
  );


  not
  g1144
  (
    n1530,
    n215
  );


  buf
  g1145
  (
    n1040,
    n526
  );


  buf
  g1146
  (
    n994,
    n212
  );


  not
  g1147
  (
    n1549,
    n349
  );


  buf
  g1148
  (
    n1072,
    n285
  );


  buf
  g1149
  (
    n1798,
    n521
  );


  not
  g1150
  (
    n1308,
    n383
  );


  not
  g1151
  (
    n1540,
    n442
  );


  buf
  g1152
  (
    n1161,
    n415
  );


  not
  g1153
  (
    n933,
    n167
  );


  buf
  g1154
  (
    n1830,
    n494
  );


  not
  g1155
  (
    n927,
    n315
  );


  not
  g1156
  (
    n1148,
    n439
  );


  not
  g1157
  (
    n699,
    n187
  );


  not
  g1158
  (
    n1839,
    n561
  );


  not
  g1159
  (
    n983,
    n419
  );


  buf
  g1160
  (
    n1378,
    n263
  );


  not
  g1161
  (
    n1564,
    n633
  );


  buf
  g1162
  (
    n1064,
    n219
  );


  buf
  g1163
  (
    n1038,
    n455
  );


  buf
  g1164
  (
    n1558,
    n436
  );


  not
  g1165
  (
    n1259,
    n640
  );


  not
  g1166
  (
    n1272,
    n564
  );


  not
  g1167
  (
    n1000,
    n516
  );


  not
  g1168
  (
    n1046,
    n389
  );


  not
  g1169
  (
    n1119,
    n159
  );


  not
  g1170
  (
    n1370,
    n164
  );


  buf
  g1171
  (
    n1548,
    n303
  );


  not
  g1172
  (
    n704,
    n193
  );


  buf
  g1173
  (
    n928,
    n419
  );


  buf
  g1174
  (
    n1694,
    n404
  );


  not
  g1175
  (
    n1372,
    n484
  );


  buf
  g1176
  (
    n1696,
    n295
  );


  not
  g1177
  (
    n1714,
    n433
  );


  not
  g1178
  (
    n1749,
    n564
  );


  buf
  g1179
  (
    n1328,
    n256
  );


  buf
  g1180
  (
    n1942,
    n635
  );


  not
  g1181
  (
    n833,
    n245
  );


  not
  g1182
  (
    n1583,
    n267
  );


  buf
  g1183
  (
    n1562,
    n190
  );


  buf
  g1184
  (
    n1736,
    n261
  );


  buf
  g1185
  (
    n1332,
    n423
  );


  buf
  g1186
  (
    n1958,
    n279
  );


  not
  g1187
  (
    n1681,
    n515
  );


  not
  g1188
  (
    n1680,
    n481
  );


  buf
  g1189
  (
    n1914,
    n610
  );


  buf
  g1190
  (
    n1743,
    n336
  );


  not
  g1191
  (
    n1663,
    n498
  );


  buf
  g1192
  (
    n1352,
    n339
  );


  not
  g1193
  (
    n843,
    n484
  );


  not
  g1194
  (
    n670,
    n285
  );


  not
  g1195
  (
    n1414,
    n372
  );


  buf
  g1196
  (
    n1527,
    n217
  );


  buf
  g1197
  (
    n945,
    n576
  );


  buf
  g1198
  (
    n1812,
    n203
  );


  not
  g1199
  (
    n858,
    n490
  );


  not
  g1200
  (
    n1608,
    n456
  );


  buf
  g1201
  (
    n810,
    n293
  );


  not
  g1202
  (
    n773,
    n304
  );


  not
  g1203
  (
    n1388,
    n304
  );


  not
  g1204
  (
    n1928,
    n590
  );


  not
  g1205
  (
    n1159,
    n367
  );


  buf
  g1206
  (
    n921,
    n300
  );


  not
  g1207
  (
    n1851,
    n177
  );


  buf
  g1208
  (
    n1896,
    n311
  );


  buf
  g1209
  (
    n1291,
    n600
  );


  not
  g1210
  (
    n1362,
    n648
  );


  buf
  g1211
  (
    n1639,
    n576
  );


  not
  g1212
  (
    n716,
    n282
  );


  buf
  g1213
  (
    n1210,
    n332
  );


  not
  g1214
  (
    n1246,
    n594
  );


  not
  g1215
  (
    n1587,
    n175
  );


  buf
  g1216
  (
    n1435,
    n470
  );


  buf
  g1217
  (
    n1020,
    n501
  );


  buf
  g1218
  (
    n1716,
    n353
  );


  buf
  g1219
  (
    n763,
    n403
  );


  buf
  g1220
  (
    n1807,
    n318
  );


  buf
  g1221
  (
    n1151,
    n181
  );


  not
  g1222
  (
    n1632,
    n211
  );


  buf
  g1223
  (
    n1400,
    n245
  );


  buf
  g1224
  (
    n1579,
    n432
  );


  buf
  g1225
  (
    n1126,
    n447
  );


  buf
  g1226
  (
    n1331,
    n522
  );


  not
  g1227
  (
    n1482,
    n489
  );


  buf
  g1228
  (
    n1243,
    n348
  );


  not
  g1229
  (
    n1768,
    n311
  );


  not
  g1230
  (
    n1221,
    n436
  );


  buf
  g1231
  (
    n932,
    n412
  );


  not
  g1232
  (
    n1846,
    n507
  );


  buf
  g1233
  (
    n1622,
    n554
  );


  buf
  g1234
  (
    n1437,
    n540
  );


  not
  g1235
  (
    n1432,
    n335
  );


  not
  g1236
  (
    n1206,
    n242
  );


  buf
  g1237
  (
    n1293,
    n563
  );


  not
  g1238
  (
    n1751,
    n389
  );


  buf
  g1239
  (
    n806,
    n315
  );


  not
  g1240
  (
    n1137,
    n241
  );


  buf
  g1241
  (
    n1023,
    n198
  );


  not
  g1242
  (
    n713,
    n263
  );


  buf
  g1243
  (
    n1852,
    n169
  );


  buf
  g1244
  (
    n1241,
    n638
  );


  buf
  g1245
  (
    n1611,
    n632
  );


  not
  g1246
  (
    n1187,
    n628
  );


  buf
  g1247
  (
    n1889,
    n553
  );


  buf
  g1248
  (
    n1506,
    n530
  );


  not
  g1249
  (
    n1837,
    n430
  );


  buf
  g1250
  (
    n1186,
    n526
  );


  buf
  g1251
  (
    n669,
    n331
  );


  not
  g1252
  (
    n1181,
    n616
  );


  not
  g1253
  (
    n1520,
    n186
  );


  not
  g1254
  (
    n1543,
    n363
  );


  not
  g1255
  (
    n1284,
    n400
  );


  not
  g1256
  (
    n1723,
    n640
  );


  not
  g1257
  (
    n1050,
    n167
  );


  buf
  g1258
  (
    n1402,
    n573
  );


  not
  g1259
  (
    n868,
    n492
  );


  buf
  g1260
  (
    n1348,
    n541
  );


  buf
  g1261
  (
    n657,
    n298
  );


  buf
  g1262
  (
    KeyWire_0_55,
    n499
  );


  buf
  g1263
  (
    n925,
    n385
  );


  not
  g1264
  (
    n1004,
    n338
  );


  not
  g1265
  (
    n1759,
    n314
  );


  buf
  g1266
  (
    n1500,
    n317
  );


  buf
  g1267
  (
    n1783,
    n266
  );


  not
  g1268
  (
    n1431,
    n170
  );


  buf
  g1269
  (
    n1665,
    n589
  );


  not
  g1270
  (
    n1227,
    n229
  );


  not
  g1271
  (
    n1016,
    n178
  );


  not
  g1272
  (
    n673,
    n503
  );


  buf
  g1273
  (
    n1082,
    n637
  );


  not
  g1274
  (
    n1375,
    n231
  );


  not
  g1275
  (
    n1970,
    n404
  );


  not
  g1276
  (
    n989,
    n275
  );


  not
  g1277
  (
    n691,
    n413
  );


  not
  g1278
  (
    n1342,
    n334
  );


  not
  g1279
  (
    n1844,
    n559
  );


  not
  g1280
  (
    n757,
    n397
  );


  not
  g1281
  (
    n781,
    n417
  );


  buf
  g1282
  (
    n1160,
    n388
  );


  buf
  g1283
  (
    n961,
    n413
  );


  not
  g1284
  (
    n970,
    n356
  );


  buf
  g1285
  (
    n1201,
    n486
  );


  not
  g1286
  (
    n968,
    n617
  );


  buf
  g1287
  (
    n1261,
    n282
  );


  not
  g1288
  (
    n1296,
    n283
  );


  not
  g1289
  (
    n1190,
    n538
  );


  buf
  g1290
  (
    n1130,
    n587
  );


  buf
  g1291
  (
    n1533,
    n345
  );


  buf
  g1292
  (
    n887,
    n418
  );


  buf
  g1293
  (
    n764,
    n520
  );


  buf
  g1294
  (
    n1832,
    n276
  );


  buf
  g1295
  (
    n1578,
    n447
  );


  buf
  g1296
  (
    n1164,
    n629
  );


  and
  g1297
  (
    n685,
    n261,
    n442
  );


  nand
  g1298
  (
    KeyWire_0_36,
    n271,
    n485
  );


  nand
  g1299
  (
    n761,
    n390,
    n339
  );


  or
  g1300
  (
    n1794,
    n573,
    n296
  );


  xor
  g1301
  (
    n1008,
    n292,
    n488
  );


  nor
  g1302
  (
    n1002,
    n362,
    n536
  );


  nand
  g1303
  (
    KeyWire_0_7,
    n589,
    n571
  );


  or
  g1304
  (
    n1888,
    n424,
    n577
  );


  xnor
  g1305
  (
    n1750,
    n318,
    n651
  );


  nand
  g1306
  (
    n675,
    n300,
    n410
  );


  or
  g1307
  (
    n770,
    n491,
    n542
  );


  or
  g1308
  (
    n1502,
    n582,
    n557
  );


  and
  g1309
  (
    n1915,
    n270,
    n449
  );


  xnor
  g1310
  (
    n1361,
    n286,
    n555
  );


  xor
  g1311
  (
    n1026,
    n335,
    n454
  );


  and
  g1312
  (
    n893,
    n343,
    n441
  );


  xor
  g1313
  (
    n1462,
    n351,
    n175
  );


  nand
  g1314
  (
    n1930,
    n267,
    n184
  );


  or
  g1315
  (
    n1764,
    n170,
    n354
  );


  nor
  g1316
  (
    n1307,
    n342,
    n417
  );


  or
  g1317
  (
    n913,
    n232,
    n348
  );


  or
  g1318
  (
    n1188,
    n326,
    n584
  );


  xor
  g1319
  (
    n1444,
    n461,
    n497
  );


  or
  g1320
  (
    n1525,
    n375,
    n245
  );


  nand
  g1321
  (
    n1131,
    n500,
    n443
  );


  xnor
  g1322
  (
    n1456,
    n474,
    n406
  );


  nor
  g1323
  (
    n1113,
    n496,
    n482
  );


  and
  g1324
  (
    n950,
    n486,
    n223
  );


  xor
  g1325
  (
    n732,
    n618,
    n605
  );


  and
  g1326
  (
    n1755,
    n192,
    n491
  );


  and
  g1327
  (
    n1394,
    n484,
    n514
  );


  xnor
  g1328
  (
    n1100,
    n633,
    n278
  );


  nor
  g1329
  (
    n1513,
    n619,
    n577
  );


  xnor
  g1330
  (
    n1473,
    n325,
    n634
  );


  xor
  g1331
  (
    n1781,
    n194,
    n303
  );


  nand
  g1332
  (
    n813,
    n223,
    n441
  );


  nor
  g1333
  (
    n1163,
    n541,
    n459
  );


  nor
  g1334
  (
    n1169,
    n583,
    n513
  );


  or
  g1335
  (
    n1917,
    n507,
    n601
  );


  xnor
  g1336
  (
    n1122,
    n506,
    n596
  );


  xor
  g1337
  (
    n1860,
    n500,
    n325
  );


  nor
  g1338
  (
    n1233,
    n249,
    n350
  );


  nand
  g1339
  (
    n655,
    n489,
    n392
  );


  xor
  g1340
  (
    n1440,
    n184,
    n529
  );


  nor
  g1341
  (
    n1031,
    n533,
    n522
  );


  or
  g1342
  (
    n1322,
    n493,
    n503
  );


  xnor
  g1343
  (
    n1806,
    n240,
    n298
  );


  nand
  g1344
  (
    n1566,
    n536,
    n262
  );


  nor
  g1345
  (
    n804,
    n255,
    n346
  );


  xnor
  g1346
  (
    n1260,
    n568,
    n162
  );


  nand
  g1347
  (
    n1672,
    n330,
    n169
  );


  xor
  g1348
  (
    n1850,
    n630,
    n251
  );


  and
  g1349
  (
    n1074,
    n600,
    n515
  );


  nor
  g1350
  (
    n1501,
    n547,
    n606
  );


  or
  g1351
  (
    n1438,
    n249,
    n649
  );


  nor
  g1352
  (
    n1979,
    n257,
    n309
  );


  nor
  g1353
  (
    KeyWire_0_24,
    n410,
    n568
  );


  xor
  g1354
  (
    n1560,
    n604,
    n408
  );


  nand
  g1355
  (
    n814,
    n532,
    n369
  );


  xnor
  g1356
  (
    n1154,
    n218,
    n575
  );


  xor
  g1357
  (
    n1336,
    n645,
    n395
  );


  and
  g1358
  (
    n1709,
    n186,
    n461
  );


  nand
  g1359
  (
    n1900,
    n334,
    n451
  );


  xnor
  g1360
  (
    n1728,
    n445,
    n503
  );


  xor
  g1361
  (
    n1058,
    n453,
    n434
  );


  and
  g1362
  (
    n1827,
    n536,
    n175
  );


  or
  g1363
  (
    n1572,
    n491,
    n476
  );


  xnor
  g1364
  (
    n1037,
    n478,
    n648
  );


  or
  g1365
  (
    n738,
    n511,
    n513
  );


  or
  g1366
  (
    n749,
    n242,
    n427
  );


  xor
  g1367
  (
    n1938,
    n243,
    n391
  );


  xnor
  g1368
  (
    n717,
    n389,
    n179
  );


  xor
  g1369
  (
    n1845,
    n159,
    n376
  );


  nor
  g1370
  (
    n1891,
    n273,
    n566
  );


  xnor
  g1371
  (
    n1032,
    n624,
    n569
  );


  nor
  g1372
  (
    n1267,
    n174,
    n220
  );


  or
  g1373
  (
    n1087,
    n408,
    n341
  );


  nand
  g1374
  (
    KeyWire_0_54,
    n441,
    n575
  );


  and
  g1375
  (
    n1199,
    n448,
    n524
  );


  nand
  g1376
  (
    n1491,
    n578,
    n182
  );


  nor
  g1377
  (
    n1317,
    n545,
    n635
  );


  nand
  g1378
  (
    n1627,
    n520,
    n507
  );


  xnor
  g1379
  (
    n1876,
    n175,
    n284
  );


  nand
  g1380
  (
    n1451,
    n327,
    n392
  );


  and
  g1381
  (
    n1796,
    n465,
    n426
  );


  xnor
  g1382
  (
    n1024,
    n468,
    n500
  );


  nor
  g1383
  (
    n1580,
    n595,
    n265
  );


  and
  g1384
  (
    n1922,
    n231,
    n631
  );


  nor
  g1385
  (
    n1285,
    n431,
    n354
  );


  xor
  g1386
  (
    n803,
    n482,
    n338
  );


  xnor
  g1387
  (
    n808,
    n374,
    n277
  );


  or
  g1388
  (
    n1408,
    n179,
    n207
  );


  xor
  g1389
  (
    n1843,
    n565,
    n185
  );


  nor
  g1390
  (
    n1595,
    n618,
    n483
  );


  xnor
  g1391
  (
    n1801,
    n308,
    n349
  );


  and
  g1392
  (
    n1453,
    n301,
    n527
  );


  nand
  g1393
  (
    n1346,
    n373,
    n159
  );


  and
  g1394
  (
    n1492,
    n547,
    n398
  );


  xnor
  g1395
  (
    n941,
    n352,
    n251
  );


  or
  g1396
  (
    n815,
    n292,
    n459
  );


  nor
  g1397
  (
    n1886,
    n177,
    n220
  );


  xor
  g1398
  (
    n1766,
    n214,
    n628
  );


  xor
  g1399
  (
    n1698,
    n369,
    n395
  );


  xor
  g1400
  (
    n962,
    n649,
    n298
  );


  xor
  g1401
  (
    n1495,
    n306,
    n466
  );


  xnor
  g1402
  (
    n881,
    n454,
    n205
  );


  nor
  g1403
  (
    n1179,
    n487,
    n425
  );


  xnor
  g1404
  (
    n1582,
    n225,
    n305
  );


  or
  g1405
  (
    n734,
    n496,
    n612
  );


  and
  g1406
  (
    n1653,
    n591,
    n429
  );


  nand
  g1407
  (
    n1777,
    n567,
    n345
  );


  xnor
  g1408
  (
    n1870,
    n222,
    n508
  );


  and
  g1409
  (
    n1908,
    n565,
    n161
  );


  and
  g1410
  (
    n1695,
    n358,
    n250
  );


  nor
  g1411
  (
    n1287,
    n269,
    n619
  );


  xor
  g1412
  (
    n1660,
    n510,
    n457
  );


  and
  g1413
  (
    n1975,
    n328,
    n294
  );


  xnor
  g1414
  (
    n1418,
    n381,
    n228
  );


  or
  g1415
  (
    n992,
    n287,
    n206
  );


  xnor
  g1416
  (
    n784,
    n620,
    n166
  );


  nand
  g1417
  (
    n1609,
    n361,
    n319
  );


  xor
  g1418
  (
    n1382,
    n285,
    n248
  );


  nor
  g1419
  (
    n1800,
    n302,
    n547
  );


  nor
  g1420
  (
    n1747,
    n457,
    n547
  );


  or
  g1421
  (
    n923,
    n197,
    n157
  );


  xor
  g1422
  (
    n1363,
    n412,
    n267
  );


  xnor
  g1423
  (
    n1692,
    n552,
    n421
  );


  xnor
  g1424
  (
    n1504,
    n447,
    n527
  );


  xnor
  g1425
  (
    n906,
    n591,
    n328
  );


  or
  g1426
  (
    n1861,
    n228,
    n301
  );


  nor
  g1427
  (
    n1767,
    n299,
    n479
  );


  nor
  g1428
  (
    n1101,
    n196,
    n602
  );


  xor
  g1429
  (
    n1503,
    n560,
    n335
  );


  xnor
  g1430
  (
    n748,
    n211,
    n230
  );


  and
  g1431
  (
    n1224,
    n326,
    n383
  );


  nand
  g1432
  (
    n1236,
    n295,
    n535
  );


  xnor
  g1433
  (
    n825,
    n355,
    n443
  );


  xnor
  g1434
  (
    n1535,
    n312,
    n468
  );


  nor
  g1435
  (
    n879,
    n384,
    n469
  );


  nor
  g1436
  (
    n729,
    n531,
    n635
  );


  xor
  g1437
  (
    n1912,
    n503,
    n592
  );


  nand
  g1438
  (
    n1268,
    n555,
    n532
  );


  xor
  g1439
  (
    n1460,
    n313,
    n523
  );


  xnor
  g1440
  (
    n1853,
    n326,
    n418
  );


  and
  g1441
  (
    n1909,
    n416,
    n405
  );


  or
  g1442
  (
    n1377,
    n229,
    n649
  );


  and
  g1443
  (
    n944,
    n505,
    n555
  );


  xor
  g1444
  (
    n1253,
    n565,
    n419
  );


  xnor
  g1445
  (
    n965,
    n511,
    n206
  );


  nand
  g1446
  (
    n1136,
    n182,
    n388
  );


  nor
  g1447
  (
    n1083,
    n348,
    n642
  );


  nor
  g1448
  (
    n693,
    n276,
    n333
  );


  or
  g1449
  (
    n755,
    n626,
    n580
  );


  and
  g1450
  (
    n1773,
    n646,
    n580
  );


  xor
  g1451
  (
    KeyWire_0_28,
    n184,
    n183
  );


  xor
  g1452
  (
    n1494,
    n173,
    n245
  );


  and
  g1453
  (
    n1333,
    n436,
    n304
  );


  xor
  g1454
  (
    n1782,
    n476,
    n279
  );


  and
  g1455
  (
    n1044,
    n168,
    n385
  );


  or
  g1456
  (
    n1536,
    n294,
    n459
  );


  and
  g1457
  (
    n1920,
    n494,
    n252
  );


  xnor
  g1458
  (
    n1195,
    n584,
    n608
  );


  xor
  g1459
  (
    n951,
    n202,
    n333
  );


  xor
  g1460
  (
    n684,
    n539,
    n519
  );


  xnor
  g1461
  (
    n1029,
    n305,
    n623
  );


  nor
  g1462
  (
    n823,
    n541,
    n199
  );


  nor
  g1463
  (
    n1165,
    n182,
    n650
  );


  xor
  g1464
  (
    n1522,
    n583,
    n620
  );


  nand
  g1465
  (
    n1257,
    n205,
    n197
  );


  xor
  g1466
  (
    n1211,
    n185,
    n518
  );


  xor
  g1467
  (
    n1787,
    n174,
    n240
  );


  and
  g1468
  (
    n794,
    n460,
    n401
  );


  nor
  g1469
  (
    n1521,
    n441,
    n478
  );


  nand
  g1470
  (
    n754,
    n622,
    n426
  );


  nor
  g1471
  (
    n658,
    n446,
    n350
  );


  or
  g1472
  (
    n1115,
    n541,
    n574
  );


  nand
  g1473
  (
    n1758,
    n579,
    n405
  );


  nand
  g1474
  (
    n1434,
    n360,
    n486
  );


  and
  g1475
  (
    n958,
    n645,
    n407
  );


  xnor
  g1476
  (
    n1193,
    n198,
    n446
  );


  nor
  g1477
  (
    n1231,
    n201,
    n352
  );


  and
  g1478
  (
    n1092,
    n202,
    n261
  );


  xor
  g1479
  (
    n1158,
    n306,
    n322
  );


  xnor
  g1480
  (
    n1961,
    n262,
    n322
  );


  xor
  g1481
  (
    n1489,
    n601,
    n345
  );


  or
  g1482
  (
    n1340,
    n650,
    n614
  );


  or
  g1483
  (
    n1965,
    n387,
    n632
  );


  xnor
  g1484
  (
    n789,
    n239,
    n309
  );


  xnor
  g1485
  (
    n1872,
    n593,
    n386
  );


  and
  g1486
  (
    n864,
    n326,
    n433
  );


  or
  g1487
  (
    n1035,
    n592,
    n562
  );


  xnor
  g1488
  (
    n910,
    n540,
    n380
  );


  nand
  g1489
  (
    n1385,
    n642,
    n256
  );


  or
  g1490
  (
    n1152,
    n279,
    n465
  );


  or
  g1491
  (
    n1700,
    n588,
    n505
  );


  nor
  g1492
  (
    n1638,
    n597,
    n161
  );


  xnor
  g1493
  (
    n795,
    n181,
    n464
  );


  or
  g1494
  (
    n1615,
    n162,
    n531
  );


  and
  g1495
  (
    n1919,
    n207,
    n588
  );


  nand
  g1496
  (
    n1039,
    n456,
    n371
  );


  and
  g1497
  (
    n1642,
    n370,
    n553
  );


  or
  g1498
  (
    n1574,
    n258,
    n239
  );


  or
  g1499
  (
    n1052,
    n471,
    n235
  );


  nand
  g1500
  (
    n1745,
    n365,
    n405
  );


  nor
  g1501
  (
    n742,
    n643,
    n615
  );


  xor
  g1502
  (
    n1945,
    n343,
    n597
  );


  nor
  g1503
  (
    n694,
    n462,
    n301
  );


  xnor
  g1504
  (
    n1468,
    n299,
    n382
  );


  and
  g1505
  (
    n1607,
    n204,
    n602
  );


  or
  g1506
  (
    n943,
    n453,
    n421
  );


  and
  g1507
  (
    n1828,
    n498,
    n595
  );


  or
  g1508
  (
    n1220,
    n232,
    n442
  );


  nor
  g1509
  (
    n1439,
    n590,
    n339
  );


  or
  g1510
  (
    KeyWire_0_14,
    n372,
    n274
  );


  xor
  g1511
  (
    n1068,
    n374,
    n259
  );


  nor
  g1512
  (
    n1881,
    n590,
    n544
  );


  xor
  g1513
  (
    n836,
    n424,
    n373
  );


  nor
  g1514
  (
    n1071,
    n190,
    n440
  );


  xor
  g1515
  (
    n1892,
    n563,
    n314
  );


  xnor
  g1516
  (
    n1866,
    n327,
    n590
  );


  xnor
  g1517
  (
    n1865,
    n248,
    n375
  );


  nor
  g1518
  (
    n1737,
    n172,
    n543
  );


  nor
  g1519
  (
    n1085,
    n386,
    n210
  );


  nand
  g1520
  (
    n1953,
    n244,
    n406
  );


  xor
  g1521
  (
    n1718,
    n238,
    n235
  );


  xor
  g1522
  (
    n1368,
    n617,
    n213
  );


  xnor
  g1523
  (
    n1628,
    n549,
    n233
  );


  xnor
  g1524
  (
    n1931,
    n418,
    n260
  );


  nor
  g1525
  (
    n839,
    n533,
    n195
  );


  nand
  g1526
  (
    n1244,
    n613,
    n364
  );


  xnor
  g1527
  (
    n1523,
    n534,
    n344
  );


  xnor
  g1528
  (
    n1575,
    n383,
    n499
  );


  nand
  g1529
  (
    n782,
    n229,
    n353
  );


  or
  g1530
  (
    n680,
    n598,
    n198
  );


  or
  g1531
  (
    n1650,
    n498,
    n572
  );


  xor
  g1532
  (
    n1661,
    n410,
    n502
  );


  nor
  g1533
  (
    n1803,
    n360,
    n168
  );


  xnor
  g1534
  (
    n1496,
    n526,
    n391
  );


  and
  g1535
  (
    n1940,
    n535,
    n414
  );


  xor
  g1536
  (
    n1180,
    n539,
    n475
  );


  nand
  g1537
  (
    KeyWire_0_51,
    n349,
    n646
  );


  nor
  g1538
  (
    n1640,
    n498,
    n572
  );


  and
  g1539
  (
    n1075,
    n228,
    n427
  );


  or
  g1540
  (
    n1693,
    n372,
    n198
  );


  nor
  g1541
  (
    n654,
    n621,
    n363
  );


  nand
  g1542
  (
    n811,
    n463,
    n521
  );


  xor
  g1543
  (
    n1943,
    n247,
    n280
  );


  and
  g1544
  (
    KeyWire_0_41,
    n410,
    n613
  );


  xnor
  g1545
  (
    n661,
    n586,
    n232
  );


  or
  g1546
  (
    n677,
    n591,
    n202
  );


  and
  g1547
  (
    n895,
    n636,
    n593
  );


  nor
  g1548
  (
    n1014,
    n451,
    n529
  );


  and
  g1549
  (
    n1637,
    n196,
    n508
  );


  xor
  g1550
  (
    n1086,
    n340,
    n268
  );


  nor
  g1551
  (
    n862,
    n174,
    n170
  );


  nor
  g1552
  (
    n1962,
    n500,
    n579
  );


  xor
  g1553
  (
    n1760,
    n188,
    n332
  );


  xnor
  g1554
  (
    n1733,
    n650,
    n407
  );


  or
  g1555
  (
    n883,
    n346,
    n358
  );


  xnor
  g1556
  (
    n1532,
    n548,
    n165
  );


  nor
  g1557
  (
    n1713,
    n516,
    n622
  );


  xor
  g1558
  (
    n946,
    n595,
    n373
  );


  nand
  g1559
  (
    n956,
    n272,
    n585
  );


  nand
  g1560
  (
    n1369,
    n376,
    n428
  );


  or
  g1561
  (
    n981,
    n390,
    n278
  );


  nor
  g1562
  (
    n1006,
    n252,
    n525
  );


  nand
  g1563
  (
    n1804,
    n171,
    n208
  );


  nand
  g1564
  (
    n1429,
    n203,
    n206
  );


  and
  g1565
  (
    n1270,
    n525,
    n266
  );


  nor
  g1566
  (
    n1950,
    n195,
    n263
  );


  nor
  g1567
  (
    n1104,
    n196,
    n478
  );


  nand
  g1568
  (
    n1297,
    n384,
    n644
  );


  xnor
  g1569
  (
    n1442,
    n489,
    n334
  );


  and
  g1570
  (
    n1515,
    n196,
    n449
  );


  and
  g1571
  (
    n1648,
    n645,
    n284
  );


  nand
  g1572
  (
    n848,
    n290,
    n351
  );


  and
  g1573
  (
    n1311,
    n336,
    n598
  );


  or
  g1574
  (
    KeyWire_0_17,
    n627,
    n501
  );


  nand
  g1575
  (
    n882,
    n412,
    n397
  );


  and
  g1576
  (
    n1902,
    n573,
    n253
  );


  and
  g1577
  (
    n831,
    n460,
    n157
  );


  xor
  g1578
  (
    n952,
    n511,
    n454
  );


  xnor
  g1579
  (
    n1670,
    n406,
    n575
  );


  and
  g1580
  (
    n690,
    n366,
    n448
  );


  xnor
  g1581
  (
    n1512,
    n176,
    n227
  );


  and
  g1582
  (
    n1339,
    n222,
    n452
  );


  or
  g1583
  (
    n1467,
    n171,
    n180
  );


  xnor
  g1584
  (
    n659,
    n378,
    n290
  );


  xor
  g1585
  (
    n1076,
    n581,
    n634
  );


  nor
  g1586
  (
    n1635,
    n210,
    n412
  );


  and
  g1587
  (
    n1746,
    n329,
    n437
  );


  xor
  g1588
  (
    n908,
    n586,
    n461
  );


  xnor
  g1589
  (
    n1923,
    n327,
    n471
  );


  or
  g1590
  (
    n822,
    n208,
    n492
  );


  nand
  g1591
  (
    n1864,
    n592,
    n256
  );


  and
  g1592
  (
    n1197,
    n312,
    n583
  );


  nand
  g1593
  (
    n1590,
    n397,
    n555
  );


  nand
  g1594
  (
    n1658,
    n449,
    n458
  );


  xor
  g1595
  (
    n991,
    n601,
    n458
  );


  nor
  g1596
  (
    n706,
    n269,
    n469
  );


  or
  g1597
  (
    n1871,
    n604,
    n371
  );


  nor
  g1598
  (
    n731,
    n423,
    n535
  );


  xor
  g1599
  (
    n1415,
    n242,
    n420
  );


  xor
  g1600
  (
    n735,
    n505,
    n188
  );


  xor
  g1601
  (
    n1704,
    n472,
    n362
  );


  nor
  g1602
  (
    n1708,
    n596,
    n445
  );


  xnor
  g1603
  (
    n1738,
    n558,
    n431
  );


  or
  g1604
  (
    n1547,
    n488,
    n299
  );


  or
  g1605
  (
    n1514,
    n163,
    n607
  );


  nor
  g1606
  (
    n1788,
    n501,
    n492
  );


  nor
  g1607
  (
    n1649,
    n281,
    n287
  );


  xor
  g1608
  (
    n1517,
    n591,
    n225
  );


  xnor
  g1609
  (
    n1705,
    n542,
    n595
  );


  nor
  g1610
  (
    n1571,
    n221,
    n639
  );


  and
  g1611
  (
    n982,
    n481,
    n641
  );


  xnor
  g1612
  (
    n1281,
    n423,
    n437
  );


  xor
  g1613
  (
    n1384,
    n435,
    n360
  );


  and
  g1614
  (
    n1329,
    n234,
    n180
  );


  and
  g1615
  (
    n1387,
    n400,
    n597
  );


  nor
  g1616
  (
    n672,
    n420,
    n435
  );


  nor
  g1617
  (
    n1808,
    n483,
    n257
  );


  xnor
  g1618
  (
    n1550,
    n419,
    n333
  );


  xnor
  g1619
  (
    n1150,
    n514,
    n574
  );


  nor
  g1620
  (
    n1407,
    n181,
    n315
  );


  nand
  g1621
  (
    n840,
    n650,
    n567
  );


  nand
  g1622
  (
    n1959,
    n559,
    n472
  );


  xor
  g1623
  (
    n1232,
    n621,
    n550
  );


  nand
  g1624
  (
    n931,
    n530,
    n637
  );


  and
  g1625
  (
    n900,
    n537,
    n492
  );


  and
  g1626
  (
    n1292,
    n570,
    n363
  );


  and
  g1627
  (
    n1392,
    n550,
    n481
  );


  and
  g1628
  (
    n664,
    n438,
    n384
  );


  xnor
  g1629
  (
    n1401,
    n521,
    n606
  );


  or
  g1630
  (
    n1599,
    n529,
    n476
  );


  nor
  g1631
  (
    n1605,
    n243,
    n223
  );


  xor
  g1632
  (
    n897,
    n265,
    n362
  );


  and
  g1633
  (
    n1073,
    n381,
    n556
  );


  xor
  g1634
  (
    n947,
    n203,
    n398
  );


  nand
  g1635
  (
    n1323,
    n374,
    n647
  );


  xor
  g1636
  (
    n1450,
    n607,
    n499
  );


  xnor
  g1637
  (
    n1603,
    n405,
    n402
  );


  and
  g1638
  (
    n1778,
    n457,
    n594
  );


  xor
  g1639
  (
    n1474,
    n178,
    n511
  );


  nor
  g1640
  (
    n1265,
    n558,
    n281
  );


  or
  g1641
  (
    n1279,
    n266,
    n408
  );


  or
  g1642
  (
    n1944,
    n359,
    n433
  );


  xnor
  g1643
  (
    KeyWire_0_31,
    n475,
    n599
  );


  xor
  g1644
  (
    n1811,
    n534,
    n333
  );


  xor
  g1645
  (
    n924,
    n345,
    n506
  );


  nor
  g1646
  (
    n1202,
    n321,
    n309
  );


  and
  g1647
  (
    n1880,
    n504,
    n559
  );


  xor
  g1648
  (
    n1620,
    n588,
    n204
  );


  nor
  g1649
  (
    n1254,
    n260,
    n435
  );


  and
  g1650
  (
    n1108,
    n413,
    n509
  );


  xor
  g1651
  (
    n1351,
    n647,
    n404
  );


  or
  g1652
  (
    n1719,
    n240,
    n370
  );


  and
  g1653
  (
    n1978,
    n630,
    n632
  );


  or
  g1654
  (
    n681,
    n524,
    n568
  );


  xnor
  g1655
  (
    n1835,
    n570,
    n275
  );


  xnor
  g1656
  (
    n1282,
    n420,
    n327
  );


  and
  g1657
  (
    n756,
    n543,
    n444
  );


  nand
  g1658
  (
    n759,
    n261,
    n554
  );


  xnor
  g1659
  (
    n851,
    n466,
    n307
  );


  xor
  g1660
  (
    n1925,
    n495,
    n311
  );


  and
  g1661
  (
    n1712,
    n309,
    n343
  );


  and
  g1662
  (
    n963,
    n368,
    n554
  );


  xnor
  g1663
  (
    n1576,
    n427,
    n450
  );


  nor
  g1664
  (
    n1121,
    n607,
    n363
  );


  or
  g1665
  (
    n1347,
    n581,
    n272
  );


  nand
  g1666
  (
    KeyWire_0_6,
    n332,
    n179
  );


  nand
  g1667
  (
    n1245,
    n235,
    n537
  );


  xor
  g1668
  (
    n1960,
    n537,
    n201
  );


  xor
  g1669
  (
    n984,
    n484,
    n618
  );


  nor
  g1670
  (
    n1761,
    n255,
    n440
  );


  and
  g1671
  (
    n1365,
    n415,
    n425
  );


  xor
  g1672
  (
    n1528,
    n209,
    n579
  );


  and
  g1673
  (
    n1927,
    n637,
    n627
  );


  xnor
  g1674
  (
    n1821,
    n166,
    n243
  );


  xnor
  g1675
  (
    n1138,
    n598,
    n246
  );


  or
  g1676
  (
    n1816,
    n614,
    n504
  );


  xnor
  g1677
  (
    n1171,
    n226,
    n460
  );


  nand
  g1678
  (
    n1051,
    n539,
    n354
  );


  and
  g1679
  (
    n1485,
    n487,
    n177
  );


  xnor
  g1680
  (
    n1657,
    n466,
    n188
  );


  nand
  g1681
  (
    n1153,
    n332,
    n262
  );


  xnor
  g1682
  (
    n747,
    n254,
    n273
  );


  and
  g1683
  (
    n1009,
    n193,
    n287
  );


  xnor
  g1684
  (
    n1371,
    n289,
    n403
  );


  or
  g1685
  (
    n1906,
    n431,
    n621
  );


  xor
  g1686
  (
    n1762,
    n633,
    n329
  );


  and
  g1687
  (
    n1183,
    n204,
    n328
  );


  xnor
  g1688
  (
    n656,
    n234,
    n158
  );


  xnor
  g1689
  (
    n1406,
    n251,
    n519
  );


  xor
  g1690
  (
    n1145,
    n341,
    n576
  );


  and
  g1691
  (
    n1519,
    n456,
    n519
  );


  or
  g1692
  (
    n1636,
    n607,
    n366
  );


  nand
  g1693
  (
    n1623,
    n229,
    n239
  );


  xnor
  g1694
  (
    n1423,
    n533,
    n446
  );


  xnor
  g1695
  (
    n1380,
    n585,
    n352
  );


  xnor
  g1696
  (
    n1887,
    n233,
    n346
  );


  nor
  g1697
  (
    n974,
    n392,
    n344
  );


  xnor
  g1698
  (
    n859,
    n258,
    n430
  );


  nor
  g1699
  (
    n1214,
    n218,
    n548
  );


  or
  g1700
  (
    n1398,
    n209,
    n451
  );


  or
  g1701
  (
    n916,
    n605,
    n212
  );


  nor
  g1702
  (
    n1107,
    n355,
    n586
  );


  xnor
  g1703
  (
    n1443,
    n580,
    n528
  );


  nor
  g1704
  (
    n802,
    n639,
    n224
  );


  or
  g1705
  (
    n662,
    n525,
    n490
  );


  nor
  g1706
  (
    n1470,
    n275,
    n380
  );


  nand
  g1707
  (
    n1885,
    n551,
    n448
  );


  or
  g1708
  (
    n739,
    n190,
    n603
  );


  nand
  g1709
  (
    n1069,
    n613,
    n493
  );


  xnor
  g1710
  (
    n1629,
    n603,
    n325
  );


  nor
  g1711
  (
    n996,
    n544,
    n176
  );


  or
  g1712
  (
    n1084,
    n169,
    n186
  );


  xnor
  g1713
  (
    n1617,
    n251,
    n556
  );


  nor
  g1714
  (
    n1455,
    n474,
    n176
  );


  nor
  g1715
  (
    n1666,
    n402,
    n296
  );


  xor
  g1716
  (
    n960,
    n460,
    n191
  );


  and
  g1717
  (
    n1884,
    n285,
    n368
  );


  nand
  g1718
  (
    n1054,
    n197,
    n244
  );


  xor
  g1719
  (
    n1786,
    n585,
    n520
  );


  and
  g1720
  (
    n679,
    n629,
    n578
  );


  nand
  g1721
  (
    n1691,
    n589,
    n158
  );


  nor
  g1722
  (
    n856,
    n416,
    n236
  );


  nand
  g1723
  (
    n1662,
    n574,
    n414
  );


  and
  g1724
  (
    n745,
    n162,
    n385
  );


  nand
  g1725
  (
    n1422,
    n612,
    n399
  );


  or
  g1726
  (
    n1304,
    n494,
    n209
  );


  and
  g1727
  (
    n1216,
    n390,
    n317
  );


  xnor
  g1728
  (
    n1167,
    n562,
    n504
  );


  or
  g1729
  (
    n1250,
    n542,
    n564
  );


  nand
  g1730
  (
    n1538,
    n571,
    n166
  );


  xor
  g1731
  (
    n986,
    n288,
    n387
  );


  xor
  g1732
  (
    n911,
    n538,
    n160
  );


  and
  g1733
  (
    n1779,
    n179,
    n362
  );


  xnor
  g1734
  (
    n1471,
    n347,
    n611
  );


  and
  g1735
  (
    n1248,
    n172,
    n614
  );


  xnor
  g1736
  (
    n849,
    n366,
    n278
  );


  xor
  g1737
  (
    n1018,
    n257,
    n546
  );


  nand
  g1738
  (
    n1634,
    n627,
    n367
  );


  xnor
  g1739
  (
    n711,
    n267,
    n414
  );


  and
  g1740
  (
    n786,
    n528,
    n629
  );


  nand
  g1741
  (
    n1321,
    n290,
    n611
  );


  nand
  g1742
  (
    n790,
    n259,
    n222
  );


  and
  g1743
  (
    n771,
    n396,
    n164
  );


  nor
  g1744
  (
    n1972,
    n401,
    n630
  );


  nor
  g1745
  (
    n964,
    n421,
    n329
  );


  xnor
  g1746
  (
    n915,
    n418,
    n324
  );


  nand
  g1747
  (
    n1079,
    n463,
    n199
  );


  xnor
  g1748
  (
    n1099,
    n255,
    n473
  );


  nand
  g1749
  (
    n1907,
    n549,
    n246
  );


  nand
  g1750
  (
    n1727,
    n361,
    n558
  );


  or
  g1751
  (
    n1869,
    n171,
    n217
  );


  or
  g1752
  (
    n692,
    n337,
    n490
  );


  xor
  g1753
  (
    n1447,
    n205,
    n355
  );


  nand
  g1754
  (
    n768,
    n477,
    n577
  );


  nand
  g1755
  (
    n1789,
    n583,
    n406
  );


  xnor
  g1756
  (
    n1081,
    n173,
    n444
  );


  and
  g1757
  (
    n1969,
    n620,
    n482
  );


  and
  g1758
  (
    n1140,
    n447,
    n214
  );


  or
  g1759
  (
    n1330,
    n399,
    n468
  );


  or
  g1760
  (
    n846,
    n514,
    n429
  );


  or
  g1761
  (
    n1488,
    n319,
    n451
  );


  xnor
  g1762
  (
    n979,
    n365,
    n282
  );


  xnor
  g1763
  (
    n710,
    n625,
    n473
  );


  xnor
  g1764
  (
    n1941,
    n344,
    n174
  );


  nand
  g1765
  (
    n1098,
    n608,
    n236
  );


  xnor
  g1766
  (
    n966,
    n291,
    n384
  );


  nor
  g1767
  (
    n1676,
    n215,
    n387
  );


  nand
  g1768
  (
    n1144,
    n314,
    n353
  );


  and
  g1769
  (
    n1541,
    n573,
    n570
  );


  nand
  g1770
  (
    n671,
    n510,
    n616
  );


  and
  g1771
  (
    n1553,
    n615,
    n636
  );


  nand
  g1772
  (
    n1552,
    n599,
    n574
  );


  xor
  g1773
  (
    n857,
    n265,
    n264
  );


  xor
  g1774
  (
    n1841,
    n543,
    n497
  );


  or
  g1775
  (
    n1954,
    n357,
    n256
  );


  xor
  g1776
  (
    n1379,
    n416,
    n227
  );


  or
  g1777
  (
    n723,
    n296,
    n348
  );


  xor
  g1778
  (
    n1364,
    n308,
    n611
  );


  xor
  g1779
  (
    n1584,
    n636,
    n340
  );


  nor
  g1780
  (
    n1524,
    n474,
    n168
  );


  nand
  g1781
  (
    n1376,
    n318,
    n365
  );


  or
  g1782
  (
    KeyWire_0_0,
    n200,
    n183
  );


  xnor
  g1783
  (
    n1070,
    n602,
    n313
  );


  and
  g1784
  (
    n1529,
    n330,
    n512
  );


  and
  g1785
  (
    n762,
    n299,
    n619
  );


  and
  g1786
  (
    n1077,
    n337,
    n539
  );


  or
  g1787
  (
    n852,
    n587,
    n527
  );


  xnor
  g1788
  (
    n1182,
    n618,
    n342
  );


  and
  g1789
  (
    n890,
    n225,
    n453
  );


  nor
  g1790
  (
    n1836,
    n394,
    n324
  );


  xnor
  g1791
  (
    n1360,
    n228,
    n411
  );


  xor
  g1792
  (
    n1563,
    n464,
    n525
  );


  or
  g1793
  (
    n1396,
    n545,
    n266
  );


  nor
  g1794
  (
    n807,
    n319,
    n631
  );


  or
  g1795
  (
    n1567,
    n490,
    n167
  );


  nor
  g1796
  (
    n1964,
    n336,
    n440
  );


  xor
  g1797
  (
    n1769,
    n471,
    n534
  );


  and
  g1798
  (
    n1859,
    n433,
    n566
  );


  nor
  g1799
  (
    n972,
    n250,
    n393
  );


  xnor
  g1800
  (
    n1170,
    n562,
    n337
  );


  xnor
  g1801
  (
    n1770,
    n626,
    n382
  );


  nand
  g1802
  (
    n730,
    n513,
    n189
  );


  xor
  g1803
  (
    n1977,
    n600,
    n502
  );


  and
  g1804
  (
    n1428,
    n611,
    n623
  );


  and
  g1805
  (
    n1955,
    n241,
    n582
  );


  xnor
  g1806
  (
    n829,
    n480,
    n599
  );


  nor
  g1807
  (
    n824,
    n522,
    n452
  );


  nor
  g1808
  (
    n816,
    n390,
    n208
  );


  xnor
  g1809
  (
    n769,
    n186,
    n623
  );


  or
  g1810
  (
    n1863,
    n620,
    n247
  );


  nand
  g1811
  (
    n1971,
    n415,
    n609
  );


  and
  g1812
  (
    n1667,
    n162,
    n203
  );


  nor
  g1813
  (
    n1062,
    n646,
    n413
  );


  nand
  g1814
  (
    n1968,
    n199,
    n268
  );


  nor
  g1815
  (
    n1089,
    n199,
    n630
  );


  xnor
  g1816
  (
    n1057,
    n594,
    n589
  );


  nor
  g1817
  (
    n959,
    n647,
    n469
  );


  or
  g1818
  (
    n1391,
    n569,
    n293
  );


  xor
  g1819
  (
    KeyWire_0_13,
    n357,
    n458
  );


  or
  g1820
  (
    n1239,
    n509,
    n520
  );


  or
  g1821
  (
    n1674,
    n457,
    n284
  );


  xor
  g1822
  (
    n1383,
    n364,
    n324
  );


  xor
  g1823
  (
    n1544,
    n338,
    n241
  );


  nand
  g1824
  (
    n1269,
    n324,
    n358
  );


  and
  g1825
  (
    n1472,
    n334,
    n517
  );


  xor
  g1826
  (
    n1554,
    n193,
    n592
  );


  xnor
  g1827
  (
    n1264,
    n296,
    n387
  );


  nand
  g1828
  (
    n1505,
    n376,
    n382
  );


  nor
  g1829
  (
    n845,
    n625,
    n359
  );


  nand
  g1830
  (
    n1283,
    n518,
    n187
  );


  xor
  g1831
  (
    n1217,
    n641,
    n598
  );


  nor
  g1832
  (
    n1739,
    n346,
    n474
  );


  and
  g1833
  (
    n878,
    n596,
    n161
  );


  or
  g1834
  (
    n1386,
    n605,
    n254
  );


  xnor
  g1835
  (
    n1055,
    n280,
    n396
  );


  xnor
  g1836
  (
    n1913,
    n160,
    n609
  );


  or
  g1837
  (
    n1720,
    n222,
    n523
  );


  or
  g1838
  (
    n1763,
    n491,
    n178
  );


  xor
  g1839
  (
    n1561,
    n638,
    n305
  );


  nor
  g1840
  (
    n1967,
    n581,
    n422
  );


  nor
  g1841
  (
    KeyWire_0_40,
    n200,
    n223
  );


  xnor
  g1842
  (
    n752,
    n385,
    n437
  );


  nor
  g1843
  (
    n1701,
    n158,
    n557
  );


  xor
  g1844
  (
    n1805,
    n339,
    n426
  );


  xor
  g1845
  (
    n809,
    n160,
    n180
  );


  and
  g1846
  (
    n1229,
    n515,
    n221
  );


  and
  g1847
  (
    n766,
    n187,
    n411
  );


  or
  g1848
  (
    n1381,
    n625,
    n168
  );


  nand
  g1849
  (
    n835,
    n378,
    n608
  );


  nor
  g1850
  (
    n1463,
    n622,
    n226
  );


  xor
  g1851
  (
    n1124,
    n454,
    n377
  );


  nand
  g1852
  (
    n1301,
    n431,
    n183
  );


  nand
  g1853
  (
    n917,
    n356,
    n483
  );


  and
  g1854
  (
    n1358,
    n651,
    n467
  );


  and
  g1855
  (
    n1633,
    n297,
    n226
  );


  and
  g1856
  (
    n1397,
    n173,
    n609
  );


  xnor
  g1857
  (
    n1724,
    n233,
    n641
  );


  xnor
  g1858
  (
    n860,
    n368,
    n401
  );


  nand
  g1859
  (
    n1306,
    n357,
    n212
  );


  xnor
  g1860
  (
    n697,
    n578,
    n178
  );


  nor
  g1861
  (
    n930,
    n248,
    n187
  );


  xor
  g1862
  (
    n1117,
    n552,
    n219
  );


  xnor
  g1863
  (
    n841,
    n563,
    n291
  );


  or
  g1864
  (
    n1481,
    n200,
    n195
  );


  nor
  g1865
  (
    n1647,
    n277,
    n578
  );


  nand
  g1866
  (
    n1334,
    n316,
    n495
  );


  xor
  g1867
  (
    n800,
    n181,
    n263
  );


  xor
  g1868
  (
    n1427,
    n493,
    n270
  );


  or
  g1869
  (
    n1929,
    n238,
    n594
  );


  nor
  g1870
  (
    n1684,
    n543,
    n310
  );


  xnor
  g1871
  (
    n1237,
    n258,
    n317
  );


  nor
  g1872
  (
    n1011,
    n497,
    n338
  );


  and
  g1873
  (
    n870,
    n238,
    n293
  );


  xnor
  g1874
  (
    n1203,
    n479,
    n276
  );


  and
  g1875
  (
    n999,
    n510,
    n540
  );


  xor
  g1876
  (
    n1410,
    n425,
    n260
  );


  xor
  g1877
  (
    n832,
    n473,
    n399
  );


  xor
  g1878
  (
    n1918,
    n556,
    n213
  );


  nor
  g1879
  (
    n788,
    n262,
    n322
  );


  xnor
  g1880
  (
    n1466,
    n445,
    n432
  );


  xor
  g1881
  (
    n1091,
    n202,
    n577
  );


  or
  g1882
  (
    n1507,
    n331,
    n305
  );


  xor
  g1883
  (
    n812,
    n271,
    n549
  );


  xor
  g1884
  (
    n1916,
    n291,
    n189
  );


  xor
  g1885
  (
    n1551,
    n201,
    n560
  );


  nor
  g1886
  (
    n935,
    n392,
    n587
  );


  xor
  g1887
  (
    n1007,
    n216,
    n271
  );


  nand
  g1888
  (
    KeyWire_0_11,
    n432,
    n396
  );


  nor
  g1889
  (
    n1271,
    n300,
    n227
  );


  nand
  g1890
  (
    n1303,
    n514,
    n601
  );


  xor
  g1891
  (
    n1555,
    n414,
    n221
  );


  and
  g1892
  (
    n1411,
    n300,
    n552
  );


  xnor
  g1893
  (
    n737,
    n584,
    n532
  );


  or
  g1894
  (
    n1956,
    n274,
    n320
  );


  and
  g1895
  (
    n797,
    n238,
    n556
  );


  xnor
  g1896
  (
    n714,
    n489,
    n527
  );


  nor
  g1897
  (
    n1890,
    n371,
    n438
  );


  and
  g1898
  (
    n1319,
    n485,
    n643
  );


  nand
  g1899
  (
    n1557,
    n395,
    n224
  );


  xor
  g1900
  (
    n1048,
    n569,
    n220
  );


  or
  g1901
  (
    n1480,
    n191,
    n597
  );


  xor
  g1902
  (
    n1596,
    n462,
    n319
  );


  nor
  g1903
  (
    n1310,
    n232,
    n217
  );


  nor
  g1904
  (
    n1177,
    n493,
    n576
  );


  and
  g1905
  (
    n1166,
    n616,
    n252
  );


  and
  g1906
  (
    n1833,
    n623,
    n302
  );


  and
  g1907
  (
    n997,
    n352,
    n158
  );


  or
  g1908
  (
    n799,
    n548,
    n535
  );


  nand
  g1909
  (
    n774,
    n330,
    n600
  );


  or
  g1910
  (
    n980,
    n422,
    n437
  );


  xnor
  g1911
  (
    n1734,
    n302,
    n439
  );


  xor
  g1912
  (
    n698,
    n312,
    n617
  );


  xor
  g1913
  (
    n1335,
    n495,
    n516
  );


  xnor
  g1914
  (
    n1172,
    n444,
    n530
  );


  nand
  g1915
  (
    n1325,
    n391,
    n302
  );


  xor
  g1916
  (
    n1374,
    n335,
    n272
  );


  and
  g1917
  (
    n1824,
    n234,
    n307
  );


  and
  g1918
  (
    n1111,
    n350,
    n180
  );


  xor
  g1919
  (
    n1280,
    n504,
    n506
  );


  nor
  g1920
  (
    n1791,
    n531,
    n280
  );


  xor
  g1921
  (
    n1819,
    n236,
    n472
  );


  and
  g1922
  (
    n1149,
    n215,
    n376
  );


  xor
  g1923
  (
    n715,
    n210,
    n221
  );


  xor
  g1924
  (
    n971,
    n517,
    n645
  );


  xnor
  g1925
  (
    n1128,
    n644,
    n341
  );


  and
  g1926
  (
    n1110,
    n477,
    n342
  );


  xor
  g1927
  (
    n1141,
    n323,
    n216
  );


  xnor
  g1928
  (
    n1120,
    n189,
    n340
  );


  xor
  g1929
  (
    n902,
    n638,
    n287
  );


  nand
  g1930
  (
    n1225,
    n409,
    n439
  );


  xor
  g1931
  (
    n820,
    n176,
    n281
  );


  and
  g1932
  (
    n914,
    n185,
    n394
  );


  or
  g1933
  (
    n903,
    n166,
    n165
  );


  or
  g1934
  (
    n1610,
    n446,
    n544
  );


  nor
  g1935
  (
    n1096,
    n278,
    n582
  );


  or
  g1936
  (
    n1933,
    n488,
    n642
  );


  nor
  g1937
  (
    n1295,
    n393,
    n375
  );


  or
  g1938
  (
    n1095,
    n355,
    n483
  );


  and
  g1939
  (
    KeyWire_0_32,
    n194,
    n276
  );


  nand
  g1940
  (
    n1262,
    n452,
    n341
  );


  nor
  g1941
  (
    n1147,
    n242,
    n548
  );


  and
  g1942
  (
    n1947,
    n361,
    n436
  );


  nor
  g1943
  (
    n1619,
    n246,
    n254
  );


  or
  g1944
  (
    n1822,
    n371,
    n427
  );


  nor
  g1945
  (
    n1105,
    n316,
    n466
  );


  xnor
  g1946
  (
    n1320,
    n331,
    n400
  );


  nand
  g1947
  (
    n787,
    n612,
    n317
  );


  xnor
  g1948
  (
    n2291,
    n824,
    n1908,
    n874,
    n929
  );


  xnor
  g1949
  (
    KeyWire_0_49,
    n1496,
    n1897,
    n1859,
    n1457
  );


  xnor
  g1950
  (
    n2203,
    n876,
    n1291,
    n1318,
    n749
  );


  and
  g1951
  (
    n2079,
    n935,
    n1180,
    n1049,
    n1161
  );


  and
  g1952
  (
    n2012,
    n1269,
    n1435,
    n1890,
    n1292
  );


  or
  g1953
  (
    n2286,
    n1284,
    n1405,
    n1498,
    n1114
  );


  nor
  g1954
  (
    n2107,
    n889,
    n1003,
    n1446,
    n1445
  );


  xnor
  g1955
  (
    n1981,
    n1896,
    n1295,
    n714,
    n1012
  );


  xor
  g1956
  (
    n2194,
    n1116,
    n716,
    n759,
    n1697
  );


  xor
  g1957
  (
    n2049,
    n1387,
    n1683,
    n1410,
    n1472
  );


  xor
  g1958
  (
    n2196,
    n1644,
    n1336,
    n989,
    n1507
  );


  xor
  g1959
  (
    n2016,
    n1040,
    n1574,
    n1538,
    n1863
  );


  nor
  g1960
  (
    n2026,
    n1335,
    n1488,
    n1137,
    n1170
  );


  and
  g1961
  (
    n2074,
    n1244,
    n1736,
    n1650,
    n1276
  );


  xnor
  g1962
  (
    n2086,
    n1717,
    n1395,
    n1018,
    n1674
  );


  nand
  g1963
  (
    n2309,
    n1767,
    n783,
    n915,
    n1786
  );


  nor
  g1964
  (
    n2181,
    n1890,
    n789,
    n822,
    n895
  );


  and
  g1965
  (
    n2158,
    n1164,
    n1583,
    n1397,
    n1352
  );


  xnor
  g1966
  (
    n2027,
    n1778,
    n1563,
    n1102,
    n1791
  );


  and
  g1967
  (
    n2224,
    n1601,
    n666,
    n1176,
    n1724
  );


  nand
  g1968
  (
    n2055,
    n1522,
    n1364,
    n1663,
    n1896
  );


  xnor
  g1969
  (
    n2285,
    n1132,
    n1867,
    n762,
    n1341
  );


  nand
  g1970
  (
    n2170,
    n1200,
    n1479,
    n1610,
    n1830
  );


  or
  g1971
  (
    n2228,
    n1258,
    n1688,
    n1464,
    n1484
  );


  xor
  g1972
  (
    n2099,
    n1667,
    n1032,
    n1356,
    n1486
  );


  and
  g1973
  (
    n2154,
    n1631,
    n966,
    n860,
    n1240
  );


  xor
  g1974
  (
    n2176,
    n1599,
    n1274,
    n1458,
    n1824
  );


  nand
  g1975
  (
    n2296,
    n774,
    n1831,
    n1721,
    n870
  );


  nor
  g1976
  (
    n2064,
    n1900,
    n1443,
    n1578,
    n829
  );


  nand
  g1977
  (
    n2255,
    n1768,
    n1803,
    n1394,
    n832
  );


  xnor
  g1978
  (
    n2248,
    n805,
    n1565,
    n1265,
    n843
  );


  nor
  g1979
  (
    n2301,
    n1266,
    n1875,
    n1454,
    n1409
  );


  or
  g1980
  (
    n2232,
    n1109,
    n1503,
    n1844,
    n1302
  );


  nor
  g1981
  (
    n2093,
    n892,
    n1866,
    n1766,
    n1852
  );


  nand
  g1982
  (
    KeyWire_0_60,
    n1230,
    n1060,
    n1306,
    n1902
  );


  and
  g1983
  (
    n2123,
    n1388,
    n907,
    n1178,
    n729
  );


  xnor
  g1984
  (
    n2008,
    n1080,
    n1905,
    n785,
    n1728
  );


  xor
  g1985
  (
    n2169,
    n1031,
    n1505,
    n1636,
    n1333
  );


  nand
  g1986
  (
    n2180,
    n1894,
    n700,
    n1797,
    n730
  );


  or
  g1987
  (
    n2076,
    n1437,
    n771,
    n695,
    n1901
  );


  or
  g1988
  (
    n2277,
    n1323,
    n1206,
    n751,
    n1466
  );


  xnor
  g1989
  (
    n2029,
    n1162,
    n1093,
    n727,
    n1615
  );


  nand
  g1990
  (
    n2097,
    n1903,
    n1662,
    n928,
    n825
  );


  xor
  g1991
  (
    n2126,
    n1304,
    n1757,
    n675,
    n1600
  );


  nand
  g1992
  (
    n2085,
    n1175,
    n1581,
    n692,
    n719
  );


  or
  g1993
  (
    n2177,
    n668,
    n1173,
    n1403,
    n992
  );


  and
  g1994
  (
    n2288,
    n1355,
    n879,
    n1770,
    n1525
  );


  and
  g1995
  (
    n2125,
    n1451,
    n859,
    n763,
    n1351
  );


  or
  g1996
  (
    n2144,
    n1900,
    n1120,
    n1847,
    n1892
  );


  xor
  g1997
  (
    n2254,
    n978,
    n1177,
    n1425,
    n669
  );


  and
  g1998
  (
    n2290,
    n953,
    n1277,
    n1231,
    n1671
  );


  nand
  g1999
  (
    n2304,
    n1582,
    n778,
    n972,
    n1798
  );


  xor
  g2000
  (
    n2303,
    n1876,
    n1755,
    n1490,
    n1400
  );


  or
  g2001
  (
    n2223,
    n1562,
    n1134,
    n1381,
    n821
  );


  xnor
  g2002
  (
    n2088,
    n1339,
    n1604,
    n1895,
    n1278
  );


  nand
  g2003
  (
    n2222,
    n1732,
    n1192,
    n856,
    n728
  );


  nor
  g2004
  (
    n2241,
    n803,
    n833,
    n1733,
    n1759
  );


  nand
  g2005
  (
    n1990,
    n1382,
    n1307,
    n1632,
    n1891
  );


  nand
  g2006
  (
    n2178,
    n1074,
    n998,
    n1868,
    n1063
  );


  nand
  g2007
  (
    KeyWire_0_58,
    n1818,
    n1532,
    n1108,
    n1096
  );


  nand
  g2008
  (
    n2221,
    n894,
    n1848,
    n896,
    n1839
  );


  xor
  g2009
  (
    n2293,
    n1150,
    n1119,
    n795,
    n1015
  );


  nor
  g2010
  (
    n2274,
    n960,
    n1907,
    n1627,
    n1890
  );


  nand
  g2011
  (
    n2077,
    n1061,
    n1414,
    n1559,
    n1398
  );


  nor
  g2012
  (
    n2242,
    n1455,
    n1342,
    n840,
    n1468
  );


  xor
  g2013
  (
    n2173,
    n1761,
    n1560,
    n1878,
    n939
  );


  xor
  g2014
  (
    n2024,
    n925,
    n1594,
    n1499,
    n1853
  );


  nand
  g2015
  (
    n2245,
    n1027,
    n1570,
    n1453,
    n1624
  );


  xnor
  g2016
  (
    n2247,
    n1477,
    n1785,
    n1422,
    n711
  );


  and
  g2017
  (
    n2106,
    n754,
    n830,
    n1584,
    n1643
  );


  xor
  g2018
  (
    n2236,
    n1190,
    n1808,
    n1429,
    n975
  );


  xnor
  g2019
  (
    n2057,
    n1201,
    n1011,
    n909,
    n997
  );


  nor
  g2020
  (
    n2002,
    n1742,
    n1285,
    n922,
    n1158
  );


  or
  g2021
  (
    n2060,
    n1704,
    n1406,
    n1151,
    n1904
  );


  xnor
  g2022
  (
    n2010,
    n1070,
    n1845,
    n942,
    n924
  );


  or
  g2023
  (
    n2163,
    n994,
    n1606,
    n1264,
    n1413
  );


  xor
  g2024
  (
    n2072,
    n1402,
    n1066,
    n796,
    n1510
  );


  xnor
  g2025
  (
    n2036,
    n1171,
    n1893,
    n706,
    n1546
  );


  xnor
  g2026
  (
    n2252,
    n1280,
    n817,
    n1494,
    n1779
  );


  xnor
  g2027
  (
    n2069,
    n722,
    n1081,
    n1370,
    n1542
  );


  xnor
  g2028
  (
    n2025,
    n903,
    n1084,
    n839,
    n1377
  );


  xnor
  g2029
  (
    n2146,
    n1692,
    n1282,
    n1816,
    n1344
  );


  xor
  g2030
  (
    n2082,
    n696,
    n950,
    n1906,
    n1589
  );


  nor
  g2031
  (
    n2298,
    n758,
    n748,
    n1521,
    n1469
  );


  nor
  g2032
  (
    n2098,
    n1545,
    n837,
    n1497,
    n1747
  );


  xnor
  g2033
  (
    KeyWire_0_29,
    n689,
    n1072,
    n1568,
    n1672
  );


  and
  g2034
  (
    n2073,
    n1218,
    n1855,
    n1054,
    n1095
  );


  and
  g2035
  (
    n2034,
    n1309,
    n697,
    n1590,
    n715
  );


  nand
  g2036
  (
    n2276,
    n1684,
    n1078,
    n717,
    n1260
  );


  xor
  g2037
  (
    n2075,
    n1726,
    n1470,
    n1567,
    n1555
  );


  and
  g2038
  (
    n2115,
    n1793,
    n1051,
    n1373,
    n1561
  );


  nor
  g2039
  (
    n2105,
    n1811,
    n1252,
    n769,
    n681
  );


  and
  g2040
  (
    n2198,
    n1639,
    n1044,
    n743,
    n1202
  );


  xor
  g2041
  (
    n2081,
    n1029,
    n1668,
    n891,
    n1204
  );


  and
  g2042
  (
    n2054,
    n1412,
    n1399,
    n677,
    n1800
  );


  or
  g2043
  (
    n2084,
    n790,
    n990,
    n1781,
    n687
  );


  and
  g2044
  (
    n2151,
    n863,
    n1769,
    n1182,
    n753
  );


  xnor
  g2045
  (
    n2188,
    n1882,
    n1118,
    n1528,
    n1357
  );


  nor
  g2046
  (
    n2240,
    n956,
    n1536,
    n1321,
    n846
  );


  nor
  g2047
  (
    n2062,
    n1149,
    n1879,
    n1439,
    n1588
  );


  and
  g2048
  (
    n2095,
    n1088,
    n1223,
    n1322,
    n1889
  );


  or
  g2049
  (
    n2227,
    n1905,
    n1383,
    n735,
    n1857
  );


  xor
  g2050
  (
    KeyWire_0_4,
    n1083,
    n1006,
    n1209,
    n1595
  );


  and
  g2051
  (
    n2130,
    n1739,
    n807,
    n1647,
    n1308
  );


  nand
  g2052
  (
    n2292,
    n921,
    n1001,
    n999,
    n1537
  );


  and
  g2053
  (
    n2257,
    n1237,
    n853,
    n1340,
    n814
  );


  xor
  g2054
  (
    n1999,
    n1310,
    n977,
    n1906,
    n1279
  );


  xor
  g2055
  (
    KeyWire_0_9,
    n1777,
    n976,
    n1622,
    n1893
  );


  xnor
  g2056
  (
    n2273,
    n1898,
    n1812,
    n890,
    n868
  );


  nor
  g2057
  (
    n2063,
    n944,
    n1609,
    n1729,
    n1191
  );


  xnor
  g2058
  (
    n2219,
    n927,
    n772,
    n1904,
    n1907
  );


  nor
  g2059
  (
    n2272,
    n750,
    n1645,
    n1106,
    n1626
  );


  xor
  g2060
  (
    n2270,
    n1901,
    n1666,
    n792,
    n1835
  );


  xnor
  g2061
  (
    n2189,
    n1030,
    n1195,
    n1085,
    n1897
  );


  xnor
  g2062
  (
    n2040,
    n1526,
    n1865,
    n1130,
    n1771
  );


  or
  g2063
  (
    n2281,
    n1564,
    n1765,
    n828,
    n1840
  );


  nor
  g2064
  (
    n2166,
    n1891,
    n1184,
    n782,
    n1207
  );


  nor
  g2065
  (
    n2131,
    n1530,
    n1159,
    n1664,
    n1428
  );


  xnor
  g2066
  (
    n2162,
    n1332,
    n664,
    n747,
    n885
  );


  and
  g2067
  (
    n2201,
    n1294,
    n898,
    n1227,
    n1144
  );


  nor
  g2068
  (
    n2266,
    n1048,
    n1432,
    n1648,
    n780
  );


  nor
  g2069
  (
    n2092,
    n1123,
    n1814,
    n1616,
    n1293
  );


  and
  g2070
  (
    n2190,
    n1050,
    n1837,
    n1376,
    n1832
  );


  or
  g2071
  (
    n2059,
    n1558,
    n1181,
    n958,
    n1541
  );


  xnor
  g2072
  (
    n2145,
    n1396,
    n951,
    n656,
    n1254
  );


  xor
  g2073
  (
    n2265,
    n1899,
    n1540,
    n733,
    n1358
  );


  nand
  g2074
  (
    n2053,
    n1238,
    n865,
    n1900,
    n1271
  );


  nand
  g2075
  (
    n2171,
    n1233,
    n1783,
    n732,
    n1107
  );


  xor
  g2076
  (
    n2235,
    n1419,
    n1598,
    n698,
    n1750
  );


  nand
  g2077
  (
    n2200,
    n1389,
    n1737,
    n1187,
    n917
  );


  xnor
  g2078
  (
    n1987,
    n850,
    n1744,
    n838,
    n670
  );


  and
  g2079
  (
    n2018,
    n1024,
    n684,
    n1903,
    n1189
  );


  xor
  g2080
  (
    n2297,
    n900,
    n1229,
    n914,
    n1008
  );


  xnor
  g2081
  (
    n2007,
    n1834,
    n1529,
    n1819,
    n1016
  );


  nand
  g2082
  (
    n2307,
    n818,
    n1679,
    n878,
    n988
  );


  nand
  g2083
  (
    n2175,
    n1901,
    n1711,
    n1034,
    n674
  );


  or
  g2084
  (
    n2259,
    n1157,
    n1891,
    n1475,
    n1270
  );


  nor
  g2085
  (
    n2037,
    n910,
    n1316,
    n1247,
    n1140
  );


  nand
  g2086
  (
    n2019,
    n1823,
    n739,
    n1092,
    n1441
  );


  xnor
  g2087
  (
    n2187,
    n979,
    n688,
    n1174,
    n1640
  );


  nand
  g2088
  (
    n2109,
    n705,
    n1301,
    n1892,
    n1139
  );


  xnor
  g2089
  (
    n2135,
    n1658,
    n1805,
    n1411,
    n963
  );


  and
  g2090
  (
    n2213,
    n1502,
    n1788,
    n931,
    n1243
  );


  nor
  g2091
  (
    n2251,
    n1415,
    n1065,
    n1421,
    n694
  );


  nand
  g2092
  (
    n2156,
    n1887,
    n848,
    n1438,
    n819
  );


  and
  g2093
  (
    n2039,
    n1773,
    n1216,
    n1706,
    n1894
  );


  xnor
  g2094
  (
    n2136,
    n712,
    n861,
    n1509,
    n679
  );


  xor
  g2095
  (
    n2102,
    n1121,
    n1602,
    n1515,
    n984
  );


  and
  g2096
  (
    n2225,
    n1557,
    n948,
    n1198,
    n1261
  );


  or
  g2097
  (
    n2041,
    n938,
    n1659,
    n1669,
    n1025
  );


  and
  g2098
  (
    n2042,
    n1099,
    n781,
    n1462,
    n835
  );


  xor
  g2099
  (
    n2138,
    n1889,
    n1348,
    n1514,
    n1607
  );


  and
  g2100
  (
    n2191,
    n1501,
    n1556,
    n1067,
    n1017
  );


  nor
  g2101
  (
    n2308,
    n1722,
    n1592,
    n1246,
    n1520
  );


  xor
  g2102
  (
    n2113,
    n1359,
    n1516,
    n1549,
    n813
  );


  xnor
  g2103
  (
    n2275,
    n881,
    n1128,
    n1143,
    n1896
  );


  xnor
  g2104
  (
    n1982,
    n798,
    n767,
    n1327,
    n1145
  );


  or
  g2105
  (
    n2080,
    n1751,
    n1311,
    n1696,
    n1211
  );


  xnor
  g2106
  (
    n2033,
    n1010,
    n682,
    n1058,
    n1380
  );


  and
  g2107
  (
    n2150,
    n1242,
    n1804,
    n1789,
    n1500
  );


  nand
  g2108
  (
    n2116,
    n1612,
    n1378,
    n1035,
    n1552
  );


  xnor
  g2109
  (
    n2078,
    n880,
    n1087,
    n1856,
    n1167
  );


  and
  g2110
  (
    n2127,
    n707,
    n1056,
    n1586,
    n737
  );


  and
  g2111
  (
    n2282,
    n1047,
    n1898,
    n726,
    n797
  );


  xnor
  g2112
  (
    n2090,
    n1343,
    n1062,
    n1891,
    n761
  );


  nand
  g2113
  (
    n2193,
    n766,
    n1219,
    n1033,
    n908
  );


  xnor
  g2114
  (
    n2133,
    n1249,
    n1892,
    n1312,
    n1360
  );


  xnor
  g2115
  (
    n2152,
    n947,
    n1543,
    n991,
    n871
  );


  xor
  g2116
  (
    n2212,
    n1708,
    n816,
    n746,
    n1478
  );


  and
  g2117
  (
    n2246,
    n1450,
    n902,
    n842,
    n1408
  );


  xnor
  g2118
  (
    n2244,
    n1743,
    n745,
    n1127,
    n1053
  );


  nor
  g2119
  (
    n2044,
    n1460,
    n844,
    n1523,
    n1677
  );


  nand
  g2120
  (
    n2035,
    n1131,
    n1548,
    n912,
    n827
  );


  and
  g2121
  (
    n2070,
    n811,
    n1257,
    n1649,
    n1727
  );


  nand
  g2122
  (
    n2047,
    n1828,
    n887,
    n1585,
    n1898
  );


  xnor
  g2123
  (
    n2231,
    n1314,
    n1021,
    n1597,
    n1183
  );


  and
  g2124
  (
    n2210,
    n1255,
    n888,
    n855,
    n701
  );


  xor
  g2125
  (
    n2195,
    n996,
    n987,
    n954,
    n1738
  );


  xnor
  g2126
  (
    n1995,
    n1262,
    n1362,
    n1901,
    n1331
  );


  nor
  g2127
  (
    n2056,
    n1880,
    n1762,
    n1713,
    n1420
  );


  nor
  g2128
  (
    n2186,
    n1375,
    n1489,
    n1512,
    n1827
  );


  xor
  g2129
  (
    n1986,
    n1579,
    n1874,
    n791,
    n1885
  );


  and
  g2130
  (
    n2114,
    n1208,
    n1678,
    n857,
    n667
  );


  nand
  g2131
  (
    n2030,
    n1416,
    n806,
    n658,
    n815
  );


  nor
  g2132
  (
    n2226,
    n1842,
    n1326,
    n1906,
    n932
  );


  or
  g2133
  (
    n2038,
    n757,
    n1372,
    n1539,
    n660
  );


  or
  g2134
  (
    n2279,
    n1605,
    n1090,
    n662,
    n1447
  );


  nor
  g2135
  (
    n2147,
    n770,
    n1210,
    n847,
    n1673
  );


  and
  g2136
  (
    n2172,
    n985,
    n1185,
    n1634,
    n1693
  );


  and
  g2137
  (
    n2209,
    n1544,
    n1653,
    n1780,
    n851
  );


  xor
  g2138
  (
    n2020,
    n1426,
    n945,
    n740,
    n1760
  );


  nor
  g2139
  (
    n2118,
    n1440,
    n1390,
    n1629,
    n1461
  );


  xnor
  g2140
  (
    n2202,
    n1101,
    n1641,
    n1655,
    n680
  );


  nor
  g2141
  (
    n2132,
    n1005,
    n1347,
    n862,
    n1487
  );


  or
  g2142
  (
    n2091,
    n1392,
    n1115,
    n1082,
    n1695
  );


  xnor
  g2143
  (
    n2052,
    n1611,
    n1775,
    n1580,
    n1113
  );


  xor
  g2144
  (
    n2048,
    n1625,
    n1635,
    n713,
    n916
  );


  nand
  g2145
  (
    n2148,
    n1069,
    n1725,
    n690,
    n1896
  );


  or
  g2146
  (
    n2153,
    n1686,
    n657,
    n1288,
    n699
  );


  or
  g2147
  (
    n2110,
    n1703,
    n672,
    n1881,
    n1897
  );


  or
  g2148
  (
    n2009,
    n1235,
    n973,
    n1334,
    n1508
  );


  or
  g2149
  (
    n2104,
    n1135,
    n1043,
    n858,
    n1506
  );


  xor
  g2150
  (
    n2295,
    n1059,
    n742,
    n1620,
    n1904
  );


  and
  g2151
  (
    n2250,
    n1434,
    n721,
    n709,
    n710
  );


  xnor
  g2152
  (
    n2214,
    n810,
    n725,
    n804,
    n1300
  );


  and
  g2153
  (
    n2262,
    n964,
    n1493,
    n1907,
    n1886
  );


  and
  g2154
  (
    n2101,
    n875,
    n845,
    n884,
    n986
  );


  or
  g2155
  (
    n2287,
    n1259,
    n799,
    n1888,
    n1825
  );


  xnor
  g2156
  (
    n2215,
    n1220,
    n760,
    n1801,
    n1905
  );


  nor
  g2157
  (
    n2117,
    n776,
    n738,
    n777,
    n1138
  );


  xnor
  g2158
  (
    n2289,
    n1367,
    n1125,
    n1795,
    n1871
  );


  nand
  g2159
  (
    n2017,
    n993,
    n1354,
    n1899,
    n661
  );


  xor
  g2160
  (
    n2229,
    n1748,
    n1752,
    n1569,
    n784
  );


  nand
  g2161
  (
    n2261,
    n1794,
    n1740,
    n1094,
    n1297
  );


  xnor
  g2162
  (
    n2128,
    n1734,
    n654,
    n1533,
    n1046
  );


  nor
  g2163
  (
    n2001,
    n802,
    n852,
    n969,
    n1710
  );


  xor
  g2164
  (
    n2179,
    n1482,
    n1872,
    n1810,
    n1110
  );


  xor
  g2165
  (
    n2263,
    n1764,
    n1052,
    n1154,
    n968
  );


  xnor
  g2166
  (
    n2208,
    n653,
    n1023,
    n1833,
    n1617
  );


  xnor
  g2167
  (
    n2159,
    n1385,
    n723,
    n1267,
    n1860
  );


  xnor
  g2168
  (
    n2230,
    n1026,
    n941,
    n801,
    n1587
  );


  and
  g2169
  (
    n2071,
    n1361,
    n1670,
    n1897,
    n1325
  );


  or
  g2170
  (
    n2067,
    n1719,
    n1554,
    n1480,
    n1452
  );


  nor
  g2171
  (
    n2032,
    n683,
    n1642,
    n961,
    n703
  );


  nor
  g2172
  (
    n2233,
    n1103,
    n1820,
    n1401,
    n1660
  );


  xnor
  g2173
  (
    n2218,
    n952,
    n1286,
    n1513,
    n1571
  );


  and
  g2174
  (
    n2161,
    n1014,
    n1345,
    n1456,
    n1898
  );


  or
  g2175
  (
    n2267,
    n1651,
    n1317,
    n794,
    n1122
  );


  or
  g2176
  (
    n2139,
    n1045,
    n1100,
    n971,
    n1272
  );


  xor
  g2177
  (
    n2141,
    n1465,
    n1806,
    n970,
    n1245
  );


  nand
  g2178
  (
    n2237,
    n1862,
    n1534,
    n1146,
    n1861
  );


  or
  g2179
  (
    n1993,
    n1654,
    n1838,
    n1687,
    n1225
  );


  nor
  g2180
  (
    n2269,
    n869,
    n893,
    n920,
    n1320
  );


  and
  g2181
  (
    n2087,
    n1036,
    n1444,
    n940,
    n897
  );


  xor
  g2182
  (
    n2050,
    n1903,
    n1199,
    n1212,
    n1826
  );


  or
  g2183
  (
    n2031,
    n1613,
    n1091,
    n1430,
    n1298
  );


  xnor
  g2184
  (
    n2249,
    n943,
    n1228,
    n1796,
    n982
  );


  and
  g2185
  (
    n2083,
    n1417,
    n1573,
    n1165,
    n1112
  );


  xor
  g2186
  (
    n2305,
    n933,
    n1013,
    n1699,
    n1694
  );


  nor
  g2187
  (
    n2205,
    n1723,
    n736,
    n1346,
    n1809
  );


  or
  g2188
  (
    n2014,
    n911,
    n663,
    n1551,
    n826
  );


  and
  g2189
  (
    n1988,
    n1903,
    n1153,
    n1904,
    n720
  );


  xnor
  g2190
  (
    n2121,
    n1776,
    n1281,
    n1064,
    n1682
  );


  nor
  g2191
  (
    n2182,
    n1661,
    n1720,
    n1111,
    n724
  );


  xnor
  g2192
  (
    n2005,
    n734,
    n1637,
    n1846,
    n1758
  );


  or
  g2193
  (
    n2197,
    n1843,
    n1215,
    n1239,
    n1000
  );


  xnor
  g2194
  (
    n2003,
    n1205,
    n1305,
    n786,
    n967
  );


  nor
  g2195
  (
    n2149,
    n1802,
    n1849,
    n1324,
    n1248
  );


  nor
  g2196
  (
    n2068,
    n1424,
    n1268,
    n1349,
    n1531
  );


  nor
  g2197
  (
    n2066,
    n918,
    n1368,
    n788,
    n1196
  );


  and
  g2198
  (
    n2119,
    n1039,
    n820,
    n1646,
    n1888
  );


  nand
  g2199
  (
    n2253,
    n1656,
    n1483,
    n1407,
    n1829
  );


  or
  g2200
  (
    n2122,
    n1902,
    n1485,
    n1675,
    n834
  );


  nor
  g2201
  (
    n2306,
    n1038,
    n1685,
    n1492,
    n1608
  );


  nand
  g2202
  (
    n2271,
    n1391,
    n1495,
    n1894,
    n1193
  );


  and
  g2203
  (
    n2216,
    n1147,
    n1700,
    n1163,
    n731
  );


  xnor
  g2204
  (
    n2011,
    n1665,
    n849,
    n744,
    n1893
  );


  or
  g2205
  (
    n2006,
    n1098,
    n995,
    n901,
    n793
  );


  xnor
  g2206
  (
    n2167,
    n1614,
    n1712,
    n708,
    n1251
  );


  nand
  g2207
  (
    n2022,
    n1869,
    n1535,
    n1787,
    n946
  );


  nand
  g2208
  (
    n2021,
    n1691,
    n1226,
    n1337,
    n1203
  );


  nor
  g2209
  (
    n2134,
    n1217,
    n1330,
    n1236,
    n764
  );


  nand
  g2210
  (
    n2278,
    n1283,
    n1873,
    n1518,
    n872
  );


  or
  g2211
  (
    n2096,
    n1633,
    n1467,
    n779,
    n1517
  );


  nand
  g2212
  (
    n2043,
    n1075,
    n809,
    n1287,
    n1524
  );


  xnor
  g2213
  (
    n2220,
    n919,
    n1681,
    n1504,
    n836
  );


  xnor
  g2214
  (
    n2294,
    n974,
    n1232,
    n691,
    n1807
  );


  nand
  g2215
  (
    n2111,
    n1055,
    n1057,
    n1519,
    n1630
  );


  xor
  g2216
  (
    n2155,
    n864,
    n1296,
    n1166,
    n1156
  );


  xor
  g2217
  (
    n2103,
    n1889,
    n1593,
    n1619,
    n1817
  );


  nand
  g2218
  (
    n2143,
    n1142,
    n1022,
    n1680,
    n1068
  );


  nor
  g2219
  (
    n2028,
    n1596,
    n1702,
    n1895,
    n655
  );


  xor
  g2220
  (
    n2284,
    n1379,
    n1547,
    n756,
    n768
  );


  or
  g2221
  (
    n2238,
    n1792,
    n1133,
    n1263,
    n1822
  );


  xnor
  g2222
  (
    n2051,
    n831,
    n1366,
    n1160,
    n1188
  );


  nand
  g2223
  (
    n2268,
    n1575,
    n1002,
    n1895,
    n1550
  );


  xor
  g2224
  (
    n2108,
    n1079,
    n676,
    n1889,
    n1716
  );


  xnor
  g2225
  (
    n2258,
    n906,
    n1117,
    n1431,
    n854
  );


  and
  g2226
  (
    n1997,
    n1384,
    n1433,
    n904,
    n1319
  );


  xor
  g2227
  (
    n2157,
    n1004,
    n1899,
    n980,
    n930
  );


  xnor
  g2228
  (
    n1996,
    n1129,
    n1353,
    n1363,
    n934
  );


  or
  g2229
  (
    n2000,
    n867,
    n1338,
    n1638,
    n1657
  );


  or
  g2230
  (
    n2192,
    n937,
    n1756,
    n1442,
    n704
  );


  and
  g2231
  (
    n2160,
    n1883,
    n1041,
    n1707,
    n1689
  );


  and
  g2232
  (
    n2094,
    n685,
    n1275,
    n1299,
    n1730
  );


  nor
  g2233
  (
    n2015,
    n1877,
    n741,
    n808,
    n1784
  );


  or
  g2234
  (
    n2243,
    n1222,
    n866,
    n1104,
    n1350
  );


  and
  g2235
  (
    n2137,
    n1086,
    n1782,
    n1315,
    n1813
  );


  and
  g2236
  (
    n2185,
    n1577,
    n1566,
    n1735,
    n959
  );


  nor
  g2237
  (
    n2300,
    n1073,
    n1527,
    n1774,
    n899
  );


  nand
  g2238
  (
    n2142,
    n1690,
    n673,
    n1019,
    n1213
  );


  nand
  g2239
  (
    n2283,
    n671,
    n1197,
    n678,
    n1841
  );


  and
  g2240
  (
    n2045,
    n1884,
    n983,
    n1404,
    n1576
  );


  nand
  g2241
  (
    n2164,
    n1042,
    n1250,
    n1448,
    n949
  );


  nor
  g2242
  (
    n2089,
    n1234,
    n775,
    n1076,
    n1221
  );


  xnor
  g2243
  (
    n2100,
    n1303,
    n755,
    n981,
    n1815
  );


  and
  g2244
  (
    n2207,
    n1890,
    n752,
    n1449,
    n1374
  );


  nor
  g2245
  (
    n2206,
    n665,
    n1459,
    n1328,
    n873
  );


  xnor
  g2246
  (
    n2129,
    n923,
    n1393,
    n1365,
    n877
  );


  or
  g2247
  (
    n1992,
    n1553,
    n1256,
    n1155,
    n1369
  );


  nor
  g2248
  (
    n2061,
    n841,
    n1194,
    n693,
    n957
  );


  and
  g2249
  (
    n2239,
    n1858,
    n1705,
    n1224,
    n1471
  );


  or
  g2250
  (
    n2211,
    n1754,
    n1701,
    n882,
    n787
  );


  xor
  g2251
  (
    n2124,
    n765,
    n1476,
    n1902,
    n1141
  );


  nand
  g2252
  (
    n2217,
    n1714,
    n1888,
    n1749,
    n1148
  );


  xor
  g2253
  (
    n1984,
    n1124,
    n1179,
    n955,
    n1718
  );


  nor
  g2254
  (
    n2299,
    n1900,
    n1864,
    n800,
    n1623
  );


  or
  g2255
  (
    n2165,
    n1603,
    n936,
    n1214,
    n812
  );


  nand
  g2256
  (
    n1998,
    n1698,
    n1289,
    n1473,
    n1572
  );


  and
  g2257
  (
    n2199,
    n1423,
    n1741,
    n1893,
    n1427
  );


  nand
  g2258
  (
    n2058,
    n905,
    n1907,
    n1772,
    n1020
  );


  and
  g2259
  (
    n1983,
    n1676,
    n1746,
    n659,
    n1474
  );


  nor
  g2260
  (
    n1994,
    n1089,
    n718,
    n1906,
    n1071
  );


  xnor
  g2261
  (
    n2264,
    n1851,
    n1821,
    n1481,
    n1436
  );


  or
  g2262
  (
    n2174,
    n1253,
    n823,
    n1591,
    n1511
  );


  or
  g2263
  (
    n2183,
    n1126,
    n1731,
    n1273,
    n1152
  );


  or
  g2264
  (
    n2256,
    n1386,
    n1491,
    n1618,
    n1136
  );


  and
  g2265
  (
    n2023,
    n773,
    n1009,
    n1899,
    n1745
  );


  nor
  g2266
  (
    n2260,
    n883,
    n1418,
    n1902,
    n1168
  );


  nand
  g2267
  (
    n1989,
    n1463,
    n1709,
    n1652,
    n1894
  );


  nor
  g2268
  (
    n2302,
    n1763,
    n1753,
    n1888,
    n886
  );


  or
  g2269
  (
    n2280,
    n1621,
    n1850,
    n965,
    n1028
  );


  and
  g2270
  (
    n1985,
    n1836,
    n1799,
    n1892,
    n926
  );


  nor
  g2271
  (
    n2065,
    n1854,
    n1313,
    n1905,
    n1628
  );


  nor
  g2272
  (
    n2046,
    n1097,
    n1037,
    n1169,
    n1105
  );


  xnor
  g2273
  (
    n2140,
    n962,
    n1371,
    n1329,
    n1241
  );


  xor
  g2274
  (
    n2004,
    n1790,
    n1870,
    n1077,
    n1290
  );


  xnor
  g2275
  (
    n2184,
    n702,
    n1007,
    n913,
    n1715
  );


  and
  g2276
  (
    n2168,
    n1172,
    n1186,
    n686,
    n1895
  );


  buf
  g2277
  (
    n2372,
    n2235
  );


  not
  g2278
  (
    n2374,
    n2075
  );


  not
  g2279
  (
    n2321,
    n2243
  );


  not
  g2280
  (
    n2327,
    n2051
  );


  not
  g2281
  (
    n2380,
    n2003
  );


  buf
  g2282
  (
    n2382,
    n2278
  );


  buf
  g2283
  (
    n2394,
    n2035
  );


  buf
  g2284
  (
    n2388,
    n2016
  );


  not
  g2285
  (
    n2371,
    n2274
  );


  not
  g2286
  (
    n2351,
    n1988
  );


  not
  g2287
  (
    n2370,
    n2131
  );


  buf
  g2288
  (
    KeyWire_0_8,
    n2183
  );


  and
  g2289
  (
    KeyWire_0_53,
    n2227,
    n2004
  );


  and
  g2290
  (
    n2389,
    n2287,
    n2086,
    n2097,
    n2053
  );


  xor
  g2291
  (
    n2342,
    n2204,
    n2029,
    n2058,
    n2065
  );


  or
  g2292
  (
    n2322,
    n2156,
    n2264,
    n2149,
    n2080
  );


  nand
  g2293
  (
    n2356,
    n2195,
    n2074,
    n2260,
    n2201
  );


  or
  g2294
  (
    n2348,
    n2008,
    n2151,
    n2114,
    n2178
  );


  or
  g2295
  (
    n2334,
    n2247,
    n2163,
    n2110,
    n2041
  );


  nand
  g2296
  (
    n2339,
    n2141,
    n2026,
    n2048,
    n2215
  );


  nor
  g2297
  (
    n2381,
    n2139,
    n2069,
    n2127,
    n1996
  );


  xor
  g2298
  (
    n2336,
    n2084,
    n2118,
    n2030,
    n2112
  );


  and
  g2299
  (
    n2383,
    n2277,
    n2211,
    n2280,
    n2055
  );


  xor
  g2300
  (
    n2393,
    n2108,
    n2023,
    n2214,
    n2095
  );


  nand
  g2301
  (
    n2367,
    n2001,
    n2135,
    n2089,
    n2076
  );


  and
  g2302
  (
    n2375,
    n2262,
    n2129,
    n2134,
    n2033
  );


  nor
  g2303
  (
    n2366,
    n2044,
    n2255,
    n2073,
    n2190
  );


  xnor
  g2304
  (
    n2319,
    n2000,
    n2162,
    n2115,
    n2085
  );


  or
  g2305
  (
    n2337,
    n2037,
    n2052,
    n2281,
    n2111
  );


  xnor
  g2306
  (
    n2346,
    n2273,
    n2094,
    n2106,
    n2144
  );


  and
  g2307
  (
    n2326,
    n2186,
    n2248,
    n2070,
    n2039
  );


  or
  g2308
  (
    n2317,
    n1984,
    n2206,
    n2254,
    n2284
  );


  xor
  g2309
  (
    n2343,
    n2205,
    n2208,
    n1998,
    n2017
  );


  nand
  g2310
  (
    n2344,
    n2050,
    n2099,
    n2068,
    n2054
  );


  and
  g2311
  (
    n2390,
    n1981,
    n2224,
    n2174,
    n2259
  );


  nor
  g2312
  (
    n2313,
    n2213,
    n2282,
    n2061,
    n2228
  );


  and
  g2313
  (
    n2345,
    n2153,
    n1987,
    n2117,
    n2167
  );


  or
  g2314
  (
    n2385,
    n2232,
    n2113,
    n2275,
    n2238
  );


  xor
  g2315
  (
    n2364,
    n2252,
    n2107,
    n2126,
    n2290
  );


  nor
  g2316
  (
    n2333,
    n2270,
    n2161,
    n2249,
    n2005
  );


  nor
  g2317
  (
    n2354,
    n2104,
    n1995,
    n2120,
    n1983
  );


  nand
  g2318
  (
    n2325,
    n1990,
    n2202,
    n2157,
    n2143
  );


  xor
  g2319
  (
    n2340,
    n2171,
    n2010,
    n1999,
    n1991
  );


  and
  g2320
  (
    n2338,
    n2216,
    n2133,
    n2142,
    n1992
  );


  or
  g2321
  (
    n2379,
    n2239,
    n2064,
    n2087,
    n2272
  );


  or
  g2322
  (
    n2330,
    n2257,
    n2203,
    n2182,
    n2226
  );


  xnor
  g2323
  (
    n2323,
    n2173,
    n2231,
    n2006,
    n2240
  );


  or
  g2324
  (
    n2324,
    n2138,
    n2036,
    n2116,
    n2196
  );


  and
  g2325
  (
    n2316,
    n2060,
    n2028,
    n2062,
    n2067
  );


  xor
  g2326
  (
    n2314,
    n2102,
    n2197,
    n2072,
    n2015
  );


  nor
  g2327
  (
    n2315,
    n2217,
    n2024,
    n2007,
    n2047
  );


  nor
  g2328
  (
    n2349,
    n2283,
    n2170,
    n2261,
    n2021
  );


  and
  g2329
  (
    n2341,
    n2210,
    n2057,
    n2014,
    n2032
  );


  nand
  g2330
  (
    n2312,
    n2091,
    n2124,
    n2098,
    n2079
  );


  xnor
  g2331
  (
    n2311,
    n2209,
    n2166,
    n2123,
    n2253
  );


  and
  g2332
  (
    n2369,
    n2176,
    n2158,
    n2137,
    n2152
  );


  nand
  g2333
  (
    n2376,
    n2212,
    n2034,
    n2221,
    n2207
  );


  nand
  g2334
  (
    n2365,
    n2130,
    n2078,
    n2031,
    n2180
  );


  nor
  g2335
  (
    n2395,
    n2159,
    n2096,
    n2245,
    n2154
  );


  nand
  g2336
  (
    n2331,
    n2147,
    n2199,
    n2194,
    n2056
  );


  xor
  g2337
  (
    n2355,
    n2092,
    n1997,
    n2244,
    n2172
  );


  nor
  g2338
  (
    n2378,
    n2230,
    n2150,
    n2038,
    n2223
  );


  and
  g2339
  (
    n2373,
    n2286,
    n2090,
    n2042,
    n1993
  );


  xnor
  g2340
  (
    n2386,
    n2105,
    n2122,
    n2266,
    n2225
  );


  xnor
  g2341
  (
    n2361,
    n2145,
    n2009,
    n2002,
    n2220
  );


  nand
  g2342
  (
    n2362,
    n2125,
    n2233,
    n2265,
    n2082
  );


  xnor
  g2343
  (
    n2360,
    n2268,
    n2018,
    n2222,
    n1986
  );


  and
  g2344
  (
    n2387,
    n2019,
    n1982,
    n2229,
    n2049
  );


  nor
  g2345
  (
    n2318,
    n2011,
    n2119,
    n2160,
    n2193
  );


  nor
  g2346
  (
    n2391,
    n2168,
    n2043,
    n2279,
    n2063
  );


  xnor
  g2347
  (
    n2352,
    n2181,
    n2198,
    n2164,
    n2200
  );


  or
  g2348
  (
    n2392,
    n2077,
    n2236,
    n2271,
    n2258
  );


  xor
  g2349
  (
    n2358,
    n2251,
    n2100,
    n2045,
    n2148
  );


  xnor
  g2350
  (
    n2396,
    n2046,
    n2013,
    n2165,
    n2155
  );


  xnor
  g2351
  (
    n2353,
    n2012,
    n2040,
    n2025,
    n2191
  );


  and
  g2352
  (
    n2384,
    n2285,
    n2269,
    n2093,
    n2066
  );


  xor
  g2353
  (
    n2368,
    n2169,
    n2140,
    n2276,
    n2121
  );


  nand
  g2354
  (
    n2347,
    n2246,
    n2234,
    n2219,
    n2088
  );


  xnor
  g2355
  (
    n2320,
    n2267,
    n2136,
    n2250,
    n2020
  );


  nand
  g2356
  (
    n2350,
    n2103,
    n2175,
    n2177,
    n2192
  );


  or
  g2357
  (
    n2359,
    n2189,
    n2109,
    n2218,
    n1989
  );


  or
  g2358
  (
    KeyWire_0_2,
    n2185,
    n2071,
    n2059,
    n2081
  );


  and
  g2359
  (
    n2328,
    n2288,
    n2256,
    n2237,
    n2101
  );


  or
  g2360
  (
    n2335,
    n1985,
    n2128,
    n2242,
    n2263
  );


  or
  g2361
  (
    n2332,
    n2027,
    n2188,
    n2179,
    n1994
  );


  and
  g2362
  (
    n2377,
    n2083,
    n2184,
    n2241,
    n2132
  );


  xnor
  g2363
  (
    n2357,
    n2289,
    n2146,
    n2022,
    n2187
  );


  not
  g2364
  (
    n2432,
    n2386
  );


  buf
  g2365
  (
    n2514,
    n1916
  );


  not
  g2366
  (
    n2460,
    n1909
  );


  not
  g2367
  (
    n2509,
    n2317
  );


  not
  g2368
  (
    n2451,
    n2361
  );


  not
  g2369
  (
    n2447,
    n2386
  );


  not
  g2370
  (
    n2433,
    n2376
  );


  buf
  g2371
  (
    n2482,
    n1915
  );


  not
  g2372
  (
    n2405,
    n2393
  );


  not
  g2373
  (
    n2516,
    n2352
  );


  buf
  g2374
  (
    n2454,
    n2344
  );


  buf
  g2375
  (
    n2471,
    n2324
  );


  buf
  g2376
  (
    n2493,
    n2396
  );


  buf
  g2377
  (
    n2461,
    n2379
  );


  buf
  g2378
  (
    n2421,
    n2391
  );


  not
  g2379
  (
    n2397,
    n2315
  );


  not
  g2380
  (
    n2499,
    n2340
  );


  not
  g2381
  (
    n2423,
    n2394
  );


  not
  g2382
  (
    n2494,
    n2358
  );


  not
  g2383
  (
    n2409,
    n2365
  );


  buf
  g2384
  (
    n2414,
    n1909
  );


  not
  g2385
  (
    n2410,
    n2395
  );


  buf
  g2386
  (
    n2453,
    n1909
  );


  buf
  g2387
  (
    n2424,
    n2363
  );


  buf
  g2388
  (
    n2466,
    n2319
  );


  not
  g2389
  (
    n2399,
    n2322
  );


  not
  g2390
  (
    n2408,
    n1913
  );


  not
  g2391
  (
    n2444,
    n1914
  );


  not
  g2392
  (
    n2449,
    n2331
  );


  buf
  g2393
  (
    n2428,
    n2349
  );


  buf
  g2394
  (
    n2434,
    n2374
  );


  buf
  g2395
  (
    n2486,
    n2391
  );


  buf
  g2396
  (
    n2440,
    n2396
  );


  buf
  g2397
  (
    n2418,
    n2316
  );


  buf
  g2398
  (
    n2400,
    n1915
  );


  not
  g2399
  (
    n2484,
    n2394
  );


  not
  g2400
  (
    n2415,
    n1916
  );


  not
  g2401
  (
    n2426,
    n2384
  );


  buf
  g2402
  (
    n2441,
    n2392
  );


  not
  g2403
  (
    n2459,
    n2390
  );


  not
  g2404
  (
    n2457,
    n2388
  );


  buf
  g2405
  (
    n2510,
    n2312
  );


  not
  g2406
  (
    n2467,
    n2390
  );


  not
  g2407
  (
    n2501,
    n2355
  );


  not
  g2408
  (
    n2480,
    n1916
  );


  buf
  g2409
  (
    KeyWire_0_56,
    n1917
  );


  not
  g2410
  (
    n2419,
    n2389
  );


  buf
  g2411
  (
    n2469,
    n1916
  );


  not
  g2412
  (
    KeyWire_0_23,
    n2390
  );


  not
  g2413
  (
    n2508,
    n2387
  );


  buf
  g2414
  (
    n2425,
    n1911
  );


  not
  g2415
  (
    n2507,
    n2386
  );


  buf
  g2416
  (
    n2462,
    n1912
  );


  not
  g2417
  (
    n2398,
    n2396
  );


  buf
  g2418
  (
    n2475,
    n1914
  );


  buf
  g2419
  (
    n2429,
    n2369
  );


  not
  g2420
  (
    n2417,
    n2350
  );


  buf
  g2421
  (
    n2427,
    n2383
  );


  buf
  g2422
  (
    n2489,
    n2326
  );


  not
  g2423
  (
    n2503,
    n2338
  );


  not
  g2424
  (
    n2517,
    n2386
  );


  buf
  g2425
  (
    n2430,
    n2389
  );


  not
  g2426
  (
    n2452,
    n2332
  );


  not
  g2427
  (
    n2479,
    n1910
  );


  buf
  g2428
  (
    n2491,
    n2395
  );


  not
  g2429
  (
    n2435,
    n2377
  );


  not
  g2430
  (
    n2443,
    n2321
  );


  buf
  g2431
  (
    n2500,
    n1914
  );


  buf
  g2432
  (
    n2437,
    n2351
  );


  buf
  g2433
  (
    n2506,
    n2390
  );


  buf
  g2434
  (
    n2442,
    n2348
  );


  not
  g2435
  (
    n2477,
    n2367
  );


  buf
  g2436
  (
    n2511,
    n2387
  );


  not
  g2437
  (
    n2456,
    n2362
  );


  buf
  g2438
  (
    n2497,
    n1910
  );


  buf
  g2439
  (
    n2518,
    n1912
  );


  buf
  g2440
  (
    n2502,
    n1911
  );


  not
  g2441
  (
    n2403,
    n2395
  );


  not
  g2442
  (
    n2487,
    n2389
  );


  not
  g2443
  (
    n2481,
    n2314
  );


  buf
  g2444
  (
    n2492,
    n2323
  );


  buf
  g2445
  (
    n2406,
    n2389
  );


  not
  g2446
  (
    n2496,
    n1917
  );


  buf
  g2447
  (
    n2445,
    n2356
  );


  buf
  g2448
  (
    n2438,
    n1910
  );


  not
  g2449
  (
    n2515,
    n1911
  );


  not
  g2450
  (
    n2490,
    n2330
  );


  not
  g2451
  (
    n2498,
    n1915
  );


  buf
  g2452
  (
    n2412,
    n2359
  );


  buf
  g2453
  (
    n2483,
    n2393
  );


  buf
  g2454
  (
    n2448,
    n2382
  );


  buf
  g2455
  (
    n2488,
    n1911
  );


  not
  g2456
  (
    n2464,
    n1917
  );


  not
  g2457
  (
    n2468,
    n2371
  );


  buf
  g2458
  (
    n2513,
    n2373
  );


  buf
  g2459
  (
    n2420,
    n2391
  );


  not
  g2460
  (
    n2465,
    n2387
  );


  not
  g2461
  (
    n2401,
    n2329
  );


  not
  g2462
  (
    n2407,
    n2337
  );


  buf
  g2463
  (
    n2512,
    n2372
  );


  buf
  g2464
  (
    n2505,
    n2381
  );


  buf
  g2465
  (
    n2478,
    n2311
  );


  not
  g2466
  (
    n2455,
    n2310
  );


  not
  g2467
  (
    n2446,
    n2325
  );


  buf
  g2468
  (
    n2439,
    n2318
  );


  not
  g2469
  (
    n2413,
    n2320
  );


  not
  g2470
  (
    n2495,
    n2380
  );


  buf
  g2471
  (
    n2436,
    n2333
  );


  not
  g2472
  (
    n2476,
    n1913
  );


  or
  g2473
  (
    n2473,
    n1908,
    n2354,
    n2346,
    n2335
  );


  and
  g2474
  (
    n2472,
    n2353,
    n2343,
    n2392
  );


  and
  g2475
  (
    n2431,
    n2313,
    n2327,
    n2370,
    n2385
  );


  nand
  g2476
  (
    n2470,
    n2392,
    n2345,
    n1912,
    n2339
  );


  xor
  g2477
  (
    n2416,
    n2341,
    n2391,
    n2360,
    n2388
  );


  xor
  g2478
  (
    n2422,
    n2395,
    n1913,
    n2385,
    n2342
  );


  nor
  g2479
  (
    n2504,
    n1915,
    n2347,
    n2394,
    n2364
  );


  xnor
  g2480
  (
    n2458,
    n1910,
    n2387,
    n2394,
    n2378
  );


  and
  g2481
  (
    n2450,
    n1917,
    n2336,
    n2375,
    n2388
  );


  nor
  g2482
  (
    n2402,
    n2357,
    n2388,
    n2334,
    n2393
  );


  and
  g2483
  (
    n2485,
    n1913,
    n2393,
    n2328,
    n2385
  );


  or
  g2484
  (
    n2474,
    n2368,
    n2385,
    n1914,
    n1912
  );


  nand
  g2485
  (
    n2411,
    n1909,
    n2366,
    n1908
  );


  not
  g2486
  (
    n2565,
    n2455
  );


  not
  g2487
  (
    n2519,
    n2426
  );


  buf
  g2488
  (
    n2563,
    n2449
  );


  not
  g2489
  (
    n2552,
    n2447
  );


  buf
  g2490
  (
    n2560,
    n2405
  );


  not
  g2491
  (
    n2549,
    n2423
  );


  buf
  g2492
  (
    n2525,
    n2414
  );


  buf
  g2493
  (
    n2528,
    n2435
  );


  not
  g2494
  (
    n2529,
    n2473
  );


  not
  g2495
  (
    n2546,
    n2474
  );


  not
  g2496
  (
    n2534,
    n2498
  );


  not
  g2497
  (
    n2537,
    n1918
  );


  buf
  g2498
  (
    n2530,
    n2462
  );


  buf
  g2499
  (
    n2536,
    n2486
  );


  xnor
  g2500
  (
    n2548,
    n2482,
    n2425
  );


  nand
  g2501
  (
    n2559,
    n1930,
    n2476,
    n2441,
    n1927
  );


  nand
  g2502
  (
    n2523,
    n2420,
    n2421,
    n1926,
    n2417
  );


  and
  g2503
  (
    n2531,
    n2501,
    n1931,
    n2492,
    n2418
  );


  xor
  g2504
  (
    n2567,
    n2439,
    n1929,
    n2406,
    n2472
  );


  or
  g2505
  (
    n2541,
    n2495,
    n1932,
    n2491,
    n1922
  );


  xor
  g2506
  (
    n2554,
    n1928,
    n2453,
    n32,
    n2463
  );


  xnor
  g2507
  (
    n2522,
    n1925,
    n2398,
    n1929,
    n1922
  );


  or
  g2508
  (
    n2571,
    n1920,
    n2440,
    n1924,
    n1931
  );


  xnor
  g2509
  (
    n2569,
    n2468,
    n2437,
    n2404,
    n2494
  );


  or
  g2510
  (
    n2526,
    n1919,
    n2475,
    n1929,
    n1922
  );


  nor
  g2511
  (
    n2538,
    n2459,
    n1929,
    n1920,
    n2467
  );


  and
  g2512
  (
    n2544,
    n1924,
    n2466,
    n1932,
    n2433
  );


  nand
  g2513
  (
    n2542,
    n2479,
    n2457,
    n1928,
    n1923
  );


  or
  g2514
  (
    n2550,
    n2431,
    n1928,
    n2470,
    n32
  );


  xor
  g2515
  (
    n2561,
    n1923,
    n2400,
    n2500,
    n2497
  );


  nand
  g2516
  (
    n2566,
    n1923,
    n2432,
    n2461,
    n2424
  );


  and
  g2517
  (
    n2558,
    n1926,
    n1925,
    n2458,
    n1920
  );


  nand
  g2518
  (
    n2557,
    n1925,
    n2412,
    n1918,
    n2427
  );


  xnor
  g2519
  (
    n2524,
    n2483,
    n2450,
    n2456,
    n2469
  );


  or
  g2520
  (
    n2532,
    n2496,
    n2480,
    n2490,
    n1926
  );


  or
  g2521
  (
    n2521,
    n2444,
    n1921,
    n2502,
    n1918
  );


  xnor
  g2522
  (
    n2564,
    n2434,
    n2448,
    n1926,
    n2416
  );


  nand
  g2523
  (
    n2533,
    n2442,
    n1932,
    n2399,
    n2499
  );


  xor
  g2524
  (
    n2535,
    n1921,
    n2413,
    n32,
    n1930
  );


  xor
  g2525
  (
    n2520,
    n2460,
    n1919,
    n2445,
    n2438
  );


  or
  g2526
  (
    n2562,
    n1919,
    n2408,
    n1923,
    n1931
  );


  nand
  g2527
  (
    n2570,
    n1927,
    n2489,
    n1919,
    n1918
  );


  or
  g2528
  (
    n2543,
    n2484,
    n1921,
    n1925,
    n2443
  );


  nand
  g2529
  (
    n2551,
    n2481,
    n2478,
    n2464,
    n2430
  );


  xor
  g2530
  (
    n2555,
    n2454,
    n2488,
    n2409,
    n2411
  );


  nor
  g2531
  (
    n2540,
    n2487,
    n1930,
    n2446
  );


  and
  g2532
  (
    n2556,
    n2465,
    n2401,
    n2485,
    n1927
  );


  and
  g2533
  (
    n2553,
    n2428,
    n1920,
    n2407,
    n1922
  );


  nor
  g2534
  (
    n2545,
    n2402,
    n2419,
    n2477,
    n2451
  );


  xor
  g2535
  (
    n2527,
    n1921,
    n2403,
    n2397,
    n2436
  );


  xor
  g2536
  (
    n2539,
    n1924,
    n1928,
    n2471,
    n2410
  );


  nor
  g2537
  (
    n2568,
    n2452,
    n1924,
    n1927,
    n2415
  );


  xor
  g2538
  (
    n2547,
    n1931,
    n2429,
    n2493,
    n2422
  );


  buf
  g2539
  (
    n2607,
    n2565
  );


  not
  g2540
  (
    n2601,
    n1942
  );


  buf
  g2541
  (
    n2578,
    n2549
  );


  buf
  g2542
  (
    n2572,
    n2565
  );


  buf
  g2543
  (
    n2575,
    n2535
  );


  buf
  g2544
  (
    n2579,
    n1941
  );


  buf
  g2545
  (
    n2586,
    n2564
  );


  not
  g2546
  (
    n2599,
    n2534
  );


  not
  g2547
  (
    n2597,
    n1935
  );


  not
  g2548
  (
    n2592,
    n1942
  );


  or
  g2549
  (
    n2591,
    n2537,
    n2566
  );


  nand
  g2550
  (
    n2577,
    n1935,
    n1936,
    n1941
  );


  or
  g2551
  (
    n2587,
    n2538,
    n1940,
    n2566,
    n2530
  );


  nand
  g2552
  (
    n2588,
    n2520,
    n2570,
    n1932,
    n2545
  );


  and
  g2553
  (
    n2589,
    n2571,
    n1938,
    n2568,
    n2529
  );


  xor
  g2554
  (
    n2602,
    n1943,
    n2568,
    n1937,
    n1934
  );


  xor
  g2555
  (
    n2603,
    n2567,
    n2523,
    n2561,
    n2557
  );


  xor
  g2556
  (
    n2598,
    n2570,
    n2555,
    n1937,
    n2569
  );


  and
  g2557
  (
    n2606,
    n2567,
    n1933,
    n2546,
    n2554
  );


  or
  g2558
  (
    n2594,
    n1933,
    n2568,
    n1940,
    n1939
  );


  nor
  g2559
  (
    n2600,
    n1940,
    n2566,
    n1933
  );


  or
  g2560
  (
    n2583,
    n2568,
    n2536,
    n2560,
    n2565
  );


  nor
  g2561
  (
    n2593,
    n2525,
    n1940,
    n2542,
    n2567
  );


  nor
  g2562
  (
    n2590,
    n2570,
    n2540,
    n2552,
    n1935
  );


  nor
  g2563
  (
    n2595,
    n1934,
    n1933,
    n1938,
    n1935
  );


  nand
  g2564
  (
    n2574,
    n1944,
    n2556,
    n2528,
    n2548
  );


  nand
  g2565
  (
    n2576,
    n2551,
    n2526,
    n2539,
    n2563
  );


  xor
  g2566
  (
    n2580,
    n2553,
    n1941,
    n2544,
    n1942
  );


  or
  g2567
  (
    n2584,
    n2570,
    n1934,
    n1943,
    n1937
  );


  nor
  g2568
  (
    n2609,
    n1943,
    n2531,
    n2571,
    n1936
  );


  and
  g2569
  (
    n2604,
    n2532,
    n2547,
    n2558,
    n1944
  );


  and
  g2570
  (
    n2596,
    n1938,
    n2533,
    n2569,
    n1941
  );


  nand
  g2571
  (
    n2581,
    n1943,
    n2541,
    n2559,
    n2527
  );


  xnor
  g2572
  (
    n2605,
    n2562,
    n2543,
    n1942,
    n1939
  );


  nand
  g2573
  (
    n2608,
    n1936,
    n1944,
    n2565,
    n2550
  );


  xnor
  g2574
  (
    n2582,
    n2521,
    n2519,
    n2524,
    n2569
  );


  nor
  g2575
  (
    n2573,
    n2567,
    n2569,
    n1934,
    n1939
  );


  xor
  g2576
  (
    n2585,
    n1938,
    n2522,
    n1939,
    n1937
  );


  or
  g2577
  (
    n2612,
    n2572,
    n1946,
    n2573
  );


  xor
  g2578
  (
    n2611,
    n1944,
    n2574,
    n1945
  );


  xnor
  g2579
  (
    n2610,
    n1946,
    n1945
  );


  or
  g2580
  (
    n2619,
    n1950,
    n1949,
    n2611,
    n1953
  );


  xor
  g2581
  (
    n2618,
    n1954,
    n1947,
    n1950,
    n2612
  );


  nand
  g2582
  (
    n2614,
    n1950,
    n2611,
    n1949
  );


  and
  g2583
  (
    n2622,
    n2612,
    n2610
  );


  xor
  g2584
  (
    n2623,
    n1947,
    n1950,
    n1955,
    n1953
  );


  nand
  g2585
  (
    n2621,
    n1954,
    n1955,
    n1951,
    n1948
  );


  or
  g2586
  (
    n2616,
    n1947,
    n1951,
    n1952
  );


  xor
  g2587
  (
    n2613,
    n2612,
    n2611,
    n1948,
    n1955
  );


  and
  g2588
  (
    n2624,
    n1951,
    n2610,
    n1954,
    n1953
  );


  or
  g2589
  (
    n2615,
    n1955,
    n2610,
    n2611,
    n1952
  );


  nor
  g2590
  (
    n2620,
    n1949,
    n1948,
    n1952,
    n1954
  );


  nand
  g2591
  (
    n2617,
    n1952,
    n1947,
    n1948,
    n1953
  );


  nor
  g2592
  (
    n2638,
    n1956,
    n1958,
    n2617,
    n1965
  );


  xor
  g2593
  (
    n2643,
    n1957,
    n1962,
    n1956,
    n1967
  );


  and
  g2594
  (
    n2639,
    n2615,
    n2616,
    n1967
  );


  xnor
  g2595
  (
    n2635,
    n2617,
    n1962,
    n1957,
    n1960
  );


  xnor
  g2596
  (
    n2632,
    n2615,
    n1963,
    n1959,
    n1956
  );


  nor
  g2597
  (
    n2641,
    n1964,
    n1963,
    n1960,
    n1961
  );


  xor
  g2598
  (
    n2629,
    n2617,
    n1959,
    n2614
  );


  nand
  g2599
  (
    n2626,
    n1964,
    n1958,
    n1963,
    n1967
  );


  nor
  g2600
  (
    n2631,
    n1962,
    n1968,
    n1965,
    n1966
  );


  nand
  g2601
  (
    n2627,
    n2613,
    n2613,
    n1966,
    n1968
  );


  nand
  g2602
  (
    n2625,
    n1965,
    n2616,
    n1970
  );


  or
  g2603
  (
    n2628,
    n1964,
    n2617,
    n1968,
    n1959
  );


  xnor
  g2604
  (
    n2644,
    n1957,
    n1960,
    n1970
  );


  xnor
  g2605
  (
    n2636,
    n2613,
    n1969,
    n1967,
    n1962
  );


  xor
  g2606
  (
    n2630,
    n1958,
    n1969,
    n1966,
    n1961
  );


  nand
  g2607
  (
    n2640,
    n2614,
    n1961,
    n1965
  );


  xnor
  g2608
  (
    n2634,
    n1956,
    n1968,
    n1966,
    n1969
  );


  nand
  g2609
  (
    n2633,
    n1963,
    n1958,
    n1957,
    n2616
  );


  and
  g2610
  (
    n2637,
    n2613,
    n1964,
    n1969,
    n1959
  );


  xor
  g2611
  (
    n2642,
    n2615,
    n2615,
    n2614,
    n1960
  );


  not
  g2612
  (
    n2646,
    n2638
  );


  not
  g2613
  (
    n2645,
    n2637
  );


  buf
  g2614
  (
    n2650,
    n2645
  );


  buf
  g2615
  (
    n2648,
    n2645
  );


  not
  g2616
  (
    n2647,
    n2645
  );


  not
  g2617
  (
    n2649,
    n2645
  );


  not
  g2618
  (
    n2654,
    n2650
  );


  not
  g2619
  (
    n2657,
    n2650
  );


  not
  g2620
  (
    n2656,
    n2648
  );


  buf
  g2621
  (
    n2658,
    n2650
  );


  not
  g2622
  (
    n2653,
    n2650
  );


  not
  g2623
  (
    n2651,
    n2647
  );


  buf
  g2624
  (
    n2652,
    n2649
  );


  not
  g2625
  (
    n2655,
    n2649
  );


  not
  g2626
  (
    n2667,
    n2653
  );


  not
  g2627
  (
    n2668,
    n2654
  );


  not
  g2628
  (
    n2671,
    n2654
  );


  buf
  g2629
  (
    n2685,
    n2655
  );


  buf
  g2630
  (
    n2675,
    n2657
  );


  not
  g2631
  (
    n2674,
    n2656
  );


  not
  g2632
  (
    n2670,
    n2654
  );


  not
  g2633
  (
    n2677,
    n2655
  );


  buf
  g2634
  (
    n2680,
    n2653
  );


  not
  g2635
  (
    n2664,
    n2652
  );


  buf
  g2636
  (
    n2661,
    n2656
  );


  not
  g2637
  (
    n2672,
    n2654
  );


  buf
  g2638
  (
    n2679,
    n2656
  );


  not
  g2639
  (
    n2676,
    n2657
  );


  not
  g2640
  (
    n2682,
    n2657
  );


  not
  g2641
  (
    n2659,
    n2657
  );


  not
  g2642
  (
    n2660,
    n2655
  );


  buf
  g2643
  (
    n2666,
    n2651
  );


  buf
  g2644
  (
    n2686,
    n2652
  );


  not
  g2645
  (
    n2662,
    n2652
  );


  not
  g2646
  (
    n2673,
    n2655
  );


  buf
  g2647
  (
    n2665,
    n2653
  );


  not
  g2648
  (
    KeyWire_0_45,
    n2656
  );


  buf
  g2649
  (
    n2669,
    n2651
  );


  buf
  g2650
  (
    n2683,
    n2653
  );


  buf
  g2651
  (
    n2684,
    n2651
  );


  not
  g2652
  (
    n2678,
    n2652
  );


  not
  g2653
  (
    n2681,
    n2651
  );


  not
  g2654
  (
    n2757,
    n2680
  );


  not
  g2655
  (
    n2744,
    n2683
  );


  buf
  g2656
  (
    n2739,
    n2686
  );


  not
  g2657
  (
    n2761,
    n2663
  );


  buf
  g2658
  (
    n2779,
    n2666
  );


  buf
  g2659
  (
    n2687,
    n2592
  );


  buf
  g2660
  (
    n2793,
    n2596
  );


  not
  g2661
  (
    n2713,
    n2662
  );


  not
  g2662
  (
    n2700,
    n2663
  );


  not
  g2663
  (
    KeyWire_0_34,
    n2597
  );


  buf
  g2664
  (
    n2755,
    n2590
  );


  buf
  g2665
  (
    n2772,
    n1971
  );


  buf
  g2666
  (
    n2749,
    n2599
  );


  not
  g2667
  (
    n2694,
    n2583
  );


  buf
  g2668
  (
    n2727,
    n1972
  );


  not
  g2669
  (
    n2737,
    n2679
  );


  buf
  g2670
  (
    n2730,
    n2603
  );


  not
  g2671
  (
    n2688,
    n2602
  );


  buf
  g2672
  (
    n2702,
    n2661
  );


  buf
  g2673
  (
    n2701,
    n2672
  );


  buf
  g2674
  (
    n2760,
    n2680
  );


  buf
  g2675
  (
    n2735,
    n2667
  );


  buf
  g2676
  (
    n2743,
    n2668
  );


  not
  g2677
  (
    n2762,
    n2676
  );


  buf
  g2678
  (
    n2721,
    n2679
  );


  buf
  g2679
  (
    n2765,
    n2669
  );


  not
  g2680
  (
    n2777,
    n2602
  );


  buf
  g2681
  (
    n2715,
    n2589
  );


  buf
  g2682
  (
    n2719,
    n2677
  );


  not
  g2683
  (
    n2724,
    n2600
  );


  not
  g2684
  (
    n2690,
    n2672
  );


  not
  g2685
  (
    n2742,
    n2599
  );


  buf
  g2686
  (
    n2795,
    n2586
  );


  buf
  g2687
  (
    n2782,
    n2591
  );


  not
  g2688
  (
    n2699,
    n2685
  );


  buf
  g2689
  (
    n2754,
    n2680
  );


  buf
  g2690
  (
    n2776,
    n2659
  );


  buf
  g2691
  (
    n2763,
    n2600
  );


  buf
  g2692
  (
    KeyWire_0_18,
    n2594
  );


  not
  g2693
  (
    n2720,
    n2601
  );


  not
  g2694
  (
    n2718,
    n2664
  );


  buf
  g2695
  (
    n2738,
    n2662
  );


  buf
  g2696
  (
    n2689,
    n2575
  );


  buf
  g2697
  (
    n2797,
    n2578
  );


  buf
  g2698
  (
    n2774,
    n2675
  );


  or
  g2699
  (
    n2787,
    n2686,
    n2681
  );


  nor
  g2700
  (
    n2704,
    n2685,
    n2603
  );


  and
  g2701
  (
    n2789,
    n2662,
    n2602
  );


  or
  g2702
  (
    n2707,
    n2674,
    n1972
  );


  xor
  g2703
  (
    n2728,
    n2668,
    n2673
  );


  nand
  g2704
  (
    n2711,
    n2660,
    n2579
  );


  and
  g2705
  (
    n2790,
    n2674,
    n2663
  );


  or
  g2706
  (
    n2784,
    n2599,
    n2678
  );


  or
  g2707
  (
    n2768,
    n1971,
    n2603
  );


  xnor
  g2708
  (
    n2692,
    n2673,
    n2682
  );


  nand
  g2709
  (
    n2722,
    n2671,
    n2666
  );


  xnor
  g2710
  (
    n2767,
    n2661,
    n2598
  );


  and
  g2711
  (
    n2708,
    n2677,
    n2678
  );


  or
  g2712
  (
    n2736,
    n1971,
    n2585
  );


  nor
  g2713
  (
    n2691,
    n2582,
    n2665
  );


  nor
  g2714
  (
    n2705,
    n2660,
    n2673
  );


  xor
  g2715
  (
    n2709,
    n2577,
    n2675
  );


  nand
  g2716
  (
    n2747,
    n2660,
    n2676
  );


  xnor
  g2717
  (
    n2791,
    n2601,
    n2666
  );


  xnor
  g2718
  (
    n2753,
    n2669,
    n2682
  );


  xnor
  g2719
  (
    n2771,
    n2675,
    n2595
  );


  xnor
  g2720
  (
    n2717,
    n2596,
    n2673
  );


  xnor
  g2721
  (
    n2792,
    n2669,
    n2681
  );


  and
  g2722
  (
    n2770,
    n2677,
    n2668
  );


  nand
  g2723
  (
    n2710,
    n2683,
    n2666
  );


  xnor
  g2724
  (
    n2729,
    n2683,
    n2674
  );


  or
  g2725
  (
    n2732,
    n2669,
    n2664
  );


  nand
  g2726
  (
    n2745,
    n2659,
    n32
  );


  or
  g2727
  (
    n2781,
    n2678,
    n2587
  );


  or
  g2728
  (
    n2693,
    n2604,
    n2580
  );


  xor
  g2729
  (
    n2778,
    n2663,
    n2678
  );


  or
  g2730
  (
    n2759,
    n2665,
    n2681
  );


  and
  g2731
  (
    KeyWire_0_3,
    n2588,
    n2676
  );


  nor
  g2732
  (
    n2712,
    n2660,
    n2603
  );


  nand
  g2733
  (
    n2756,
    n2596,
    n1973
  );


  or
  g2734
  (
    n2695,
    n2684,
    n2584
  );


  xor
  g2735
  (
    n2783,
    n2596,
    n2671
  );


  not
  g2736
  (
    n2788,
    n2601
  );


  and
  g2737
  (
    n2697,
    n2684,
    n2664
  );


  or
  g2738
  (
    n2740,
    n2682,
    n2671
  );


  nand
  g2739
  (
    n2746,
    n2598,
    n2665
  );


  or
  g2740
  (
    n2703,
    n2681,
    n2599
  );


  xor
  g2741
  (
    n2734,
    n2661,
    n2670
  );


  xor
  g2742
  (
    n2785,
    n2597,
    n2686
  );


  xor
  g2743
  (
    n2769,
    n2674,
    n2685
  );


  xor
  g2744
  (
    n2731,
    n2593,
    n2581
  );


  xnor
  g2745
  (
    n2698,
    n2598,
    n2604
  );


  xnor
  g2746
  (
    n2716,
    n1971,
    n2667
  );


  and
  g2747
  (
    n2750,
    n2668,
    n2670
  );


  and
  g2748
  (
    n2766,
    n2665,
    n2671
  );


  nor
  g2749
  (
    n2714,
    n2675,
    n2677
  );


  and
  g2750
  (
    n2780,
    n2679,
    n2670
  );


  or
  g2751
  (
    n2796,
    n2685,
    n2604
  );


  nand
  g2752
  (
    n2786,
    n2670,
    n2661
  );


  or
  g2753
  (
    n2733,
    n1972,
    n2602
  );


  and
  g2754
  (
    n2752,
    n2672,
    n2600
  );


  and
  g2755
  (
    n2758,
    n2598,
    n2667
  );


  nor
  g2756
  (
    n2748,
    n2684,
    n1972
  );


  or
  g2757
  (
    n2696,
    n2600,
    n2682
  );


  and
  g2758
  (
    n2741,
    n2676,
    n2679
  );


  nor
  g2759
  (
    n2725,
    n2667,
    n2680
  );


  nand
  g2760
  (
    n2773,
    n2597,
    n2604
  );


  nor
  g2761
  (
    n2723,
    n2672,
    n2684
  );


  xnor
  g2762
  (
    n2775,
    n2659,
    n2597
  );


  and
  g2763
  (
    n2751,
    n2576,
    n2659
  );


  xnor
  g2764
  (
    n2764,
    n2686,
    n2683
  );


  xor
  g2765
  (
    n2794,
    n2664,
    n2662
  );


  xor
  g2766
  (
    n2808,
    n2718,
    n2688,
    n2709,
    n2703
  );


  or
  g2767
  (
    n2805,
    n2739,
    n2726,
    n2734,
    n2729
  );


  xor
  g2768
  (
    n2801,
    n2733,
    n2736,
    n2735,
    n2693
  );


  xnor
  g2769
  (
    n2809,
    n2710,
    n2707,
    n2716,
    n2719
  );


  nand
  g2770
  (
    n2812,
    n2694,
    n2698,
    n2723,
    n2690
  );


  xnor
  g2771
  (
    n2799,
    n2717,
    n2720,
    n2732,
    n2699
  );


  nor
  g2772
  (
    n2806,
    n2738,
    n2737,
    n2706,
    n2701
  );


  nand
  g2773
  (
    n2804,
    n2742,
    n2712,
    n2724,
    n2728
  );


  xor
  g2774
  (
    n2800,
    n2689,
    n2687,
    n2715,
    n2705
  );


  xor
  g2775
  (
    n2802,
    n2741,
    n2695,
    n2725,
    n2704
  );


  nand
  g2776
  (
    n2807,
    n2740,
    n2714,
    n2700,
    n2730
  );


  xnor
  g2777
  (
    n2810,
    n2713,
    n2697,
    n2708,
    n2727
  );


  or
  g2778
  (
    n2811,
    n2721,
    n2722,
    n2702,
    n2731
  );


  xnor
  g2779
  (
    n2803,
    n2691,
    n2696,
    n2692,
    n2711
  );


  or
  g2780
  (
    n2827,
    n1976,
    n1973,
    n2621
  );


  xnor
  g2781
  (
    n2837,
    n2300,
    n2303,
    n2301,
    n2292
  );


  xnor
  g2782
  (
    n2825,
    n2621,
    n2571,
    n2807,
    n2809
  );


  or
  g2783
  (
    n2830,
    n2297,
    n2811,
    n2643,
    n2808
  );


  or
  g2784
  (
    n2826,
    n2810,
    n652,
    n1975,
    n2624
  );


  nor
  g2785
  (
    n2834,
    n2808,
    n2571,
    n2622,
    n2618
  );


  xnor
  g2786
  (
    n2840,
    n2812,
    n2622,
    n2517,
    n2646
  );


  xor
  g2787
  (
    n2835,
    n2810,
    n2620,
    n1975,
    n2623
  );


  or
  g2788
  (
    n2829,
    n2619,
    n2619,
    n2620,
    n2644
  );


  nor
  g2789
  (
    n2821,
    n1974,
    n2621,
    n2298,
    n2296
  );


  xor
  g2790
  (
    n2824,
    n2806,
    n2516,
    n2304,
    n2622
  );


  xnor
  g2791
  (
    n2816,
    n2646,
    n1974,
    n2809,
    n2512
  );


  or
  g2792
  (
    n2815,
    n2503,
    n1976,
    n2804,
    n2646
  );


  and
  g2793
  (
    KeyWire_0_47,
    n651,
    n2506,
    n2812,
    n2513
  );


  xor
  g2794
  (
    n2820,
    n2624,
    n2807,
    n652,
    n2623
  );


  nand
  g2795
  (
    n2819,
    n2517,
    n2803,
    n2622,
    n2811
  );


  and
  g2796
  (
    n2838,
    n2641,
    n2811,
    n2295,
    n1974
  );


  nor
  g2797
  (
    n2836,
    n2812,
    n2805,
    n2619,
    n2504
  );


  nor
  g2798
  (
    n2832,
    n1973,
    n2810,
    n2809,
    n2293
  );


  xor
  g2799
  (
    n2818,
    n2808,
    n1975,
    n2646,
    n1974
  );


  and
  g2800
  (
    n2841,
    n2507,
    n2514,
    n2618,
    n2802
  );


  xor
  g2801
  (
    n2823,
    n1975,
    n2618,
    n2517,
    n2623
  );


  nor
  g2802
  (
    n2833,
    n2302,
    n2801,
    n2515,
    n2799
  );


  xor
  g2803
  (
    n2839,
    n2619,
    n2811,
    n2510,
    n2809
  );


  nor
  g2804
  (
    n2842,
    n2509,
    n2810,
    n2505,
    n2511
  );


  or
  g2805
  (
    n2822,
    n2800,
    n2620,
    n652,
    n2623
  );


  or
  g2806
  (
    n2817,
    n1976,
    n2620,
    n1973,
    n2621
  );


  nand
  g2807
  (
    n2814,
    n2639,
    n652,
    n2508,
    n2299
  );


  xor
  g2808
  (
    n2813,
    n2640,
    n2812,
    n2808,
    n2291
  );


  xnor
  g2809
  (
    n2828,
    n2618,
    n2642,
    n2294,
    n1976
  );


  buf
  g2810
  (
    n2845,
    n2823
  );


  buf
  g2811
  (
    n2843,
    n2824
  );


  buf
  g2812
  (
    n2844,
    n2825
  );


  not
  g2813
  (
    n2846,
    n2826
  );


  not
  g2814
  (
    n2850,
    n2846
  );


  buf
  g2815
  (
    n2852,
    n2843
  );


  not
  g2816
  (
    n2853,
    n2844
  );


  not
  g2817
  (
    n2848,
    n2845
  );


  not
  g2818
  (
    n2847,
    n2846
  );


  buf
  g2819
  (
    n2849,
    n2845
  );


  not
  g2820
  (
    n2854,
    n2846
  );


  buf
  g2821
  (
    n2851,
    n2846
  );


  not
  g2822
  (
    n2855,
    n2849
  );


  buf
  g2823
  (
    n2856,
    n2848
  );


  buf
  g2824
  (
    n2860,
    n2854
  );


  buf
  g2825
  (
    n2858,
    n2852
  );


  nand
  g2826
  (
    n2859,
    n2850,
    n2853
  );


  xor
  g2827
  (
    n2857,
    n2851,
    n2847
  );


  nor
  g2828
  (
    n2861,
    n2745,
    n1978,
    n1977
  );


  xor
  g2829
  (
    n2863,
    n2750,
    n1978,
    n1977
  );


  nand
  g2830
  (
    n2867,
    n2753,
    n2752,
    n2859,
    n2855
  );


  nor
  g2831
  (
    n2864,
    n2860,
    n1979,
    n2858,
    n2749
  );


  xor
  g2832
  (
    n2866,
    n2748,
    n2746,
    n2743,
    n1979
  );


  nor
  g2833
  (
    n2865,
    n2751,
    n2860,
    n2744,
    n2857
  );


  or
  g2834
  (
    n2862,
    n1977,
    n1978,
    n2856,
    n2747
  );


  buf
  g2835
  (
    n2873,
    n2863
  );


  buf
  g2836
  (
    n2872,
    n2864
  );


  not
  g2837
  (
    n2874,
    n2865
  );


  not
  g2838
  (
    n2870,
    n2866
  );


  buf
  g2839
  (
    n2869,
    n2862
  );


  buf
  g2840
  (
    n2868,
    n2866
  );


  buf
  g2841
  (
    n2875,
    n2861
  );


  not
  g2842
  (
    n2871,
    n2866
  );


  xnor
  g2843
  (
    n2881,
    n2868,
    n2776,
    n2755,
    n2756
  );


  xor
  g2844
  (
    n2883,
    n2769,
    n2869,
    n2868,
    n2760
  );


  nand
  g2845
  (
    n2878,
    n2305,
    n2759,
    n2772,
    n2758
  );


  and
  g2846
  (
    n2886,
    n2762,
    n2773,
    n2766,
    n2779
  );


  xor
  g2847
  (
    n2880,
    n2868,
    n2770,
    n2764,
    n2783
  );


  nand
  g2848
  (
    n2876,
    n2757,
    n2869,
    n2870,
    n2754
  );


  nand
  g2849
  (
    n2882,
    n2785,
    n2781,
    n2774,
    n2782
  );


  or
  g2850
  (
    n2885,
    n2870,
    n2768,
    n2777,
    n2771
  );


  or
  g2851
  (
    n2877,
    n2869,
    n2767,
    n2784,
    n2778
  );


  xor
  g2852
  (
    n2879,
    n2763,
    n2775,
    n2870,
    n2868
  );


  nand
  g2853
  (
    n2884,
    n2765,
    n2761,
    n2869,
    n2780
  );


  buf
  g2854
  (
    n2916,
    n2879
  );


  buf
  g2855
  (
    n2918,
    n2882
  );


  buf
  g2856
  (
    n2906,
    n2794
  );


  buf
  g2857
  (
    n2917,
    n2605
  );


  buf
  g2858
  (
    n2905,
    n2883
  );


  not
  g2859
  (
    n2896,
    n2881
  );


  not
  g2860
  (
    n2893,
    n2798
  );


  not
  g2861
  (
    n2924,
    n2880
  );


  not
  g2862
  (
    n2914,
    n1980
  );


  buf
  g2863
  (
    n2889,
    n2796
  );


  not
  g2864
  (
    n2911,
    n2605
  );


  buf
  g2865
  (
    n2915,
    n1979
  );


  not
  g2866
  (
    n2921,
    n2879
  );


  not
  g2867
  (
    n2888,
    n2884
  );


  not
  g2868
  (
    n2920,
    n2798
  );


  not
  g2869
  (
    n2913,
    n2842
  );


  not
  g2870
  (
    n2890,
    n2886
  );


  not
  g2871
  (
    n2909,
    n2840
  );


  not
  g2872
  (
    n2898,
    n2786
  );


  nor
  g2873
  (
    n2903,
    n2877,
    n2396,
    n2882
  );


  nand
  g2874
  (
    n2900,
    n2879,
    n2306,
    n2791
  );


  or
  g2875
  (
    n2923,
    n2876,
    n2877,
    n2885
  );


  nor
  g2876
  (
    n2901,
    n2788,
    n2787,
    n2307,
    n2879
  );


  nor
  g2877
  (
    n2908,
    n2885,
    n2886,
    n2309,
    n2827
  );


  xnor
  g2878
  (
    n2899,
    n2829,
    n2831,
    n2835,
    n2832
  );


  xor
  g2879
  (
    n2897,
    n2886,
    n2881,
    n2797,
    n2606
  );


  xor
  g2880
  (
    KeyWire_0_52,
    n2883,
    n2798,
    n2830,
    n2792
  );


  or
  g2881
  (
    n2910,
    n2839,
    n2605,
    n2885,
    n2876
  );


  nand
  g2882
  (
    n2907,
    n2876,
    n2878,
    n2606
  );


  xnor
  g2883
  (
    n2919,
    n2795,
    n2828,
    n2878,
    n2883
  );


  xnor
  g2884
  (
    n2904,
    n2841,
    n2836,
    n2605,
    n2606
  );


  nand
  g2885
  (
    n2902,
    n2877,
    n2882,
    n2880
  );


  xnor
  g2886
  (
    n2892,
    n2834,
    n2790,
    n2884,
    n2883
  );


  nand
  g2887
  (
    n2895,
    n2798,
    n2789,
    n2876,
    n2837
  );


  xnor
  g2888
  (
    n2912,
    n2886,
    n2884,
    n2881,
    n2880
  );


  nor
  g2889
  (
    n2891,
    n2878,
    n2793,
    n2838,
    n2885
  );


  xor
  g2890
  (
    n2887,
    n2517,
    n2308,
    n2884,
    n2880
  );


  nand
  g2891
  (
    n2894,
    n2833,
    n2878,
    n2881,
    n1979
  );


  and
  g2892
  (
    n2934,
    n2889,
    n2891,
    n2892,
    n2895
  );


  or
  g2893
  (
    n2927,
    n2887,
    n2889,
    n2893
  );


  xor
  g2894
  (
    n2929,
    n2887,
    n2895,
    n2889,
    n2892
  );


  nor
  g2895
  (
    n2933,
    n2891,
    n2888,
    n2893,
    n2897
  );


  or
  g2896
  (
    n2931,
    n2896,
    n2896,
    n2891,
    n2888
  );


  and
  g2897
  (
    n2935,
    n2893,
    n2895,
    n2892,
    n2894
  );


  nand
  g2898
  (
    n2926,
    n2894,
    n2890,
    n2897,
    n2895
  );


  xnor
  g2899
  (
    n2930,
    n2896,
    n2888,
    n2892,
    n2897
  );


  xnor
  g2900
  (
    n2932,
    n2893,
    n2896,
    n2894,
    n2887
  );


  nand
  g2901
  (
    n2928,
    n2887,
    n2890,
    n2894
  );


  and
  g2902
  (
    n2925,
    n2891,
    n2890,
    n2897,
    n2888
  );


  buf
  g2903
  (
    n2936,
    n1980
  );


  buf
  g2904
  (
    n2937,
    n1980
  );


  nor
  g2905
  (
    n2938,
    n2925,
    n2926,
    n1980,
    n2927
  );


  nand
  g2906
  (
    n2941,
    n2607,
    n2608
  );


  nand
  g2907
  (
    n2942,
    n2608,
    n2938,
    n2609,
    n2607
  );


  xnor
  g2908
  (
    n2939,
    n2609,
    n2607,
    n2938,
    n2936
  );


  and
  g2909
  (
    n2940,
    n2937,
    n2607,
    n2609
  );


  not
  g2910
  (
    n2944,
    n2939
  );


  not
  g2911
  (
    n2947,
    n2941
  );


  buf
  g2912
  (
    n2943,
    n2942
  );


  buf
  g2913
  (
    n2948,
    n2942
  );


  buf
  g2914
  (
    n2946,
    n2942
  );


  not
  g2915
  (
    n2950,
    n2942
  );


  buf
  g2916
  (
    n2945,
    n2941
  );


  not
  g2917
  (
    n2949,
    n2940
  );


  not
  g2918
  (
    n2971,
    n2902
  );


  buf
  g2919
  (
    n2957,
    n2902
  );


  not
  g2920
  (
    n2964,
    n2943
  );


  buf
  g2921
  (
    n2978,
    n2871
  );


  not
  g2922
  (
    n2955,
    n2900
  );


  xnor
  g2923
  (
    n2961,
    n2871,
    n2935,
    n2930,
    n2901
  );


  and
  g2924
  (
    n2963,
    n2874,
    n2902,
    n2948,
    n2898
  );


  nor
  g2925
  (
    n2966,
    n2900,
    n2950,
    n2944,
    n2898
  );


  nand
  g2926
  (
    n2965,
    n2949,
    n2948,
    n2932,
    n2875
  );


  or
  g2927
  (
    n2958,
    n2903,
    n2944,
    n2945,
    n2905
  );


  xnor
  g2928
  (
    n2959,
    n2875,
    n2904,
    n2872
  );


  nand
  g2929
  (
    n2956,
    n2904,
    n2901,
    n2949,
    n2872
  );


  and
  g2930
  (
    n2975,
    n2904,
    n2873,
    n2899
  );


  or
  g2931
  (
    n2976,
    n2905,
    n2949,
    n2873,
    n2906
  );


  and
  g2932
  (
    n2951,
    n2658,
    n2872,
    n2903,
    n2947
  );


  or
  g2933
  (
    n2972,
    n2518,
    n2933,
    n2899,
    n2943
  );


  and
  g2934
  (
    n2968,
    n2875,
    n2928,
    n2931,
    n2871
  );


  nand
  g2935
  (
    n2954,
    n2949,
    n2946,
    n2948,
    n2658
  );


  or
  g2936
  (
    n2962,
    n2906,
    n2944,
    n2867
  );


  nand
  g2937
  (
    n2977,
    n2624,
    n2870,
    n2874,
    n2929
  );


  and
  g2938
  (
    n2982,
    n2946,
    n2950,
    n2947,
    n2906
  );


  xnor
  g2939
  (
    n2953,
    n2658,
    n2898,
    n2944,
    n2875
  );


  xnor
  g2940
  (
    n2979,
    n2943,
    n2873,
    n2945,
    n2905
  );


  nor
  g2941
  (
    n2970,
    n2907,
    n2871,
    n2873,
    n2899
  );


  and
  g2942
  (
    n2952,
    n2900,
    n2947,
    n2867,
    n2906
  );


  xnor
  g2943
  (
    n2969,
    n2947,
    n2950,
    n2518,
    n2658
  );


  nor
  g2944
  (
    n2973,
    n2518,
    n2948,
    n2943,
    n2901
  );


  or
  g2945
  (
    n2967,
    n2867,
    n2945,
    n2872,
    n2900
  );


  xor
  g2946
  (
    n2960,
    n2903,
    n2518,
    n2905,
    n2901
  );


  nor
  g2947
  (
    n2981,
    n2902,
    n2946,
    n2874
  );


  xor
  g2948
  (
    n2974,
    n2950,
    n2945,
    n2874,
    n2866
  );


  xor
  g2949
  (
    n2980,
    n2934,
    n2898,
    n2903,
    n2624
  );


  xnor
  g2950
  (
    n3013,
    n2924,
    n2981,
    n2977,
    n2922
  );


  and
  g2951
  (
    n3011,
    n2964,
    n2977,
    n2973,
    n2917
  );


  or
  g2952
  (
    n2998,
    n2979,
    n2968,
    n2921,
    n2967
  );


  and
  g2953
  (
    n2987,
    n2919,
    n2978,
    n2951,
    n2923
  );


  and
  g2954
  (
    n3004,
    n2971,
    n2907,
    n2913,
    n2914
  );


  or
  g2955
  (
    n2996,
    n2917,
    n2919,
    n2909,
    n2970
  );


  nor
  g2956
  (
    n2988,
    n2914,
    n2907,
    n2954,
    n2916
  );


  nand
  g2957
  (
    n2991,
    n2974,
    n2966,
    n2921
  );


  and
  g2958
  (
    n3001,
    n2923,
    n2976,
    n2970,
    n2977
  );


  nand
  g2959
  (
    n2985,
    n2963,
    n2955,
    n2919,
    n2914
  );


  and
  g2960
  (
    n2997,
    n2982,
    n2971,
    n2910,
    n2973
  );


  nand
  g2961
  (
    n3016,
    n2965,
    n2965,
    n2920,
    n2966
  );


  xnor
  g2962
  (
    n3018,
    n2980,
    n2962,
    n2975,
    n2978
  );


  xnor
  g2963
  (
    n2999,
    n2964,
    n2918,
    n2967,
    n2916
  );


  nand
  g2964
  (
    KeyWire_0_27,
    n2965,
    n2972,
    n2974,
    n2968
  );


  xnor
  g2965
  (
    n2986,
    n2968,
    n2923,
    n2913,
    n2953
  );


  xnor
  g2966
  (
    n2995,
    n2974,
    n2915,
    n2970,
    n2961
  );


  xor
  g2967
  (
    n3003,
    n2971,
    n2911,
    n2917,
    n2921
  );


  nand
  g2968
  (
    n3021,
    n2975,
    n2974,
    n2972,
    n2916
  );


  nor
  g2969
  (
    n3014,
    n2959,
    n2979,
    n2910,
    n2915
  );


  xor
  g2970
  (
    n2992,
    n2924,
    n2907,
    n2981,
    n2982
  );


  and
  g2971
  (
    n3008,
    n2969,
    n2977,
    n2914,
    n2918
  );


  or
  g2972
  (
    n3019,
    n2909,
    n2972,
    n2966,
    n2912
  );


  xnor
  g2973
  (
    n2983,
    n2964,
    n2910,
    n2913,
    n2915
  );


  or
  g2974
  (
    n3002,
    n2972,
    n2912,
    n2980,
    n2969
  );


  nor
  g2975
  (
    n3015,
    n2917,
    n2975,
    n2908,
    n2976
  );


  nand
  g2976
  (
    n3012,
    n2921,
    n2919,
    n2969,
    n2960
  );


  nand
  g2977
  (
    n3010,
    n2967,
    n2923,
    n2908,
    n2975
  );


  xnor
  g2978
  (
    n2994,
    n2909,
    n2976,
    n2912,
    n2981
  );


  nand
  g2979
  (
    n2989,
    n2969,
    n2922,
    n2958,
    n2924
  );


  xor
  g2980
  (
    n3007,
    n2973,
    n2911,
    n2908,
    n2968
  );


  and
  g2981
  (
    n3022,
    n2982,
    n2956,
    n2979,
    n2967
  );


  and
  g2982
  (
    n3017,
    n2965,
    n2970,
    n2978
  );


  or
  g2983
  (
    n3006,
    n2920,
    n2920,
    n2913,
    n2976
  );


  nand
  g2984
  (
    n3020,
    n2920,
    n2922,
    n2952,
    n2982
  );


  nor
  g2985
  (
    KeyWire_0_46,
    n2909,
    n2908,
    n2957,
    n2911
  );


  nand
  g2986
  (
    n2984,
    n2979,
    n2964,
    n2980
  );


  xor
  g2987
  (
    n2990,
    n2924,
    n2922,
    n2910,
    n2918
  );


  or
  g2988
  (
    n2993,
    n2973,
    n2916,
    n2911,
    n2918
  );


  nor
  g2989
  (
    n3005,
    n2981,
    n2971,
    n2912,
    n2915
  );


  and
  g2990
  (
    n3030,
    n3002,
    n2983,
    n3014,
    n3000
  );


  or
  g2991
  (
    n3027,
    n3010,
    n3006,
    n3011,
    n2985
  );


  nand
  g2992
  (
    n3026,
    n3007,
    n2994,
    n3015,
    n2992
  );


  nor
  g2993
  (
    n3029,
    n3020,
    n2984,
    n3016,
    n2991
  );


  nor
  g2994
  (
    n3028,
    n3005,
    n2993,
    n2995,
    n3021
  );


  xor
  g2995
  (
    n3025,
    n3018,
    n2998,
    n2997,
    n2999
  );


  nor
  g2996
  (
    n3024,
    n2986,
    n2996,
    n2988,
    n3004
  );


  xor
  g2997
  (
    n3023,
    n3003,
    n3009,
    n2987,
    n3017
  );


  or
  g2998
  (
    n3032,
    n3019,
    n2990,
    n3022,
    n3001
  );


  nand
  g2999
  (
    n3031,
    n3013,
    n3008,
    n3012,
    n2989
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1454,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1882,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n2363,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n2706,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n2120,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n554,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n741,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1840,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n2329,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n2234,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n429,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1312,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n445,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n702,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1814,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1618,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n322,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n922,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n2798,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n783,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1389,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1425,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n498,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n2404,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1465,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n1910,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n255,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n3009,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n1356,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1991,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n830,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n665,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n863,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n634,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n2726,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n720,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1196,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n325,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n133,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n937,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n1897,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n1752,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n35,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n447,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n70,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n2663,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n3000,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n2831,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1017,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n2204,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n397,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n1219,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n2922,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n2310,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n837,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n1594,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n2463,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n541,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n2013,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n514,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n2112,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n793,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n798,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n1702,
    KeyNOTWire_0_63
  );


endmodule

