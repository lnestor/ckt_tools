// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_103 written by SynthGen on 2021/04/05 11:08:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_103 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1024, n1017, n1020, n1012, n1008, n1005, n1025, n1016,
 n1007, n1027, n1011, n1026, n1031, n1023, n1003, n1014,
 n1021, n1019, n1009, n1028, n1013, n1006, n1001, n1002,
 n1015, n1022, n1032, n1018, n1004, n1029, n1010, n1030);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1024, n1017, n1020, n1012, n1008, n1005, n1025, n1016,
 n1007, n1027, n1011, n1026, n1031, n1023, n1003, n1014,
 n1021, n1019, n1009, n1028, n1013, n1006, n1001, n1002,
 n1015, n1022, n1032, n1018, n1004, n1029, n1010, n1030;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000;

not  g0 (n145, n6);
not  g1 (n34, n16);
not  g2 (n160, n23);
not  g3 (n157, n24);
buf  g4 (n131, n10);
not  g5 (n147, n17);
not  g6 (n45, n22);
not  g7 (n59, n6);
not  g8 (n117, n11);
buf  g9 (n62, n4);
not  g10 (n115, n4);
not  g11 (n119, n26);
buf  g12 (n77, n9);
buf  g13 (n42, n32);
not  g14 (n100, n32);
buf  g15 (n54, n3);
not  g16 (n101, n27);
buf  g17 (n57, n13);
not  g18 (n134, n31);
not  g19 (n116, n1);
buf  g20 (n123, n8);
buf  g21 (n105, n26);
buf  g22 (n152, n6);
not  g23 (n83, n9);
buf  g24 (n149, n3);
not  g25 (n60, n15);
buf  g26 (n78, n18);
buf  g27 (n108, n2);
buf  g28 (n88, n4);
buf  g29 (n70, n3);
buf  g30 (n144, n14);
buf  g31 (n67, n28);
buf  g32 (n53, n11);
buf  g33 (n76, n2);
not  g34 (n107, n12);
not  g35 (n95, n25);
buf  g36 (n151, n28);
not  g37 (n73, n15);
not  g38 (n143, n2);
not  g39 (n137, n31);
buf  g40 (n75, n8);
buf  g41 (n159, n16);
not  g42 (n154, n5);
not  g43 (n85, n7);
not  g44 (n113, n30);
buf  g45 (n132, n26);
not  g46 (n71, n8);
buf  g47 (n94, n23);
not  g48 (n81, n6);
buf  g49 (n99, n30);
buf  g50 (n40, n21);
buf  g51 (n148, n29);
not  g52 (n66, n27);
buf  g53 (n140, n30);
buf  g54 (n47, n22);
not  g55 (n96, n20);
buf  g56 (n43, n21);
not  g57 (n102, n9);
not  g58 (n86, n32);
buf  g59 (n139, n16);
buf  g60 (n61, n22);
not  g61 (n52, n22);
buf  g62 (n38, n5);
not  g63 (n93, n5);
not  g64 (n121, n31);
not  g65 (n36, n28);
buf  g66 (n135, n25);
buf  g67 (n138, n24);
not  g68 (n82, n20);
not  g69 (n87, n12);
buf  g70 (n124, n5);
buf  g71 (n63, n21);
not  g72 (n158, n14);
not  g73 (n58, n19);
not  g74 (n39, n15);
buf  g75 (n103, n13);
buf  g76 (n110, n27);
buf  g77 (n129, n11);
not  g78 (n79, n17);
not  g79 (n56, n19);
not  g80 (n48, n17);
not  g81 (n127, n13);
buf  g82 (n114, n2);
buf  g83 (n155, n25);
buf  g84 (n89, n8);
not  g85 (n128, n1);
not  g86 (n133, n15);
not  g87 (n122, n13);
not  g88 (n141, n9);
not  g89 (n118, n12);
buf  g90 (n55, n19);
buf  g91 (n37, n10);
buf  g92 (n35, n31);
buf  g93 (n156, n28);
buf  g94 (n92, n1);
not  g95 (n64, n23);
not  g96 (n65, n16);
buf  g97 (n84, n24);
buf  g98 (n130, n27);
buf  g99 (n142, n12);
buf  g100 (n146, n18);
not  g101 (n44, n14);
buf  g102 (n72, n18);
buf  g103 (n90, n7);
buf  g104 (n91, n7);
not  g105 (n126, n29);
buf  g106 (n150, n26);
not  g107 (n112, n1);
buf  g108 (n68, n23);
buf  g109 (n33, n21);
not  g110 (n120, n18);
not  g111 (n74, n20);
buf  g112 (n51, n19);
buf  g113 (n97, n20);
buf  g114 (n46, n11);
not  g115 (n98, n30);
not  g116 (n111, n4);
not  g117 (n109, n10);
not  g118 (n69, n25);
buf  g119 (n80, n29);
buf  g120 (n125, n17);
buf  g121 (n41, n32);
not  g122 (n106, n7);
not  g123 (n153, n10);
not  g124 (n104, n14);
buf  g125 (n49, n3);
buf  g126 (n136, n29);
not  g127 (n50, n24);
not  g128 (n294, n69);
buf  g129 (n394, n75);
not  g130 (n419, n112);
buf  g131 (n300, n86);
buf  g132 (n386, n125);
buf  g133 (n440, n112);
buf  g134 (n485, n54);
buf  g135 (n420, n78);
not  g136 (n410, n120);
not  g137 (n208, n55);
buf  g138 (n472, n44);
buf  g139 (n436, n85);
not  g140 (n296, n85);
buf  g141 (n343, n118);
buf  g142 (n185, n54);
buf  g143 (n166, n77);
buf  g144 (n198, n123);
not  g145 (n334, n70);
not  g146 (n355, n69);
not  g147 (n243, n74);
buf  g148 (n517, n50);
buf  g149 (n191, n60);
not  g150 (n525, n60);
buf  g151 (n324, n81);
not  g152 (n384, n105);
buf  g153 (n400, n52);
buf  g154 (n427, n40);
buf  g155 (n459, n93);
not  g156 (n426, n105);
buf  g157 (n197, n71);
buf  g158 (n399, n112);
buf  g159 (n402, n35);
buf  g160 (n524, n34);
buf  g161 (n377, n74);
not  g162 (n266, n126);
buf  g163 (n206, n51);
buf  g164 (n240, n104);
buf  g165 (n454, n44);
buf  g166 (n391, n83);
not  g167 (n409, n88);
not  g168 (n477, n39);
not  g169 (n467, n80);
not  g170 (n456, n94);
not  g171 (n278, n83);
not  g172 (n265, n64);
buf  g173 (n232, n80);
not  g174 (n313, n73);
not  g175 (n257, n68);
buf  g176 (n530, n102);
not  g177 (n230, n90);
not  g178 (n496, n39);
not  g179 (n482, n68);
not  g180 (n203, n108);
buf  g181 (n209, n109);
not  g182 (n455, n45);
not  g183 (n210, n53);
buf  g184 (n255, n86);
buf  g185 (n319, n47);
not  g186 (n219, n120);
not  g187 (n483, n50);
not  g188 (n336, n86);
not  g189 (n171, n88);
not  g190 (n441, n79);
buf  g191 (n533, n51);
buf  g192 (n186, n88);
buf  g193 (n487, n37);
not  g194 (n228, n82);
not  g195 (n292, n87);
not  g196 (n174, n103);
not  g197 (n451, n81);
not  g198 (n452, n107);
buf  g199 (n453, n66);
not  g200 (n225, n63);
not  g201 (n463, n118);
buf  g202 (n307, n51);
buf  g203 (n254, n76);
buf  g204 (n505, n117);
buf  g205 (n393, n47);
buf  g206 (n162, n56);
not  g207 (n489, n114);
not  g208 (n405, n116);
not  g209 (n207, n111);
buf  g210 (n433, n54);
buf  g211 (n305, n107);
not  g212 (n301, n43);
buf  g213 (n202, n115);
not  g214 (n424, n52);
not  g215 (n273, n95);
buf  g216 (n371, n71);
not  g217 (n217, n87);
not  g218 (n309, n75);
buf  g219 (n416, n121);
buf  g220 (n182, n91);
buf  g221 (n249, n103);
buf  g222 (n381, n96);
buf  g223 (n318, n50);
not  g224 (n513, n111);
not  g225 (n490, n34);
buf  g226 (n281, n58);
buf  g227 (n368, n110);
not  g228 (n448, n55);
buf  g229 (n346, n97);
not  g230 (n479, n104);
buf  g231 (n168, n105);
buf  g232 (n231, n55);
buf  g233 (n508, n47);
not  g234 (n260, n36);
buf  g235 (n366, n114);
not  g236 (n196, n49);
buf  g237 (n442, n48);
buf  g238 (n507, n46);
buf  g239 (n434, n110);
buf  g240 (n311, n108);
buf  g241 (n261, n59);
not  g242 (n302, n71);
not  g243 (n241, n50);
buf  g244 (n474, n92);
buf  g245 (n491, n38);
buf  g246 (n326, n73);
not  g247 (n445, n61);
not  g248 (n526, n38);
buf  g249 (n187, n54);
not  g250 (n520, n105);
not  g251 (n527, n106);
buf  g252 (n439, n62);
buf  g253 (n329, n120);
not  g254 (n389, n123);
not  g255 (n361, n120);
buf  g256 (n413, n41);
buf  g257 (n415, n70);
buf  g258 (n330, n97);
buf  g259 (n365, n95);
buf  g260 (n164, n121);
not  g261 (n481, n124);
not  g262 (n170, n34);
buf  g263 (n169, n41);
not  g264 (n447, n63);
buf  g265 (n475, n40);
buf  g266 (n519, n77);
buf  g267 (n175, n108);
buf  g268 (n308, n84);
not  g269 (n165, n61);
not  g270 (n180, n119);
buf  g271 (n177, n68);
buf  g272 (n529, n89);
buf  g273 (n504, n96);
not  g274 (n316, n113);
buf  g275 (n204, n84);
not  g276 (n473, n35);
buf  g277 (n417, n72);
not  g278 (n512, n36);
not  g279 (n471, n64);
not  g280 (n468, n117);
not  g281 (n276, n65);
buf  g282 (n268, n35);
not  g283 (n431, n75);
not  g284 (n235, n98);
buf  g285 (n347, n69);
buf  g286 (n429, n103);
buf  g287 (n299, n42);
buf  g288 (n214, n125);
buf  g289 (n398, n56);
not  g290 (n488, n109);
not  g291 (n353, n107);
buf  g292 (n248, n80);
buf  g293 (n161, n71);
not  g294 (n205, n125);
buf  g295 (n221, n80);
buf  g296 (n360, n91);
buf  g297 (n211, n40);
buf  g298 (n279, n59);
buf  g299 (n460, n95);
not  g300 (n335, n33);
buf  g301 (n457, n94);
buf  g302 (n163, n100);
not  g303 (n262, n63);
not  g304 (n523, n122);
not  g305 (n500, n45);
not  g306 (n181, n96);
not  g307 (n184, n124);
not  g308 (n531, n83);
not  g309 (n291, n92);
buf  g310 (n282, n97);
buf  g311 (n341, n113);
not  g312 (n224, n123);
buf  g313 (n369, n42);
buf  g314 (n303, n53);
not  g315 (n408, n62);
buf  g316 (n338, n58);
buf  g317 (n325, n42);
buf  g318 (n256, n106);
not  g319 (n193, n61);
buf  g320 (n277, n35);
not  g321 (n321, n81);
buf  g322 (n480, n116);
not  g323 (n484, n78);
buf  g324 (n342, n58);
not  g325 (n345, n39);
not  g326 (n317, n45);
buf  g327 (n287, n73);
not  g328 (n444, n49);
not  g329 (n357, n109);
buf  g330 (n465, n116);
not  g331 (n229, n74);
buf  g332 (n476, n99);
buf  g333 (n242, n51);
buf  g334 (n337, n45);
buf  g335 (n446, n79);
not  g336 (n437, n76);
buf  g337 (n315, n37);
buf  g338 (n364, n91);
not  g339 (n327, n101);
not  g340 (n497, n101);
not  g341 (n449, n56);
buf  g342 (n323, n100);
buf  g343 (n173, n46);
not  g344 (n201, n84);
buf  g345 (n199, n81);
buf  g346 (n502, n76);
buf  g347 (n397, n44);
buf  g348 (n227, n94);
not  g349 (n438, n92);
buf  g350 (n322, n79);
buf  g351 (n295, n62);
not  g352 (n352, n48);
not  g353 (n430, n66);
buf  g354 (n470, n59);
buf  g355 (n403, n70);
buf  g356 (n216, n98);
not  g357 (n274, n75);
buf  g358 (n469, n118);
not  g359 (n250, n85);
not  g360 (n267, n92);
not  g361 (n306, n119);
not  g362 (n220, n82);
buf  g363 (n414, n83);
not  g364 (n379, n43);
not  g365 (n226, n115);
buf  g366 (n354, n62);
not  g367 (n239, n72);
not  g368 (n466, n111);
buf  g369 (n298, n73);
buf  g370 (n392, n104);
buf  g371 (n189, n78);
buf  g372 (n516, n47);
not  g373 (n461, n67);
not  g374 (n501, n112);
buf  g375 (n304, n41);
buf  g376 (n290, n122);
buf  g377 (n506, n102);
not  g378 (n511, n123);
not  g379 (n222, n43);
not  g380 (n258, n98);
buf  g381 (n494, n91);
buf  g382 (n532, n39);
buf  g383 (n200, n90);
not  g384 (n422, n61);
not  g385 (n331, n33);
not  g386 (n167, n38);
not  g387 (n358, n57);
not  g388 (n339, n113);
buf  g389 (n406, n84);
not  g390 (n236, n121);
not  g391 (n458, n102);
not  g392 (n275, n100);
not  g393 (n411, n89);
not  g394 (n396, n49);
buf  g395 (n432, n57);
not  g396 (n362, n89);
buf  g397 (n499, n85);
not  g398 (n401, n98);
not  g399 (n218, n41);
not  g400 (n518, n57);
buf  g401 (n376, n34);
buf  g402 (n493, n33);
not  g403 (n348, n65);
buf  g404 (n359, n117);
buf  g405 (n374, n82);
not  g406 (n350, n101);
not  g407 (n510, n53);
buf  g408 (n450, n67);
not  g409 (n522, n63);
buf  g410 (n195, n104);
buf  g411 (n407, n64);
buf  g412 (n314, n72);
not  g413 (n503, n36);
not  g414 (n367, n90);
buf  g415 (n247, n118);
buf  g416 (n344, n76);
buf  g417 (n190, n37);
buf  g418 (n269, n67);
not  g419 (n382, n113);
not  g420 (n509, n124);
buf  g421 (n237, n43);
not  g422 (n478, n52);
not  g423 (n443, n89);
buf  g424 (n349, n88);
not  g425 (n213, n114);
not  g426 (n263, n101);
buf  g427 (n312, n102);
not  g428 (n390, n111);
buf  g429 (n244, n56);
not  g430 (n515, n79);
not  g431 (n223, n59);
buf  g432 (n259, n49);
buf  g433 (n245, n36);
buf  g434 (n412, n93);
not  g435 (n383, n93);
buf  g436 (n428, n97);
not  g437 (n387, n99);
not  g438 (n351, n38);
buf  g439 (n404, n106);
not  g440 (n283, n99);
buf  g441 (n514, n107);
buf  g442 (n238, n60);
buf  g443 (n425, n86);
buf  g444 (n297, n60);
not  g445 (n320, n55);
not  g446 (n192, n33);
buf  g447 (n421, n53);
buf  g448 (n233, n65);
buf  g449 (n464, n66);
buf  g450 (n418, n70);
buf  g451 (n179, n67);
buf  g452 (n264, n69);
buf  g453 (n176, n46);
not  g454 (n521, n100);
buf  g455 (n378, n64);
not  g456 (n251, n65);
buf  g457 (n486, n99);
not  g458 (n172, n77);
not  g459 (n373, n124);
buf  g460 (n272, n48);
not  g461 (n385, n58);
buf  g462 (n286, n93);
not  g463 (n310, n74);
not  g464 (n188, n37);
not  g465 (n375, n96);
buf  g466 (n372, n78);
not  g467 (n356, n115);
buf  g468 (n332, n122);
not  g469 (n212, n77);
not  g470 (n183, n109);
not  g471 (n328, n82);
buf  g472 (n462, n103);
not  g473 (n340, n72);
not  g474 (n423, n119);
buf  g475 (n495, n90);
buf  g476 (n363, n42);
buf  g477 (n252, n115);
buf  g478 (n498, n108);
not  g479 (n388, n48);
buf  g480 (n370, n95);
buf  g481 (n246, n52);
not  g482 (n253, n46);
not  g483 (n178, n68);
buf  g484 (n215, n121);
not  g485 (n395, n40);
not  g486 (n270, n114);
not  g487 (n380, n119);
buf  g488 (n280, n94);
not  g489 (n293, n117);
buf  g490 (n271, n110);
buf  g491 (n288, n106);
buf  g492 (n234, n125);
not  g493 (n492, n44);
not  g494 (n289, n110);
not  g495 (n528, n87);
not  g496 (n194, n87);
not  g497 (n435, n57);
buf  g498 (n285, n116);
buf  g499 (n333, n122);
not  g500 (n284, n66);
not  g501 (n541, n164);
buf  g502 (n540, n167);
not  g503 (n537, n168);
buf  g504 (n538, n166);
not  g505 (n539, n163);
buf  g506 (n543, n161);
buf  g507 (n546, n161);
not  g508 (n535, n162);
buf  g509 (n542, n165);
not  g510 (n544, n164);
buf  g511 (n547, n162);
not  g512 (n536, n167);
not  g513 (n545, n163);
not  g514 (n534, n165);
buf  g515 (n548, n166);
buf  g516 (n567, n538);
not  g517 (n556, n174);
buf  g518 (n580, n548);
not  g519 (n561, n182);
not  g520 (n557, n169);
not  g521 (n563, n179);
not  g522 (n569, n176);
buf  g523 (n553, n175);
not  g524 (n559, n172);
buf  g525 (n554, n180);
not  g526 (n555, n547);
not  g527 (n571, n537);
not  g528 (n570, n548);
not  g529 (n565, n534);
not  g530 (n562, n540);
not  g531 (n578, n543);
buf  g532 (n551, n178);
buf  g533 (n568, n539);
buf  g534 (n566, n176);
not  g535 (n579, n539);
nor  g536 (n573, n538, n544);
xnor g537 (n576, n177, n171);
nor  g538 (n577, n179, n548, n182, n541);
nand g539 (n549, n536, n543, n546, n169);
and  g540 (n572, n168, n535, n546, n183);
xnor g541 (n564, n545, n175, n180, n542);
nand g542 (n550, n540, n171, n184, n534);
xor  g543 (n558, n173, n542, n181, n537);
and  g544 (n574, n170, n544, n545, n173);
nor  g545 (n560, n178, n174, n172, n177);
xnor g546 (n552, n183, n170, n541, n547);
xor  g547 (n575, n535, n181, n547, n536);
not  g548 (n581, n159);
xnor g549 (n617, n552, n129, n155);
or   g550 (n599, n550, n142, n137, n575);
nand g551 (n628, n566, n158, n141);
nand g552 (n586, n556, n128, n155, n159);
and  g553 (n615, n566, n577, n155, n130);
xnor g554 (n601, n131, n156, n569, n149);
or   g555 (n610, n127, n144, n568, n135);
and  g556 (n627, n571, n159, n134, n140);
or   g557 (n597, n576, n137, n160, n141);
xor  g558 (n611, n148, n145, n144, n132);
nor  g559 (n593, n553, n145, n160, n127);
nand g560 (n607, n568, n138, n145, n126);
and  g561 (n620, n148, n147, n570, n150);
xor  g562 (n624, n156, n128, n126, n555);
or   g563 (n591, n154, n157, n142, n143);
nand g564 (n588, n129, n153, n133, n132);
xor  g565 (n613, n146, n561, n152, n136);
xnor g566 (n606, n142, n133, n129, n562);
xnor g567 (n623, n151, n141, n549, n564);
xor  g568 (n585, n133, n560, n134, n137);
xnor g569 (n582, n572, n158, n580, n154);
xor  g570 (n618, n574, n138, n139, n145);
and  g571 (n603, n141, n140, n142, n557);
nor  g572 (n609, n136, n134, n135, n578);
xnor g573 (n600, n577, n148, n132, n147);
xnor g574 (n592, n149, n127, n152, n130);
and  g575 (n604, n128, n576, n151, n156);
nor  g576 (n583, n150, n155, n580, n579);
xnor g577 (n608, n135, n565, n156, n184);
xor  g578 (n621, n154, n157, n132, n128);
nand g579 (n612, n143, n554, n579, n152);
or   g580 (n622, n149, n139, n151, n129);
xnor g581 (n614, n127, n147, n572, n139);
xnor g582 (n598, n570, n131, n159, n573);
nor  g583 (n596, n138, n146, n126, n143);
or   g584 (n626, n569, n144, n150, n130);
nand g585 (n594, n136, n157, n151, n160);
and  g586 (n616, n563, n130, n551, n131);
nand g587 (n590, n148, n137, n135, n147);
nand g588 (n625, n140, n157, n153, n138);
xor  g589 (n602, n160, n149, n131, n559);
or   g590 (n584, n152, n140, n578, n136);
or   g591 (n605, n139, n158, n571, n146);
xnor g592 (n589, n153, n134, n150, n567);
xnor g593 (n595, n153, n133, n573, n558);
nand g594 (n587, n567, n574, n143, n575);
xor  g595 (n619, n144, n146, n154, n565);
xnor g596 (n769, n246, n428, n285, n279);
or   g597 (n807, n249, n304, n417, n289);
nand g598 (n638, n618, n430, n582, n213);
xnor g599 (n698, n584, n315, n330, n269);
xnor g600 (n675, n380, n276, n364, n351);
and  g601 (n810, n235, n411, n372, n207);
nand g602 (n713, n607, n367, n281, n604);
xnor g603 (n781, n602, n616, n322, n598);
nor  g604 (n652, n432, n325, n233, n625);
xor  g605 (n804, n311, n605, n410, n398);
xnor g606 (n635, n384, n241, n599, n219);
xor  g607 (n703, n366, n308, n397, n215);
and  g608 (n637, n365, n396, n298, n336);
nand g609 (n738, n286, n323, n599, n400);
xor  g610 (n646, n185, n599, n387, n275);
xor  g611 (n733, n618, n276, n262, n408);
and  g612 (n661, n369, n423, n601, n387);
nand g613 (n654, n370, n583, n622, n595);
or   g614 (n741, n194, n215, n195, n427);
xor  g615 (n672, n399, n396, n258, n381);
nand g616 (n650, n360, n626, n384, n590);
nand g617 (n789, n366, n610, n585, n321);
nor  g618 (n792, n415, n204, n342, n594);
nor  g619 (n712, n244, n353, n200, n434);
nand g620 (n772, n191, n597, n598, n217);
or   g621 (n734, n279, n299, n600, n388);
and  g622 (n724, n375, n585, n384, n425);
xor  g623 (n719, n257, n186, n342, n359);
nand g624 (n693, n374, n592, n431, n195);
or   g625 (n641, n381, n583, n267, n404);
and  g626 (n817, n592, n240, n190, n365);
and  g627 (n697, n604, n373, n418, n627);
and  g628 (n629, n412, n613, n312, n232);
and  g629 (n707, n263, n229, n372, n391);
and  g630 (n680, n583, n305, n319, n626);
nand g631 (n720, n619, n264, n205, n227);
and  g632 (n791, n380, n308, n406, n203);
nand g633 (n717, n303, n602, n407, n283);
nand g634 (n784, n258, n600, n259, n589);
nand g635 (n808, n313, n188, n289, n285);
nand g636 (n761, n290, n298, n251, n382);
xnor g637 (n766, n593, n619, n340, n364);
or   g638 (n640, n601, n352, n241, n323);
xor  g639 (n630, n286, n620, n347, n189);
nor  g640 (n705, n331, n593, n261, n390);
xor  g641 (n658, n603, n261, n226, n628);
or   g642 (n753, n204, n584, n231, n617);
xnor g643 (n800, n604, n292, n376, n277);
xnor g644 (n685, n387, n350, n347, n222);
nand g645 (n806, n581, n628, n357, n615);
xor  g646 (n731, n344, n349, n332, n328);
nor  g647 (n696, n220, n314, n300, n252);
or   g648 (n775, n586, n595, n296, n307);
nand g649 (n732, n605, n398, n217, n371);
xor  g650 (n748, n197, n612, n594, n221);
nor  g651 (n760, n366, n362, n211, n301);
or   g652 (n715, n233, n268, n248, n198);
and  g653 (n673, n250, n414, n325, n318);
nor  g654 (n723, n212, n346, n419, n402);
and  g655 (n657, n412, n196, n343, n424);
or   g656 (n721, n304, n327, n382, n256);
or   g657 (n643, n311, n202, n406, n234);
nor  g658 (n710, n411, n297, n612, n310);
nand g659 (n659, n592, n377, n238, n405);
nor  g660 (n754, n395, n380, n605, n581);
nor  g661 (n815, n602, n627, n225, n592);
xnor g662 (n737, n385, n274, n346, n378);
and  g663 (n729, n374, n389, n350, n257);
nor  g664 (n633, n255, n609, n269, n359);
nor  g665 (n662, n400, n209, n392, n388);
xor  g666 (n704, n418, n191, n622, n400);
nor  g667 (n681, n406, n272, n337, n609);
nand g668 (n780, n596, n369, n589, n317);
nor  g669 (n726, n193, n405, n208, n293);
xnor g670 (n798, n256, n377, n619, n620);
and  g671 (n758, n421, n322, n231, n288);
nand g672 (n634, n588, n420, n303, n423);
xnor g673 (n777, n266, n333, n409, n582);
nor  g674 (n788, n615, n302, n608, n382);
xnor g675 (n639, n392, n416, n225, n355);
or   g676 (n631, n420, n594, n338, n324);
nor  g677 (n664, n607, n265, n414, n356);
and  g678 (n799, n287, n616, n393, n606);
xor  g679 (n674, n343, n432, n429, n365);
and  g680 (n790, n388, n613, n394, n620);
or   g681 (n725, n430, n309, n591, n194);
xnor g682 (n689, n584, n598, n372, n317);
nor  g683 (n809, n604, n273, n216, n211);
or   g684 (n677, n422, n236, n377, n265);
nand g685 (n679, n198, n358, n433, n383);
nand g686 (n711, n368, n610, n586, n402);
nor  g687 (n779, n354, n618, n282, n208);
and  g688 (n814, n209, n623, n610, n606);
or   g689 (n805, n207, n294, n245, n266);
or   g690 (n671, n228, n214, n426, n353);
and  g691 (n682, n363, n316, n603, n282);
nor  g692 (n651, n415, n627, n288, n407);
xor  g693 (n813, n583, n228, n597, n186);
xnor g694 (n770, n232, n330, n428, n414);
xnor g695 (n797, n433, n200, n278, n367);
nand g696 (n655, n223, n354, n416, n375);
and  g697 (n660, n373, n326, n584, n293);
and  g698 (n776, n267, n609, n251, n332);
or   g699 (n708, n335, n612, n352, n296);
nand g700 (n714, n242, n421, n596, n606);
or   g701 (n632, n320, n320, n334, n329);
nor  g702 (n668, n611, n341, n614, n393);
xor  g703 (n676, n386, n397, n588, n624);
nand g704 (n745, n621, n626, n284, n402);
nor  g705 (n653, n278, n187, n290, n299);
nor  g706 (n678, n240, n237, n202, n341);
nand g707 (n752, n610, n585, n606, n259);
and  g708 (n730, n219, n218, n328, n415);
nor  g709 (n644, n254, n313, n431, n335);
xnor g710 (n787, n339, n295, n268, n427);
xor  g711 (n667, n595, n603, n427, n401);
and  g712 (n706, n395, n601, n401, n591);
nor  g713 (n656, n331, n622, n260, n394);
xor  g714 (n716, n242, n221, n581, n397);
nor  g715 (n783, n621, n376, n389, n197);
xor  g716 (n767, n609, n375, n587, n403);
nor  g717 (n666, n612, n611, n422, n613);
nor  g718 (n701, n420, n588, n607, n625);
or   g719 (n649, n199, n424, n274, n615);
and  g720 (n751, n410, n391, n411, n602);
nor  g721 (n687, n409, n199, n196, n315);
and  g722 (n749, n409, n374, n404, n306);
xor  g723 (n768, n300, n270, n364, n206);
nand g724 (n816, n255, n595, n403, n370);
xor  g725 (n794, n248, n359, n246, n422);
nor  g726 (n759, n203, n367, n608, n403);
nand g727 (n718, n386, n318, n433, n614);
xor  g728 (n819, n376, n430, n625, n390);
xnor g729 (n699, n624, n357, n312, n192);
and  g730 (n728, n361, n247, n249, n244);
and  g731 (n636, n291, n434, n586, n316);
or   g732 (n691, n396, n226, n611, n287);
xnor g733 (n818, n368, n608, n336, n213);
xnor g734 (n688, n424, n253, n413, n306);
nor  g735 (n756, n363, n271, n264, n398);
nor  g736 (n695, n239, n192, n385, n338);
and  g737 (n742, n210, n379, n227, n371);
nand g738 (n743, n250, n408, n597, n613);
xor  g739 (n744, n628, n624, n247, n205);
nand g740 (n771, n294, n302, n324, n627);
xnor g741 (n642, n238, n301, n356, n587);
nand g742 (n665, n389, n607, n224, n235);
xnor g743 (n801, n337, n399, n410, n412);
xnor g744 (n750, n307, n230, n617, n297);
nand g745 (n663, n596, n582, n429, n349);
nor  g746 (n786, n426, n362, n358, n621);
and  g747 (n692, n236, n345, n419, n416);
nand g748 (n647, n405, n587, n362, n378);
xnor g749 (n709, n624, n622, n214, n587);
xnor g750 (n782, n329, n421, n189, n237);
and  g751 (n735, n425, n590, n361, n355);
or   g752 (n785, n601, n585, n253, n210);
xor  g753 (n736, n586, n385, n188, n399);
xnor g754 (n702, n611, n270, n190, n383);
or   g755 (n796, n185, n392, n426, n321);
nand g756 (n669, n419, n619, n348, n394);
nor  g757 (n802, n272, n277, n594, n361);
xnor g758 (n757, n623, n327, n284, n617);
xor  g759 (n765, n326, n234, n360, n589);
or   g760 (n811, n423, n391, n281, n222);
nand g761 (n694, n379, n310, n344, n616);
nor  g762 (n773, n589, n223, n368, n252);
xor  g763 (n727, n407, n254, n360, n401);
nand g764 (n739, n614, n220, n620, n370);
xnor g765 (n755, n418, n597, n334, n340);
xor  g766 (n686, n600, n305, n617, n603);
nor  g767 (n700, n333, n596, n363, n588);
nand g768 (n763, n206, n230, n605, n386);
xnor g769 (n803, n431, n623, n591, n593);
and  g770 (n684, n383, n201, n291, n273);
nor  g771 (n670, n309, n615, n351, n339);
nand g772 (n820, n600, n239, n187, n413);
or   g773 (n648, n369, n280, n582, n621);
nor  g774 (n762, n245, n590, n432, n358);
or   g775 (n778, n314, n243, n260, n425);
nor  g776 (n690, n608, n591, n614, n628);
and  g777 (n812, n345, n373, n283, n381);
xnor g778 (n747, n417, n201, n395, n616);
nor  g779 (n795, n393, n229, n428, n275);
xnor g780 (n645, n271, n348, n599, n408);
or   g781 (n774, n263, n593, n598, n378);
and  g782 (n764, n404, n623, n371, n581);
or   g783 (n793, n379, n417, n413, n390);
nor  g784 (n746, n280, n216, n590, n224);
and  g785 (n683, n429, n212, n292, n625);
nand g786 (n740, n243, n295, n218, n618);
nand g787 (n722, n626, n262, n319, n193);
nor  g788 (n889, n450, n446, n680);
xnor g789 (n896, n751, n694, n723, n481);
and  g790 (n870, n479, n631, n688, n441);
nand g791 (n895, n482, n443, n752, n731);
xor  g792 (n869, n746, n466, n739, n747);
and  g793 (n863, n658, n467, n719, n718);
xnor g794 (n891, n482, n459, n455, n726);
xnor g795 (n829, n676, n467, n719, n705);
xnor g796 (n872, n703, n634, n444, n708);
and  g797 (n883, n475, n737, n705, n460);
or   g798 (n834, n749, n752, n739, n717);
xor  g799 (n821, n468, n730, n448, n669);
nor  g800 (n842, n469, n648, n735, n477);
nor  g801 (n843, n724, n629, n445, n704);
xnor g802 (n901, n753, n654, n438, n732);
nand g803 (n904, n464, n722, n652, n483);
nand g804 (n899, n714, n468, n734, n445);
nand g805 (n850, n711, n650, n447, n693);
xor  g806 (n890, n734, n730, n703, n738);
nand g807 (n897, n720, n461, n463, n671);
nor  g808 (n825, n720, n436, n651, n449);
nand g809 (n846, n732, n691, n684, n456);
xnor g810 (n868, n642, n667, n710, n466);
nand g811 (n884, n443, n449, n715, n462);
nor  g812 (n903, n481, n461, n701, n483);
or   g813 (n855, n662, n750, n475, n471);
nand g814 (n854, n630, n451, n440, n458);
nand g815 (n865, n702, n485, n456, n447);
xnor g816 (n885, n673, n687, n458, n663);
or   g817 (n822, n641, n744, n476, n735);
xnor g818 (n827, n450, n701, n467, n440);
nor  g819 (n849, n710, n683, n745, n460);
xor  g820 (n881, n713, n475, n738, n472);
and  g821 (n877, n485, n736, n465, n453);
nor  g822 (n898, n706, n477, n714, n677);
nand g823 (n873, n440, n480, n674, n449);
and  g824 (n862, n453, n653, n479, n438);
xnor g825 (n864, n468, n640, n482, n462);
nor  g826 (n875, n457, n479, n435, n713);
nand g827 (n857, n721, n476, n463, n692);
nor  g828 (n847, n478, n733, n698, n633);
xnor g829 (n838, n726, n477, n462, n459);
and  g830 (n878, n457, n478, n473, n731);
xor  g831 (n826, n472, n454, n727, n723);
and  g832 (n893, n465, n753, n736, n439);
xor  g833 (n876, n451, n724, n708, n452);
xnor g834 (n880, n712, n469, n484, n747);
and  g835 (n882, n469, n750, n727, n442);
and  g836 (n874, n670, n453, n452, n743);
nand g837 (n839, n434, n473, n446, n741);
xnor g838 (n900, n480, n438, n442, n660);
xnor g839 (n871, n442, n483, n685, n718);
nor  g840 (n886, n455, n444, n644, n668);
nor  g841 (n894, n435, n729, n452, n679);
nand g842 (n833, n649, n743, n472, n484);
xor  g843 (n841, n655, n721, n446, n742);
xnor g844 (n844, n725, n740, n733, n456);
xnor g845 (n830, n672, n437, n457);
xor  g846 (n858, n441, n448, n635);
or   g847 (n848, n450, n439, n666, n711);
nand g848 (n860, n741, n725, n704, n455);
xor  g849 (n832, n436, n484, n678, n461);
xor  g850 (n879, n745, n435, n746, n458);
and  g851 (n835, n700, n695, n699, n643);
nand g852 (n866, n696, n751, n485, n445);
and  g853 (n837, n645, n690, n709, n451);
nor  g854 (n853, n647, n748, n636, n664);
or   g855 (n824, n470, n480, n682, n689);
nand g856 (n861, n742, n439, n748, n728);
nand g857 (n840, n675, n471, n459, n470);
xor  g858 (n888, n481, n637, n646, n717);
and  g859 (n836, n436, n656, n447, n702);
xnor g860 (n828, n737, n698, n638, n639);
nor  g861 (n823, n709, n686, n470, n454);
xnor g862 (n845, n699, n749, n478, n632);
or   g863 (n892, n707, n716, n657);
xor  g864 (n859, n661, n715, n441, n722);
nor  g865 (n831, n444, n463, n465, n460);
xnor g866 (n867, n476, n473, n740, n474);
nand g867 (n851, n700, n437, n454, n659);
xor  g868 (n856, n471, n706, n474, n665);
or   g869 (n852, n707, n466, n697, n474);
and  g870 (n887, n728, n712, n729, n681);
nor  g871 (n902, n744, n464, n443);
nand g872 (n928, n767, n755, n889, n757);
and  g873 (n930, n842, n761, n859, n825);
nor  g874 (n927, n757, n759, n892, n832);
or   g875 (n920, n755, n847, n831, n769);
and  g876 (n907, n871, n764, n767, n844);
nor  g877 (n919, n770, n861, n766, n875);
nor  g878 (n931, n874, n860, n835, n754);
xnor g879 (n915, n756, n821, n771, n853);
nand g880 (n916, n758, n893, n837, n888);
xnor g881 (n911, n851, n858, n823, n824);
and  g882 (n932, n879, n840, n882, n761);
nor  g883 (n908, n893, n770, n829, n890);
or   g884 (n914, n870, n872, n856, n852);
xnor g885 (n912, n830, n892, n839, n854);
nor  g886 (n922, n841, n869, n876, n765);
nand g887 (n923, n862, n887, n891, n769);
nor  g888 (n921, n754, n891, n836, n762);
or   g889 (n909, n765, n877, n885, n886);
xnor g890 (n910, n846, n771, n822, n867);
xnor g891 (n925, n855, n766, n880, n884);
and  g892 (n918, n843, n760, n865, n763);
or   g893 (n905, n826, n764, n827, n834);
or   g894 (n906, n863, n828, n768, n838);
xnor g895 (n913, n878, n848, n868, n759);
nand g896 (n917, n756, n763, n768, n864);
nor  g897 (n929, n849, n845, n760, n833);
xor  g898 (n926, n873, n883, n850, n758);
xor  g899 (n924, n881, n866, n762, n857);
or   g900 (n959, n908, n526, n900, n508);
and  g901 (n980, n490, n507, n906, n504);
or   g902 (n952, n913, n533, n490, n512);
and  g903 (n943, n898, n488, n503, n904);
xnor g904 (n937, n487, n498, n497);
and  g905 (n957, n785, n531, n528, n506);
xor  g906 (n999, n530, n488, n912, n780);
or   g907 (n1000, n905, n511, n489, n932);
nor  g908 (n998, n775, n932, n505, n780);
or   g909 (n987, n517, n486, n903, n495);
and  g910 (n949, n921, n492, n923);
nor  g911 (n939, n782, n516, n925, n928);
nand g912 (n990, n521, n513, n508, n533);
or   g913 (n965, n899, n924, n919, n529);
xor  g914 (n934, n500, n514, n789, n907);
nand g915 (n981, n509, n533, n492, n503);
nand g916 (n935, n510, n906, n777, n496);
nor  g917 (n984, n914, n529, n526, n496);
and  g918 (n995, n532, n530, n510, n494);
nand g919 (n960, n929, n923, n527, n517);
or   g920 (n955, n911, n529, n774, n511);
or   g921 (n977, n500, n501, n927, n907);
nand g922 (n988, n521, n912, n896, n498);
xnor g923 (n974, n897, n782, n909, n775);
xnor g924 (n972, n510, n491, n928, n895);
nand g925 (n953, n506, n788, n524, n523);
and  g926 (n950, n489, n486, n505, n904);
xnor g927 (n954, n911, n908, n515, n790);
xor  g928 (n975, n518, n897, n773, n772);
nand g929 (n970, n926, n504, n919, n520);
and  g930 (n986, n895, n777, n493, n931);
or   g931 (n961, n930, n527, n913, n524);
xnor g932 (n942, n503, n926, n514, n778);
and  g933 (n940, n516, n917, n920, n929);
and  g934 (n936, n920, n531, n916, n491);
nand g935 (n951, n776, n786, n523);
nor  g936 (n946, n921, n488, n525);
and  g937 (n976, n783, n512, n894, n778);
nor  g938 (n982, n495, n511, n521, n513);
nor  g939 (n997, n784, n910, n520, n519);
xor  g940 (n947, n502, n519, n513, n495);
and  g941 (n978, n528, n517, n507, n518);
xor  g942 (n962, n499, n499, n494, n903);
nor  g943 (n979, n506, n779, n531, n923);
or   g944 (n983, n505, n902, n523, n772);
or   g945 (n969, n925, n931, n501, n526);
nor  g946 (n985, n779, n783, n929, n532);
xor  g947 (n996, n930, n785, n901, n902);
xor  g948 (n948, n915, n916, n930, n918);
or   g949 (n989, n784, n905, n787, n781);
and  g950 (n992, n900, n932, n776, n787);
or   g951 (n964, n774, n924, n490, n527);
or   g952 (n994, n493, n520, n512, n927);
nor  g953 (n973, n910, n922, n491, n516);
or   g954 (n967, n508, n493, n486, n918);
and  g955 (n971, n926, n494, n928, n922);
or   g956 (n956, n530, n509, n524, n489);
nand g957 (n968, n525, n502, n915, n522);
xnor g958 (n933, n497, n788, n515, n773);
nand g959 (n938, n790, n924, n500, n921);
and  g960 (n945, n497, n899, n528, n532);
nor  g961 (n963, n931, n894, n917, n927);
and  g962 (n966, n914, n518, n507, n909);
and  g963 (n991, n781, n509, n499, n901);
or   g964 (n958, n487, n487, n496, n898);
nand g965 (n941, n925, n922, n502, n789);
xor  g966 (n944, n522, n896, n504, n515);
nor  g967 (n993, n514, n522, n501, n519);
nor  g968 (n1001, n958, n808, n977, n798);
xor  g969 (n1020, n991, n986, n818, n972);
and  g970 (n1017, n955, n808, n959, n935);
xor  g971 (n1021, n957, n966, n814, n968);
xnor g972 (n1010, n794, n797, n796, n814);
or   g973 (n1004, n953, n817, n940, n795);
and  g974 (n1008, n799, n795, n811, n796);
and  g975 (n1002, n792, n815, n818, n987);
or   g976 (n1030, n800, n807, n819, n944);
xnor g977 (n1019, n943, n812, n952, n817);
or   g978 (n1024, n996, n806, n976, n961);
xor  g979 (n1032, n1000, n819, n992, n820);
and  g980 (n1011, n933, n791, n816, n970);
or   g981 (n1003, n979, n969, n975, n806);
and  g982 (n1016, n960, n948, n815, n978);
nand g983 (n1023, n994, n988, n809, n813);
xor  g984 (n1014, n956, n934, n983, n985);
and  g985 (n1025, n981, n938, n945, n995);
nand g986 (n1007, n941, n816, n980, n802);
or   g987 (n1029, n813, n947, n982, n792);
and  g988 (n1027, n964, n974, n967, n807);
and  g989 (n1015, n803, n793, n794);
or   g990 (n1026, n800, n803, n950, n999);
xor  g991 (n1009, n809, n939, n810, n984);
xor  g992 (n1018, n954, n804, n942, n812);
or   g993 (n1022, n998, n805, n971, n997);
or   g994 (n1006, n965, n799, n949, n990);
or   g995 (n1012, n937, n820, n804, n798);
or   g996 (n1031, n802, n811, n801, n791);
and  g997 (n1013, n797, n951, n989, n962);
and  g998 (n1005, n993, n963, n801, n946);
xnor g999 (n1028, n805, n973, n810, n936);
endmodule
