

module Stat_2000_228
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n171,
  n167,
  n123,
  n79,
  n155,
  n85,
  n185,
  n132,
  n195,
  n179,
  n93,
  n162,
  n108,
  n151,
  n176,
  n191,
  n1881,
  n2025,
  n2021,
  n2020,
  n2019,
  n2023,
  n2027,
  n2022,
  n2028,
  n2032,
  n2031,
  n2026,
  n2029,
  n2024,
  n2030,
  n2018
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n171;output n167;output n123;output n79;output n155;output n85;output n185;output n132;output n195;output n179;output n93;output n162;output n108;output n151;output n176;output n191;output n1881;output n2025;output n2021;output n2020;output n2019;output n2023;output n2027;output n2022;output n2028;output n2032;output n2031;output n2026;output n2029;output n2024;output n2030;output n2018;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n80;wire n81;wire n82;wire n83;wire n84;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n152;wire n153;wire n154;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n163;wire n164;wire n165;wire n166;wire n168;wire n169;wire n170;wire n172;wire n173;wire n174;wire n175;wire n177;wire n178;wire n180;wire n181;wire n182;wire n183;wire n184;wire n186;wire n187;wire n188;wire n189;wire n190;wire n192;wire n193;wire n194;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n34,
    n16
  );


  buf
  g1
  (
    n40,
    n18
  );


  buf
  g2
  (
    n35,
    n13
  );


  buf
  g3
  (
    n41,
    n4
  );


  buf
  g4
  (
    n33,
    n8
  );


  buf
  g5
  (
    n39,
    n1
  );


  nor
  g6
  (
    n37,
    n5,
    n15,
    n9,
    n3
  );


  nand
  g7
  (
    n36,
    n12,
    n17,
    n11,
    n7
  );


  xnor
  g8
  (
    n38,
    n14,
    n2,
    n10,
    n6
  );


  not
  g9
  (
    n54,
    n41
  );


  not
  g10
  (
    n66,
    n34
  );


  buf
  g11
  (
    n47,
    n22
  );


  buf
  g12
  (
    n42,
    n21
  );


  not
  g13
  (
    n59,
    n36
  );


  not
  g14
  (
    n63,
    n35
  );


  buf
  g15
  (
    n65,
    n34
  );


  not
  g16
  (
    n56,
    n41
  );


  buf
  g17
  (
    n45,
    n40
  );


  buf
  g18
  (
    n68,
    n23
  );


  not
  g19
  (
    n75,
    n33
  );


  not
  g20
  (
    n64,
    n37
  );


  buf
  g21
  (
    n51,
    n35
  );


  buf
  g22
  (
    KeyWire_0_3,
    n37
  );


  buf
  g23
  (
    n46,
    n20
  );


  buf
  g24
  (
    n62,
    n39
  );


  not
  g25
  (
    n77,
    n39
  );


  buf
  g26
  (
    n58,
    n40
  );


  not
  g27
  (
    n76,
    n36
  );


  not
  g28
  (
    n55,
    n39
  );


  not
  g29
  (
    n61,
    n24
  );


  buf
  g30
  (
    n57,
    n33
  );


  buf
  g31
  (
    n44,
    n38
  );


  not
  g32
  (
    n49,
    n33
  );


  not
  g33
  (
    n74,
    n38
  );


  not
  g34
  (
    n70,
    n37
  );


  not
  g35
  (
    n71,
    n40
  );


  not
  g36
  (
    n50,
    n34
  );


  not
  g37
  (
    n67,
    n36
  );


  not
  g38
  (
    n53,
    n35
  );


  not
  g39
  (
    n69,
    n33
  );


  not
  g40
  (
    n43,
    n38
  );


  buf
  g41
  (
    n60,
    n37
  );


  xor
  g42
  (
    n52,
    n35,
    n41,
    n38
  );


  nor
  g43
  (
    n73,
    n19,
    n40,
    n36
  );


  and
  g44
  (
    n48,
    n34,
    n39,
    n41
  );


  not
  g45
  (
    n133,
    n44
  );


  buf
  g46
  (
    n103,
    n45
  );


  not
  g47
  (
    n119,
    n45
  );


  not
  g48
  (
    n190,
    n69
  );


  not
  g49
  (
    n172,
    n68
  );


  buf
  g50
  (
    n95,
    n68
  );


  buf
  g51
  (
    n171,
    n52
  );


  buf
  g52
  (
    n123,
    n57
  );


  not
  g53
  (
    n164,
    n69
  );


  buf
  g54
  (
    n122,
    n71
  );


  buf
  g55
  (
    n170,
    n44
  );


  not
  g56
  (
    n174,
    n58
  );


  not
  g57
  (
    n145,
    n53
  );


  buf
  g58
  (
    n96,
    n44
  );


  not
  g59
  (
    n173,
    n46
  );


  buf
  g60
  (
    n79,
    n64
  );


  not
  g61
  (
    n108,
    n51
  );


  buf
  g62
  (
    n168,
    n45
  );


  not
  g63
  (
    n140,
    n47
  );


  buf
  g64
  (
    n126,
    n49
  );


  not
  g65
  (
    n193,
    n56
  );


  buf
  g66
  (
    n151,
    n57
  );


  buf
  g67
  (
    n106,
    n55
  );


  buf
  g68
  (
    n118,
    n58
  );


  not
  g69
  (
    n86,
    n71
  );


  buf
  g70
  (
    n182,
    n47
  );


  not
  g71
  (
    n180,
    n71
  );


  buf
  g72
  (
    n185,
    n46
  );


  buf
  g73
  (
    n128,
    n63
  );


  buf
  g74
  (
    n196,
    n60
  );


  buf
  g75
  (
    n167,
    n53
  );


  not
  g76
  (
    n110,
    n42
  );


  buf
  g77
  (
    n152,
    n63
  );


  buf
  g78
  (
    n139,
    n65
  );


  buf
  g79
  (
    n127,
    n47
  );


  buf
  g80
  (
    n99,
    n53
  );


  not
  g81
  (
    n163,
    n44
  );


  buf
  g82
  (
    n112,
    n64
  );


  buf
  g83
  (
    n194,
    n67
  );


  buf
  g84
  (
    n154,
    n51
  );


  not
  g85
  (
    n121,
    n53
  );


  not
  g86
  (
    n138,
    n56
  );


  buf
  g87
  (
    n83,
    n43
  );


  buf
  g88
  (
    n82,
    n59
  );


  not
  g89
  (
    n197,
    n55
  );


  buf
  g90
  (
    n176,
    n50
  );


  buf
  g91
  (
    n160,
    n60
  );


  buf
  g92
  (
    n192,
    n60
  );


  not
  g93
  (
    n179,
    n68
  );


  buf
  g94
  (
    n129,
    n56
  );


  buf
  g95
  (
    n120,
    n61
  );


  not
  g96
  (
    n148,
    n55
  );


  buf
  g97
  (
    n161,
    n58
  );


  buf
  g98
  (
    n81,
    n54
  );


  not
  g99
  (
    n195,
    n58
  );


  buf
  g100
  (
    n84,
    n57
  );


  not
  g101
  (
    n125,
    n50
  );


  not
  g102
  (
    n155,
    n43
  );


  not
  g103
  (
    n98,
    n70
  );


  not
  g104
  (
    n94,
    n50
  );


  buf
  g105
  (
    n141,
    n62
  );


  not
  g106
  (
    n159,
    n66
  );


  buf
  g107
  (
    n113,
    n43
  );


  not
  g108
  (
    n115,
    n45
  );


  buf
  g109
  (
    n91,
    n50
  );


  buf
  g110
  (
    n135,
    n52
  );


  buf
  g111
  (
    n189,
    n48
  );


  not
  g112
  (
    n178,
    n49
  );


  not
  g113
  (
    n100,
    n71
  );


  not
  g114
  (
    n175,
    n59
  );


  buf
  g115
  (
    n184,
    n67
  );


  buf
  g116
  (
    n105,
    n49
  );


  buf
  g117
  (
    n111,
    n43
  );


  buf
  g118
  (
    n87,
    n51
  );


  not
  g119
  (
    n109,
    n69
  );


  not
  g120
  (
    n134,
    n65
  );


  not
  g121
  (
    n102,
    n61
  );


  buf
  g122
  (
    n116,
    n46
  );


  not
  g123
  (
    n198,
    n54
  );


  not
  g124
  (
    n166,
    n52
  );


  not
  g125
  (
    n188,
    n66
  );


  not
  g126
  (
    n137,
    n65
  );


  buf
  g127
  (
    n130,
    n61
  );


  buf
  g128
  (
    n101,
    n68
  );


  buf
  g129
  (
    n78,
    n55
  );


  not
  g130
  (
    KeyWire_0_31,
    n49
  );


  buf
  g131
  (
    n149,
    n48
  );


  buf
  g132
  (
    n93,
    n59
  );


  buf
  g133
  (
    n165,
    n48
  );


  not
  g134
  (
    n183,
    n61
  );


  not
  g135
  (
    n124,
    n66
  );


  buf
  g136
  (
    n186,
    n54
  );


  not
  g137
  (
    n88,
    n51
  );


  not
  g138
  (
    n80,
    n63
  );


  buf
  g139
  (
    n92,
    n42
  );


  not
  g140
  (
    n143,
    n62
  );


  buf
  g141
  (
    n132,
    n72
  );


  not
  g142
  (
    n90,
    n52
  );


  buf
  g143
  (
    n157,
    n59
  );


  not
  g144
  (
    n104,
    n42
  );


  not
  g145
  (
    n147,
    n66
  );


  not
  g146
  (
    n156,
    n47
  );


  not
  g147
  (
    n169,
    n65
  );


  not
  g148
  (
    KeyWire_0_10,
    n69
  );


  not
  g149
  (
    n153,
    n64
  );


  buf
  g150
  (
    n187,
    n70
  );


  not
  g151
  (
    n89,
    n67
  );


  not
  g152
  (
    n191,
    n60
  );


  buf
  g153
  (
    n150,
    n62
  );


  not
  g154
  (
    n97,
    n64
  );


  buf
  g155
  (
    n131,
    n48
  );


  buf
  g156
  (
    n162,
    n63
  );


  buf
  g157
  (
    n117,
    n70
  );


  buf
  g158
  (
    n181,
    n42
  );


  buf
  g159
  (
    n85,
    n54
  );


  not
  g160
  (
    n177,
    n46
  );


  buf
  g161
  (
    n114,
    n56
  );


  not
  g162
  (
    n158,
    n57
  );


  buf
  g163
  (
    n142,
    n70
  );


  not
  g164
  (
    n136,
    n67
  );


  not
  g165
  (
    n107,
    n62
  );


  not
  g166
  (
    n208,
    n155
  );


  not
  g167
  (
    n257,
    n122
  );


  not
  g168
  (
    n238,
    n177
  );


  not
  g169
  (
    n400,
    n140
  );


  buf
  g170
  (
    n388,
    n163
  );


  not
  g171
  (
    n381,
    n158
  );


  buf
  g172
  (
    n317,
    n180
  );


  buf
  g173
  (
    n409,
    n156
  );


  not
  g174
  (
    n382,
    n162
  );


  buf
  g175
  (
    n345,
    n172
  );


  not
  g176
  (
    n337,
    n168
  );


  not
  g177
  (
    n313,
    n139
  );


  buf
  g178
  (
    n407,
    n188
  );


  not
  g179
  (
    n362,
    n143
  );


  not
  g180
  (
    n380,
    n152
  );


  not
  g181
  (
    n339,
    n181
  );


  buf
  g182
  (
    n360,
    n162
  );


  buf
  g183
  (
    n268,
    n157
  );


  buf
  g184
  (
    n295,
    n78
  );


  not
  g185
  (
    n338,
    n184
  );


  buf
  g186
  (
    n386,
    n173
  );


  buf
  g187
  (
    n371,
    n129
  );


  not
  g188
  (
    n403,
    n191
  );


  buf
  g189
  (
    n209,
    n126
  );


  not
  g190
  (
    n349,
    n176
  );


  not
  g191
  (
    n287,
    n187
  );


  buf
  g192
  (
    n301,
    n99
  );


  not
  g193
  (
    n264,
    n158
  );


  not
  g194
  (
    n391,
    n164
  );


  not
  g195
  (
    n366,
    n165
  );


  not
  g196
  (
    n274,
    n191
  );


  buf
  g197
  (
    n325,
    n179
  );


  not
  g198
  (
    n385,
    n178
  );


  buf
  g199
  (
    n297,
    n183
  );


  buf
  g200
  (
    n379,
    n106
  );


  buf
  g201
  (
    n378,
    n188
  );


  buf
  g202
  (
    n342,
    n138
  );


  buf
  g203
  (
    n254,
    n136
  );


  buf
  g204
  (
    n229,
    n150
  );


  buf
  g205
  (
    n341,
    n112
  );


  not
  g206
  (
    n377,
    n174
  );


  not
  g207
  (
    n402,
    n187
  );


  buf
  g208
  (
    n411,
    n152
  );


  buf
  g209
  (
    n279,
    n148
  );


  buf
  g210
  (
    n405,
    n145
  );


  buf
  g211
  (
    n364,
    n172
  );


  buf
  g212
  (
    n260,
    n176
  );


  not
  g213
  (
    n240,
    n184
  );


  buf
  g214
  (
    n284,
    n181
  );


  not
  g215
  (
    n305,
    n144
  );


  buf
  g216
  (
    n415,
    n169
  );


  buf
  g217
  (
    n414,
    n167
  );


  buf
  g218
  (
    n256,
    n95
  );


  not
  g219
  (
    n370,
    n132
  );


  buf
  g220
  (
    n273,
    n147
  );


  not
  g221
  (
    n335,
    n157
  );


  not
  g222
  (
    n350,
    n182
  );


  buf
  g223
  (
    n223,
    n153
  );


  buf
  g224
  (
    n401,
    n190
  );


  buf
  g225
  (
    n231,
    n130
  );


  buf
  g226
  (
    n340,
    n103
  );


  buf
  g227
  (
    n214,
    n150
  );


  buf
  g228
  (
    n320,
    n144
  );


  not
  g229
  (
    n315,
    n118
  );


  not
  g230
  (
    n418,
    n174
  );


  not
  g231
  (
    n314,
    n96
  );


  buf
  g232
  (
    n404,
    n164
  );


  buf
  g233
  (
    n237,
    n171
  );


  not
  g234
  (
    n354,
    n111
  );


  buf
  g235
  (
    n259,
    n140
  );


  not
  g236
  (
    KeyWire_0_30,
    n113
  );


  buf
  g237
  (
    n303,
    n191
  );


  not
  g238
  (
    n351,
    n115
  );


  not
  g239
  (
    n316,
    n177
  );


  buf
  g240
  (
    n406,
    n183
  );


  not
  g241
  (
    n361,
    n143
  );


  buf
  g242
  (
    n389,
    n149
  );


  not
  g243
  (
    n251,
    n135
  );


  not
  g244
  (
    n291,
    n92
  );


  buf
  g245
  (
    n225,
    n186
  );


  buf
  g246
  (
    n226,
    n142
  );


  buf
  g247
  (
    n282,
    n190
  );


  not
  g248
  (
    n278,
    n189
  );


  buf
  g249
  (
    n227,
    n180
  );


  not
  g250
  (
    n236,
    n147
  );


  buf
  g251
  (
    n250,
    n181
  );


  not
  g252
  (
    n272,
    n152
  );


  not
  g253
  (
    n333,
    n123
  );


  buf
  g254
  (
    n365,
    n189
  );


  not
  g255
  (
    n343,
    n100
  );


  not
  g256
  (
    n252,
    n82
  );


  buf
  g257
  (
    n275,
    n154
  );


  not
  g258
  (
    n373,
    n119
  );


  buf
  g259
  (
    n294,
    n131
  );


  buf
  g260
  (
    n393,
    n182
  );


  not
  g261
  (
    n416,
    n141
  );


  buf
  g262
  (
    KeyWire_0_20,
    n91
  );


  not
  g263
  (
    n412,
    n94
  );


  buf
  g264
  (
    n392,
    n79
  );


  buf
  g265
  (
    n258,
    n162
  );


  not
  g266
  (
    n263,
    n168
  );


  not
  g267
  (
    n306,
    n81
  );


  buf
  g268
  (
    n283,
    n124
  );


  not
  g269
  (
    n336,
    n167
  );


  not
  g270
  (
    n300,
    n183
  );


  buf
  g271
  (
    n348,
    n127
  );


  not
  g272
  (
    n290,
    n88
  );


  not
  g273
  (
    n218,
    n173
  );


  not
  g274
  (
    n255,
    n133
  );


  buf
  g275
  (
    KeyWire_0_21,
    n145
  );


  buf
  g276
  (
    n245,
    n169
  );


  buf
  g277
  (
    n212,
    n182
  );


  not
  g278
  (
    n244,
    n155
  );


  not
  g279
  (
    n281,
    n163
  );


  buf
  g280
  (
    n397,
    n110
  );


  buf
  g281
  (
    n285,
    n109
  );


  not
  g282
  (
    n277,
    n178
  );


  buf
  g283
  (
    n230,
    n143
  );


  not
  g284
  (
    n280,
    n159
  );


  not
  g285
  (
    n249,
    n186
  );


  not
  g286
  (
    n233,
    n132
  );


  buf
  g287
  (
    n266,
    n137
  );


  not
  g288
  (
    n201,
    n185
  );


  not
  g289
  (
    n286,
    n150
  );


  buf
  g290
  (
    n248,
    n136
  );


  buf
  g291
  (
    KeyWire_0_23,
    n189
  );


  buf
  g292
  (
    n328,
    n97
  );


  buf
  g293
  (
    n307,
    n187
  );


  buf
  g294
  (
    n359,
    n182
  );


  buf
  g295
  (
    n396,
    n104
  );


  buf
  g296
  (
    n367,
    n146
  );


  not
  g297
  (
    n352,
    n166
  );


  not
  g298
  (
    n289,
    n156
  );


  buf
  g299
  (
    n347,
    n161
  );


  not
  g300
  (
    n213,
    n85
  );


  buf
  g301
  (
    n265,
    n139
  );


  buf
  g302
  (
    n410,
    n166
  );


  buf
  g303
  (
    n221,
    n151
  );


  buf
  g304
  (
    n200,
    n128
  );


  not
  g305
  (
    n242,
    n145
  );


  not
  g306
  (
    n363,
    n169
  );


  not
  g307
  (
    n222,
    n183
  );


  not
  g308
  (
    n206,
    n138
  );


  not
  g309
  (
    n271,
    n173
  );


  buf
  g310
  (
    n235,
    n181
  );


  not
  g311
  (
    n298,
    n93
  );


  not
  g312
  (
    n304,
    n178
  );


  not
  g313
  (
    n383,
    n154
  );


  buf
  g314
  (
    n394,
    n186
  );


  buf
  g315
  (
    n330,
    n163
  );


  not
  g316
  (
    n199,
    n170
  );


  not
  g317
  (
    n220,
    n151
  );


  buf
  g318
  (
    n353,
    n134
  );


  buf
  g319
  (
    n376,
    n135
  );


  not
  g320
  (
    n357,
    n146
  );


  buf
  g321
  (
    n358,
    n146
  );


  buf
  g322
  (
    n413,
    n172
  );


  not
  g323
  (
    n207,
    n148
  );


  not
  g324
  (
    n375,
    n137
  );


  buf
  g325
  (
    n368,
    n105
  );


  not
  g326
  (
    n374,
    n171
  );


  buf
  g327
  (
    n323,
    n141
  );


  buf
  g328
  (
    n204,
    n89
  );


  buf
  g329
  (
    n417,
    n161
  );


  buf
  g330
  (
    n395,
    n141
  );


  not
  g331
  (
    n205,
    n121
  );


  not
  g332
  (
    n369,
    n170
  );


  not
  g333
  (
    n217,
    n153
  );


  buf
  g334
  (
    n293,
    n191
  );


  buf
  g335
  (
    n246,
    n167
  );


  not
  g336
  (
    n312,
    n185
  );


  not
  g337
  (
    n267,
    n139
  );


  buf
  g338
  (
    n276,
    n179
  );


  buf
  g339
  (
    n310,
    n160
  );


  buf
  g340
  (
    n329,
    n166
  );


  not
  g341
  (
    n387,
    n134
  );


  not
  g342
  (
    n210,
    n185
  );


  not
  g343
  (
    n419,
    n114
  );


  not
  g344
  (
    n322,
    n83
  );


  not
  g345
  (
    n292,
    n157
  );


  buf
  g346
  (
    n202,
    n132
  );


  buf
  g347
  (
    n356,
    n117
  );


  buf
  g348
  (
    n319,
    n187
  );


  buf
  g349
  (
    n332,
    n185
  );


  not
  g350
  (
    n228,
    n138
  );


  buf
  g351
  (
    n390,
    n142
  );


  not
  g352
  (
    n234,
    n168
  );


  buf
  g353
  (
    n355,
    n186
  );


  buf
  g354
  (
    n219,
    n177
  );


  not
  g355
  (
    n215,
    n142
  );


  buf
  g356
  (
    n299,
    n188
  );


  buf
  g357
  (
    n331,
    n87
  );


  buf
  g358
  (
    n203,
    n120
  );


  buf
  g359
  (
    n334,
    n133
  );


  buf
  g360
  (
    n372,
    n90
  );


  buf
  g361
  (
    n232,
    n108
  );


  not
  g362
  (
    n296,
    n140
  );


  or
  g363
  (
    n253,
    n134,
    n84
  );


  or
  g364
  (
    n321,
    n116,
    n160
  );


  xor
  g365
  (
    n239,
    n180,
    n133
  );


  and
  g366
  (
    n302,
    n151,
    n149
  );


  nand
  g367
  (
    n309,
    n155,
    n156
  );


  or
  g368
  (
    n224,
    n125,
    n107
  );


  nor
  g369
  (
    n262,
    n160,
    n171
  );


  and
  g370
  (
    n270,
    n175,
    n80
  );


  or
  g371
  (
    n247,
    n170,
    n101
  );


  and
  g372
  (
    n398,
    n102,
    n153
  );


  and
  g373
  (
    n216,
    n165,
    n184
  );


  nand
  g374
  (
    n243,
    n158,
    n159
  );


  nand
  g375
  (
    n344,
    n175,
    n164
  );


  nand
  g376
  (
    n211,
    n188,
    n86
  );


  and
  g377
  (
    n346,
    n190,
    n159
  );


  or
  g378
  (
    n399,
    n189,
    n136
  );


  xor
  g379
  (
    n308,
    n149,
    n184
  );


  xor
  g380
  (
    n318,
    n137,
    n175
  );


  xor
  g381
  (
    n241,
    n144,
    n148
  );


  nor
  g382
  (
    n269,
    n161,
    n135
  );


  xnor
  g383
  (
    n408,
    n147,
    n165
  );


  nor
  g384
  (
    n261,
    n179,
    n154
  );


  nand
  g385
  (
    n324,
    n176,
    n190
  );


  xnor
  g386
  (
    n327,
    n98,
    n174
  );


  buf
  g387
  (
    n421,
    n200
  );


  buf
  g388
  (
    n420,
    n199
  );


  xnor
  g389
  (
    n422,
    n203,
    n204
  );


  buf
  g390
  (
    n424,
    n420
  );


  nand
  g391
  (
    n423,
    n202,
    n201,
    n420,
    n205
  );


  not
  g392
  (
    n431,
    n421
  );


  not
  g393
  (
    n432,
    n423
  );


  nor
  g394
  (
    n425,
    n194,
    n192
  );


  xor
  g395
  (
    n434,
    n194,
    n194,
    n195,
    n424
  );


  xnor
  g396
  (
    n430,
    n195,
    n194,
    n422,
    n192
  );


  xor
  g397
  (
    n433,
    n423,
    n424,
    n421,
    n193
  );


  and
  g398
  (
    n429,
    n424,
    n72,
    n192,
    n422
  );


  or
  g399
  (
    n428,
    n192,
    n421,
    n193,
    n423
  );


  or
  g400
  (
    n426,
    n207,
    n193,
    n72,
    n206
  );


  xnor
  g401
  (
    n427,
    n424,
    n420,
    n423,
    n193
  );


  not
  g402
  (
    n446,
    n429
  );


  not
  g403
  (
    n437,
    n434
  );


  buf
  g404
  (
    n438,
    n425
  );


  buf
  g405
  (
    n447,
    n209
  );


  not
  g406
  (
    n442,
    n433
  );


  not
  g407
  (
    n435,
    n432
  );


  buf
  g408
  (
    n444,
    n434
  );


  buf
  g409
  (
    n450,
    n208
  );


  not
  g410
  (
    KeyWire_0_16,
    n426
  );


  not
  g411
  (
    n439,
    n431
  );


  not
  g412
  (
    n440,
    n427
  );


  not
  g413
  (
    n445,
    n433
  );


  not
  g414
  (
    n441,
    n431
  );


  buf
  g415
  (
    n443,
    n428
  );


  not
  g416
  (
    n448,
    n434
  );


  xor
  g417
  (
    n449,
    n430,
    n434,
    n432
  );


  not
  g418
  (
    n505,
    n437
  );


  not
  g419
  (
    n491,
    n281
  );


  buf
  g420
  (
    n470,
    n288
  );


  not
  g421
  (
    n458,
    n251
  );


  not
  g422
  (
    n509,
    n210
  );


  not
  g423
  (
    n494,
    n440
  );


  not
  g424
  (
    n464,
    n435
  );


  buf
  g425
  (
    n480,
    n435
  );


  buf
  g426
  (
    n453,
    n440
  );


  not
  g427
  (
    n475,
    n217
  );


  buf
  g428
  (
    n457,
    n256
  );


  not
  g429
  (
    n460,
    n219
  );


  not
  g430
  (
    n476,
    n223
  );


  not
  g431
  (
    n498,
    n261
  );


  buf
  g432
  (
    n504,
    n439
  );


  buf
  g433
  (
    n487,
    n257
  );


  not
  g434
  (
    n513,
    n284
  );


  buf
  g435
  (
    n486,
    n450
  );


  buf
  g436
  (
    n484,
    n275
  );


  buf
  g437
  (
    n506,
    n266
  );


  buf
  g438
  (
    n461,
    n216
  );


  not
  g439
  (
    n485,
    n233
  );


  buf
  g440
  (
    n496,
    n436
  );


  buf
  g441
  (
    n463,
    n269
  );


  not
  g442
  (
    n472,
    n213
  );


  buf
  g443
  (
    n503,
    n446
  );


  not
  g444
  (
    KeyWire_0_7,
    n447
  );


  buf
  g445
  (
    n490,
    n232
  );


  not
  g446
  (
    n467,
    n265
  );


  buf
  g447
  (
    n454,
    n450
  );


  buf
  g448
  (
    n512,
    n259
  );


  buf
  g449
  (
    n474,
    n221
  );


  buf
  g450
  (
    n492,
    n264
  );


  buf
  g451
  (
    n452,
    n228
  );


  not
  g452
  (
    n469,
    n446
  );


  buf
  g453
  (
    n488,
    n443
  );


  xnor
  g454
  (
    n499,
    n220,
    n446
  );


  and
  g455
  (
    n471,
    n444,
    n244,
    n242,
    n279
  );


  and
  g456
  (
    n514,
    n282,
    n436,
    n246,
    n241
  );


  xnor
  g457
  (
    n500,
    n253,
    n212,
    n442,
    n247
  );


  nand
  g458
  (
    n478,
    n445,
    n290,
    n278,
    n287
  );


  nand
  g459
  (
    n473,
    n448,
    n444,
    n249,
    n263
  );


  xnor
  g460
  (
    n462,
    n449,
    n445,
    n254,
    n273
  );


  nor
  g461
  (
    n497,
    n214,
    n450,
    n243,
    n211
  );


  nor
  g462
  (
    n455,
    n238,
    n435,
    n443,
    n449
  );


  nand
  g463
  (
    n468,
    n268,
    n240,
    n235,
    n234
  );


  nand
  g464
  (
    n456,
    n448,
    n439,
    n437,
    n231
  );


  or
  g465
  (
    n502,
    n449,
    n280,
    n436,
    n262
  );


  or
  g466
  (
    n479,
    n446,
    n435,
    n229,
    n450
  );


  or
  g467
  (
    n466,
    n255,
    n445,
    n225,
    n443
  );


  nand
  g468
  (
    n508,
    n441,
    n270,
    n239,
    n224
  );


  nand
  g469
  (
    n481,
    n250,
    n448,
    n442,
    n258
  );


  nand
  g470
  (
    n482,
    n267,
    n222,
    n272,
    n441
  );


  xor
  g471
  (
    n501,
    n438,
    n277,
    n248,
    n439
  );


  nand
  g472
  (
    n477,
    n230,
    n218,
    n289,
    n443
  );


  nand
  g473
  (
    n507,
    n444,
    n447,
    n276,
    n215
  );


  xnor
  g474
  (
    n510,
    n245,
    n437,
    n438,
    n252
  );


  xnor
  g475
  (
    n511,
    n438,
    n442,
    n285,
    n226
  );


  xnor
  g476
  (
    n493,
    n227,
    n447,
    n440,
    n439
  );


  xnor
  g477
  (
    n451,
    n441,
    n440,
    n286,
    n442
  );


  nand
  g478
  (
    n459,
    n448,
    n283,
    n437,
    n291
  );


  nor
  g479
  (
    n489,
    n237,
    n271,
    n274,
    n260
  );


  nor
  g480
  (
    n495,
    n447,
    n445,
    n436,
    n236
  );


  xor
  g481
  (
    n483,
    n444,
    n441,
    n438,
    n449
  );


  buf
  g482
  (
    n584,
    n461
  );


  not
  g483
  (
    n580,
    n496
  );


  not
  g484
  (
    n682,
    n497
  );


  buf
  g485
  (
    n628,
    n452
  );


  not
  g486
  (
    n743,
    n454
  );


  not
  g487
  (
    n708,
    n457
  );


  not
  g488
  (
    n659,
    n496
  );


  buf
  g489
  (
    n548,
    n468
  );


  not
  g490
  (
    n531,
    n475
  );


  not
  g491
  (
    n732,
    n513
  );


  buf
  g492
  (
    n720,
    n471
  );


  buf
  g493
  (
    n748,
    n477
  );


  not
  g494
  (
    n701,
    n488
  );


  buf
  g495
  (
    n677,
    n507
  );


  buf
  g496
  (
    n590,
    n26
  );


  not
  g497
  (
    n712,
    n466
  );


  buf
  g498
  (
    n621,
    n73
  );


  buf
  g499
  (
    n650,
    n469
  );


  buf
  g500
  (
    n671,
    n504
  );


  not
  g501
  (
    n752,
    n494
  );


  not
  g502
  (
    n691,
    n197
  );


  buf
  g503
  (
    n747,
    n460
  );


  buf
  g504
  (
    n601,
    n462
  );


  buf
  g505
  (
    n526,
    n456
  );


  buf
  g506
  (
    n704,
    n511
  );


  not
  g507
  (
    KeyWire_0_17,
    n462
  );


  buf
  g508
  (
    n751,
    n478
  );


  not
  g509
  (
    n600,
    n490
  );


  not
  g510
  (
    n521,
    n453
  );


  buf
  g511
  (
    n658,
    n507
  );


  not
  g512
  (
    n577,
    n196
  );


  buf
  g513
  (
    n594,
    n505
  );


  not
  g514
  (
    KeyWire_0_15,
    n451
  );


  buf
  g515
  (
    n766,
    n492
  );


  buf
  g516
  (
    n690,
    n296
  );


  buf
  g517
  (
    n755,
    n460
  );


  buf
  g518
  (
    n663,
    n494
  );


  buf
  g519
  (
    n554,
    n508
  );


  not
  g520
  (
    n759,
    n498
  );


  not
  g521
  (
    n637,
    n482
  );


  buf
  g522
  (
    n745,
    n488
  );


  buf
  g523
  (
    n608,
    n489
  );


  not
  g524
  (
    n611,
    n489
  );


  buf
  g525
  (
    n726,
    n484
  );


  not
  g526
  (
    n674,
    n464
  );


  buf
  g527
  (
    n614,
    n452
  );


  not
  g528
  (
    n763,
    n472
  );


  not
  g529
  (
    n733,
    n511
  );


  buf
  g530
  (
    n542,
    n506
  );


  buf
  g531
  (
    n762,
    n514
  );


  buf
  g532
  (
    n685,
    n479
  );


  buf
  g533
  (
    n588,
    n502
  );


  not
  g534
  (
    n676,
    n492
  );


  buf
  g535
  (
    n769,
    n473
  );


  not
  g536
  (
    n758,
    n74
  );


  not
  g537
  (
    n686,
    n506
  );


  buf
  g538
  (
    n620,
    n196
  );


  not
  g539
  (
    n656,
    n498
  );


  not
  g540
  (
    n666,
    n491
  );


  not
  g541
  (
    n592,
    n455
  );


  buf
  g542
  (
    n753,
    n77
  );


  buf
  g543
  (
    n524,
    n491
  );


  not
  g544
  (
    n717,
    n497
  );


  not
  g545
  (
    n591,
    n466
  );


  buf
  g546
  (
    n523,
    n503
  );


  buf
  g547
  (
    n578,
    n510
  );


  buf
  g548
  (
    n606,
    n465
  );


  buf
  g549
  (
    n736,
    n466
  );


  not
  g550
  (
    n557,
    n484
  );


  buf
  g551
  (
    n573,
    n74
  );


  buf
  g552
  (
    n665,
    n491
  );


  buf
  g553
  (
    n599,
    n489
  );


  buf
  g554
  (
    n532,
    n198
  );


  not
  g555
  (
    n718,
    n421
  );


  not
  g556
  (
    n630,
    n504
  );


  not
  g557
  (
    n567,
    n479
  );


  buf
  g558
  (
    n527,
    n300
  );


  buf
  g559
  (
    n749,
    n454
  );


  not
  g560
  (
    n569,
    n466
  );


  buf
  g561
  (
    n731,
    n453
  );


  not
  g562
  (
    n741,
    n505
  );


  buf
  g563
  (
    n538,
    n77
  );


  buf
  g564
  (
    n604,
    n459
  );


  buf
  g565
  (
    n655,
    n495
  );


  buf
  g566
  (
    n638,
    n506
  );


  not
  g567
  (
    n668,
    n486
  );


  buf
  g568
  (
    n727,
    n472
  );


  buf
  g569
  (
    n565,
    n485
  );


  not
  g570
  (
    n681,
    n488
  );


  buf
  g571
  (
    n647,
    n294
  );


  buf
  g572
  (
    n556,
    n198
  );


  not
  g573
  (
    n767,
    n483
  );


  not
  g574
  (
    n667,
    n299
  );


  not
  g575
  (
    n724,
    n76
  );


  buf
  g576
  (
    n645,
    n470
  );


  not
  g577
  (
    n518,
    n76
  );


  buf
  g578
  (
    n729,
    n503
  );


  buf
  g579
  (
    n610,
    n487
  );


  not
  g580
  (
    n641,
    n496
  );


  buf
  g581
  (
    n546,
    n302
  );


  not
  g582
  (
    n642,
    n508
  );


  not
  g583
  (
    n694,
    n480
  );


  buf
  g584
  (
    n636,
    n499
  );


  not
  g585
  (
    n547,
    n197
  );


  buf
  g586
  (
    n684,
    n474
  );


  not
  g587
  (
    n707,
    n458
  );


  not
  g588
  (
    n539,
    n306
  );


  not
  g589
  (
    n673,
    n297
  );


  buf
  g590
  (
    n583,
    n501
  );


  buf
  g591
  (
    n689,
    n461
  );


  not
  g592
  (
    n649,
    n455
  );


  not
  g593
  (
    n617,
    n512
  );


  buf
  g594
  (
    n644,
    n514
  );


  not
  g595
  (
    n536,
    n474
  );


  not
  g596
  (
    n533,
    n485
  );


  buf
  g597
  (
    n643,
    n463
  );


  buf
  g598
  (
    n549,
    n460
  );


  buf
  g599
  (
    n715,
    n77
  );


  buf
  g600
  (
    n657,
    n462
  );


  not
  g601
  (
    n560,
    n25
  );


  not
  g602
  (
    n744,
    n506
  );


  buf
  g603
  (
    n570,
    n504
  );


  not
  g604
  (
    n670,
    n451
  );


  not
  g605
  (
    n582,
    n30
  );


  buf
  g606
  (
    n597,
    n480
  );


  buf
  g607
  (
    n624,
    n459
  );


  not
  g608
  (
    n697,
    n75
  );


  not
  g609
  (
    n678,
    n74
  );


  buf
  g610
  (
    n563,
    n510
  );


  not
  g611
  (
    n571,
    n196
  );


  not
  g612
  (
    n739,
    n463
  );


  buf
  g613
  (
    n593,
    n492
  );


  not
  g614
  (
    n705,
    n76
  );


  not
  g615
  (
    n756,
    n498
  );


  buf
  g616
  (
    n723,
    n469
  );


  buf
  g617
  (
    n738,
    n455
  );


  buf
  g618
  (
    n535,
    n31
  );


  not
  g619
  (
    n566,
    n29
  );


  buf
  g620
  (
    n559,
    n502
  );


  buf
  g621
  (
    n740,
    n453
  );


  not
  g622
  (
    n648,
    n490
  );


  not
  g623
  (
    n646,
    n484
  );


  not
  g624
  (
    n537,
    n511
  );


  not
  g625
  (
    n765,
    n477
  );


  not
  g626
  (
    n576,
    n463
  );


  not
  g627
  (
    n725,
    n197
  );


  buf
  g628
  (
    n639,
    n482
  );


  not
  g629
  (
    n688,
    n512
  );


  not
  g630
  (
    n735,
    n514
  );


  buf
  g631
  (
    n700,
    n481
  );


  not
  g632
  (
    n669,
    n464
  );


  not
  g633
  (
    n710,
    n464
  );


  not
  g634
  (
    n564,
    n303
  );


  buf
  g635
  (
    n616,
    n467
  );


  buf
  g636
  (
    n661,
    n451
  );


  buf
  g637
  (
    n579,
    n514
  );


  not
  g638
  (
    n693,
    n476
  );


  buf
  g639
  (
    n633,
    n493
  );


  not
  g640
  (
    n517,
    n198
  );


  buf
  g641
  (
    n581,
    n474
  );


  buf
  g642
  (
    n562,
    n195
  );


  not
  g643
  (
    n619,
    n509
  );


  not
  g644
  (
    n631,
    n468
  );


  not
  g645
  (
    n703,
    n472
  );


  not
  g646
  (
    n520,
    n507
  );


  buf
  g647
  (
    n585,
    n493
  );


  buf
  g648
  (
    n683,
    n451
  );


  not
  g649
  (
    n530,
    n293
  );


  not
  g650
  (
    n522,
    n483
  );


  not
  g651
  (
    n589,
    n472
  );


  buf
  g652
  (
    n768,
    n461
  );


  buf
  g653
  (
    n696,
    n490
  );


  buf
  g654
  (
    n629,
    n478
  );


  not
  g655
  (
    n680,
    n475
  );


  buf
  g656
  (
    n626,
    n295
  );


  buf
  g657
  (
    n764,
    n479
  );


  not
  g658
  (
    KeyWire_0_9,
    n508
  );


  buf
  g659
  (
    n596,
    n501
  );


  not
  g660
  (
    n692,
    n478
  );


  not
  g661
  (
    n706,
    n498
  );


  not
  g662
  (
    n528,
    n505
  );


  not
  g663
  (
    n730,
    n500
  );


  buf
  g664
  (
    n544,
    n458
  );


  not
  g665
  (
    n519,
    n477
  );


  not
  g666
  (
    n558,
    n463
  );


  not
  g667
  (
    n550,
    n494
  );


  buf
  g668
  (
    n714,
    n509
  );


  buf
  g669
  (
    n553,
    n28
  );


  not
  g670
  (
    n555,
    n467
  );


  not
  g671
  (
    n746,
    n454
  );


  not
  g672
  (
    n603,
    n492
  );


  buf
  g673
  (
    n653,
    n465
  );


  not
  g674
  (
    n545,
    n483
  );


  not
  g675
  (
    n607,
    n304
  );


  buf
  g676
  (
    n515,
    n486
  );


  not
  g677
  (
    n612,
    n481
  );


  not
  g678
  (
    n575,
    n195
  );


  buf
  g679
  (
    n716,
    n292
  );


  buf
  g680
  (
    n742,
    n74
  );


  buf
  g681
  (
    n672,
    n457
  );


  not
  g682
  (
    n618,
    n196
  );


  buf
  g683
  (
    n634,
    n453
  );


  not
  g684
  (
    n587,
    n307
  );


  not
  g685
  (
    n721,
    n458
  );


  buf
  g686
  (
    n675,
    n512
  );


  not
  g687
  (
    n737,
    n470
  );


  not
  g688
  (
    n602,
    n456
  );


  buf
  g689
  (
    n761,
    n476
  );


  buf
  g690
  (
    n719,
    n301
  );


  not
  g691
  (
    n695,
    n461
  );


  not
  g692
  (
    n609,
    n481
  );


  buf
  g693
  (
    n652,
    n500
  );


  buf
  g694
  (
    n529,
    n470
  );


  buf
  g695
  (
    n702,
    n499
  );


  buf
  g696
  (
    n598,
    n471
  );


  buf
  g697
  (
    n728,
    n464
  );


  not
  g698
  (
    n574,
    n459
  );


  buf
  g699
  (
    n568,
    n494
  );


  buf
  g700
  (
    n664,
    n197
  );


  not
  g701
  (
    n709,
    n502
  );


  not
  g702
  (
    n713,
    n75
  );


  not
  g703
  (
    n534,
    n476
  );


  buf
  g704
  (
    n572,
    n32
  );


  not
  g705
  (
    n516,
    n298
  );


  not
  g706
  (
    n595,
    n452
  );


  not
  g707
  (
    n734,
    n473
  );


  buf
  g708
  (
    n622,
    n480
  );


  buf
  g709
  (
    n561,
    n467
  );


  buf
  g710
  (
    n760,
    n456
  );


  not
  g711
  (
    n698,
    n485
  );


  not
  g712
  (
    KeyWire_0_2,
    n481
  );


  not
  g713
  (
    n640,
    n478
  );


  not
  g714
  (
    n632,
    n460
  );


  not
  g715
  (
    n651,
    n487
  );


  buf
  g716
  (
    n750,
    n487
  );


  buf
  g717
  (
    n754,
    n77
  );


  nor
  g718
  (
    n541,
    n469,
    n73,
    n491,
    n510
  );


  xor
  g719
  (
    n722,
    n507,
    n465,
    n497,
    n76
  );


  and
  g720
  (
    n551,
    n198,
    n482,
    n496,
    n465
  );


  and
  g721
  (
    n615,
    n475,
    n493,
    n497,
    n508
  );


  xor
  g722
  (
    n699,
    n489,
    n468,
    n471,
    n73
  );


  or
  g723
  (
    n552,
    n474,
    n488,
    n469,
    n485
  );


  xor
  g724
  (
    n654,
    n483,
    n495,
    n500,
    n499
  );


  nor
  g725
  (
    n543,
    n454,
    n495,
    n467,
    n502
  );


  or
  g726
  (
    n586,
    n484,
    n505,
    n459,
    n493
  );


  and
  g727
  (
    n540,
    n305,
    n504,
    n455,
    n513
  );


  nand
  g728
  (
    n613,
    n476,
    n475,
    n470,
    n452
  );


  xor
  g729
  (
    n627,
    n509,
    n501,
    n457,
    n495
  );


  nand
  g730
  (
    n687,
    n500,
    n511,
    n75,
    n513
  );


  nor
  g731
  (
    n711,
    n468,
    n473,
    n509
  );


  xnor
  g732
  (
    n770,
    n27,
    n501,
    n513,
    n458
  );


  nor
  g733
  (
    n757,
    n490,
    n487,
    n480,
    n503
  );


  nand
  g734
  (
    n660,
    n482,
    n512,
    n462,
    n72
  );


  or
  g735
  (
    n625,
    n75,
    n503,
    n479,
    n457
  );


  nand
  g736
  (
    n679,
    n73,
    n486,
    n471,
    n477
  );


  xnor
  g737
  (
    n605,
    n456,
    n486,
    n499,
    n510
  );


  and
  g738
  (
    n814,
    n664,
    n577,
    n599,
    n589
  );


  or
  g739
  (
    n772,
    n659,
    n656,
    n592,
    n572
  );


  or
  g740
  (
    n846,
    n576,
    n546,
    n557,
    n640
  );


  nor
  g741
  (
    n789,
    n665,
    n629,
    n660,
    n645
  );


  xnor
  g742
  (
    n825,
    n645,
    n646,
    n606,
    n627
  );


  xnor
  g743
  (
    n829,
    n549,
    n678,
    n614,
    n599
  );


  xnor
  g744
  (
    n833,
    n588,
    n680,
    n641,
    n645
  );


  and
  g745
  (
    n811,
    n605,
    n663,
    n638,
    n578
  );


  nand
  g746
  (
    n838,
    n667,
    n609,
    n642,
    n659
  );


  nor
  g747
  (
    n845,
    n600,
    n657,
    n635,
    n546
  );


  or
  g748
  (
    n824,
    n616,
    n647,
    n661,
    n615
  );


  xnor
  g749
  (
    n837,
    n578,
    n636,
    n610,
    n543
  );


  xor
  g750
  (
    n802,
    n531,
    n673,
    n627,
    n643
  );


  nand
  g751
  (
    n859,
    n677,
    n555,
    n628,
    n660
  );


  xor
  g752
  (
    n827,
    n667,
    n575,
    n675,
    n567
  );


  and
  g753
  (
    n832,
    n606,
    n653,
    n676,
    n658
  );


  and
  g754
  (
    n819,
    n672,
    n683,
    n678,
    n625
  );


  or
  g755
  (
    n790,
    n582,
    n576,
    n640,
    n631
  );


  or
  g756
  (
    n848,
    n654,
    n683,
    n670,
    n647
  );


  xor
  g757
  (
    n803,
    n662,
    n592,
    n556,
    n617
  );


  xor
  g758
  (
    n776,
    n550,
    n581,
    n594,
    n674
  );


  xnor
  g759
  (
    n796,
    n672,
    n601,
    n535,
    n551
  );


  nor
  g760
  (
    n852,
    n574,
    n593,
    n634,
    n644
  );


  nor
  g761
  (
    n795,
    n623,
    n668,
    n665,
    n515
  );


  and
  g762
  (
    n786,
    n560,
    n611,
    n521,
    n631
  );


  and
  g763
  (
    n821,
    n655,
    n641,
    n632,
    n616
  );


  xor
  g764
  (
    n783,
    n663,
    n524,
    n664,
    n613
  );


  nand
  g765
  (
    n847,
    n666,
    n552,
    n637,
    n580
  );


  and
  g766
  (
    n851,
    n607,
    n646,
    n632,
    n667
  );


  nand
  g767
  (
    n843,
    n598,
    n680,
    n679,
    n668
  );


  or
  g768
  (
    n773,
    n675,
    n650,
    n555,
    n534
  );


  nand
  g769
  (
    n777,
    n542,
    n647,
    n575,
    n635
  );


  xor
  g770
  (
    n807,
    n650,
    n639,
    n536,
    n652
  );


  and
  g771
  (
    n808,
    n570,
    n649,
    n594,
    n603
  );


  and
  g772
  (
    n775,
    n622,
    n671,
    n602,
    n583
  );


  nand
  g773
  (
    n817,
    n516,
    n564,
    n658,
    n597
  );


  or
  g774
  (
    n840,
    n584,
    n624,
    n556,
    n526
  );


  nand
  g775
  (
    n809,
    n527,
    n583,
    n625,
    n681
  );


  and
  g776
  (
    n850,
    n591,
    n669,
    n637,
    n642
  );


  xnor
  g777
  (
    n815,
    n655,
    n618,
    n681,
    n653
  );


  nor
  g778
  (
    n805,
    n644,
    n619,
    n682,
    n591
  );


  xor
  g779
  (
    n813,
    n581,
    n651,
    n654,
    n630
  );


  xor
  g780
  (
    n780,
    n657,
    n551,
    n607,
    n666
  );


  xor
  g781
  (
    n856,
    n611,
    n661,
    n680,
    n672
  );


  and
  g782
  (
    n828,
    n520,
    n610,
    n590,
    n585
  );


  xnor
  g783
  (
    n812,
    n668,
    n571,
    n646,
    n638
  );


  xor
  g784
  (
    n800,
    n544,
    n532,
    n614,
    n540
  );


  or
  g785
  (
    n781,
    n544,
    n655,
    n571,
    n609
  );


  xor
  g786
  (
    n853,
    n673,
    n604,
    n552,
    n559
  );


  nor
  g787
  (
    n834,
    n587,
    n605,
    n600,
    n678
  );


  nand
  g788
  (
    n836,
    n585,
    n563,
    n548,
    n619
  );


  xnor
  g789
  (
    n835,
    n626,
    n561,
    n517,
    n656
  );


  or
  g790
  (
    n782,
    n558,
    n622,
    n665,
    n580
  );


  nor
  g791
  (
    n854,
    n559,
    n621,
    n582,
    n670
  );


  xor
  g792
  (
    n842,
    n567,
    n620,
    n653,
    n577
  );


  xor
  g793
  (
    n793,
    n553,
    n633,
    n597,
    n523
  );


  xnor
  g794
  (
    KeyWire_0_6,
    n574,
    n545,
    n664,
    n643
  );


  xor
  g795
  (
    n788,
    n543,
    n595,
    n530,
    n658
  );


  xor
  g796
  (
    n787,
    n661,
    n677,
    n671
  );


  xnor
  g797
  (
    n822,
    n539,
    n626,
    n595,
    n637
  );


  and
  g798
  (
    n831,
    n548,
    n640,
    n615,
    n598
  );


  xnor
  g799
  (
    n816,
    n562,
    n650,
    n612
  );


  xnor
  g800
  (
    n844,
    n654,
    n589,
    n676,
    n620
  );


  and
  g801
  (
    n820,
    n679,
    n558,
    n549,
    n525
  );


  xnor
  g802
  (
    n826,
    n648,
    n670,
    n561,
    n566
  );


  xnor
  g803
  (
    n797,
    n519,
    n638,
    n533,
    n604
  );


  nand
  g804
  (
    n771,
    n584,
    n569,
    n590,
    n565
  );


  xnor
  g805
  (
    n857,
    n586,
    n643,
    n662,
    n679
  );


  xnor
  g806
  (
    n841,
    n677,
    n579,
    n565,
    n596
  );


  nand
  g807
  (
    n791,
    n621,
    n550,
    n663,
    n656
  );


  nor
  g808
  (
    n778,
    n639,
    n676,
    n596,
    n659
  );


  nand
  g809
  (
    n784,
    n568,
    n675,
    n613,
    n674
  );


  xor
  g810
  (
    n810,
    n562,
    n674,
    n518,
    n573
  );


  nand
  g811
  (
    n855,
    n648,
    n566,
    n560,
    n537
  );


  and
  g812
  (
    n839,
    n634,
    n554,
    n657,
    n617
  );


  xnor
  g813
  (
    n858,
    n660,
    n669,
    n545,
    n636
  );


  nor
  g814
  (
    n830,
    n587,
    n579,
    n608,
    n651
  );


  and
  g815
  (
    n823,
    n602,
    n623,
    n569,
    n529
  );


  xor
  g816
  (
    n801,
    n563,
    n593,
    n564,
    n642
  );


  xnor
  g817
  (
    n804,
    n633,
    n681,
    n662,
    n644
  );


  nand
  g818
  (
    n794,
    n648,
    n573,
    n641,
    n628
  );


  xnor
  g819
  (
    n792,
    n554,
    n528,
    n639,
    n557
  );


  nor
  g820
  (
    n785,
    n541,
    n649,
    n682,
    n586
  );


  nand
  g821
  (
    n779,
    n547,
    n652,
    n629,
    n588
  );


  xnor
  g822
  (
    n818,
    n624,
    n553,
    n572,
    n669
  );


  xor
  g823
  (
    n799,
    n608,
    n649,
    n603,
    n568
  );


  xor
  g824
  (
    n806,
    n538,
    n682,
    n601,
    n547
  );


  nand
  g825
  (
    n798,
    n651,
    n666,
    n522,
    n570
  );


  and
  g826
  (
    n849,
    n652,
    n618,
    n673,
    n630
  );


  or
  g827
  (
    n891,
    n778,
    n765,
    n780,
    n718
  );


  nand
  g828
  (
    n927,
    n767,
    n745,
    n759,
    n746
  );


  and
  g829
  (
    n937,
    n758,
    n738,
    n753,
    n685
  );


  nor
  g830
  (
    n944,
    n728,
    n718,
    n757,
    n733
  );


  xor
  g831
  (
    n881,
    n733,
    n836,
    n710,
    n776
  );


  nand
  g832
  (
    n864,
    n759,
    n784,
    n812,
    n746
  );


  nand
  g833
  (
    n870,
    n769,
    n722,
    n843,
    n810
  );


  xnor
  g834
  (
    n893,
    n760,
    n709,
    n773,
    n761
  );


  nand
  g835
  (
    n939,
    n714,
    n758,
    n838,
    n696
  );


  or
  g836
  (
    n863,
    n737,
    n749,
    n699,
    n734
  );


  and
  g837
  (
    n933,
    n837,
    n716,
    n723,
    n727
  );


  nor
  g838
  (
    n875,
    n804,
    n754,
    n697,
    n309
  );


  or
  g839
  (
    n925,
    n732,
    n701,
    n690,
    n809
  );


  nor
  g840
  (
    n890,
    n792,
    n744,
    n757,
    n716
  );


  xor
  g841
  (
    n922,
    n684,
    n855,
    n768,
    n737
  );


  xnor
  g842
  (
    n926,
    n714,
    n739,
    n732,
    n684
  );


  xnor
  g843
  (
    n935,
    n715,
    n777,
    n689,
    n736
  );


  xor
  g844
  (
    n869,
    n730,
    n689,
    n684,
    n758
  );


  xor
  g845
  (
    n880,
    n719,
    n748,
    n761,
    n750
  );


  xnor
  g846
  (
    n874,
    n841,
    n731,
    n692,
    n723
  );


  nand
  g847
  (
    n934,
    n852,
    n807,
    n785,
    n741
  );


  and
  g848
  (
    n919,
    n728,
    n765,
    n693,
    n831
  );


  nand
  g849
  (
    n887,
    n787,
    n729,
    n786,
    n707
  );


  xor
  g850
  (
    n883,
    n751,
    n742,
    n781,
    n805
  );


  or
  g851
  (
    n915,
    n693,
    n760,
    n772,
    n733
  );


  and
  g852
  (
    n888,
    n739,
    n740,
    n700,
    n686
  );


  nand
  g853
  (
    n886,
    n690,
    n706,
    n711,
    n695
  );


  xnor
  g854
  (
    n945,
    n710,
    n706,
    n794,
    n725
  );


  and
  g855
  (
    n866,
    n767,
    n692,
    n730,
    n683
  );


  xnor
  g856
  (
    n892,
    n691,
    n720,
    n749,
    n840
  );


  nor
  g857
  (
    n900,
    n705,
    n716,
    n751,
    n760
  );


  nand
  g858
  (
    n860,
    n842,
    n709,
    n820,
    n705
  );


  and
  g859
  (
    KeyWire_0_12,
    n698,
    n797,
    n802,
    n769
  );


  xor
  g860
  (
    n914,
    n795,
    n755,
    n791,
    n308
  );


  and
  g861
  (
    KeyWire_0_27,
    n700,
    n696,
    n762,
    n705
  );


  xnor
  g862
  (
    n907,
    n721,
    n821,
    n726,
    n708
  );


  xor
  g863
  (
    n876,
    n701,
    n762,
    n738,
    n686
  );


  xor
  g864
  (
    n889,
    n731,
    n717,
    n694,
    n713
  );


  nor
  g865
  (
    n868,
    n720,
    n763,
    n728,
    n813
  );


  xor
  g866
  (
    n912,
    n846,
    n719,
    n691,
    n844
  );


  nand
  g867
  (
    n862,
    n694,
    n729,
    n828,
    n847
  );


  nor
  g868
  (
    n931,
    n718,
    n747,
    n775,
    n713
  );


  and
  g869
  (
    n923,
    n732,
    n708,
    n712,
    n721
  );


  nor
  g870
  (
    n896,
    n762,
    n737,
    n720,
    n695
  );


  nand
  g871
  (
    n905,
    n688,
    n736,
    n750
  );


  or
  g872
  (
    n930,
    n761,
    n722,
    n738,
    n825
  );


  nor
  g873
  (
    n936,
    n699,
    n752,
    n696,
    n735
  );


  xnor
  g874
  (
    n942,
    n814,
    n744,
    n709,
    n751
  );


  or
  g875
  (
    n909,
    n748,
    n796,
    n764,
    n707
  );


  and
  g876
  (
    n885,
    n726,
    n687,
    n702,
    n723
  );


  xor
  g877
  (
    n941,
    n856,
    n755,
    n770,
    n753
  );


  xnor
  g878
  (
    n917,
    n815,
    n685,
    n703,
    n694
  );


  and
  g879
  (
    n871,
    n745,
    n734,
    n853,
    n727
  );


  nor
  g880
  (
    n882,
    n789,
    n806,
    n755,
    n748
  );


  xor
  g881
  (
    n918,
    n747,
    n727,
    n746,
    n744
  );


  xor
  g882
  (
    n867,
    n801,
    n749,
    n690,
    n702
  );


  nand
  g883
  (
    n899,
    n754,
    n712,
    n756,
    n835
  );


  nor
  g884
  (
    n940,
    n717,
    n817,
    n800,
    n730
  );


  nor
  g885
  (
    n943,
    n703,
    n763,
    n857,
    n745
  );


  xor
  g886
  (
    n910,
    n700,
    n743,
    n689,
    n783
  );


  nand
  g887
  (
    n895,
    n767,
    n724,
    n829,
    n729
  );


  nor
  g888
  (
    n947,
    n803,
    n743,
    n739,
    n687
  );


  xnor
  g889
  (
    n894,
    n717,
    n808,
    n747,
    n713
  );


  xor
  g890
  (
    n921,
    n698,
    n798,
    n764,
    n845
  );


  nand
  g891
  (
    n884,
    n714,
    n704,
    n706,
    n830
  );


  xnor
  g892
  (
    n865,
    n691,
    n768,
    n763,
    n698
  );


  xnor
  g893
  (
    n916,
    n740,
    n759,
    n811,
    n766
  );


  and
  g894
  (
    n913,
    n799,
    n771,
    n743,
    n725
  );


  nor
  g895
  (
    n898,
    n833,
    n742,
    n816,
    n858
  );


  nand
  g896
  (
    n902,
    n765,
    n752,
    n715,
    n768
  );


  nand
  g897
  (
    n932,
    n697,
    n711,
    n753,
    n721
  );


  xor
  g898
  (
    n911,
    n707,
    n699,
    n782,
    n686
  );


  or
  g899
  (
    n938,
    n710,
    n724,
    n793,
    n708
  );


  xnor
  g900
  (
    n861,
    n726,
    n766,
    n764,
    n701
  );


  or
  g901
  (
    n873,
    n823,
    n822,
    n849,
    n754
  );


  and
  g902
  (
    n904,
    n824,
    n834,
    n687,
    n854
  );


  nor
  g903
  (
    n872,
    n779,
    n756,
    n725,
    n851
  );


  and
  g904
  (
    n924,
    n715,
    n688,
    n741,
    n736
  );


  xnor
  g905
  (
    n877,
    n719,
    n770,
    n826,
    n704
  );


  nand
  g906
  (
    n878,
    n766,
    n819,
    n695,
    n769
  );


  xnor
  g907
  (
    n946,
    n688,
    n790,
    n774,
    n818
  );


  and
  g908
  (
    n879,
    n703,
    n685,
    n735
  );


  or
  g909
  (
    n897,
    n722,
    n832,
    n697,
    n742
  );


  xor
  g910
  (
    n929,
    n740,
    n724,
    n712,
    n693
  );


  and
  g911
  (
    n901,
    n752,
    n692,
    n770,
    n704
  );


  xnor
  g912
  (
    n906,
    n788,
    n757,
    n850,
    n702
  );


  nor
  g913
  (
    n903,
    n839,
    n756,
    n848,
    n827
  );


  nand
  g914
  (
    n928,
    n734,
    n711,
    n731,
    n741
  );


  nor
  g915
  (
    n948,
    n863,
    n887
  );


  xor
  g916
  (
    n966,
    n312,
    n913,
    n906,
    n864
  );


  nor
  g917
  (
    n955,
    n903,
    n893,
    n920,
    n871
  );


  or
  g918
  (
    n954,
    n899,
    n869,
    n884,
    n859
  );


  xnor
  g919
  (
    n950,
    n877,
    n892,
    n888,
    n919
  );


  nand
  g920
  (
    n951,
    n911,
    n894,
    n881,
    n323
  );


  or
  g921
  (
    n959,
    n311,
    n918,
    n862,
    n880
  );


  xnor
  g922
  (
    n949,
    n872,
    n319,
    n313,
    n909
  );


  nor
  g923
  (
    n953,
    n905,
    n898,
    n895,
    n901
  );


  xor
  g924
  (
    n956,
    n883,
    n916,
    n890,
    n912
  );


  or
  g925
  (
    n952,
    n318,
    n882,
    n878,
    n907
  );


  xnor
  g926
  (
    n962,
    n876,
    n897,
    n896,
    n873
  );


  or
  g927
  (
    n964,
    n868,
    n885,
    n886,
    n910
  );


  xnor
  g928
  (
    n957,
    n317,
    n320,
    n875,
    n321
  );


  xnor
  g929
  (
    n963,
    n325,
    n915,
    n914,
    n902
  );


  nand
  g930
  (
    n960,
    n314,
    n917,
    n879,
    n860
  );


  xor
  g931
  (
    n958,
    n900,
    n866,
    n324,
    n889
  );


  and
  g932
  (
    n961,
    n316,
    n865,
    n867,
    n908
  );


  or
  g933
  (
    n965,
    n874,
    n891,
    n315,
    n310
  );


  or
  g934
  (
    n967,
    n322,
    n861,
    n904,
    n870
  );


  or
  g935
  (
    n973,
    n939,
    n926,
    n921,
    n944
  );


  xor
  g936
  (
    n969,
    n923,
    n942,
    n966,
    n954
  );


  xnor
  g937
  (
    n979,
    n966,
    n934,
    n940
  );


  xnor
  g938
  (
    n981,
    n963,
    n967,
    n941,
    n929
  );


  nor
  g939
  (
    n983,
    n939,
    n937,
    n944,
    n943
  );


  and
  g940
  (
    n989,
    n931,
    n965,
    n944,
    n938
  );


  nand
  g941
  (
    n970,
    n941,
    n936,
    n937,
    n924
  );


  xnor
  g942
  (
    n978,
    n947,
    n950,
    n967,
    n946
  );


  or
  g943
  (
    n984,
    n927,
    n930,
    n962,
    n964
  );


  and
  g944
  (
    n971,
    n956,
    n943,
    n959,
    n935
  );


  xnor
  g945
  (
    n976,
    n942,
    n960,
    n945,
    n941
  );


  xor
  g946
  (
    n988,
    n939,
    n957,
    n925,
    n947
  );


  xnor
  g947
  (
    n987,
    n939,
    n935,
    n933,
    n945
  );


  or
  g948
  (
    n986,
    n937,
    n949,
    n936,
    n935
  );


  and
  g949
  (
    n975,
    n943,
    n936,
    n945,
    n938
  );


  or
  g950
  (
    n982,
    n951,
    n932,
    n946
  );


  or
  g951
  (
    n968,
    n953,
    n938,
    n946
  );


  xnor
  g952
  (
    n972,
    n922,
    n941,
    n948,
    n952
  );


  and
  g953
  (
    n985,
    n928,
    n961,
    n942,
    n936
  );


  or
  g954
  (
    n977,
    n937,
    n947,
    n944,
    n945
  );


  nor
  g955
  (
    n974,
    n935,
    n940,
    n947,
    n958
  );


  xor
  g956
  (
    n980,
    n940,
    n955,
    n942,
    n943
  );


  not
  g957
  (
    n1069,
    n974
  );


  buf
  g958
  (
    n1053,
    n970
  );


  buf
  g959
  (
    n1008,
    n986
  );


  buf
  g960
  (
    n1034,
    n975
  );


  buf
  g961
  (
    n1006,
    n980
  );


  buf
  g962
  (
    n1022,
    n979
  );


  buf
  g963
  (
    n1000,
    n972
  );


  buf
  g964
  (
    n1050,
    n972
  );


  buf
  g965
  (
    n1031,
    n974
  );


  not
  g966
  (
    n1068,
    n974
  );


  buf
  g967
  (
    n998,
    n980
  );


  buf
  g968
  (
    n1035,
    n986
  );


  buf
  g969
  (
    n1057,
    n968
  );


  buf
  g970
  (
    KeyWire_0_19,
    n988
  );


  buf
  g971
  (
    n1064,
    n968
  );


  not
  g972
  (
    n1047,
    n982
  );


  buf
  g973
  (
    n994,
    n971
  );


  not
  g974
  (
    n1012,
    n980
  );


  buf
  g975
  (
    n1045,
    n976
  );


  buf
  g976
  (
    n1071,
    n978
  );


  buf
  g977
  (
    n1015,
    n985
  );


  not
  g978
  (
    n1017,
    n969
  );


  not
  g979
  (
    n1032,
    n973
  );


  not
  g980
  (
    n1016,
    n982
  );


  not
  g981
  (
    n992,
    n986
  );


  buf
  g982
  (
    n1048,
    n983
  );


  not
  g983
  (
    n1063,
    n976
  );


  buf
  g984
  (
    n1067,
    n983
  );


  not
  g985
  (
    n1043,
    n978
  );


  buf
  g986
  (
    n1058,
    n982
  );


  not
  g987
  (
    n1036,
    n987
  );


  buf
  g988
  (
    n1028,
    n987
  );


  not
  g989
  (
    n990,
    n971
  );


  buf
  g990
  (
    n1054,
    n987
  );


  not
  g991
  (
    n1023,
    n986
  );


  buf
  g992
  (
    n1051,
    n985
  );


  buf
  g993
  (
    n996,
    n981
  );


  buf
  g994
  (
    n1007,
    n981
  );


  not
  g995
  (
    n1070,
    n968
  );


  not
  g996
  (
    KeyWire_0_11,
    n983
  );


  not
  g997
  (
    n1049,
    n982
  );


  buf
  g998
  (
    n999,
    n972
  );


  buf
  g999
  (
    n1030,
    n979
  );


  buf
  g1000
  (
    n991,
    n970
  );


  buf
  g1001
  (
    n1065,
    n973
  );


  buf
  g1002
  (
    n1005,
    n975
  );


  buf
  g1003
  (
    KeyWire_0_24,
    n975
  );


  not
  g1004
  (
    n1044,
    n326
  );


  not
  g1005
  (
    n1042,
    n978
  );


  not
  g1006
  (
    n1025,
    n977
  );


  not
  g1007
  (
    n1018,
    n974
  );


  buf
  g1008
  (
    n1062,
    n971
  );


  not
  g1009
  (
    n993,
    n968
  );


  not
  g1010
  (
    n1060,
    n969
  );


  buf
  g1011
  (
    n1038,
    n984
  );


  not
  g1012
  (
    n1014,
    n977
  );


  buf
  g1013
  (
    n1001,
    n988
  );


  buf
  g1014
  (
    n1046,
    n977
  );


  buf
  g1015
  (
    n1013,
    n978
  );


  not
  g1016
  (
    n1021,
    n973
  );


  buf
  g1017
  (
    n1026,
    n981
  );


  buf
  g1018
  (
    n1024,
    n969
  );


  not
  g1019
  (
    n1002,
    n973
  );


  not
  g1020
  (
    n1009,
    n977
  );


  buf
  g1021
  (
    n1029,
    n969
  );


  not
  g1022
  (
    n1059,
    n971
  );


  buf
  g1023
  (
    n995,
    n970
  );


  not
  g1024
  (
    n1020,
    n984
  );


  not
  g1025
  (
    n1019,
    n980
  );


  not
  g1026
  (
    n1039,
    n976
  );


  not
  g1027
  (
    n997,
    n976
  );


  buf
  g1028
  (
    n1052,
    n970
  );


  not
  g1029
  (
    n1004,
    n984
  );


  not
  g1030
  (
    n1041,
    n327
  );


  buf
  g1031
  (
    n1037,
    n981
  );


  not
  g1032
  (
    n1011,
    n979
  );


  not
  g1033
  (
    n1027,
    n979
  );


  not
  g1034
  (
    n1033,
    n987
  );


  buf
  g1035
  (
    n1055,
    n972
  );


  buf
  g1036
  (
    n1003,
    n975
  );


  not
  g1037
  (
    n1010,
    n985
  );


  nand
  g1038
  (
    n1066,
    n983,
    n984
  );


  not
  g1039
  (
    n1072,
    n1005
  );


  not
  g1040
  (
    n1077,
    n1025
  );


  not
  g1041
  (
    n1094,
    n1007
  );


  buf
  g1042
  (
    n1086,
    n1009
  );


  not
  g1043
  (
    n1134,
    n1028
  );


  buf
  g1044
  (
    n1107,
    n1025
  );


  not
  g1045
  (
    n1127,
    n336
  );


  not
  g1046
  (
    n1113,
    n1026
  );


  not
  g1047
  (
    n1073,
    n1015
  );


  buf
  g1048
  (
    n1089,
    n1028
  );


  buf
  g1049
  (
    n1117,
    n1023
  );


  buf
  g1050
  (
    n1088,
    n1011
  );


  not
  g1051
  (
    n1110,
    n1007
  );


  not
  g1052
  (
    n1091,
    n1019
  );


  not
  g1053
  (
    n1135,
    n338
  );


  not
  g1054
  (
    n1114,
    n988
  );


  buf
  g1055
  (
    n1112,
    n1007
  );


  buf
  g1056
  (
    n1078,
    n1018
  );


  buf
  g1057
  (
    n1100,
    n1008
  );


  not
  g1058
  (
    n1121,
    n1024
  );


  not
  g1059
  (
    n1079,
    n1015
  );


  not
  g1060
  (
    n1109,
    n1027
  );


  not
  g1061
  (
    n1075,
    n1017
  );


  not
  g1062
  (
    n1129,
    n1012
  );


  buf
  g1063
  (
    n1074,
    n989
  );


  not
  g1064
  (
    n1098,
    n1017
  );


  not
  g1065
  (
    n1092,
    n337
  );


  buf
  g1066
  (
    n1095,
    n1011
  );


  not
  g1067
  (
    n1083,
    n1012
  );


  not
  g1068
  (
    n1103,
    n1022
  );


  not
  g1069
  (
    n1093,
    n1022
  );


  not
  g1070
  (
    n1124,
    n331
  );


  buf
  g1071
  (
    n1118,
    n1006
  );


  not
  g1072
  (
    n1106,
    n1016
  );


  buf
  g1073
  (
    n1097,
    n1009
  );


  buf
  g1074
  (
    n1130,
    n1021
  );


  not
  g1075
  (
    n1101,
    n339
  );


  buf
  g1076
  (
    n1082,
    n1008
  );


  not
  g1077
  (
    n1105,
    n1027
  );


  buf
  g1078
  (
    n1115,
    n1014
  );


  not
  g1079
  (
    n1080,
    n988
  );


  not
  g1080
  (
    n1119,
    n1026
  );


  not
  g1081
  (
    n1120,
    n1019
  );


  not
  g1082
  (
    n1111,
    n1024
  );


  buf
  g1083
  (
    n1132,
    n335
  );


  not
  g1084
  (
    n1102,
    n333
  );


  buf
  g1085
  (
    n1099,
    n1022
  );


  buf
  g1086
  (
    n1123,
    n340
  );


  buf
  g1087
  (
    n1104,
    n1026
  );


  not
  g1088
  (
    n1085,
    n1013
  );


  buf
  g1089
  (
    n1084,
    n330
  );


  not
  g1090
  (
    n1087,
    n1028
  );


  not
  g1091
  (
    n1122,
    n1008
  );


  buf
  g1092
  (
    n1125,
    n1015
  );


  nand
  g1093
  (
    n1076,
    n1020,
    n1013
  );


  xnor
  g1094
  (
    n1090,
    n1027,
    n1010
  );


  xnor
  g1095
  (
    n1096,
    n1011,
    n1009,
    n1016,
    n341
  );


  nand
  g1096
  (
    n1133,
    n1014,
    n1020,
    n1021
  );


  xnor
  g1097
  (
    n1081,
    n1018,
    n1029,
    n1023,
    n1010
  );


  or
  g1098
  (
    n1116,
    n1014,
    n989,
    n332,
    n1010
  );


  xor
  g1099
  (
    n1126,
    n1017,
    n1023,
    n1019,
    n1018
  );


  xor
  g1100
  (
    n1131,
    n1012,
    n1013,
    n334,
    n328
  );


  xor
  g1101
  (
    n1128,
    n1016,
    n342,
    n329,
    n1024
  );


  xnor
  g1102
  (
    n1108,
    n1020,
    n1025,
    n989
  );


  buf
  g1103
  (
    n1216,
    n1096
  );


  buf
  g1104
  (
    n1278,
    n1117
  );


  buf
  g1105
  (
    n1371,
    n1099
  );


  buf
  g1106
  (
    n1212,
    n1110
  );


  not
  g1107
  (
    n1148,
    n1125
  );


  not
  g1108
  (
    n1230,
    n1054
  );


  buf
  g1109
  (
    n1286,
    n1101
  );


  buf
  g1110
  (
    n1391,
    n1095
  );


  buf
  g1111
  (
    n1307,
    n1043
  );


  buf
  g1112
  (
    n1163,
    n1066
  );


  not
  g1113
  (
    n1143,
    n1134
  );


  not
  g1114
  (
    n1218,
    n1115
  );


  not
  g1115
  (
    n1138,
    n1090
  );


  buf
  g1116
  (
    n1352,
    n1063
  );


  not
  g1117
  (
    n1267,
    n1091
  );


  not
  g1118
  (
    n1388,
    n1072
  );


  buf
  g1119
  (
    n1320,
    n1098
  );


  buf
  g1120
  (
    n1187,
    n1061
  );


  buf
  g1121
  (
    n1289,
    n1116
  );


  not
  g1122
  (
    n1231,
    n1064
  );


  buf
  g1123
  (
    n1275,
    n1089
  );


  not
  g1124
  (
    n1342,
    n1118
  );


  buf
  g1125
  (
    n1324,
    n1100
  );


  buf
  g1126
  (
    n1246,
    n1103
  );


  buf
  g1127
  (
    n1260,
    n1080
  );


  not
  g1128
  (
    n1338,
    n1084
  );


  not
  g1129
  (
    n1377,
    n1075
  );


  not
  g1130
  (
    n1271,
    n1087
  );


  not
  g1131
  (
    n1169,
    n1077
  );


  buf
  g1132
  (
    n1345,
    n1133
  );


  not
  g1133
  (
    n1259,
    n1128
  );


  not
  g1134
  (
    n1217,
    n1083
  );


  not
  g1135
  (
    n1195,
    n1065
  );


  not
  g1136
  (
    n1257,
    n1049
  );


  not
  g1137
  (
    n1334,
    n1029
  );


  not
  g1138
  (
    n1379,
    n1129
  );


  buf
  g1139
  (
    n1319,
    n1067
  );


  buf
  g1140
  (
    n1198,
    n1069
  );


  buf
  g1141
  (
    KeyWire_0_25,
    n1111
  );


  not
  g1142
  (
    n1165,
    n1075
  );


  buf
  g1143
  (
    n1242,
    n1085
  );


  not
  g1144
  (
    n1375,
    n1105
  );


  not
  g1145
  (
    n1317,
    n1128
  );


  not
  g1146
  (
    n1144,
    n1106
  );


  buf
  g1147
  (
    n1224,
    n1132
  );


  not
  g1148
  (
    n1177,
    n1069
  );


  not
  g1149
  (
    n1327,
    n1070
  );


  buf
  g1150
  (
    n1347,
    n1083
  );


  not
  g1151
  (
    n1350,
    n1081
  );


  buf
  g1152
  (
    n1321,
    n1097
  );


  buf
  g1153
  (
    n1378,
    n1124
  );


  buf
  g1154
  (
    n1182,
    n1042
  );


  not
  g1155
  (
    n1383,
    n1091
  );


  not
  g1156
  (
    n1213,
    n1114
  );


  buf
  g1157
  (
    n1190,
    n1109
  );


  not
  g1158
  (
    n1156,
    n1088
  );


  buf
  g1159
  (
    n1263,
    n1093
  );


  buf
  g1160
  (
    n1185,
    n1060
  );


  buf
  g1161
  (
    n1237,
    n1032
  );


  not
  g1162
  (
    n1358,
    n1033
  );


  not
  g1163
  (
    n1316,
    n1099
  );


  not
  g1164
  (
    n1179,
    n1085
  );


  not
  g1165
  (
    n1219,
    n1046
  );


  not
  g1166
  (
    n1174,
    n1055
  );


  not
  g1167
  (
    n1244,
    n1131
  );


  buf
  g1168
  (
    n1243,
    n1110
  );


  not
  g1169
  (
    n1227,
    n1096
  );


  buf
  g1170
  (
    n1290,
    n1093
  );


  buf
  g1171
  (
    n1204,
    n1064
  );


  not
  g1172
  (
    n1239,
    n1033
  );


  buf
  g1173
  (
    n1283,
    n1045
  );


  not
  g1174
  (
    n1149,
    n1036
  );


  buf
  g1175
  (
    n1329,
    n1065
  );


  buf
  g1176
  (
    n1344,
    n1109
  );


  buf
  g1177
  (
    n1184,
    n1125
  );


  buf
  g1178
  (
    n1155,
    n1056
  );


  not
  g1179
  (
    n1372,
    n1107
  );


  buf
  g1180
  (
    n1252,
    n1115
  );


  not
  g1181
  (
    n1340,
    n1107
  );


  not
  g1182
  (
    n1390,
    n1094
  );


  buf
  g1183
  (
    n1168,
    n1057
  );


  not
  g1184
  (
    n1296,
    n1134
  );


  not
  g1185
  (
    n1364,
    n1096
  );


  buf
  g1186
  (
    n1308,
    n1030
  );


  not
  g1187
  (
    n1247,
    n1035
  );


  not
  g1188
  (
    n1311,
    n1124
  );


  not
  g1189
  (
    n1199,
    n1101
  );


  not
  g1190
  (
    n1203,
    n1073
  );


  not
  g1191
  (
    n1282,
    n1082
  );


  not
  g1192
  (
    n1233,
    n1047
  );


  buf
  g1193
  (
    n1147,
    n1111
  );


  buf
  g1194
  (
    n1200,
    n1054
  );


  not
  g1195
  (
    n1336,
    n1077
  );


  not
  g1196
  (
    n1280,
    n1127
  );


  not
  g1197
  (
    n1245,
    n1112
  );


  not
  g1198
  (
    KeyWire_0_29,
    n1105
  );


  not
  g1199
  (
    n1248,
    n1050
  );


  buf
  g1200
  (
    n1380,
    n1127
  );


  buf
  g1201
  (
    n1370,
    n1073
  );


  not
  g1202
  (
    n1140,
    n1115
  );


  buf
  g1203
  (
    n1258,
    n1086
  );


  buf
  g1204
  (
    n1303,
    n1031
  );


  not
  g1205
  (
    n1356,
    n1029
  );


  not
  g1206
  (
    n1226,
    n1045
  );


  not
  g1207
  (
    n1173,
    n1112
  );


  not
  g1208
  (
    KeyWire_0_5,
    n1061
  );


  buf
  g1209
  (
    n1207,
    n1074
  );


  not
  g1210
  (
    n1305,
    n1084
  );


  not
  g1211
  (
    n1285,
    n1121
  );


  not
  g1212
  (
    n1254,
    n1117
  );


  not
  g1213
  (
    n1201,
    n1042
  );


  not
  g1214
  (
    n1152,
    n1123
  );


  buf
  g1215
  (
    n1297,
    n1114
  );


  buf
  g1216
  (
    n1314,
    n1031
  );


  not
  g1217
  (
    n1181,
    n1079
  );


  not
  g1218
  (
    n1274,
    n1127
  );


  buf
  g1219
  (
    n1145,
    n1118
  );


  not
  g1220
  (
    n1310,
    n1122
  );


  not
  g1221
  (
    n1295,
    n1076
  );


  not
  g1222
  (
    n1313,
    n1097
  );


  buf
  g1223
  (
    n1291,
    n1089
  );


  not
  g1224
  (
    n1272,
    n1083
  );


  buf
  g1225
  (
    n1229,
    n1082
  );


  buf
  g1226
  (
    n1360,
    n1051
  );


  not
  g1227
  (
    n1381,
    n1041
  );


  not
  g1228
  (
    n1193,
    n1076
  );


  not
  g1229
  (
    n1157,
    n1109
  );


  buf
  g1230
  (
    n1228,
    n1089
  );


  buf
  g1231
  (
    n1359,
    n1049
  );


  buf
  g1232
  (
    n1170,
    n1078
  );


  not
  g1233
  (
    n1137,
    n1135
  );


  not
  g1234
  (
    n1172,
    n1078
  );


  buf
  g1235
  (
    n1374,
    n1053
  );


  buf
  g1236
  (
    n1269,
    n1038
  );


  not
  g1237
  (
    n1234,
    n1126
  );


  buf
  g1238
  (
    n1273,
    n1095
  );


  buf
  g1239
  (
    n1264,
    n1051
  );


  not
  g1240
  (
    n1365,
    n1044
  );


  buf
  g1241
  (
    n1222,
    n1135
  );


  buf
  g1242
  (
    n1196,
    n1075
  );


  not
  g1243
  (
    n1176,
    n1052
  );


  not
  g1244
  (
    n1141,
    n1084
  );


  not
  g1245
  (
    n1387,
    n1091
  );


  not
  g1246
  (
    n1266,
    n1033
  );


  buf
  g1247
  (
    n1343,
    n1066
  );


  not
  g1248
  (
    n1232,
    n1102
  );


  buf
  g1249
  (
    n1241,
    n1104
  );


  buf
  g1250
  (
    n1349,
    n1034
  );


  not
  g1251
  (
    n1180,
    n1050
  );


  not
  g1252
  (
    n1281,
    n1122
  );


  not
  g1253
  (
    n1151,
    n1054
  );


  not
  g1254
  (
    n1209,
    n1087
  );


  not
  g1255
  (
    n1178,
    n1047
  );


  buf
  g1256
  (
    n1205,
    n349
  );


  buf
  g1257
  (
    n1315,
    n344
  );


  not
  g1258
  (
    n1253,
    n1102
  );


  not
  g1259
  (
    n1183,
    n1094
  );


  buf
  g1260
  (
    n1136,
    n1100
  );


  buf
  g1261
  (
    n1197,
    n1098
  );


  not
  g1262
  (
    n1366,
    n1107
  );


  not
  g1263
  (
    n1382,
    n1039
  );


  buf
  g1264
  (
    n1146,
    n1103
  );


  not
  g1265
  (
    n1223,
    n1058
  );


  buf
  g1266
  (
    n1309,
    n1059
  );


  buf
  g1267
  (
    n1322,
    n1061
  );


  not
  g1268
  (
    n1154,
    n1059
  );


  buf
  g1269
  (
    n1357,
    n1104
  );


  buf
  g1270
  (
    n1348,
    n1072
  );


  buf
  g1271
  (
    n1268,
    n1058
  );


  buf
  g1272
  (
    n1368,
    n1073
  );


  not
  g1273
  (
    n1206,
    n1128
  );


  buf
  g1274
  (
    n1256,
    n1081
  );


  not
  g1275
  (
    n1188,
    n1116
  );


  buf
  g1276
  (
    n1270,
    n1043
  );


  buf
  g1277
  (
    n1159,
    n1086
  );


  buf
  g1278
  (
    n1214,
    n1102
  );


  not
  g1279
  (
    n1367,
    n1063
  );


  not
  g1280
  (
    n1335,
    n1052
  );


  not
  g1281
  (
    n1300,
    n1090
  );


  buf
  g1282
  (
    n1162,
    n1035
  );


  buf
  g1283
  (
    n1220,
    n1133
  );


  buf
  g1284
  (
    n1221,
    n1067
  );


  not
  g1285
  (
    n1384,
    n1069
  );


  buf
  g1286
  (
    n1279,
    n1119
  );


  not
  g1287
  (
    n1353,
    n1041
  );


  buf
  g1288
  (
    n1277,
    n1056
  );


  not
  g1289
  (
    n1208,
    n1113
  );


  buf
  g1290
  (
    n1331,
    n1120
  );


  not
  g1291
  (
    n1328,
    n1130
  );


  not
  g1292
  (
    n1301,
    n1062
  );


  not
  g1293
  (
    n1158,
    n1096
  );


  not
  g1294
  (
    n1330,
    n1129
  );


  buf
  g1295
  (
    n1139,
    n1115
  );


  buf
  g1296
  (
    n1189,
    n1132
  );


  buf
  g1297
  (
    n1255,
    n1129
  );


  buf
  g1298
  (
    n1302,
    n1072
  );


  buf
  g1299
  (
    n1351,
    n1077
  );


  buf
  g1300
  (
    n1293,
    n1100
  );


  buf
  g1301
  (
    n1164,
    n1112
  );


  not
  g1302
  (
    n1265,
    n1118
  );


  buf
  g1303
  (
    n1153,
    n1128
  );


  not
  g1304
  (
    n1261,
    n1070
  );


  buf
  g1305
  (
    n1171,
    n1050
  );


  not
  g1306
  (
    n1341,
    n1068
  );


  buf
  g1307
  (
    n1262,
    n1119
  );


  not
  g1308
  (
    n1211,
    n1106
  );


  not
  g1309
  (
    n1373,
    n1126
  );


  buf
  g1310
  (
    n1376,
    n1060
  );


  not
  g1311
  (
    n1160,
    n1101
  );


  not
  g1312
  (
    n1210,
    n1088
  );


  buf
  g1313
  (
    n1304,
    n1068
  );


  and
  g1314
  (
    n1249,
    n1082,
    n1117,
    n1121,
    n1056
  );


  or
  g1315
  (
    n1276,
    n1103,
    n1037,
    n1074,
    n1092
  );


  or
  g1316
  (
    n1332,
    n1053,
    n1118,
    n1130,
    n1037
  );


  and
  g1317
  (
    n1385,
    n1078,
    n1055,
    n1119,
    n1080
  );


  nand
  g1318
  (
    n1215,
    n1058,
    n1075,
    n1040,
    n1120
  );


  nand
  g1319
  (
    n1288,
    n1094,
    n1130,
    n1102,
    n1105
  );


  xnor
  g1320
  (
    n1362,
    n1100,
    n1106,
    n1066,
    n1120
  );


  and
  g1321
  (
    n1251,
    n1089,
    n1080,
    n1062
  );


  xor
  g1322
  (
    n1363,
    n1114,
    n1135,
    n1036,
    n1133
  );


  nor
  g1323
  (
    n1337,
    n1063,
    n1076,
    n1123,
    n1065
  );


  xnor
  g1324
  (
    n1150,
    n1072,
    n1104,
    n1051,
    n1068
  );


  and
  g1325
  (
    n1292,
    n1041,
    n1122,
    n1107,
    n1095
  );


  nor
  g1326
  (
    n1339,
    n1113,
    n1124,
    n1049,
    n1104
  );


  nand
  g1327
  (
    KeyWire_0_22,
    n1081,
    n1090,
    n1101,
    n1126
  );


  and
  g1328
  (
    n1238,
    n1048,
    n1032,
    n1079,
    n1123
  );


  xnor
  g1329
  (
    n1192,
    n1125,
    n1133,
    n1074,
    n1099
  );


  nand
  g1330
  (
    n1225,
    n1038,
    n1052,
    n1122,
    n1108
  );


  nand
  g1331
  (
    n1312,
    n1126,
    n1036,
    n1046,
    n343
  );


  and
  g1332
  (
    n1240,
    n1135,
    n1079,
    n1123,
    n1076
  );


  nand
  g1333
  (
    n1202,
    n347,
    n1073,
    n1132,
    n1092
  );


  and
  g1334
  (
    n1298,
    n345,
    n1087,
    n1117,
    n1039
  );


  xor
  g1335
  (
    n1323,
    n1034,
    n1044,
    n1071,
    n1113
  );


  nor
  g1336
  (
    n1299,
    n1047,
    n1044,
    n1053,
    n1091
  );


  xor
  g1337
  (
    n1333,
    n1090,
    n1111,
    n1098
  );


  xor
  g1338
  (
    n1287,
    n1116,
    n1094,
    n1105,
    n1030
  );


  nand
  g1339
  (
    n1236,
    n1092,
    n1083,
    n1037,
    n1125
  );


  nor
  g1340
  (
    n1191,
    n1132,
    n1110,
    n1098,
    n1086
  );


  xnor
  g1341
  (
    n1294,
    n1067,
    n346,
    n1062,
    n1042
  );


  nand
  g1342
  (
    n1326,
    n1088,
    n1046,
    n1035,
    n1134
  );


  xnor
  g1343
  (
    n1161,
    n1131,
    n1070,
    n1059,
    n1093
  );


  nand
  g1344
  (
    n1306,
    n1130,
    n1131,
    n1127,
    n1129
  );


  or
  g1345
  (
    n1325,
    n1119,
    n1030,
    n1057,
    n1124
  );


  nand
  g1346
  (
    n1318,
    n1064,
    n1108,
    n1040,
    n1048
  );


  nor
  g1347
  (
    n1284,
    n1110,
    n1108,
    n1121,
    n1116
  );


  xor
  g1348
  (
    n1250,
    n1131,
    n1097,
    n1114,
    n1071
  );


  nor
  g1349
  (
    n1166,
    n1109,
    n1031,
    n1055,
    n1074
  );


  or
  g1350
  (
    n1354,
    n1086,
    n1103,
    n1040,
    n1071
  );


  or
  g1351
  (
    n1389,
    n1081,
    n1079,
    n1034,
    n1106
  );


  and
  g1352
  (
    n1235,
    n1120,
    n1108,
    n1112,
    n1060
  );


  and
  g1353
  (
    n1369,
    n1048,
    n1088,
    n1078,
    n1057
  );


  xor
  g1354
  (
    n1346,
    n1121,
    n1092,
    n1093,
    n1087
  );


  xnor
  g1355
  (
    n1361,
    n1099,
    n1082,
    n1084,
    n1085
  );


  xor
  g1356
  (
    n1186,
    n1097,
    n1077,
    n1032,
    n1095
  );


  nand
  g1357
  (
    n1175,
    n1039,
    n1038,
    n348,
    n1085
  );


  or
  g1358
  (
    n1355,
    n1045,
    n1043,
    n1134,
    n1113
  );


  buf
  g1359
  (
    n1619,
    n1188
  );


  buf
  g1360
  (
    n1432,
    n1253
  );


  buf
  g1361
  (
    n1451,
    n355
  );


  not
  g1362
  (
    n1509,
    n1165
  );


  buf
  g1363
  (
    n1581,
    n1190
  );


  buf
  g1364
  (
    n1430,
    n1247
  );


  not
  g1365
  (
    n1563,
    n1171
  );


  not
  g1366
  (
    n1543,
    n1169
  );


  not
  g1367
  (
    n1478,
    n1259
  );


  not
  g1368
  (
    n1403,
    n1196
  );


  buf
  g1369
  (
    n1453,
    n1147
  );


  not
  g1370
  (
    n1602,
    n1226
  );


  not
  g1371
  (
    n1491,
    n1178
  );


  not
  g1372
  (
    n1573,
    n1212
  );


  not
  g1373
  (
    n1426,
    n1252
  );


  not
  g1374
  (
    KeyWire_0_14,
    n1247
  );


  not
  g1375
  (
    n1544,
    n1249
  );


  not
  g1376
  (
    n1497,
    n1235
  );


  not
  g1377
  (
    n1500,
    n1245
  );


  buf
  g1378
  (
    n1548,
    n357
  );


  buf
  g1379
  (
    n1537,
    n1198
  );


  not
  g1380
  (
    n1607,
    n1243
  );


  buf
  g1381
  (
    n1501,
    n360
  );


  not
  g1382
  (
    n1610,
    n1220
  );


  buf
  g1383
  (
    n1618,
    n1189
  );


  buf
  g1384
  (
    n1542,
    n1200
  );


  buf
  g1385
  (
    n1489,
    n1240
  );


  buf
  g1386
  (
    n1617,
    n1238
  );


  not
  g1387
  (
    n1605,
    n1237
  );


  not
  g1388
  (
    n1530,
    n1237
  );


  not
  g1389
  (
    n1458,
    n1234
  );


  not
  g1390
  (
    n1446,
    n1140
  );


  not
  g1391
  (
    n1541,
    n1211
  );


  buf
  g1392
  (
    n1608,
    n1244
  );


  not
  g1393
  (
    n1567,
    n1181
  );


  buf
  g1394
  (
    n1601,
    n1261
  );


  buf
  g1395
  (
    n1551,
    n1193
  );


  buf
  g1396
  (
    n1565,
    n1240
  );


  not
  g1397
  (
    n1571,
    n1233
  );


  not
  g1398
  (
    n1622,
    n1159
  );


  buf
  g1399
  (
    n1477,
    n1164
  );


  not
  g1400
  (
    n1480,
    n1202
  );


  buf
  g1401
  (
    n1427,
    n1163
  );


  buf
  g1402
  (
    n1433,
    n1258
  );


  buf
  g1403
  (
    n1612,
    n354
  );


  not
  g1404
  (
    KeyWire_0_4,
    n1245
  );


  buf
  g1405
  (
    n1419,
    n1208
  );


  buf
  g1406
  (
    n1452,
    n1245
  );


  not
  g1407
  (
    n1596,
    n1225
  );


  buf
  g1408
  (
    n1492,
    n1248
  );


  not
  g1409
  (
    n1519,
    n1254
  );


  buf
  g1410
  (
    n1598,
    n1260
  );


  buf
  g1411
  (
    n1396,
    n1242
  );


  buf
  g1412
  (
    n1431,
    n1251
  );


  buf
  g1413
  (
    n1514,
    n1258
  );


  not
  g1414
  (
    n1400,
    n1237
  );


  not
  g1415
  (
    n1597,
    n1236
  );


  not
  g1416
  (
    n1465,
    n1243
  );


  buf
  g1417
  (
    KeyWire_0_8,
    n1256
  );


  not
  g1418
  (
    n1599,
    n1161
  );


  buf
  g1419
  (
    n1429,
    n1235
  );


  not
  g1420
  (
    n1402,
    n1139
  );


  buf
  g1421
  (
    n1423,
    n1233
  );


  buf
  g1422
  (
    n1553,
    n1246
  );


  buf
  g1423
  (
    n1437,
    n1243
  );


  buf
  g1424
  (
    n1606,
    n1260
  );


  not
  g1425
  (
    n1549,
    n1234
  );


  buf
  g1426
  (
    n1439,
    n1173
  );


  not
  g1427
  (
    n1523,
    n351
  );


  buf
  g1428
  (
    n1576,
    n1207
  );


  not
  g1429
  (
    n1592,
    n1166
  );


  not
  g1430
  (
    n1524,
    n1194
  );


  not
  g1431
  (
    n1444,
    n1255
  );


  buf
  g1432
  (
    n1448,
    n1249
  );


  buf
  g1433
  (
    n1466,
    n1247
  );


  not
  g1434
  (
    n1482,
    n1239
  );


  buf
  g1435
  (
    n1474,
    n1255
  );


  not
  g1436
  (
    n1572,
    n1265
  );


  not
  g1437
  (
    n1533,
    n361
  );


  buf
  g1438
  (
    n1407,
    n1251
  );


  not
  g1439
  (
    n1447,
    n1197
  );


  not
  g1440
  (
    n1529,
    n1255
  );


  not
  g1441
  (
    n1593,
    n358
  );


  not
  g1442
  (
    n1463,
    n1246
  );


  buf
  g1443
  (
    n1539,
    n1154
  );


  not
  g1444
  (
    n1595,
    n363
  );


  not
  g1445
  (
    n1578,
    n1231
  );


  buf
  g1446
  (
    n1411,
    n1260
  );


  buf
  g1447
  (
    n1410,
    n1249
  );


  not
  g1448
  (
    n1546,
    n1256
  );


  buf
  g1449
  (
    n1487,
    n1215
  );


  not
  g1450
  (
    n1393,
    n1146
  );


  not
  g1451
  (
    n1461,
    n1251
  );


  buf
  g1452
  (
    n1414,
    n1182
  );


  buf
  g1453
  (
    n1434,
    n1264
  );


  not
  g1454
  (
    n1417,
    n1137
  );


  buf
  g1455
  (
    n1496,
    n1218
  );


  buf
  g1456
  (
    n1580,
    n1261
  );


  not
  g1457
  (
    n1609,
    n1176
  );


  not
  g1458
  (
    n1424,
    n1254
  );


  not
  g1459
  (
    n1504,
    n1250
  );


  not
  g1460
  (
    n1600,
    n1236
  );


  not
  g1461
  (
    n1604,
    n1209
  );


  buf
  g1462
  (
    n1512,
    n1232
  );


  buf
  g1463
  (
    n1525,
    n1241
  );


  buf
  g1464
  (
    n1591,
    n1232
  );


  buf
  g1465
  (
    n1413,
    n356
  );


  not
  g1466
  (
    n1594,
    n1236
  );


  buf
  g1467
  (
    n1513,
    n1155
  );


  not
  g1468
  (
    n1457,
    n1203
  );


  buf
  g1469
  (
    n1449,
    n1239
  );


  buf
  g1470
  (
    n1527,
    n1247
  );


  buf
  g1471
  (
    n1558,
    n1236
  );


  not
  g1472
  (
    n1586,
    n1252
  );


  not
  g1473
  (
    n1412,
    n1235
  );


  buf
  g1474
  (
    n1590,
    n1253
  );


  not
  g1475
  (
    n1468,
    n1205
  );


  buf
  g1476
  (
    n1577,
    n1259
  );


  not
  g1477
  (
    n1568,
    n1240
  );


  not
  g1478
  (
    n1493,
    n1244
  );


  not
  g1479
  (
    n1462,
    n1149
  );


  buf
  g1480
  (
    n1584,
    n1258
  );


  buf
  g1481
  (
    n1416,
    n1249
  );


  not
  g1482
  (
    n1475,
    n1162
  );


  buf
  g1483
  (
    n1589,
    n1227
  );


  buf
  g1484
  (
    n1560,
    n1253
  );


  not
  g1485
  (
    n1455,
    n1246
  );


  not
  g1486
  (
    n1615,
    n1263
  );


  buf
  g1487
  (
    n1483,
    n1250
  );


  not
  g1488
  (
    n1522,
    n1248
  );


  buf
  g1489
  (
    n1405,
    n1261
  );


  not
  g1490
  (
    n1579,
    n1233
  );


  not
  g1491
  (
    n1516,
    n1256
  );


  not
  g1492
  (
    n1435,
    n1242
  );


  buf
  g1493
  (
    n1505,
    n1145
  );


  buf
  g1494
  (
    n1570,
    n1251
  );


  buf
  g1495
  (
    n1566,
    n1229
  );


  buf
  g1496
  (
    n1479,
    n1232
  );


  buf
  g1497
  (
    n1404,
    n1259
  );


  buf
  g1498
  (
    n1518,
    n1252
  );


  not
  g1499
  (
    n1561,
    n1257
  );


  buf
  g1500
  (
    n1456,
    n1167
  );


  buf
  g1501
  (
    n1394,
    n1241
  );


  not
  g1502
  (
    n1555,
    n1234
  );


  not
  g1503
  (
    n1472,
    n1213
  );


  not
  g1504
  (
    n1526,
    n1183
  );


  not
  g1505
  (
    n1420,
    n1144
  );


  buf
  g1506
  (
    n1502,
    n1258
  );


  not
  g1507
  (
    n1445,
    n1238
  );


  not
  g1508
  (
    n1507,
    n1235
  );


  not
  g1509
  (
    n1556,
    n1244
  );


  buf
  g1510
  (
    n1488,
    n1259
  );


  buf
  g1511
  (
    n1397,
    n1240
  );


  buf
  g1512
  (
    n1392,
    n359
  );


  not
  g1513
  (
    n1481,
    n1185
  );


  not
  g1514
  (
    n1422,
    n1168
  );


  not
  g1515
  (
    n1498,
    n1241
  );


  buf
  g1516
  (
    n1587,
    n1257
  );


  not
  g1517
  (
    n1517,
    n1180
  );


  buf
  g1518
  (
    n1464,
    n1237
  );


  buf
  g1519
  (
    n1614,
    n1187
  );


  buf
  g1520
  (
    n1460,
    n1262
  );


  buf
  g1521
  (
    n1409,
    n1222
  );


  not
  g1522
  (
    n1510,
    n1228
  );


  buf
  g1523
  (
    n1442,
    n350
  );


  not
  g1524
  (
    n1620,
    n1256
  );


  buf
  g1525
  (
    n1440,
    n1210
  );


  buf
  g1526
  (
    n1521,
    n1191
  );


  not
  g1527
  (
    n1511,
    n1232
  );


  not
  g1528
  (
    n1470,
    n1246
  );


  buf
  g1529
  (
    n1611,
    n1223
  );


  buf
  g1530
  (
    KeyWire_0_0,
    n1221
  );


  not
  g1531
  (
    n1603,
    n1170
  );


  not
  g1532
  (
    n1515,
    n1219
  );


  buf
  g1533
  (
    n1441,
    n1184
  );


  not
  g1534
  (
    n1421,
    n1172
  );


  buf
  g1535
  (
    n1534,
    n1204
  );


  not
  g1536
  (
    n1613,
    n1239
  );


  buf
  g1537
  (
    n1574,
    n1179
  );


  buf
  g1538
  (
    n1471,
    n1262
  );


  buf
  g1539
  (
    n1499,
    n1242
  );


  buf
  g1540
  (
    n1535,
    n1138
  );


  not
  g1541
  (
    n1469,
    n1206
  );


  buf
  g1542
  (
    n1528,
    n352
  );


  buf
  g1543
  (
    n1508,
    n1216
  );


  buf
  g1544
  (
    n1408,
    n1231
  );


  not
  g1545
  (
    n1520,
    n1245
  );


  buf
  g1546
  (
    n1531,
    n1195
  );


  not
  g1547
  (
    n1506,
    n1142
  );


  not
  g1548
  (
    n1552,
    n1262
  );


  not
  g1549
  (
    n1554,
    n1264
  );


  not
  g1550
  (
    n1490,
    n1152
  );


  not
  g1551
  (
    n1557,
    n1239
  );


  buf
  g1552
  (
    n1486,
    n1158
  );


  not
  g1553
  (
    n1415,
    n1248
  );


  not
  g1554
  (
    n1616,
    n1263
  );


  not
  g1555
  (
    n1473,
    n1157
  );


  not
  g1556
  (
    n1575,
    n1263
  );


  not
  g1557
  (
    n1569,
    n1243
  );


  buf
  g1558
  (
    n1401,
    n362
  );


  not
  g1559
  (
    n1585,
    n1250
  );


  buf
  g1560
  (
    n1588,
    n1252
  );


  not
  g1561
  (
    n1425,
    n1255
  );


  buf
  g1562
  (
    n1485,
    n1192
  );


  buf
  g1563
  (
    n1582,
    n1186
  );


  not
  g1564
  (
    n1495,
    n1233
  );


  not
  g1565
  (
    n1467,
    n1141
  );


  not
  g1566
  (
    n1536,
    n1254
  );


  buf
  g1567
  (
    n1550,
    n353
  );


  not
  g1568
  (
    n1562,
    n1214
  );


  buf
  g1569
  (
    n1459,
    n1262
  );


  not
  g1570
  (
    n1436,
    n1160
  );


  buf
  g1571
  (
    n1494,
    n1199
  );


  not
  g1572
  (
    n1418,
    n1153
  );


  not
  g1573
  (
    n1621,
    n1224
  );


  buf
  g1574
  (
    n1443,
    n1201
  );


  buf
  g1575
  (
    n1540,
    n1244
  );


  not
  g1576
  (
    n1484,
    n1260
  );


  buf
  g1577
  (
    n1547,
    n1217
  );


  not
  g1578
  (
    n1450,
    n1254
  );


  buf
  g1579
  (
    n1406,
    n1174
  );


  not
  g1580
  (
    n1438,
    n1263
  );


  not
  g1581
  (
    n1538,
    n1250
  );


  not
  g1582
  (
    n1559,
    n1242
  );


  not
  g1583
  (
    n1476,
    n1248
  );


  nand
  g1584
  (
    n1532,
    n1175,
    n1150
  );


  nand
  g1585
  (
    n1395,
    n1261,
    n1234
  );


  nand
  g1586
  (
    n1545,
    n1151,
    n1238,
    n1264,
    n1143
  );


  xnor
  g1587
  (
    n1399,
    n1230,
    n1177,
    n1156,
    n1264
  );


  xor
  g1588
  (
    n1583,
    n1257,
    n1257,
    n1241,
    n1231
  );


  nor
  g1589
  (
    n1503,
    n1148,
    n1231,
    n1253,
    n1238
  );


  or
  g1590
  (
    n1693,
    n1526,
    n1268,
    n1338,
    n1481
  );


  and
  g1591
  (
    n1788,
    n1474,
    n1412,
    n1484,
    n1602
  );


  xnor
  g1592
  (
    n1913,
    n1551,
    n1311,
    n1354,
    n1519
  );


  nand
  g1593
  (
    n1896,
    n1291,
    n1470,
    n1341,
    n1563
  );


  and
  g1594
  (
    n1868,
    n1554,
    n1275,
    n1387,
    n1331
  );


  or
  g1595
  (
    n1837,
    n1560,
    n1375,
    n1420,
    n1305
  );


  nor
  g1596
  (
    n1630,
    n1491,
    n1339,
    n1575,
    n1498
  );


  xnor
  g1597
  (
    n1875,
    n1497,
    n1348,
    n1520,
    n1317
  );


  xor
  g1598
  (
    n1838,
    n1385,
    n1314,
    n1366,
    n1562
  );


  nor
  g1599
  (
    n1820,
    n1325,
    n1300,
    n1430,
    n1606
  );


  xor
  g1600
  (
    n1877,
    n1379,
    n1391,
    n1618,
    n1367
  );


  nand
  g1601
  (
    n1794,
    n1602,
    n1602,
    n1500,
    n1485
  );


  xor
  g1602
  (
    n1674,
    n1303,
    n1265,
    n1604,
    n1611
  );


  and
  g1603
  (
    n1886,
    n1612,
    n1325,
    n1584,
    n1546
  );


  xor
  g1604
  (
    n1745,
    n1359,
    n1363,
    n1600,
    n1464
  );


  xnor
  g1605
  (
    n1668,
    n1491,
    n1574,
    n1611,
    n1474
  );


  and
  g1606
  (
    n1735,
    n1275,
    n1276,
    n1545,
    n1293
  );


  xnor
  g1607
  (
    n1811,
    n1337,
    n1287,
    n1504,
    n1272
  );


  nand
  g1608
  (
    n1878,
    n1268,
    n1267,
    n1553,
    n1481
  );


  nor
  g1609
  (
    n1832,
    n1329,
    n1313,
    n1521,
    n1361
  );


  and
  g1610
  (
    n1881,
    n1507,
    n1517,
    n1322,
    n1548
  );


  nand
  g1611
  (
    n1836,
    n1524,
    n1389,
    n1394,
    n1364
  );


  nand
  g1612
  (
    n1712,
    n1533,
    n1539,
    n1605,
    n1603
  );


  xor
  g1613
  (
    n1769,
    n1396,
    n1568,
    n1341,
    n1300
  );


  or
  g1614
  (
    n1902,
    n1577,
    n1370,
    n1539,
    n1468
  );


  xnor
  g1615
  (
    n1815,
    n1522,
    n1493,
    n1289,
    n1363
  );


  and
  g1616
  (
    n1892,
    n1360,
    n1448,
    n1593,
    n1318
  );


  and
  g1617
  (
    n1824,
    n1517,
    n1374,
    n1537,
    n1318
  );


  xor
  g1618
  (
    n1831,
    n1364,
    n1306,
    n1496,
    n1367
  );


  nor
  g1619
  (
    n1817,
    n1533,
    n1315,
    n1542,
    n1444
  );


  and
  g1620
  (
    n1812,
    n1280,
    n1340,
    n1349,
    n1507
  );


  xnor
  g1621
  (
    n1797,
    n1513,
    n1548,
    n1589,
    n1294
  );


  xor
  g1622
  (
    n1864,
    n1277,
    n1345,
    n1336,
    n1293
  );


  and
  g1623
  (
    n1854,
    n1332,
    n1525,
    n1500,
    n1350
  );


  nor
  g1624
  (
    n1917,
    n1284,
    n1549,
    n1422,
    n1476
  );


  xor
  g1625
  (
    n1867,
    n1433,
    n1537,
    n1293,
    n1490
  );


  or
  g1626
  (
    n1677,
    n1353,
    n1333,
    n1573,
    n1460
  );


  nor
  g1627
  (
    n1907,
    n1384,
    n1588,
    n1480,
    n1544
  );


  nor
  g1628
  (
    n1773,
    n1303,
    n1487,
    n1373,
    n1520
  );


  and
  g1629
  (
    n1887,
    n1531,
    n1542,
    n1370,
    n1316
  );


  or
  g1630
  (
    n1623,
    n1596,
    n1595,
    n1533,
    n1495
  );


  xnor
  g1631
  (
    n1792,
    n1494,
    n1328,
    n1414,
    n1386
  );


  and
  g1632
  (
    n1781,
    n1306,
    n1510,
    n1330,
    n1604
  );


  nor
  g1633
  (
    n1921,
    n1300,
    n1597,
    n1330,
    n1511
  );


  nand
  g1634
  (
    n1888,
    n1478,
    n1337,
    n1329,
    n1302
  );


  nor
  g1635
  (
    n1874,
    n1486,
    n1532,
    n1527,
    n1310
  );


  nor
  g1636
  (
    n1903,
    n1364,
    n1291,
    n1616,
    n1524
  );


  nor
  g1637
  (
    n1732,
    n1512,
    n1368,
    n1379,
    n369
  );


  or
  g1638
  (
    n1829,
    n1369,
    n1376,
    n1419,
    n1478
  );


  nor
  g1639
  (
    n1810,
    n1521,
    n1571,
    n1316,
    n1382
  );


  or
  g1640
  (
    n1636,
    n1360,
    n1607,
    n1592,
    n1534
  );


  or
  g1641
  (
    n1755,
    n1509,
    n1598,
    n1559,
    n1451
  );


  xor
  g1642
  (
    n1871,
    n1369,
    n1499,
    n1310,
    n1356
  );


  nand
  g1643
  (
    n1624,
    n1609,
    n1476,
    n1359,
    n1502
  );


  or
  g1644
  (
    n1870,
    n1520,
    n1597,
    n1584,
    n1619
  );


  xor
  g1645
  (
    n1653,
    n1385,
    n1567,
    n1508,
    n1564
  );


  nand
  g1646
  (
    n1840,
    n1273,
    n1355,
    n1323,
    n367
  );


  xnor
  g1647
  (
    n1747,
    n1556,
    n1456,
    n1382,
    n1322
  );


  or
  g1648
  (
    n1716,
    n1567,
    n1325,
    n1519,
    n1551
  );


  and
  g1649
  (
    n1642,
    n1499,
    n1429,
    n1288,
    n1572
  );


  nor
  g1650
  (
    n1908,
    n1489,
    n1437,
    n1323,
    n1458
  );


  and
  g1651
  (
    n1651,
    n1610,
    n1265,
    n1552,
    n1378
  );


  nor
  g1652
  (
    n1628,
    n1290,
    n1613,
    n1474,
    n1536
  );


  and
  g1653
  (
    n1650,
    n1513,
    n1285,
    n1478,
    n1598
  );


  xor
  g1654
  (
    n1713,
    n1292,
    n1503,
    n1365,
    n1528
  );


  xnor
  g1655
  (
    n1640,
    n1276,
    n1371,
    n1515,
    n1593
  );


  and
  g1656
  (
    n1690,
    n1570,
    n1388,
    n1615,
    n1299
  );


  xnor
  g1657
  (
    n1647,
    n1526,
    n1525,
    n1566,
    n1295
  );


  nor
  g1658
  (
    n1779,
    n1324,
    n1296,
    n1438,
    n1523
  );


  or
  g1659
  (
    n1809,
    n1343,
    n1471,
    n1435,
    n1485
  );


  nor
  g1660
  (
    n1826,
    n1352,
    n1320,
    n1335,
    n1541
  );


  and
  g1661
  (
    n1872,
    n1557,
    n1389,
    n1380,
    n1361
  );


  or
  g1662
  (
    n1783,
    n1356,
    n1543,
    n1424,
    n1308
  );


  nand
  g1663
  (
    n1789,
    n1542,
    n1380,
    n1536,
    n1587
  );


  nand
  g1664
  (
    n1782,
    n1280,
    n1298,
    n1616,
    n1408
  );


  nand
  g1665
  (
    n1834,
    n1488,
    n1517,
    n1545,
    n1341
  );


  nand
  g1666
  (
    n1849,
    n1565,
    n1338,
    n1374,
    n1426
  );


  nand
  g1667
  (
    n1744,
    n1584,
    n1501,
    n1619,
    n1340
  );


  nand
  g1668
  (
    n1825,
    n1336,
    n1599,
    n1295,
    n1535
  );


  or
  g1669
  (
    n1727,
    n1365,
    n1364,
    n1535,
    n1519
  );


  nand
  g1670
  (
    n1785,
    n1362,
    n1489,
    n1571,
    n1514
  );


  xor
  g1671
  (
    n1759,
    n1585,
    n1347,
    n1540,
    n1552
  );


  or
  g1672
  (
    n1778,
    n1610,
    n1561,
    n1578,
    n1551
  );


  nand
  g1673
  (
    n1710,
    n1447,
    n1281,
    n1277,
    n1316
  );


  or
  g1674
  (
    n1859,
    n1359,
    n371,
    n1479,
    n1543
  );


  and
  g1675
  (
    n1906,
    n1488,
    n1549,
    n1266,
    n1368
  );


  xor
  g1676
  (
    n1711,
    n1615,
    n1327,
    n1538,
    n1553
  );


  or
  g1677
  (
    n1659,
    n1506,
    n1393,
    n1572,
    n1286
  );


  xnor
  g1678
  (
    n1865,
    n1303,
    n1485,
    n1612
  );


  xor
  g1679
  (
    n1791,
    n1352,
    n1511,
    n1578,
    n1282
  );


  xnor
  g1680
  (
    n1863,
    n1372,
    n1617,
    n1309,
    n1330
  );


  and
  g1681
  (
    n1723,
    n1490,
    n1530,
    n1298,
    n1406
  );


  or
  g1682
  (
    n1814,
    n1559,
    n1622,
    n1476,
    n1333
  );


  or
  g1683
  (
    n1691,
    n1600,
    n1617,
    n1523,
    n1335
  );


  xnor
  g1684
  (
    n1858,
    n1579,
    n1449,
    n1363,
    n1309
  );


  xor
  g1685
  (
    n1746,
    n1302,
    n1554,
    n1606,
    n1348
  );


  or
  g1686
  (
    n1784,
    n1583,
    n1269,
    n1266,
    n1280
  );


  and
  g1687
  (
    n1680,
    n1301,
    n1288,
    n1498,
    n1289
  );


  nand
  g1688
  (
    n1638,
    n1373,
    n1494,
    n1577,
    n1550
  );


  nor
  g1689
  (
    n1920,
    n1605,
    n1497,
    n1366,
    n1294
  );


  and
  g1690
  (
    n1635,
    n1547,
    n1316,
    n1540,
    n1322
  );


  nor
  g1691
  (
    n1830,
    n1381,
    n1320,
    n1527,
    n1290
  );


  nand
  g1692
  (
    n1757,
    n1599,
    n1280,
    n1314,
    n1335
  );


  xnor
  g1693
  (
    n1856,
    n1598,
    n1294,
    n1480,
    n1482
  );


  xor
  g1694
  (
    n1804,
    n1440,
    n1389,
    n1397,
    n1381
  );


  or
  g1695
  (
    n1800,
    n1488,
    n1290,
    n1487,
    n1585
  );


  and
  g1696
  (
    n1704,
    n1492,
    n1524,
    n1274,
    n1387
  );


  nor
  g1697
  (
    n1740,
    n1285,
    n1328,
    n1564,
    n1486
  );


  and
  g1698
  (
    n1669,
    n1382,
    n1502,
    n1555,
    n1588
  );


  or
  g1699
  (
    n1823,
    n1583,
    n1510,
    n1473,
    n1508
  );


  nand
  g1700
  (
    n1717,
    n1273,
    n1605,
    n1452,
    n1613
  );


  or
  g1701
  (
    n1673,
    n1513,
    n1446,
    n1481,
    n1610
  );


  nor
  g1702
  (
    n1822,
    n1362,
    n1529,
    n1391,
    n1497
  );


  or
  g1703
  (
    n1894,
    n1577,
    n1274,
    n1475,
    n1354
  );


  xnor
  g1704
  (
    n1689,
    n1270,
    n1339,
    n1287,
    n1332
  );


  nand
  g1705
  (
    n1861,
    n1308,
    n1486,
    n1279,
    n1411
  );


  nand
  g1706
  (
    n1764,
    n1590,
    n1369,
    n1317,
    n1307
  );


  nand
  g1707
  (
    n1686,
    n1483,
    n1352,
    n1292,
    n1326
  );


  or
  g1708
  (
    n1909,
    n1512,
    n1342,
    n1320,
    n1356
  );


  and
  g1709
  (
    n1775,
    n1383,
    n1529,
    n1489,
    n1455
  );


  or
  g1710
  (
    n1733,
    n1479,
    n1297,
    n1354,
    n1385
  );


  xnor
  g1711
  (
    n1687,
    n1551,
    n1591,
    n1621,
    n1345
  );


  and
  g1712
  (
    n1632,
    n1281,
    n1326,
    n1603,
    n1334
  );


  xor
  g1713
  (
    n1667,
    n1311,
    n1283,
    n1450,
    n1563
  );


  and
  g1714
  (
    n1649,
    n1496,
    n1331,
    n1519,
    n1423
  );


  xor
  g1715
  (
    n1911,
    n1528,
    n1611,
    n1431,
    n1548
  );


  nand
  g1716
  (
    n1664,
    n1384,
    n1384,
    n1383,
    n1522
  );


  xnor
  g1717
  (
    n1898,
    n1344,
    n372,
    n1579,
    n1549
  );


  nor
  g1718
  (
    n1679,
    n1283,
    n1307,
    n1555
  );


  or
  g1719
  (
    n1682,
    n1388,
    n1327,
    n1361,
    n1272
  );


  nor
  g1720
  (
    n1641,
    n1602,
    n1284,
    n1606,
    n1434
  );


  xnor
  g1721
  (
    n1726,
    n1413,
    n1580,
    n1587,
    n1582
  );


  or
  g1722
  (
    n1637,
    n1588,
    n1578,
    n1586,
    n1620
  );


  xnor
  g1723
  (
    n1683,
    n1608,
    n1531,
    n1491,
    n1365
  );


  or
  g1724
  (
    n1827,
    n1338,
    n1360,
    n1307,
    n1301
  );


  or
  g1725
  (
    n1758,
    n1404,
    n1463,
    n1540,
    n1277
  );


  or
  g1726
  (
    n1633,
    n1321,
    n1613,
    n1340,
    n1620
  );


  xor
  g1727
  (
    n1890,
    n1622,
    n1328,
    n1594,
    n1612
  );


  nor
  g1728
  (
    n1786,
    n1507,
    n1331,
    n1547,
    n1606
  );


  and
  g1729
  (
    n1706,
    n1569,
    n1590,
    n1576,
    n1328
  );


  nand
  g1730
  (
    n1699,
    n1350,
    n1284,
    n1358,
    n1576
  );


  and
  g1731
  (
    n1644,
    n1592,
    n1570,
    n1421,
    n1571
  );


  xnor
  g1732
  (
    n1833,
    n1516,
    n1586,
    n1510,
    n1351
  );


  nand
  g1733
  (
    n1737,
    n364,
    n1526,
    n1269,
    n1579
  );


  nand
  g1734
  (
    n1627,
    n1617,
    n1531,
    n1554,
    n1568
  );


  and
  g1735
  (
    n1793,
    n1326,
    n1275,
    n1613,
    n1566
  );


  nand
  g1736
  (
    n1852,
    n1289,
    n370,
    n1319,
    n1473
  );


  xnor
  g1737
  (
    n1860,
    n1580,
    n1387,
    n1554,
    n1608
  );


  nor
  g1738
  (
    n1884,
    n1267,
    n1599,
    n1488,
    n1335
  );


  and
  g1739
  (
    n1893,
    n1357,
    n1371,
    n1288,
    n1370
  );


  nand
  g1740
  (
    n1660,
    n1418,
    n1494,
    n1392,
    n1506
  );


  and
  g1741
  (
    KeyWire_0_28,
    n1523,
    n1492,
    n1585,
    n1603
  );


  and
  g1742
  (
    n1626,
    n1571,
    n1525,
    n1275,
    n1614
  );


  and
  g1743
  (
    n1912,
    n1363,
    n1337,
    n1386,
    n1368
  );


  and
  g1744
  (
    n1767,
    n1534,
    n1477,
    n1398,
    n1299
  );


  xnor
  g1745
  (
    n1648,
    n1534,
    n1278,
    n1304,
    n1544
  );


  xor
  g1746
  (
    n1678,
    n1482,
    n1536,
    n1319,
    n1461
  );


  nor
  g1747
  (
    n1806,
    n1555,
    n1565,
    n1405,
    n1545
  );


  or
  g1748
  (
    n1770,
    n1337,
    n1614,
    n1284,
    n1292
  );


  xor
  g1749
  (
    n1821,
    n1268,
    n1544,
    n1546,
    n1569
  );


  xor
  g1750
  (
    n1857,
    n1282,
    n1593,
    n1563,
    n1339
  );


  nand
  g1751
  (
    n1801,
    n1575,
    n1298,
    n373,
    n1526
  );


  or
  g1752
  (
    n1748,
    n1378,
    n1480,
    n1271,
    n1321
  );


  or
  g1753
  (
    n1695,
    n1385,
    n1507,
    n1291,
    n1546
  );


  nand
  g1754
  (
    n1658,
    n1417,
    n1380,
    n1332,
    n1605
  );


  xnor
  g1755
  (
    n1899,
    n1561,
    n1567,
    n1536,
    n1436
  );


  xor
  g1756
  (
    n1772,
    n1503,
    n1357,
    n1298,
    n1479
  );


  nor
  g1757
  (
    n1803,
    n1480,
    n1391,
    n1472,
    n1518
  );


  nand
  g1758
  (
    n1625,
    n1287,
    n1306,
    n1273,
    n1379
  );


  nor
  g1759
  (
    n1692,
    n1296,
    n1537,
    n1395,
    n1308
  );


  xnor
  g1760
  (
    n1910,
    n1557,
    n1555,
    n1384,
    n1614
  );


  nand
  g1761
  (
    n1805,
    n1410,
    n1515,
    n1309,
    n1378
  );


  xnor
  g1762
  (
    n1853,
    n1343,
    n1365,
    n1353,
    n1574
  );


  or
  g1763
  (
    n1718,
    n1318,
    n1348,
    n1390,
    n1388
  );


  or
  g1764
  (
    n1841,
    n1487,
    n1370,
    n1553,
    n1591
  );


  nand
  g1765
  (
    n1734,
    n1301,
    n1469,
    n1346,
    n1505
  );


  xnor
  g1766
  (
    n1904,
    n1283,
    n1399,
    n1509,
    n1336
  );


  or
  g1767
  (
    n1869,
    n1512,
    n1522,
    n1356,
    n1415
  );


  xnor
  g1768
  (
    n1846,
    n1317,
    n1351,
    n1401,
    n1497
  );


  xor
  g1769
  (
    n1905,
    n1596,
    n1327,
    n1390,
    n1382
  );


  and
  g1770
  (
    n1676,
    n1301,
    n1443,
    n1574,
    n1565
  );


  nand
  g1771
  (
    n1796,
    n1501,
    n1490,
    n1362,
    n1582
  );


  or
  g1772
  (
    n1891,
    n1539,
    n1303,
    n1556,
    n1492
  );


  or
  g1773
  (
    n1802,
    n1582,
    n1513,
    n1479,
    n1386
  );


  and
  g1774
  (
    n1787,
    n1359,
    n1285,
    n1336,
    n1333
  );


  or
  g1775
  (
    n1760,
    n1375,
    n1445,
    n1373,
    n1618
  );


  and
  g1776
  (
    n1728,
    n1386,
    n1596,
    n1518,
    n1566
  );


  or
  g1777
  (
    n1666,
    n1407,
    n1278,
    n1274,
    n1383
  );


  and
  g1778
  (
    n1901,
    n1441,
    n1532,
    n1582,
    n1286
  );


  nor
  g1779
  (
    n1742,
    n1279,
    n1521,
    n1381,
    n1427
  );


  xnor
  g1780
  (
    n1662,
    n1538,
    n1387,
    n1311,
    n1617
  );


  nand
  g1781
  (
    n1697,
    n1531,
    n1330,
    n1457,
    n1353
  );


  xor
  g1782
  (
    n1708,
    n1490,
    n1305,
    n1473,
    n1565
  );


  xnor
  g1783
  (
    n1656,
    n1402,
    n1541,
    n1297
  );


  and
  g1784
  (
    n1866,
    n1529,
    n1281,
    n1380,
    n1343
  );


  nor
  g1785
  (
    n1774,
    n1331,
    n1272,
    n1491,
    n1376
  );


  xnor
  g1786
  (
    n1701,
    n1270,
    n1558,
    n1292,
    n1604
  );


  xor
  g1787
  (
    n1882,
    n1508,
    n1268,
    n1496,
    n1266
  );


  xor
  g1788
  (
    n1780,
    n1620,
    n1312,
    n1501,
    n1345
  );


  or
  g1789
  (
    n1762,
    n1552,
    n1534,
    n1358,
    n1500
  );


  and
  g1790
  (
    n1639,
    n1279,
    n1310,
    n1484,
    n1285
  );


  nand
  g1791
  (
    n1725,
    n1622,
    n1287,
    n1289,
    n1590
  );


  xor
  g1792
  (
    n1655,
    n1338,
    n1346,
    n1515,
    n1477
  );


  nor
  g1793
  (
    n1895,
    n1557,
    n1311,
    n1495,
    n1508
  );


  or
  g1794
  (
    n1634,
    n1358,
    n1622,
    n1377,
    n1597
  );


  and
  g1795
  (
    n1761,
    n1562,
    n1509,
    n1494,
    n1271
  );


  and
  g1796
  (
    n1646,
    n1581,
    n1532,
    n1616,
    n1278
  );


  xnor
  g1797
  (
    n1883,
    n1344,
    n1472,
    n1390,
    n1299
  );


  xor
  g1798
  (
    n1724,
    n1425,
    n1620,
    n1383,
    n1556
  );


  and
  g1799
  (
    n1684,
    n1327,
    n1367,
    n1504,
    n1598
  );


  xor
  g1800
  (
    n1808,
    n1375,
    n1389,
    n1594,
    n1496
  );


  xnor
  g1801
  (
    n1671,
    n1544,
    n1282,
    n1558,
    n1353
  );


  nor
  g1802
  (
    KeyWire_0_1,
    n1590,
    n1269,
    n1320,
    n1564
  );


  nor
  g1803
  (
    n1915,
    n1304,
    n1315,
    n1374,
    n1269
  );


  xnor
  g1804
  (
    n1722,
    n1483,
    n1314,
    n1512,
    n1621
  );


  or
  g1805
  (
    n1862,
    n1607,
    n1500,
    n1409,
    n1344
  );


  xnor
  g1806
  (
    n1750,
    n1334,
    n1439,
    n1472,
    n1522
  );


  xor
  g1807
  (
    n1731,
    n1329,
    n1616,
    n1581,
    n1350
  );


  xnor
  g1808
  (
    n1698,
    n1332,
    n1375,
    n1614,
    n1538
  );


  and
  g1809
  (
    n1652,
    n1563,
    n1505,
    n1486,
    n1454
  );


  and
  g1810
  (
    n1700,
    n1604,
    n1505,
    n1482,
    n1349
  );


  and
  g1811
  (
    n1672,
    n1591,
    n1334,
    n1323,
    n1266
  );


  or
  g1812
  (
    n1657,
    n1302,
    n1305,
    n1615,
    n1543
  );


  xnor
  g1813
  (
    n1795,
    n1372,
    n1351,
    n1560,
    n1428
  );


  nand
  g1814
  (
    n1848,
    n1510,
    n1343,
    n1502,
    n1552
  );


  nand
  g1815
  (
    n1729,
    n1495,
    n1575,
    n1530,
    n1376
  );


  nor
  g1816
  (
    n1876,
    n1342,
    n1267,
    n1294,
    n1503
  );


  or
  g1817
  (
    n1816,
    n1579,
    n1352,
    n1586,
    n1346
  );


  xnor
  g1818
  (
    n1665,
    n1379,
    n1473,
    n1334,
    n1592
  );


  and
  g1819
  (
    n1736,
    n1347,
    n1477,
    n1546,
    n1573
  );


  and
  g1820
  (
    n1741,
    n1442,
    n1564,
    n1273,
    n1478
  );


  xnor
  g1821
  (
    n1818,
    n1276,
    n1369,
    n1588,
    n1591
  );


  nand
  g1822
  (
    n1900,
    n1342,
    n1485,
    n1550,
    n1530
  );


  xnor
  g1823
  (
    n1765,
    n1374,
    n1371,
    n1511,
    n1475
  );


  xor
  g1824
  (
    n1855,
    n1378,
    n1315,
    n1313,
    n1271
  );


  or
  g1825
  (
    n1753,
    n1279,
    n1344,
    n1560,
    n1592
  );


  nand
  g1826
  (
    n1790,
    n1283,
    n1539,
    n1483,
    n1535
  );


  xor
  g1827
  (
    n1719,
    n1558,
    n1368,
    n1282,
    n1308
  );


  nand
  g1828
  (
    KeyWire_0_13,
    n1270,
    n1530,
    n1573,
    n1492
  );


  xor
  g1829
  (
    n1661,
    n1274,
    n1608,
    n1366,
    n1495
  );


  xor
  g1830
  (
    n1807,
    n1572,
    n1499,
    n1381,
    n1319
  );


  nor
  g1831
  (
    n1670,
    n1366,
    n1569,
    n1589,
    n1306
  );


  nand
  g1832
  (
    n1702,
    n1573,
    n1516,
    n1351,
    n1545
  );


  nor
  g1833
  (
    n1751,
    n1499,
    n1560,
    n1589,
    n1265
  );


  xnor
  g1834
  (
    n1776,
    n1619,
    n1618,
    n1373,
    n1360
  );


  nor
  g1835
  (
    n1922,
    n1583,
    n1559,
    n1345,
    n1277
  );


  nand
  g1836
  (
    n1715,
    n1487,
    n1553,
    n1538,
    n1290
  );


  and
  g1837
  (
    n1766,
    n1558,
    n1540,
    n1270,
    n1587
  );


  xnor
  g1838
  (
    n1847,
    n1475,
    n1509,
    n1514,
    n1453
  );


  nor
  g1839
  (
    n1916,
    n1583,
    n1482,
    n1295,
    n1416
  );


  and
  g1840
  (
    n1842,
    n1589,
    n1483,
    n1346,
    n1501
  );


  or
  g1841
  (
    n1756,
    n1567,
    n1391,
    n1619,
    n1576
  );


  and
  g1842
  (
    n1631,
    n1465,
    n1504,
    n1610,
    n1286
  );


  nand
  g1843
  (
    n1813,
    n1521,
    n1596,
    n1498,
    n1340
  );


  xnor
  g1844
  (
    n1873,
    n1593,
    n1325,
    n1355,
    n1520
  );


  xnor
  g1845
  (
    n1771,
    n1304,
    n1580,
    n1476,
    n1302
  );


  xor
  g1846
  (
    n1763,
    n1309,
    n1601,
    n1524,
    n1312
  );


  xnor
  g1847
  (
    n1663,
    n1548,
    n1299,
    n1537,
    n1295
  );


  and
  g1848
  (
    n1675,
    n1527,
    n1600,
    n1475,
    n1533
  );


  or
  g1849
  (
    n1918,
    n1529,
    n1609,
    n1572,
    n1506
  );


  xor
  g1850
  (
    n1749,
    n1341,
    n1547,
    n1317,
    n1300
  );


  xnor
  g1851
  (
    n1654,
    n1611,
    n1324,
    n1608,
    n1581
  );


  nor
  g1852
  (
    n1681,
    n1276,
    n1550,
    n1350,
    n1377
  );


  xor
  g1853
  (
    n1897,
    n1291,
    n1594,
    n1550,
    n1367
  );


  or
  g1854
  (
    n1643,
    n1549,
    n1355,
    n1333,
    n1621
  );


  or
  g1855
  (
    n1879,
    n1388,
    n1618,
    n1577,
    n1484
  );


  or
  g1856
  (
    n1919,
    n1324,
    n1587,
    n1371,
    n1466
  );


  xnor
  g1857
  (
    n1743,
    n1527,
    n1570,
    n1575,
    n1377
  );


  nand
  g1858
  (
    n1880,
    n1481,
    n1321,
    n1514,
    n1296
  );


  nand
  g1859
  (
    n1694,
    n1586,
    n1493,
    n368,
    n1319
  );


  xor
  g1860
  (
    n1696,
    n1601,
    n1516,
    n1597,
    n1324
  );


  nand
  g1861
  (
    n1752,
    n1584,
    n1505,
    n1503,
    n1568
  );


  or
  g1862
  (
    n1889,
    n1357,
    n1502,
    n1474,
    n1272
  );


  nor
  g1863
  (
    n1709,
    n1288,
    n1318,
    n1523,
    n1312
  );


  or
  g1864
  (
    n1828,
    n1312,
    n1516,
    n1390,
    n1498
  );


  and
  g1865
  (
    n1914,
    n1528,
    n1484,
    n1562,
    n1347
  );


  or
  g1866
  (
    n1629,
    n1281,
    n1326,
    n1315,
    n1403
  );


  and
  g1867
  (
    n1850,
    n1517,
    n1329,
    n1467,
    n1615
  );


  or
  g1868
  (
    n1843,
    n1322,
    n1601,
    n1293,
    n1504
  );


  nor
  g1869
  (
    n1799,
    n1532,
    n1566,
    n1543,
    n1377
  );


  and
  g1870
  (
    n1839,
    n1580,
    n1305,
    n1541,
    n1362
  );


  xnor
  g1871
  (
    n1845,
    n1607,
    n1557,
    n1547,
    n1574
  );


  nor
  g1872
  (
    n1705,
    n1518,
    n1585,
    n1493,
    n1515
  );


  and
  g1873
  (
    n1714,
    n1576,
    n1493,
    n1462,
    n1562
  );


  or
  g1874
  (
    n1721,
    n365,
    n1349,
    n1600,
    n1314
  );


  or
  g1875
  (
    n1685,
    n1528,
    n1286,
    n1313,
    n1357
  );


  xor
  g1876
  (
    n1707,
    n1347,
    n1304,
    n1594,
    n1518
  );


  xnor
  g1877
  (
    n1730,
    n1372,
    n1535,
    n1595,
    n1489
  );


  nand
  g1878
  (
    n1645,
    n1339,
    n1432,
    n1541,
    n1578
  );


  xnor
  g1879
  (
    n1835,
    n1376,
    n1570,
    n1607,
    n1569
  );


  or
  g1880
  (
    n1688,
    n1477,
    n1342,
    n1581,
    n366
  );


  or
  g1881
  (
    n1844,
    n1278,
    n1354,
    n1267,
    n1321
  );


  and
  g1882
  (
    n1768,
    n1595,
    n1511,
    n1542,
    n1561
  );


  or
  g1883
  (
    n1777,
    n1323,
    n1361,
    n1556,
    n1621
  );


  nand
  g1884
  (
    n1738,
    n1514,
    n1601,
    n1609,
    n1595
  );


  and
  g1885
  (
    n1720,
    n1561,
    n1459,
    n1525,
    n1297
  );


  nor
  g1886
  (
    n1703,
    n1355,
    n1310,
    n1568,
    n1271
  );


  and
  g1887
  (
    n1851,
    n1603,
    n1599,
    n1559,
    n1372
  );


  xor
  g1888
  (
    n1754,
    n1400,
    n1348,
    n1609,
    n1358
  );


  or
  g1889
  (
    n1739,
    n1296,
    n1349,
    n1313,
    n1506
  );


  nor
  g1890
  (
    n1964,
    n1894,
    n1785,
    n1880,
    n1729
  );


  or
  g1891
  (
    n1952,
    n1764,
    n1651,
    n1781,
    n1702
  );


  and
  g1892
  (
    n1949,
    n1867,
    n1794,
    n1878,
    n1918
  );


  xnor
  g1893
  (
    n1995,
    n377,
    n1828,
    n1630,
    n1837
  );


  or
  g1894
  (
    n1955,
    n1649,
    n1628,
    n1638,
    n1779
  );


  nand
  g1895
  (
    n1948,
    n1920,
    n1788,
    n1732,
    n1802
  );


  xnor
  g1896
  (
    n1934,
    n1667,
    n1865,
    n1790,
    n1727
  );


  nor
  g1897
  (
    n1987,
    n1869,
    n1858,
    n1758,
    n1848
  );


  or
  g1898
  (
    KeyWire_0_18,
    n1754,
    n1910,
    n1634,
    n1637
  );


  xnor
  g1899
  (
    n1939,
    n1705,
    n1711,
    n1908,
    n1666
  );


  nand
  g1900
  (
    n1969,
    n1716,
    n1806,
    n1812,
    n1752
  );


  or
  g1901
  (
    n1966,
    n1825,
    n1680,
    n1726,
    n1783
  );


  xnor
  g1902
  (
    n1980,
    n1690,
    n1818,
    n1652,
    n1743
  );


  nand
  g1903
  (
    n1959,
    n1853,
    n1738,
    n1744,
    n1919
  );


  xnor
  g1904
  (
    n1942,
    n1887,
    n1792,
    n1870,
    n1898
  );


  xnor
  g1905
  (
    n1994,
    n1762,
    n1826,
    n1766,
    n1677
  );


  xor
  g1906
  (
    n1978,
    n375,
    n1760,
    n1856,
    n1733
  );


  nor
  g1907
  (
    n1946,
    n1907,
    n1770,
    n1750,
    n1805
  );


  xor
  g1908
  (
    n1940,
    n1842,
    n1647,
    n1903,
    n1681
  );


  or
  g1909
  (
    n1975,
    n1710,
    n1787,
    n1684,
    n1661
  );


  xor
  g1910
  (
    n1933,
    n1852,
    n1778,
    n1724,
    n1854
  );


  xor
  g1911
  (
    n1953,
    n1849,
    n1776,
    n1696,
    n1698
  );


  xnor
  g1912
  (
    n1972,
    n1753,
    n1694,
    n1780,
    n1832
  );


  nand
  g1913
  (
    n1974,
    n1713,
    n1759,
    n1746,
    n1701
  );


  nor
  g1914
  (
    n1923,
    n1817,
    n1909,
    n1768,
    n1742
  );


  nand
  g1915
  (
    n1929,
    n1905,
    n1821,
    n1723,
    n1749
  );


  or
  g1916
  (
    n1992,
    n1755,
    n1761,
    n1829,
    n1922
  );


  xnor
  g1917
  (
    n1986,
    n1917,
    n1889,
    n1674,
    n1665
  );


  xor
  g1918
  (
    n1963,
    n1739,
    n1731,
    n1714,
    n1659
  );


  nand
  g1919
  (
    n1941,
    n1860,
    n1657,
    n1914,
    n1655
  );


  xnor
  g1920
  (
    n1979,
    n1844,
    n1686,
    n1786,
    n1673
  );


  xnor
  g1921
  (
    n1945,
    n1735,
    n1804,
    n1662,
    n1866
  );


  nand
  g1922
  (
    n1982,
    n1693,
    n1757,
    n1900,
    n1672
  );


  xnor
  g1923
  (
    n1951,
    n1648,
    n1808,
    n1650,
    n1915
  );


  nand
  g1924
  (
    n1927,
    n1669,
    n1774,
    n1748,
    n1633
  );


  xnor
  g1925
  (
    n1962,
    n1751,
    n1820,
    n1916,
    n1895
  );


  or
  g1926
  (
    n1997,
    n1911,
    n1901,
    n1885,
    n1830
  );


  and
  g1927
  (
    n1938,
    n376,
    n1797,
    n1697,
    n1839
  );


  or
  g1928
  (
    n1936,
    n1707,
    n1730,
    n1678,
    n1721
  );


  or
  g1929
  (
    n1932,
    n1827,
    n1789,
    n1857,
    n1741
  );


  or
  g1930
  (
    n1931,
    n1831,
    n1841,
    n1879,
    n1913
  );


  nand
  g1931
  (
    n1958,
    n1893,
    n1799,
    n1663,
    n1784
  );


  xor
  g1932
  (
    n1954,
    n1765,
    n1692,
    n1708,
    n1888
  );


  nand
  g1933
  (
    n1977,
    n1855,
    n1921,
    n1801,
    n1896
  );


  xor
  g1934
  (
    n1950,
    n1631,
    n1899,
    n1712,
    n1834
  );


  and
  g1935
  (
    n1996,
    n1656,
    n1660,
    n1793,
    n1683
  );


  nand
  g1936
  (
    n1971,
    n1875,
    n1704,
    n1771,
    n1717
  );


  xor
  g1937
  (
    n1983,
    n1636,
    n1640,
    n1881,
    n1819
  );


  or
  g1938
  (
    n1988,
    n1736,
    n1809,
    n1777,
    n1864
  );


  nor
  g1939
  (
    n1967,
    n1644,
    n1737,
    n1836,
    n1679
  );


  and
  g1940
  (
    n1981,
    n1691,
    n1671,
    n1775,
    n1675
  );


  xnor
  g1941
  (
    n1956,
    n1873,
    n1845,
    n1811,
    n1646
  );


  and
  g1942
  (
    n1973,
    n1654,
    n1807,
    n1700,
    n1709
  );


  nand
  g1943
  (
    n1985,
    n1629,
    n1840,
    n1670,
    n1877
  );


  and
  g1944
  (
    n1957,
    n1699,
    n1624,
    n1816,
    n1862
  );


  or
  g1945
  (
    n1937,
    n1688,
    n378,
    n1782,
    n1815
  );


  or
  g1946
  (
    n1924,
    n1823,
    n1703,
    n1813,
    n1810
  );


  or
  g1947
  (
    n1944,
    n1706,
    n1838,
    n1668,
    n1747
  );


  or
  g1948
  (
    n1984,
    n1798,
    n1874,
    n1861,
    n1847
  );


  or
  g1949
  (
    n1965,
    n1803,
    n1883,
    n1627,
    n1645
  );


  xor
  g1950
  (
    n1935,
    n1814,
    n1626,
    n1664,
    n1859
  );


  nor
  g1951
  (
    n1925,
    n1685,
    n1851,
    n1871,
    n1734
  );


  xor
  g1952
  (
    n1976,
    n1740,
    n1897,
    n1850,
    n1722
  );


  or
  g1953
  (
    n1993,
    n1822,
    n1687,
    n1868,
    n1641
  );


  xnor
  g1954
  (
    n1991,
    n1720,
    n1689,
    n1695,
    n1763
  );


  nor
  g1955
  (
    n1970,
    n1772,
    n1846,
    n1902,
    n1791
  );


  nor
  g1956
  (
    n1990,
    n1796,
    n1639,
    n1718,
    n1912
  );


  xor
  g1957
  (
    n1998,
    n1643,
    n1835,
    n1725,
    n1635
  );


  or
  g1958
  (
    n1926,
    n1653,
    n1769,
    n1892,
    n1800
  );


  xor
  g1959
  (
    n1960,
    n1745,
    n1863,
    n1773,
    n1767
  );


  xnor
  g1960
  (
    n1968,
    n1682,
    n1886,
    n1891,
    n1795
  );


  or
  g1961
  (
    n1943,
    n1843,
    n1906,
    n1676,
    n1632
  );


  xor
  g1962
  (
    n1930,
    n1824,
    n1876,
    n1715,
    n1884
  );


  or
  g1963
  (
    n1947,
    n1728,
    n1756,
    n1625,
    n1890
  );


  and
  g1964
  (
    n1961,
    n1882,
    n1658,
    n1833,
    n1904
  );


  and
  g1965
  (
    n1989,
    n1642,
    n1719,
    n1872,
    n374
  );


  nor
  g1966
  (
    n2002,
    n1962,
    n1995,
    n1989,
    n1946
  );


  nand
  g1967
  (
    n2004,
    n1956,
    n1935,
    n1950,
    n1963
  );


  or
  g1968
  (
    n2015,
    n1966,
    n1985,
    n1933,
    n1955
  );


  nor
  g1969
  (
    n2017,
    n1993,
    n1972,
    n1960,
    n1930
  );


  xor
  g1970
  (
    n2000,
    n1937,
    n1976,
    n1988,
    n1926
  );


  xnor
  g1971
  (
    n2013,
    n1969,
    n1984,
    n1941,
    n1982
  );


  nand
  g1972
  (
    KeyWire_0_26,
    n1991,
    n1942,
    n1997,
    n1990
  );


  xor
  g1973
  (
    n2006,
    n1944,
    n1928,
    n1964,
    n1952
  );


  nor
  g1974
  (
    n2003,
    n1974,
    n1939,
    n1938,
    n1965
  );


  and
  g1975
  (
    n2010,
    n1975,
    n1970,
    n1980,
    n1929
  );


  nand
  g1976
  (
    n2001,
    n1957,
    n1967,
    n1953,
    n1925
  );


  or
  g1977
  (
    n2011,
    n1961,
    n1940,
    n1959,
    n1992
  );


  nor
  g1978
  (
    n2014,
    n1994,
    n1948,
    n1943,
    n1978
  );


  xor
  g1979
  (
    n2007,
    n1934,
    n1949,
    n1983,
    n1958
  );


  nand
  g1980
  (
    n2016,
    n1947,
    n1927,
    n1932,
    n1986
  );


  and
  g1981
  (
    n2008,
    n1979,
    n1998,
    n1945,
    n1954
  );


  or
  g1982
  (
    n1999,
    n1996,
    n1951,
    n1923,
    n1924
  );


  xnor
  g1983
  (
    n2009,
    n1971,
    n1968,
    n1931,
    n1977
  );


  xor
  g1984
  (
    n2012,
    n1981,
    n1973,
    n1987,
    n1936
  );


  or
  g1985
  (
    n2025,
    n2003,
    n398,
    n383,
    n2005
  );


  and
  g1986
  (
    n2018,
    n2008,
    n2016,
    n385,
    n388
  );


  xnor
  g1987
  (
    n2027,
    n399,
    n395,
    n380,
    n2009
  );


  or
  g1988
  (
    n2028,
    n386,
    n396,
    n387,
    n2007
  );


  nor
  g1989
  (
    n2029,
    n2002,
    n2015,
    n408,
    n389
  );


  xnor
  g1990
  (
    n2023,
    n404,
    n401,
    n2000,
    n391
  );


  or
  g1991
  (
    n2030,
    n381,
    n2006,
    n2014,
    n1999
  );


  nor
  g1992
  (
    n2019,
    n418,
    n405,
    n397,
    n407
  );


  or
  g1993
  (
    n2031,
    n382,
    n379,
    n2013,
    n394
  );


  nand
  g1994
  (
    n2032,
    n406,
    n393,
    n415,
    n410
  );


  and
  g1995
  (
    n2022,
    n412,
    n400,
    n2011,
    n413
  );


  or
  g1996
  (
    n2021,
    n416,
    n384,
    n2004,
    n2001
  );


  nand
  g1997
  (
    n2026,
    n390,
    n402,
    n2010,
    n392
  );


  nor
  g1998
  (
    n2020,
    n419,
    n2017,
    n409,
    n2012
  );


  and
  g1999
  (
    n2024,
    n414,
    n417,
    n411,
    n403
  );


  xnor
  KeyGate_0_0
  (
    n1428,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1798,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n635,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n72,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1454,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1167,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n774,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n465,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1398,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n623,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n146,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1061,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n920,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1885,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1564,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n525,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n436,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n662,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n1928,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1040,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n384,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n326,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1386,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n288,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1056,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1194,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n2005,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n908,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1819,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1142,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n311,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n144,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


