

module Stat_4000_402
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n3750,
  n3884,
  n3879,
  n3922,
  n3921,
  n3912,
  n3913,
  n3926,
  n3918,
  n3919,
  n3917,
  n3920,
  n3914,
  n3924,
  n3982,
  n3981,
  n3992,
  n3996,
  n3985,
  n3987,
  n3991,
  n3984,
  n3990,
  n3988,
  n3995,
  n3989,
  n3993,
  n3986,
  n3994,
  n4031,
  n4030,
  n4032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n3750;output n3884;output n3879;output n3922;output n3921;output n3912;output n3913;output n3926;output n3918;output n3919;output n3917;output n3920;output n3914;output n3924;output n3982;output n3981;output n3992;output n3996;output n3985;output n3987;output n3991;output n3984;output n3990;output n3988;output n3995;output n3989;output n3993;output n3986;output n3994;output n4031;output n4030;output n4032;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire n3011;wire n3012;wire n3013;wire n3014;wire n3015;wire n3016;wire n3017;wire n3018;wire n3019;wire n3020;wire n3021;wire n3022;wire n3023;wire n3024;wire n3025;wire n3026;wire n3027;wire n3028;wire n3029;wire n3030;wire n3031;wire n3032;wire n3033;wire n3034;wire n3035;wire n3036;wire n3037;wire n3038;wire n3039;wire n3040;wire n3041;wire n3042;wire n3043;wire n3044;wire n3045;wire n3046;wire n3047;wire n3048;wire n3049;wire n3050;wire n3051;wire n3052;wire n3053;wire n3054;wire n3055;wire n3056;wire n3057;wire n3058;wire n3059;wire n3060;wire n3061;wire n3062;wire n3063;wire n3064;wire n3065;wire n3066;wire n3067;wire n3068;wire n3069;wire n3070;wire n3071;wire n3072;wire n3073;wire n3074;wire n3075;wire n3076;wire n3077;wire n3078;wire n3079;wire n3080;wire n3081;wire n3082;wire n3083;wire n3084;wire n3085;wire n3086;wire n3087;wire n3088;wire n3089;wire n3090;wire n3091;wire n3092;wire n3093;wire n3094;wire n3095;wire n3096;wire n3097;wire n3098;wire n3099;wire n3100;wire n3101;wire n3102;wire n3103;wire n3104;wire n3105;wire n3106;wire n3107;wire n3108;wire n3109;wire n3110;wire n3111;wire n3112;wire n3113;wire n3114;wire n3115;wire n3116;wire n3117;wire n3118;wire n3119;wire n3120;wire n3121;wire n3122;wire n3123;wire n3124;wire n3125;wire n3126;wire n3127;wire n3128;wire n3129;wire n3130;wire n3131;wire n3132;wire n3133;wire n3134;wire n3135;wire n3136;wire n3137;wire n3138;wire n3139;wire n3140;wire n3141;wire n3142;wire n3143;wire n3144;wire n3145;wire n3146;wire n3147;wire n3148;wire n3149;wire n3150;wire n3151;wire n3152;wire n3153;wire n3154;wire n3155;wire n3156;wire n3157;wire n3158;wire n3159;wire n3160;wire n3161;wire n3162;wire n3163;wire n3164;wire n3165;wire n3166;wire n3167;wire n3168;wire n3169;wire n3170;wire n3171;wire n3172;wire n3173;wire n3174;wire n3175;wire n3176;wire n3177;wire n3178;wire n3179;wire n3180;wire n3181;wire n3182;wire n3183;wire n3184;wire n3185;wire n3186;wire n3187;wire n3188;wire n3189;wire n3190;wire n3191;wire n3192;wire n3193;wire n3194;wire n3195;wire n3196;wire n3197;wire n3198;wire n3199;wire n3200;wire n3201;wire n3202;wire n3203;wire n3204;wire n3205;wire n3206;wire n3207;wire n3208;wire n3209;wire n3210;wire n3211;wire n3212;wire n3213;wire n3214;wire n3215;wire n3216;wire n3217;wire n3218;wire n3219;wire n3220;wire n3221;wire n3222;wire n3223;wire n3224;wire n3225;wire n3226;wire n3227;wire n3228;wire n3229;wire n3230;wire n3231;wire n3232;wire n3233;wire n3234;wire n3235;wire n3236;wire n3237;wire n3238;wire n3239;wire n3240;wire n3241;wire n3242;wire n3243;wire n3244;wire n3245;wire n3246;wire n3247;wire n3248;wire n3249;wire n3250;wire n3251;wire n3252;wire n3253;wire n3254;wire n3255;wire n3256;wire n3257;wire n3258;wire n3259;wire n3260;wire n3261;wire n3262;wire n3263;wire n3264;wire n3265;wire n3266;wire n3267;wire n3268;wire n3269;wire n3270;wire n3271;wire n3272;wire n3273;wire n3274;wire n3275;wire n3276;wire n3277;wire n3278;wire n3279;wire n3280;wire n3281;wire n3282;wire n3283;wire n3284;wire n3285;wire n3286;wire n3287;wire n3288;wire n3289;wire n3290;wire n3291;wire n3292;wire n3293;wire n3294;wire n3295;wire n3296;wire n3297;wire n3298;wire n3299;wire n3300;wire n3301;wire n3302;wire n3303;wire n3304;wire n3305;wire n3306;wire n3307;wire n3308;wire n3309;wire n3310;wire n3311;wire n3312;wire n3313;wire n3314;wire n3315;wire n3316;wire n3317;wire n3318;wire n3319;wire n3320;wire n3321;wire n3322;wire n3323;wire n3324;wire n3325;wire n3326;wire n3327;wire n3328;wire n3329;wire n3330;wire n3331;wire n3332;wire n3333;wire n3334;wire n3335;wire n3336;wire n3337;wire n3338;wire n3339;wire n3340;wire n3341;wire n3342;wire n3343;wire n3344;wire n3345;wire n3346;wire n3347;wire n3348;wire n3349;wire n3350;wire n3351;wire n3352;wire n3353;wire n3354;wire n3355;wire n3356;wire n3357;wire n3358;wire n3359;wire n3360;wire n3361;wire n3362;wire n3363;wire n3364;wire n3365;wire n3366;wire n3367;wire n3368;wire n3369;wire n3370;wire n3371;wire n3372;wire n3373;wire n3374;wire n3375;wire n3376;wire n3377;wire n3378;wire n3379;wire n3380;wire n3381;wire n3382;wire n3383;wire n3384;wire n3385;wire n3386;wire n3387;wire n3388;wire n3389;wire n3390;wire n3391;wire n3392;wire n3393;wire n3394;wire n3395;wire n3396;wire n3397;wire n3398;wire n3399;wire n3400;wire n3401;wire n3402;wire n3403;wire n3404;wire n3405;wire n3406;wire n3407;wire n3408;wire n3409;wire n3410;wire n3411;wire n3412;wire n3413;wire n3414;wire n3415;wire n3416;wire n3417;wire n3418;wire n3419;wire n3420;wire n3421;wire n3422;wire n3423;wire n3424;wire n3425;wire n3426;wire n3427;wire n3428;wire n3429;wire n3430;wire n3431;wire n3432;wire n3433;wire n3434;wire n3435;wire n3436;wire n3437;wire n3438;wire n3439;wire n3440;wire n3441;wire n3442;wire n3443;wire n3444;wire n3445;wire n3446;wire n3447;wire n3448;wire n3449;wire n3450;wire n3451;wire n3452;wire n3453;wire n3454;wire n3455;wire n3456;wire n3457;wire n3458;wire n3459;wire n3460;wire n3461;wire n3462;wire n3463;wire n3464;wire n3465;wire n3466;wire n3467;wire n3468;wire n3469;wire n3470;wire n3471;wire n3472;wire n3473;wire n3474;wire n3475;wire n3476;wire n3477;wire n3478;wire n3479;wire n3480;wire n3481;wire n3482;wire n3483;wire n3484;wire n3485;wire n3486;wire n3487;wire n3488;wire n3489;wire n3490;wire n3491;wire n3492;wire n3493;wire n3494;wire n3495;wire n3496;wire n3497;wire n3498;wire n3499;wire n3500;wire n3501;wire n3502;wire n3503;wire n3504;wire n3505;wire n3506;wire n3507;wire n3508;wire n3509;wire n3510;wire n3511;wire n3512;wire n3513;wire n3514;wire n3515;wire n3516;wire n3517;wire n3518;wire n3519;wire n3520;wire n3521;wire n3522;wire n3523;wire n3524;wire n3525;wire n3526;wire n3527;wire n3528;wire n3529;wire n3530;wire n3531;wire n3532;wire n3533;wire n3534;wire n3535;wire n3536;wire n3537;wire n3538;wire n3539;wire n3540;wire n3541;wire n3542;wire n3543;wire n3544;wire n3545;wire n3546;wire n3547;wire n3548;wire n3549;wire n3550;wire n3551;wire n3552;wire n3553;wire n3554;wire n3555;wire n3556;wire n3557;wire n3558;wire n3559;wire n3560;wire n3561;wire n3562;wire n3563;wire n3564;wire n3565;wire n3566;wire n3567;wire n3568;wire n3569;wire n3570;wire n3571;wire n3572;wire n3573;wire n3574;wire n3575;wire n3576;wire n3577;wire n3578;wire n3579;wire n3580;wire n3581;wire n3582;wire n3583;wire n3584;wire n3585;wire n3586;wire n3587;wire n3588;wire n3589;wire n3590;wire n3591;wire n3592;wire n3593;wire n3594;wire n3595;wire n3596;wire n3597;wire n3598;wire n3599;wire n3600;wire n3601;wire n3602;wire n3603;wire n3604;wire n3605;wire n3606;wire n3607;wire n3608;wire n3609;wire n3610;wire n3611;wire n3612;wire n3613;wire n3614;wire n3615;wire n3616;wire n3617;wire n3618;wire n3619;wire n3620;wire n3621;wire n3622;wire n3623;wire n3624;wire n3625;wire n3626;wire n3627;wire n3628;wire n3629;wire n3630;wire n3631;wire n3632;wire n3633;wire n3634;wire n3635;wire n3636;wire n3637;wire n3638;wire n3639;wire n3640;wire n3641;wire n3642;wire n3643;wire n3644;wire n3645;wire n3646;wire n3647;wire n3648;wire n3649;wire n3650;wire n3651;wire n3652;wire n3653;wire n3654;wire n3655;wire n3656;wire n3657;wire n3658;wire n3659;wire n3660;wire n3661;wire n3662;wire n3663;wire n3664;wire n3665;wire n3666;wire n3667;wire n3668;wire n3669;wire n3670;wire n3671;wire n3672;wire n3673;wire n3674;wire n3675;wire n3676;wire n3677;wire n3678;wire n3679;wire n3680;wire n3681;wire n3682;wire n3683;wire n3684;wire n3685;wire n3686;wire n3687;wire n3688;wire n3689;wire n3690;wire n3691;wire n3692;wire n3693;wire n3694;wire n3695;wire n3696;wire n3697;wire n3698;wire n3699;wire n3700;wire n3701;wire n3702;wire n3703;wire n3704;wire n3705;wire n3706;wire n3707;wire n3708;wire n3709;wire n3710;wire n3711;wire n3712;wire n3713;wire n3714;wire n3715;wire n3716;wire n3717;wire n3718;wire n3719;wire n3720;wire n3721;wire n3722;wire n3723;wire n3724;wire n3725;wire n3726;wire n3727;wire n3728;wire n3729;wire n3730;wire n3731;wire n3732;wire n3733;wire n3734;wire n3735;wire n3736;wire n3737;wire n3738;wire n3739;wire n3740;wire n3741;wire n3742;wire n3743;wire n3744;wire n3745;wire n3746;wire n3747;wire n3748;wire n3749;wire n3751;wire n3752;wire n3753;wire n3754;wire n3755;wire n3756;wire n3757;wire n3758;wire n3759;wire n3760;wire n3761;wire n3762;wire n3763;wire n3764;wire n3765;wire n3766;wire n3767;wire n3768;wire n3769;wire n3770;wire n3771;wire n3772;wire n3773;wire n3774;wire n3775;wire n3776;wire n3777;wire n3778;wire n3779;wire n3780;wire n3781;wire n3782;wire n3783;wire n3784;wire n3785;wire n3786;wire n3787;wire n3788;wire n3789;wire n3790;wire n3791;wire n3792;wire n3793;wire n3794;wire n3795;wire n3796;wire n3797;wire n3798;wire n3799;wire n3800;wire n3801;wire n3802;wire n3803;wire n3804;wire n3805;wire n3806;wire n3807;wire n3808;wire n3809;wire n3810;wire n3811;wire n3812;wire n3813;wire n3814;wire n3815;wire n3816;wire n3817;wire n3818;wire n3819;wire n3820;wire n3821;wire n3822;wire n3823;wire n3824;wire n3825;wire n3826;wire n3827;wire n3828;wire n3829;wire n3830;wire n3831;wire n3832;wire n3833;wire n3834;wire n3835;wire n3836;wire n3837;wire n3838;wire n3839;wire n3840;wire n3841;wire n3842;wire n3843;wire n3844;wire n3845;wire n3846;wire n3847;wire n3848;wire n3849;wire n3850;wire n3851;wire n3852;wire n3853;wire n3854;wire n3855;wire n3856;wire n3857;wire n3858;wire n3859;wire n3860;wire n3861;wire n3862;wire n3863;wire n3864;wire n3865;wire n3866;wire n3867;wire n3868;wire n3869;wire n3870;wire n3871;wire n3872;wire n3873;wire n3874;wire n3875;wire n3876;wire n3877;wire n3878;wire n3880;wire n3881;wire n3882;wire n3883;wire n3885;wire n3886;wire n3887;wire n3888;wire n3889;wire n3890;wire n3891;wire n3892;wire n3893;wire n3894;wire n3895;wire n3896;wire n3897;wire n3898;wire n3899;wire n3900;wire n3901;wire n3902;wire n3903;wire n3904;wire n3905;wire n3906;wire n3907;wire n3908;wire n3909;wire n3910;wire n3911;wire n3915;wire n3916;wire n3923;wire n3925;wire n3927;wire n3928;wire n3929;wire n3930;wire n3931;wire n3932;wire n3933;wire n3934;wire n3935;wire n3936;wire n3937;wire n3938;wire n3939;wire n3940;wire n3941;wire n3942;wire n3943;wire n3944;wire n3945;wire n3946;wire n3947;wire n3948;wire n3949;wire n3950;wire n3951;wire n3952;wire n3953;wire n3954;wire n3955;wire n3956;wire n3957;wire n3958;wire n3959;wire n3960;wire n3961;wire n3962;wire n3963;wire n3964;wire n3965;wire n3966;wire n3967;wire n3968;wire n3969;wire n3970;wire n3971;wire n3972;wire n3973;wire n3974;wire n3975;wire n3976;wire n3977;wire n3978;wire n3979;wire n3980;wire n3983;wire n3997;wire n3998;wire n3999;wire n4000;wire n4001;wire n4002;wire n4003;wire n4004;wire n4005;wire n4006;wire n4007;wire n4008;wire n4009;wire n4010;wire n4011;wire n4012;wire n4013;wire n4014;wire n4015;wire n4016;wire n4017;wire n4018;wire n4019;wire n4020;wire n4021;wire n4022;wire n4023;wire n4024;wire n4025;wire n4026;wire n4027;wire n4028;wire n4029;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n156,
    n32
  );


  buf
  g1
  (
    n87,
    n8
  );


  buf
  g2
  (
    n119,
    n10
  );


  not
  g3
  (
    n88,
    n11
  );


  not
  g4
  (
    n41,
    n7
  );


  buf
  g5
  (
    n58,
    n22
  );


  not
  g6
  (
    n134,
    n3
  );


  buf
  g7
  (
    n104,
    n30
  );


  not
  g8
  (
    n64,
    n20
  );


  not
  g9
  (
    n154,
    n21
  );


  not
  g10
  (
    n85,
    n28
  );


  not
  g11
  (
    n48,
    n5
  );


  buf
  g12
  (
    n128,
    n32
  );


  not
  g13
  (
    n94,
    n18
  );


  not
  g14
  (
    n69,
    n6
  );


  buf
  g15
  (
    n149,
    n16
  );


  not
  g16
  (
    n114,
    n6
  );


  buf
  g17
  (
    n135,
    n29
  );


  not
  g18
  (
    n144,
    n17
  );


  buf
  g19
  (
    n72,
    n20
  );


  buf
  g20
  (
    n99,
    n5
  );


  buf
  g21
  (
    n146,
    n4
  );


  buf
  g22
  (
    n147,
    n29
  );


  not
  g23
  (
    n118,
    n2
  );


  not
  g24
  (
    n120,
    n31
  );


  not
  g25
  (
    n49,
    n32
  );


  not
  g26
  (
    n92,
    n16
  );


  buf
  g27
  (
    n122,
    n6
  );


  buf
  g28
  (
    n65,
    n24
  );


  not
  g29
  (
    n39,
    n25
  );


  buf
  g30
  (
    n59,
    n11
  );


  buf
  g31
  (
    n38,
    n24
  );


  buf
  g32
  (
    n62,
    n24
  );


  not
  g33
  (
    n133,
    n18
  );


  not
  g34
  (
    n117,
    n7
  );


  not
  g35
  (
    n155,
    n29
  );


  not
  g36
  (
    n74,
    n19
  );


  buf
  g37
  (
    n121,
    n23
  );


  buf
  g38
  (
    n159,
    n8
  );


  not
  g39
  (
    n53,
    n14
  );


  not
  g40
  (
    n66,
    n27
  );


  buf
  g41
  (
    n97,
    n27
  );


  not
  g42
  (
    n110,
    n8
  );


  not
  g43
  (
    n145,
    n5
  );


  buf
  g44
  (
    n130,
    n26
  );


  buf
  g45
  (
    n56,
    n13
  );


  buf
  g46
  (
    n109,
    n31
  );


  buf
  g47
  (
    n127,
    n7
  );


  not
  g48
  (
    n140,
    n27
  );


  not
  g49
  (
    n116,
    n9
  );


  not
  g50
  (
    n153,
    n12
  );


  buf
  g51
  (
    n141,
    n21
  );


  not
  g52
  (
    n79,
    n9
  );


  buf
  g53
  (
    n158,
    n9
  );


  buf
  g54
  (
    n46,
    n17
  );


  buf
  g55
  (
    n40,
    n15
  );


  not
  g56
  (
    n96,
    n28
  );


  not
  g57
  (
    n45,
    n3
  );


  buf
  g58
  (
    n106,
    n16
  );


  not
  g59
  (
    n150,
    n12
  );


  not
  g60
  (
    n131,
    n23
  );


  not
  g61
  (
    n35,
    n28
  );


  not
  g62
  (
    n44,
    n16
  );


  buf
  g63
  (
    n107,
    n14
  );


  not
  g64
  (
    n86,
    n1
  );


  not
  g65
  (
    n105,
    n4
  );


  not
  g66
  (
    n36,
    n22
  );


  not
  g67
  (
    n42,
    n13
  );


  buf
  g68
  (
    n126,
    n22
  );


  not
  g69
  (
    n34,
    n30
  );


  buf
  g70
  (
    n148,
    n21
  );


  buf
  g71
  (
    n47,
    n22
  );


  not
  g72
  (
    n90,
    n25
  );


  not
  g73
  (
    n68,
    n4
  );


  buf
  g74
  (
    n137,
    n7
  );


  not
  g75
  (
    n33,
    n24
  );


  not
  g76
  (
    n95,
    n3
  );


  buf
  g77
  (
    n73,
    n19
  );


  not
  g78
  (
    n51,
    n13
  );


  buf
  g79
  (
    n83,
    n25
  );


  not
  g80
  (
    n143,
    n13
  );


  buf
  g81
  (
    n123,
    n17
  );


  not
  g82
  (
    n81,
    n4
  );


  not
  g83
  (
    n60,
    n6
  );


  not
  g84
  (
    n152,
    n9
  );


  not
  g85
  (
    n52,
    n12
  );


  not
  g86
  (
    n71,
    n26
  );


  not
  g87
  (
    n103,
    n11
  );


  not
  g88
  (
    n84,
    n20
  );


  buf
  g89
  (
    n111,
    n19
  );


  not
  g90
  (
    n112,
    n30
  );


  not
  g91
  (
    n78,
    n10
  );


  not
  g92
  (
    n113,
    n25
  );


  not
  g93
  (
    n43,
    n15
  );


  buf
  g94
  (
    n139,
    n19
  );


  buf
  g95
  (
    n91,
    n27
  );


  not
  g96
  (
    n76,
    n18
  );


  buf
  g97
  (
    n93,
    n15
  );


  not
  g98
  (
    n124,
    n10
  );


  not
  g99
  (
    n57,
    n20
  );


  buf
  g100
  (
    n70,
    n2
  );


  buf
  g101
  (
    n132,
    n31
  );


  buf
  g102
  (
    n102,
    n14
  );


  not
  g103
  (
    n54,
    n5
  );


  buf
  g104
  (
    n160,
    n17
  );


  not
  g105
  (
    n98,
    n14
  );


  buf
  g106
  (
    n55,
    n26
  );


  buf
  g107
  (
    n142,
    n21
  );


  not
  g108
  (
    n138,
    n3
  );


  buf
  g109
  (
    n115,
    n12
  );


  buf
  g110
  (
    n77,
    n28
  );


  not
  g111
  (
    n63,
    n18
  );


  not
  g112
  (
    n136,
    n2
  );


  not
  g113
  (
    n80,
    n26
  );


  buf
  g114
  (
    n101,
    n23
  );


  buf
  g115
  (
    n129,
    n1
  );


  buf
  g116
  (
    n151,
    n31
  );


  not
  g117
  (
    n61,
    n23
  );


  buf
  g118
  (
    n67,
    n1
  );


  buf
  g119
  (
    n82,
    n10
  );


  not
  g120
  (
    n89,
    n32
  );


  buf
  g121
  (
    n157,
    n2
  );


  buf
  g122
  (
    n108,
    n11
  );


  not
  g123
  (
    n37,
    n1
  );


  buf
  g124
  (
    n100,
    n15
  );


  not
  g125
  (
    n50,
    n8
  );


  buf
  g126
  (
    n75,
    n29
  );


  buf
  g127
  (
    n125,
    n30
  );


  not
  g128
  (
    n386,
    n141
  );


  not
  g129
  (
    n521,
    n112
  );


  not
  g130
  (
    n325,
    n47
  );


  not
  g131
  (
    n404,
    n81
  );


  buf
  g132
  (
    n387,
    n38
  );


  not
  g133
  (
    n458,
    n120
  );


  buf
  g134
  (
    n168,
    n66
  );


  buf
  g135
  (
    n343,
    n84
  );


  not
  g136
  (
    n527,
    n99
  );


  buf
  g137
  (
    n487,
    n141
  );


  not
  g138
  (
    n600,
    n149
  );


  not
  g139
  (
    n226,
    n128
  );


  buf
  g140
  (
    n162,
    n159
  );


  buf
  g141
  (
    n503,
    n43
  );


  buf
  g142
  (
    n353,
    n124
  );


  buf
  g143
  (
    n562,
    n126
  );


  buf
  g144
  (
    n219,
    n81
  );


  buf
  g145
  (
    n258,
    n113
  );


  not
  g146
  (
    n557,
    n72
  );


  not
  g147
  (
    n582,
    n144
  );


  not
  g148
  (
    n260,
    n153
  );


  not
  g149
  (
    n237,
    n47
  );


  not
  g150
  (
    n516,
    n155
  );


  buf
  g151
  (
    n351,
    n82
  );


  buf
  g152
  (
    n310,
    n133
  );


  buf
  g153
  (
    n267,
    n33
  );


  not
  g154
  (
    n482,
    n68
  );


  buf
  g155
  (
    n463,
    n121
  );


  not
  g156
  (
    n427,
    n96
  );


  buf
  g157
  (
    n502,
    n133
  );


  not
  g158
  (
    n259,
    n149
  );


  buf
  g159
  (
    n570,
    n41
  );


  not
  g160
  (
    n576,
    n86
  );


  buf
  g161
  (
    n672,
    n82
  );


  buf
  g162
  (
    n640,
    n154
  );


  buf
  g163
  (
    n435,
    n145
  );


  not
  g164
  (
    n328,
    n46
  );


  buf
  g165
  (
    n432,
    n126
  );


  buf
  g166
  (
    n323,
    n138
  );


  not
  g167
  (
    n255,
    n92
  );


  buf
  g168
  (
    n401,
    n73
  );


  not
  g169
  (
    n541,
    n147
  );


  buf
  g170
  (
    n249,
    n134
  );


  buf
  g171
  (
    n395,
    n43
  );


  not
  g172
  (
    n359,
    n130
  );


  not
  g173
  (
    n641,
    n42
  );


  buf
  g174
  (
    n397,
    n84
  );


  buf
  g175
  (
    n410,
    n61
  );


  not
  g176
  (
    n306,
    n98
  );


  not
  g177
  (
    n592,
    n136
  );


  buf
  g178
  (
    n468,
    n80
  );


  buf
  g179
  (
    n302,
    n106
  );


  not
  g180
  (
    n202,
    n95
  );


  buf
  g181
  (
    n301,
    n82
  );


  buf
  g182
  (
    n304,
    n45
  );


  not
  g183
  (
    n393,
    n117
  );


  buf
  g184
  (
    n519,
    n121
  );


  buf
  g185
  (
    n256,
    n39
  );


  buf
  g186
  (
    n426,
    n102
  );


  not
  g187
  (
    n480,
    n145
  );


  not
  g188
  (
    n244,
    n104
  );


  buf
  g189
  (
    n455,
    n70
  );


  buf
  g190
  (
    n470,
    n74
  );


  buf
  g191
  (
    n217,
    n107
  );


  buf
  g192
  (
    n645,
    n77
  );


  not
  g193
  (
    n383,
    n115
  );


  not
  g194
  (
    n424,
    n120
  );


  not
  g195
  (
    n370,
    n117
  );


  buf
  g196
  (
    n634,
    n149
  );


  buf
  g197
  (
    n291,
    n145
  );


  not
  g198
  (
    n510,
    n109
  );


  not
  g199
  (
    n668,
    n80
  );


  buf
  g200
  (
    n170,
    n151
  );


  not
  g201
  (
    n529,
    n158
  );


  not
  g202
  (
    n218,
    n38
  );


  not
  g203
  (
    n329,
    n63
  );


  buf
  g204
  (
    n484,
    n79
  );


  not
  g205
  (
    n501,
    n137
  );


  not
  g206
  (
    n282,
    n53
  );


  buf
  g207
  (
    n284,
    n116
  );


  not
  g208
  (
    n409,
    n64
  );


  not
  g209
  (
    n615,
    n153
  );


  buf
  g210
  (
    n561,
    n122
  );


  not
  g211
  (
    n415,
    n115
  );


  buf
  g212
  (
    n498,
    n140
  );


  not
  g213
  (
    n209,
    n151
  );


  not
  g214
  (
    n220,
    n98
  );


  not
  g215
  (
    n621,
    n91
  );


  buf
  g216
  (
    n382,
    n78
  );


  not
  g217
  (
    n192,
    n59
  );


  buf
  g218
  (
    n188,
    n55
  );


  buf
  g219
  (
    n210,
    n34
  );


  not
  g220
  (
    n368,
    n111
  );


  not
  g221
  (
    n273,
    n152
  );


  not
  g222
  (
    n491,
    n65
  );


  buf
  g223
  (
    n476,
    n69
  );


  not
  g224
  (
    n546,
    n160
  );


  buf
  g225
  (
    n405,
    n84
  );


  buf
  g226
  (
    n474,
    n34
  );


  buf
  g227
  (
    n337,
    n131
  );


  buf
  g228
  (
    n173,
    n136
  );


  buf
  g229
  (
    n224,
    n111
  );


  buf
  g230
  (
    n591,
    n53
  );


  buf
  g231
  (
    n646,
    n100
  );


  not
  g232
  (
    n315,
    n119
  );


  not
  g233
  (
    n185,
    n118
  );


  buf
  g234
  (
    n272,
    n157
  );


  buf
  g235
  (
    n614,
    n44
  );


  buf
  g236
  (
    n268,
    n150
  );


  not
  g237
  (
    n633,
    n104
  );


  buf
  g238
  (
    n664,
    n160
  );


  not
  g239
  (
    n593,
    n67
  );


  not
  g240
  (
    n590,
    n105
  );


  not
  g241
  (
    n264,
    n59
  );


  not
  g242
  (
    n183,
    n103
  );


  not
  g243
  (
    n605,
    n64
  );


  buf
  g244
  (
    n396,
    n45
  );


  not
  g245
  (
    n620,
    n126
  );


  not
  g246
  (
    n342,
    n140
  );


  not
  g247
  (
    n610,
    n153
  );


  buf
  g248
  (
    n367,
    n123
  );


  buf
  g249
  (
    n438,
    n44
  );


  not
  g250
  (
    n241,
    n56
  );


  buf
  g251
  (
    n622,
    n56
  );


  buf
  g252
  (
    n652,
    n33
  );


  buf
  g253
  (
    n662,
    n96
  );


  not
  g254
  (
    n371,
    n99
  );


  buf
  g255
  (
    n230,
    n57
  );


  buf
  g256
  (
    n511,
    n108
  );


  not
  g257
  (
    n626,
    n106
  );


  not
  g258
  (
    n603,
    n100
  );


  buf
  g259
  (
    n618,
    n93
  );


  not
  g260
  (
    n366,
    n41
  );


  not
  g261
  (
    n655,
    n106
  );


  buf
  g262
  (
    n317,
    n57
  );


  not
  g263
  (
    n481,
    n159
  );


  buf
  g264
  (
    n670,
    n152
  );


  not
  g265
  (
    n171,
    n45
  );


  buf
  g266
  (
    n617,
    n154
  );


  not
  g267
  (
    n178,
    n113
  );


  buf
  g268
  (
    n240,
    n84
  );


  not
  g269
  (
    n214,
    n75
  );


  not
  g270
  (
    n245,
    n86
  );


  buf
  g271
  (
    n642,
    n62
  );


  buf
  g272
  (
    n669,
    n146
  );


  not
  g273
  (
    n475,
    n102
  );


  buf
  g274
  (
    n335,
    n49
  );


  buf
  g275
  (
    n212,
    n70
  );


  buf
  g276
  (
    n186,
    n50
  );


  not
  g277
  (
    n316,
    n42
  );


  buf
  g278
  (
    n211,
    n89
  );


  not
  g279
  (
    n454,
    n118
  );


  buf
  g280
  (
    n189,
    n33
  );


  buf
  g281
  (
    n281,
    n117
  );


  not
  g282
  (
    n198,
    n158
  );


  not
  g283
  (
    n201,
    n74
  );


  not
  g284
  (
    n336,
    n142
  );


  not
  g285
  (
    n638,
    n72
  );


  buf
  g286
  (
    n456,
    n71
  );


  not
  g287
  (
    n307,
    n62
  );


  buf
  g288
  (
    n653,
    n108
  );


  buf
  g289
  (
    n538,
    n87
  );


  not
  g290
  (
    n631,
    n61
  );


  buf
  g291
  (
    n577,
    n63
  );


  buf
  g292
  (
    n195,
    n135
  );


  buf
  g293
  (
    n563,
    n134
  );


  not
  g294
  (
    n449,
    n131
  );


  buf
  g295
  (
    n632,
    n146
  );


  buf
  g296
  (
    n313,
    n157
  );


  not
  g297
  (
    n453,
    n141
  );


  not
  g298
  (
    n190,
    n43
  );


  buf
  g299
  (
    n191,
    n142
  );


  buf
  g300
  (
    n263,
    n142
  );


  not
  g301
  (
    n554,
    n36
  );


  not
  g302
  (
    n347,
    n48
  );


  buf
  g303
  (
    n450,
    n103
  );


  buf
  g304
  (
    n479,
    n61
  );


  buf
  g305
  (
    n630,
    n90
  );


  buf
  g306
  (
    n276,
    n110
  );


  buf
  g307
  (
    n445,
    n73
  );


  not
  g308
  (
    n251,
    n109
  );


  not
  g309
  (
    n526,
    n144
  );


  not
  g310
  (
    n536,
    n128
  );


  not
  g311
  (
    n492,
    n54
  );


  not
  g312
  (
    n609,
    n62
  );


  buf
  g313
  (
    n571,
    n116
  );


  buf
  g314
  (
    n231,
    n45
  );


  buf
  g315
  (
    n585,
    n65
  );


  not
  g316
  (
    n277,
    n147
  );


  not
  g317
  (
    n583,
    n66
  );


  not
  g318
  (
    n373,
    n107
  );


  buf
  g319
  (
    n514,
    n152
  );


  buf
  g320
  (
    n419,
    n47
  );


  buf
  g321
  (
    n459,
    n40
  );


  buf
  g322
  (
    n352,
    n42
  );


  buf
  g323
  (
    n391,
    n56
  );


  not
  g324
  (
    n362,
    n83
  );


  buf
  g325
  (
    n250,
    n97
  );


  buf
  g326
  (
    n385,
    n102
  );


  buf
  g327
  (
    n208,
    n61
  );


  buf
  g328
  (
    n176,
    n140
  );


  not
  g329
  (
    n627,
    n95
  );


  buf
  g330
  (
    n493,
    n96
  );


  buf
  g331
  (
    n346,
    n134
  );


  not
  g332
  (
    n232,
    n146
  );


  buf
  g333
  (
    n660,
    n150
  );


  not
  g334
  (
    n650,
    n115
  );


  not
  g335
  (
    n205,
    n128
  );


  not
  g336
  (
    n528,
    n46
  );


  buf
  g337
  (
    n381,
    n155
  );


  not
  g338
  (
    n206,
    n153
  );


  buf
  g339
  (
    n547,
    n90
  );


  not
  g340
  (
    n579,
    n131
  );


  buf
  g341
  (
    n215,
    n50
  );


  buf
  g342
  (
    n629,
    n148
  );


  buf
  g343
  (
    n242,
    n124
  );


  buf
  g344
  (
    n418,
    n54
  );


  buf
  g345
  (
    n166,
    n85
  );


  buf
  g346
  (
    n525,
    n125
  );


  buf
  g347
  (
    n384,
    n139
  );


  buf
  g348
  (
    n169,
    n133
  );


  not
  g349
  (
    n471,
    n83
  );


  buf
  g350
  (
    n334,
    n94
  );


  buf
  g351
  (
    n535,
    n118
  );


  buf
  g352
  (
    n239,
    n104
  );


  buf
  g353
  (
    n513,
    n81
  );


  not
  g354
  (
    n661,
    n52
  );


  buf
  g355
  (
    n507,
    n69
  );


  not
  g356
  (
    n565,
    n158
  );


  buf
  g357
  (
    n540,
    n68
  );


  not
  g358
  (
    n278,
    n89
  );


  buf
  g359
  (
    n270,
    n75
  );


  buf
  g360
  (
    n442,
    n86
  );


  buf
  g361
  (
    n515,
    n59
  );


  buf
  g362
  (
    n196,
    n130
  );


  buf
  g363
  (
    n477,
    n72
  );


  buf
  g364
  (
    n604,
    n110
  );


  not
  g365
  (
    n443,
    n48
  );


  buf
  g366
  (
    n567,
    n33
  );


  not
  g367
  (
    n457,
    n119
  );


  buf
  g368
  (
    n420,
    n125
  );


  buf
  g369
  (
    n663,
    n77
  );


  not
  g370
  (
    n286,
    n160
  );


  not
  g371
  (
    n539,
    n38
  );


  buf
  g372
  (
    n564,
    n101
  );


  not
  g373
  (
    n625,
    n34
  );


  buf
  g374
  (
    n437,
    n124
  );


  not
  g375
  (
    n376,
    n99
  );


  buf
  g376
  (
    n413,
    n129
  );


  not
  g377
  (
    n506,
    n103
  );


  not
  g378
  (
    n187,
    n54
  );


  not
  g379
  (
    n324,
    n53
  );


  buf
  g380
  (
    n560,
    n94
  );


  buf
  g381
  (
    n594,
    n121
  );


  not
  g382
  (
    n303,
    n137
  );


  not
  g383
  (
    n222,
    n129
  );


  buf
  g384
  (
    n364,
    n141
  );


  not
  g385
  (
    n300,
    n143
  );


  buf
  g386
  (
    n283,
    n88
  );


  not
  g387
  (
    n573,
    n88
  );


  not
  g388
  (
    n164,
    n62
  );


  buf
  g389
  (
    n466,
    n114
  );


  not
  g390
  (
    n262,
    n79
  );


  not
  g391
  (
    n483,
    n79
  );


  buf
  g392
  (
    n327,
    n97
  );


  buf
  g393
  (
    n665,
    n60
  );


  buf
  g394
  (
    n428,
    n101
  );


  not
  g395
  (
    n568,
    n37
  );


  buf
  g396
  (
    n549,
    n95
  );


  buf
  g397
  (
    n265,
    n120
  );


  not
  g398
  (
    n531,
    n112
  );


  buf
  g399
  (
    n586,
    n77
  );


  buf
  g400
  (
    n490,
    n131
  );


  buf
  g401
  (
    n271,
    n80
  );


  not
  g402
  (
    n509,
    n73
  );


  buf
  g403
  (
    n274,
    n91
  );


  not
  g404
  (
    n326,
    n66
  );


  buf
  g405
  (
    n414,
    n157
  );


  buf
  g406
  (
    n207,
    n156
  );


  buf
  g407
  (
    n165,
    n78
  );


  buf
  g408
  (
    n223,
    n74
  );


  not
  g409
  (
    n377,
    n100
  );


  buf
  g410
  (
    n299,
    n93
  );


  not
  g411
  (
    n447,
    n156
  );


  not
  g412
  (
    n279,
    n100
  );


  not
  g413
  (
    n394,
    n111
  );


  buf
  g414
  (
    n321,
    n132
  );


  not
  g415
  (
    n446,
    n55
  );


  buf
  g416
  (
    n553,
    n49
  );


  not
  g417
  (
    n365,
    n159
  );


  not
  g418
  (
    n194,
    n122
  );


  buf
  g419
  (
    n497,
    n35
  );


  buf
  g420
  (
    n294,
    n87
  );


  buf
  g421
  (
    n524,
    n37
  );


  buf
  g422
  (
    n275,
    n50
  );


  buf
  g423
  (
    n460,
    n123
  );


  not
  g424
  (
    n597,
    n88
  );


  buf
  g425
  (
    n318,
    n36
  );


  buf
  g426
  (
    n587,
    n39
  );


  buf
  g427
  (
    n289,
    n51
  );


  buf
  g428
  (
    n486,
    n109
  );


  buf
  g429
  (
    n234,
    n51
  );


  buf
  g430
  (
    n656,
    n78
  );


  buf
  g431
  (
    n462,
    n64
  );


  buf
  g432
  (
    n292,
    n41
  );


  not
  g433
  (
    n236,
    n57
  );


  buf
  g434
  (
    n545,
    n92
  );


  not
  g435
  (
    n623,
    n75
  );


  not
  g436
  (
    n379,
    n91
  );


  not
  g437
  (
    n344,
    n99
  );


  buf
  g438
  (
    n312,
    n107
  );


  not
  g439
  (
    n174,
    n146
  );


  buf
  g440
  (
    n374,
    n135
  );


  buf
  g441
  (
    n649,
    n155
  );


  buf
  g442
  (
    n216,
    n156
  );


  not
  g443
  (
    n494,
    n53
  );


  not
  g444
  (
    n602,
    n150
  );


  not
  g445
  (
    n651,
    n143
  );


  buf
  g446
  (
    n402,
    n157
  );


  not
  g447
  (
    n555,
    n50
  );


  not
  g448
  (
    n425,
    n101
  );


  buf
  g449
  (
    n512,
    n90
  );


  not
  g450
  (
    n473,
    n69
  );


  not
  g451
  (
    n430,
    n137
  );


  not
  g452
  (
    n363,
    n122
  );


  buf
  g453
  (
    n197,
    n119
  );


  not
  g454
  (
    n422,
    n69
  );


  buf
  g455
  (
    n348,
    n136
  );


  buf
  g456
  (
    n578,
    n75
  );


  buf
  g457
  (
    n532,
    n51
  );


  buf
  g458
  (
    n261,
    n80
  );


  buf
  g459
  (
    n180,
    n158
  );


  not
  g460
  (
    n350,
    n136
  );


  buf
  g461
  (
    n406,
    n134
  );


  buf
  g462
  (
    n588,
    n144
  );


  not
  g463
  (
    n247,
    n40
  );


  not
  g464
  (
    n297,
    n124
  );


  buf
  g465
  (
    n530,
    n140
  );


  not
  g466
  (
    n671,
    n101
  );


  not
  g467
  (
    n647,
    n56
  );


  buf
  g468
  (
    n248,
    n48
  );


  buf
  g469
  (
    n558,
    n105
  );


  not
  g470
  (
    n411,
    n132
  );


  buf
  g471
  (
    n559,
    n113
  );


  buf
  g472
  (
    n360,
    n96
  );


  not
  g473
  (
    n666,
    n154
  );


  not
  g474
  (
    n552,
    n102
  );


  not
  g475
  (
    n581,
    n76
  );


  buf
  g476
  (
    n574,
    n155
  );


  buf
  g477
  (
    n569,
    n154
  );


  not
  g478
  (
    n499,
    n85
  );


  not
  g479
  (
    n254,
    n64
  );


  buf
  g480
  (
    n575,
    n123
  );


  buf
  g481
  (
    n508,
    n130
  );


  buf
  g482
  (
    n416,
    n72
  );


  buf
  g483
  (
    n612,
    n119
  );


  not
  g484
  (
    n252,
    n98
  );


  not
  g485
  (
    n203,
    n148
  );


  buf
  g486
  (
    n182,
    n129
  );


  buf
  g487
  (
    n534,
    n48
  );


  buf
  g488
  (
    n338,
    n41
  );


  buf
  g489
  (
    n355,
    n121
  );


  buf
  g490
  (
    n533,
    n127
  );


  not
  g491
  (
    n333,
    n127
  );


  not
  g492
  (
    n167,
    n143
  );


  not
  g493
  (
    n608,
    n52
  );


  not
  g494
  (
    n319,
    n40
  );


  not
  g495
  (
    n434,
    n135
  );


  not
  g496
  (
    n330,
    n58
  );


  buf
  g497
  (
    n628,
    n67
  );


  buf
  g498
  (
    n472,
    n148
  );


  buf
  g499
  (
    n358,
    n83
  );


  not
  g500
  (
    n407,
    n43
  );


  buf
  g501
  (
    n421,
    n150
  );


  buf
  g502
  (
    n175,
    n114
  );


  not
  g503
  (
    n580,
    n104
  );


  buf
  g504
  (
    n667,
    n93
  );


  buf
  g505
  (
    n452,
    n138
  );


  not
  g506
  (
    n643,
    n125
  );


  buf
  g507
  (
    n606,
    n138
  );


  not
  g508
  (
    n349,
    n35
  );


  not
  g509
  (
    n163,
    n46
  );


  not
  g510
  (
    n305,
    n94
  );


  not
  g511
  (
    n495,
    n38
  );


  not
  g512
  (
    n522,
    n44
  );


  not
  g513
  (
    n193,
    n60
  );


  not
  g514
  (
    n172,
    n44
  );


  not
  g515
  (
    n253,
    n139
  );


  not
  g516
  (
    n357,
    n156
  );


  buf
  g517
  (
    n266,
    n118
  );


  buf
  g518
  (
    n441,
    n71
  );


  buf
  g519
  (
    n496,
    n68
  );


  not
  g520
  (
    n465,
    n66
  );


  not
  g521
  (
    n431,
    n98
  );


  not
  g522
  (
    n285,
    n58
  );


  not
  g523
  (
    n644,
    n36
  );


  buf
  g524
  (
    n398,
    n42
  );


  buf
  g525
  (
    n439,
    n142
  );


  not
  g526
  (
    n584,
    n132
  );


  buf
  g527
  (
    n200,
    n87
  );


  not
  g528
  (
    n448,
    n105
  );


  buf
  g529
  (
    n451,
    n132
  );


  not
  g530
  (
    n635,
    n145
  );


  buf
  g531
  (
    n369,
    n74
  );


  buf
  g532
  (
    n340,
    n127
  );


  not
  g533
  (
    n469,
    n108
  );


  not
  g534
  (
    n619,
    n77
  );


  buf
  g535
  (
    n380,
    n79
  );


  buf
  g536
  (
    n596,
    n147
  );


  buf
  g537
  (
    n478,
    n97
  );


  buf
  g538
  (
    n399,
    n65
  );


  not
  g539
  (
    n280,
    n111
  );


  not
  g540
  (
    n372,
    n60
  );


  buf
  g541
  (
    n296,
    n57
  );


  buf
  g542
  (
    n269,
    n93
  );


  buf
  g543
  (
    n235,
    n71
  );


  buf
  g544
  (
    n225,
    n51
  );


  not
  g545
  (
    n311,
    n137
  );


  buf
  g546
  (
    n485,
    n113
  );


  not
  g547
  (
    n436,
    n91
  );


  buf
  g548
  (
    n572,
    n114
  );


  buf
  g549
  (
    n598,
    n125
  );


  buf
  g550
  (
    n589,
    n92
  );


  buf
  g551
  (
    n551,
    n133
  );


  buf
  g552
  (
    n227,
    n130
  );


  not
  g553
  (
    n339,
    n55
  );


  buf
  g554
  (
    n293,
    n92
  );


  not
  g555
  (
    n520,
    n106
  );


  buf
  g556
  (
    n658,
    n159
  );


  buf
  g557
  (
    n566,
    n126
  );


  not
  g558
  (
    n636,
    n116
  );


  buf
  g559
  (
    n550,
    n138
  );


  not
  g560
  (
    n378,
    n109
  );


  buf
  g561
  (
    n309,
    n73
  );


  buf
  g562
  (
    n204,
    n116
  );


  buf
  g563
  (
    n177,
    n112
  );


  buf
  g564
  (
    n517,
    n94
  );


  buf
  g565
  (
    n341,
    n135
  );


  buf
  g566
  (
    n537,
    n58
  );


  buf
  g567
  (
    n213,
    n148
  );


  buf
  g568
  (
    n607,
    n63
  );


  not
  g569
  (
    n657,
    n59
  );


  buf
  g570
  (
    n354,
    n35
  );


  buf
  g571
  (
    n298,
    n86
  );


  not
  g572
  (
    n556,
    n107
  );


  buf
  g573
  (
    n199,
    n78
  );


  buf
  g574
  (
    n542,
    n55
  );


  buf
  g575
  (
    n489,
    n128
  );


  buf
  g576
  (
    n639,
    n70
  );


  buf
  g577
  (
    n659,
    n144
  );


  not
  g578
  (
    n179,
    n89
  );


  not
  g579
  (
    n221,
    n47
  );


  not
  g580
  (
    n161,
    n63
  );


  not
  g581
  (
    n308,
    n108
  );


  not
  g582
  (
    n595,
    n39
  );


  buf
  g583
  (
    n184,
    n35
  );


  buf
  g584
  (
    n464,
    n112
  );


  buf
  g585
  (
    n403,
    n143
  );


  not
  g586
  (
    n433,
    n115
  );


  not
  g587
  (
    n637,
    n52
  );


  buf
  g588
  (
    n488,
    n110
  );


  buf
  g589
  (
    n388,
    n147
  );


  buf
  g590
  (
    n288,
    n149
  );


  buf
  g591
  (
    n228,
    n95
  );


  not
  g592
  (
    n500,
    n127
  );


  not
  g593
  (
    n611,
    n117
  );


  buf
  g594
  (
    n412,
    n90
  );


  not
  g595
  (
    n601,
    n114
  );


  buf
  g596
  (
    n389,
    n87
  );


  buf
  g597
  (
    n599,
    n82
  );


  not
  g598
  (
    n314,
    n122
  );


  not
  g599
  (
    n518,
    n71
  );


  not
  g600
  (
    n408,
    n103
  );


  not
  g601
  (
    n544,
    n40
  );


  buf
  g602
  (
    n356,
    n152
  );


  not
  g603
  (
    n504,
    n139
  );


  not
  g604
  (
    n345,
    n123
  );


  buf
  g605
  (
    n461,
    n129
  );


  buf
  g606
  (
    n243,
    n81
  );


  not
  g607
  (
    n400,
    n70
  );


  not
  g608
  (
    n417,
    n39
  );


  buf
  g609
  (
    n616,
    n151
  );


  buf
  g610
  (
    n320,
    n49
  );


  buf
  g611
  (
    n613,
    n97
  );


  not
  g612
  (
    n543,
    n83
  );


  buf
  g613
  (
    n390,
    n68
  );


  not
  g614
  (
    n444,
    n34
  );


  buf
  g615
  (
    n295,
    n67
  );


  not
  g616
  (
    n429,
    n105
  );


  buf
  g617
  (
    n233,
    n67
  );


  not
  g618
  (
    n440,
    n36
  );


  not
  g619
  (
    n505,
    n120
  );


  not
  g620
  (
    n654,
    n89
  );


  not
  g621
  (
    n287,
    n160
  );


  buf
  g622
  (
    n423,
    n60
  );


  buf
  g623
  (
    n246,
    n54
  );


  not
  g624
  (
    n229,
    n49
  );


  not
  g625
  (
    n290,
    n37
  );


  not
  g626
  (
    n467,
    n151
  );


  not
  g627
  (
    n322,
    n76
  );


  not
  g628
  (
    n257,
    n76
  );


  not
  g629
  (
    n331,
    n76
  );


  not
  g630
  (
    n648,
    n46
  );


  buf
  g631
  (
    n624,
    n52
  );


  not
  g632
  (
    n238,
    n58
  );


  buf
  g633
  (
    n548,
    n139
  );


  not
  g634
  (
    n332,
    n110
  );


  buf
  g635
  (
    n181,
    n85
  );


  not
  g636
  (
    n375,
    n85
  );


  buf
  g637
  (
    n392,
    n88
  );


  not
  g638
  (
    n523,
    n37
  );


  not
  g639
  (
    n361,
    n65
  );


  not
  g640
  (
    n716,
    n183
  );


  buf
  g641
  (
    n1383,
    n171
  );


  buf
  g642
  (
    n1289,
    n226
  );


  not
  g643
  (
    n1430,
    n387
  );


  not
  g644
  (
    n1584,
    n422
  );


  not
  g645
  (
    n727,
    n569
  );


  not
  g646
  (
    n1060,
    n551
  );


  buf
  g647
  (
    n1598,
    n566
  );


  buf
  g648
  (
    n675,
    n592
  );


  buf
  g649
  (
    n987,
    n610
  );


  buf
  g650
  (
    n1394,
    n178
  );


  not
  g651
  (
    n1151,
    n613
  );


  buf
  g652
  (
    n1145,
    n199
  );


  not
  g653
  (
    n998,
    n162
  );


  not
  g654
  (
    n1277,
    n258
  );


  buf
  g655
  (
    n1220,
    n340
  );


  buf
  g656
  (
    n1555,
    n335
  );


  not
  g657
  (
    n1556,
    n307
  );


  not
  g658
  (
    n1483,
    n193
  );


  not
  g659
  (
    n1650,
    n323
  );


  buf
  g660
  (
    n856,
    n559
  );


  buf
  g661
  (
    n1272,
    n510
  );


  not
  g662
  (
    n1647,
    n658
  );


  not
  g663
  (
    n1102,
    n603
  );


  buf
  g664
  (
    n903,
    n653
  );


  buf
  g665
  (
    n677,
    n559
  );


  not
  g666
  (
    n674,
    n565
  );


  not
  g667
  (
    n682,
    n288
  );


  not
  g668
  (
    n843,
    n185
  );


  buf
  g669
  (
    n842,
    n315
  );


  not
  g670
  (
    n868,
    n206
  );


  buf
  g671
  (
    n1138,
    n221
  );


  not
  g672
  (
    n1152,
    n513
  );


  buf
  g673
  (
    n1523,
    n264
  );


  buf
  g674
  (
    n1494,
    n249
  );


  not
  g675
  (
    n1520,
    n332
  );


  not
  g676
  (
    n1617,
    n182
  );


  not
  g677
  (
    n1292,
    n568
  );


  buf
  g678
  (
    n1173,
    n519
  );


  not
  g679
  (
    n1499,
    n666
  );


  not
  g680
  (
    n887,
    n298
  );


  not
  g681
  (
    n1249,
    n191
  );


  buf
  g682
  (
    n1517,
    n460
  );


  not
  g683
  (
    n1595,
    n519
  );


  buf
  g684
  (
    n1620,
    n204
  );


  buf
  g685
  (
    n996,
    n175
  );


  buf
  g686
  (
    n1615,
    n366
  );


  buf
  g687
  (
    n730,
    n409
  );


  not
  g688
  (
    n696,
    n488
  );


  not
  g689
  (
    n934,
    n355
  );


  buf
  g690
  (
    n1099,
    n431
  );


  buf
  g691
  (
    n1259,
    n178
  );


  buf
  g692
  (
    n1509,
    n650
  );


  buf
  g693
  (
    n1547,
    n649
  );


  buf
  g694
  (
    n1548,
    n255
  );


  not
  g695
  (
    n1126,
    n593
  );


  not
  g696
  (
    n764,
    n534
  );


  not
  g697
  (
    n1117,
    n252
  );


  not
  g698
  (
    n1330,
    n667
  );


  buf
  g699
  (
    n1658,
    n196
  );


  buf
  g700
  (
    n1422,
    n186
  );


  not
  g701
  (
    n834,
    n295
  );


  not
  g702
  (
    n1589,
    n275
  );


  not
  g703
  (
    n1542,
    n470
  );


  not
  g704
  (
    n1618,
    n668
  );


  buf
  g705
  (
    n1592,
    n482
  );


  buf
  g706
  (
    n1124,
    n491
  );


  not
  g707
  (
    n959,
    n574
  );


  buf
  g708
  (
    n1680,
    n402
  );


  not
  g709
  (
    n1263,
    n203
  );


  buf
  g710
  (
    n1527,
    n316
  );


  buf
  g711
  (
    n1367,
    n304
  );


  not
  g712
  (
    n992,
    n177
  );


  buf
  g713
  (
    n1171,
    n526
  );


  buf
  g714
  (
    n1135,
    n230
  );


  buf
  g715
  (
    n732,
    n396
  );


  not
  g716
  (
    n1036,
    n310
  );


  buf
  g717
  (
    n1382,
    n448
  );


  buf
  g718
  (
    n1233,
    n179
  );


  not
  g719
  (
    n1101,
    n456
  );


  buf
  g720
  (
    n1341,
    n493
  );


  not
  g721
  (
    n809,
    n507
  );


  buf
  g722
  (
    n1626,
    n528
  );


  buf
  g723
  (
    n1693,
    n667
  );


  not
  g724
  (
    n1578,
    n397
  );


  not
  g725
  (
    n1378,
    n580
  );


  buf
  g726
  (
    n704,
    n306
  );


  buf
  g727
  (
    n1427,
    n659
  );


  not
  g728
  (
    n821,
    n375
  );


  not
  g729
  (
    n1420,
    n197
  );


  buf
  g730
  (
    n1004,
    n211
  );


  buf
  g731
  (
    n1601,
    n316
  );


  not
  g732
  (
    n1683,
    n277
  );


  not
  g733
  (
    n708,
    n326
  );


  buf
  g734
  (
    n1561,
    n490
  );


  buf
  g735
  (
    n781,
    n404
  );


  not
  g736
  (
    n1304,
    n619
  );


  buf
  g737
  (
    n961,
    n462
  );


  not
  g738
  (
    n819,
    n301
  );


  buf
  g739
  (
    n1157,
    n660
  );


  not
  g740
  (
    n744,
    n434
  );


  not
  g741
  (
    n1055,
    n315
  );


  buf
  g742
  (
    n1400,
    n350
  );


  not
  g743
  (
    n806,
    n242
  );


  buf
  g744
  (
    n837,
    n396
  );


  buf
  g745
  (
    n1264,
    n499
  );


  buf
  g746
  (
    n988,
    n411
  );


  not
  g747
  (
    n1319,
    n585
  );


  buf
  g748
  (
    n1566,
    n442
  );


  not
  g749
  (
    n1597,
    n560
  );


  buf
  g750
  (
    n1031,
    n246
  );


  not
  g751
  (
    n1487,
    n397
  );


  buf
  g752
  (
    n736,
    n470
  );


  not
  g753
  (
    n1014,
    n463
  );


  buf
  g754
  (
    n920,
    n467
  );


  not
  g755
  (
    n770,
    n478
  );


  not
  g756
  (
    n869,
    n337
  );


  not
  g757
  (
    n765,
    n613
  );


  not
  g758
  (
    n811,
    n398
  );


  not
  g759
  (
    n972,
    n407
  );


  buf
  g760
  (
    n1488,
    n581
  );


  buf
  g761
  (
    n1112,
    n182
  );


  buf
  g762
  (
    n1021,
    n188
  );


  buf
  g763
  (
    n800,
    n274
  );


  buf
  g764
  (
    n1491,
    n431
  );


  not
  g765
  (
    n928,
    n258
  );


  not
  g766
  (
    n1666,
    n397
  );


  not
  g767
  (
    n854,
    n600
  );


  buf
  g768
  (
    n1078,
    n385
  );


  buf
  g769
  (
    n1245,
    n336
  );


  not
  g770
  (
    n1602,
    n212
  );


  not
  g771
  (
    n1200,
    n554
  );


  not
  g772
  (
    n991,
    n220
  );


  not
  g773
  (
    n912,
    n376
  );


  buf
  g774
  (
    n796,
    n196
  );


  not
  g775
  (
    n1235,
    n582
  );


  buf
  g776
  (
    n805,
    n359
  );


  not
  g777
  (
    n1415,
    n401
  );


  not
  g778
  (
    n939,
    n484
  );


  not
  g779
  (
    n820,
    n257
  );


  buf
  g780
  (
    n703,
    n635
  );


  not
  g781
  (
    n1396,
    n399
  );


  not
  g782
  (
    n835,
    n425
  );


  buf
  g783
  (
    n1244,
    n286
  );


  not
  g784
  (
    n1406,
    n289
  );


  buf
  g785
  (
    n1283,
    n589
  );


  buf
  g786
  (
    n898,
    n598
  );


  not
  g787
  (
    n1239,
    n466
  );


  buf
  g788
  (
    n1194,
    n618
  );


  buf
  g789
  (
    n1552,
    n481
  );


  buf
  g790
  (
    n876,
    n497
  );


  buf
  g791
  (
    n890,
    n232
  );


  not
  g792
  (
    n1034,
    n181
  );


  buf
  g793
  (
    n1252,
    n205
  );


  not
  g794
  (
    n1366,
    n421
  );


  not
  g795
  (
    n1623,
    n496
  );


  not
  g796
  (
    n1389,
    n393
  );


  not
  g797
  (
    n795,
    n231
  );


  buf
  g798
  (
    n1388,
    n476
  );


  buf
  g799
  (
    n1166,
    n646
  );


  buf
  g800
  (
    n1248,
    n192
  );


  not
  g801
  (
    n1596,
    n504
  );


  not
  g802
  (
    n713,
    n435
  );


  buf
  g803
  (
    n1624,
    n271
  );


  buf
  g804
  (
    n1111,
    n549
  );


  buf
  g805
  (
    n892,
    n249
  );


  not
  g806
  (
    n1510,
    n486
  );


  not
  g807
  (
    n1211,
    n219
  );


  buf
  g808
  (
    n1441,
    n592
  );


  buf
  g809
  (
    n1333,
    n261
  );


  buf
  g810
  (
    n1678,
    n652
  );


  not
  g811
  (
    n1350,
    n298
  );


  buf
  g812
  (
    n709,
    n174
  );


  not
  g813
  (
    n1237,
    n590
  );


  buf
  g814
  (
    n980,
    n346
  );


  not
  g815
  (
    n1403,
    n177
  );


  not
  g816
  (
    n838,
    n169
  );


  not
  g817
  (
    n1652,
    n633
  );


  buf
  g818
  (
    n1477,
    n605
  );


  not
  g819
  (
    n1358,
    n477
  );


  buf
  g820
  (
    n1116,
    n175
  );


  buf
  g821
  (
    n1230,
    n555
  );


  not
  g822
  (
    n1447,
    n439
  );


  not
  g823
  (
    n1240,
    n165
  );


  not
  g824
  (
    n1671,
    n351
  );


  buf
  g825
  (
    n1435,
    n280
  );


  not
  g826
  (
    n1522,
    n327
  );


  buf
  g827
  (
    n1250,
    n629
  );


  not
  g828
  (
    n702,
    n222
  );


  buf
  g829
  (
    n1218,
    n556
  );


  buf
  g830
  (
    n1635,
    n323
  );


  not
  g831
  (
    n1466,
    n528
  );


  buf
  g832
  (
    n1069,
    n203
  );


  not
  g833
  (
    n1397,
    n292
  );


  buf
  g834
  (
    n719,
    n620
  );


  not
  g835
  (
    n1037,
    n264
  );


  not
  g836
  (
    n1191,
    n518
  );


  buf
  g837
  (
    n683,
    n604
  );


  buf
  g838
  (
    n1576,
    n250
  );


  not
  g839
  (
    n1500,
    n563
  );


  buf
  g840
  (
    n1558,
    n332
  );


  buf
  g841
  (
    n865,
    n552
  );


  not
  g842
  (
    n1046,
    n650
  );


  not
  g843
  (
    n687,
    n645
  );


  not
  g844
  (
    n1007,
    n580
  );


  not
  g845
  (
    n1337,
    n530
  );


  not
  g846
  (
    n1075,
    n434
  );


  buf
  g847
  (
    n699,
    n513
  );


  not
  g848
  (
    n1327,
    n430
  );


  buf
  g849
  (
    n1316,
    n317
  );


  not
  g850
  (
    n1176,
    n507
  );


  buf
  g851
  (
    n1362,
    n508
  );


  not
  g852
  (
    n977,
    n545
  );


  not
  g853
  (
    n1651,
    n406
  );


  buf
  g854
  (
    n1442,
    n555
  );


  buf
  g855
  (
    n726,
    n368
  );


  buf
  g856
  (
    n1275,
    n471
  );


  not
  g857
  (
    n1005,
    n452
  );


  buf
  g858
  (
    n1554,
    n328
  );


  not
  g859
  (
    n1674,
    n621
  );


  not
  g860
  (
    n864,
    n601
  );


  buf
  g861
  (
    n1656,
    n460
  );


  buf
  g862
  (
    n1467,
    n366
  );


  not
  g863
  (
    n1550,
    n419
  );


  buf
  g864
  (
    n1290,
    n639
  );


  not
  g865
  (
    n1519,
    n374
  );


  buf
  g866
  (
    n799,
    n480
  );


  not
  g867
  (
    n1481,
    n578
  );


  not
  g868
  (
    n1332,
    n240
  );


  not
  g869
  (
    n1073,
    n632
  );


  not
  g870
  (
    n1460,
    n186
  );


  not
  g871
  (
    n739,
    n441
  );


  not
  g872
  (
    n1204,
    n326
  );


  not
  g873
  (
    n1322,
    n296
  );


  not
  g874
  (
    n871,
    n292
  );


  buf
  g875
  (
    n1056,
    n633
  );


  buf
  g876
  (
    n1374,
    n339
  );


  buf
  g877
  (
    n841,
    n345
  );


  buf
  g878
  (
    n943,
    n549
  );


  buf
  g879
  (
    n701,
    n541
  );


  not
  g880
  (
    n1132,
    n266
  );


  buf
  g881
  (
    n1213,
    n589
  );


  not
  g882
  (
    n966,
    n631
  );


  not
  g883
  (
    n1456,
    n402
  );


  not
  g884
  (
    n907,
    n252
  );


  buf
  g885
  (
    n1521,
    n592
  );


  buf
  g886
  (
    n1604,
    n438
  );


  buf
  g887
  (
    n1190,
    n227
  );


  buf
  g888
  (
    n738,
    n400
  );


  buf
  g889
  (
    n722,
    n562
  );


  buf
  g890
  (
    n844,
    n188
  );


  buf
  g891
  (
    n1365,
    n330
  );


  not
  g892
  (
    n794,
    n450
  );


  buf
  g893
  (
    n1405,
    n276
  );


  buf
  g894
  (
    n1480,
    n367
  );


  not
  g895
  (
    n1359,
    n236
  );


  buf
  g896
  (
    n906,
    n498
  );


  not
  g897
  (
    n1090,
    n504
  );


  not
  g898
  (
    n1318,
    n343
  );


  not
  g899
  (
    n1310,
    n357
  );


  not
  g900
  (
    n1114,
    n665
  );


  not
  g901
  (
    n983,
    n666
  );


  buf
  g902
  (
    n822,
    n479
  );


  buf
  g903
  (
    n1431,
    n643
  );


  buf
  g904
  (
    n1507,
    n640
  );


  not
  g905
  (
    n1475,
    n582
  );


  not
  g906
  (
    n1363,
    n661
  );


  buf
  g907
  (
    n973,
    n282
  );


  not
  g908
  (
    n974,
    n500
  );


  buf
  g909
  (
    n1170,
    n517
  );


  not
  g910
  (
    n1209,
    n465
  );


  not
  g911
  (
    n1028,
    n625
  );


  buf
  g912
  (
    n897,
    n200
  );


  buf
  g913
  (
    n1098,
    n505
  );


  buf
  g914
  (
    n862,
    n577
  );


  not
  g915
  (
    n1454,
    n296
  );


  not
  g916
  (
    n1413,
    n316
  );


  buf
  g917
  (
    n1120,
    n475
  );


  not
  g918
  (
    n1172,
    n577
  );


  not
  g919
  (
    n882,
    n446
  );


  buf
  g920
  (
    n1670,
    n487
  );


  buf
  g921
  (
    n1089,
    n372
  );


  not
  g922
  (
    n1013,
    n247
  );


  buf
  g923
  (
    n1043,
    n558
  );


  buf
  g924
  (
    n1096,
    n359
  );


  buf
  g925
  (
    n1395,
    n223
  );


  buf
  g926
  (
    n1594,
    n425
  );


  not
  g927
  (
    n1381,
    n514
  );


  buf
  g928
  (
    n1352,
    n449
  );


  not
  g929
  (
    n923,
    n243
  );


  buf
  g930
  (
    n1305,
    n332
  );


  buf
  g931
  (
    n1546,
    n403
  );


  buf
  g932
  (
    n904,
    n163
  );


  not
  g933
  (
    n1251,
    n553
  );


  buf
  g934
  (
    n1531,
    n461
  );


  buf
  g935
  (
    n913,
    n333
  );


  not
  g936
  (
    n1052,
    n453
  );


  buf
  g937
  (
    n1147,
    n172
  );


  buf
  g938
  (
    n916,
    n574
  );


  not
  g939
  (
    n1539,
    n170
  );


  buf
  g940
  (
    n1492,
    n243
  );


  not
  g941
  (
    n1223,
    n627
  );


  buf
  g942
  (
    n824,
    n481
  );


  not
  g943
  (
    n1679,
    n281
  );


  not
  g944
  (
    n1082,
    n358
  );


  buf
  g945
  (
    n1154,
    n509
  );


  not
  g946
  (
    n958,
    n253
  );


  not
  g947
  (
    n1479,
    n348
  );


  not
  g948
  (
    n1439,
    n631
  );


  buf
  g949
  (
    n1309,
    n228
  );


  not
  g950
  (
    n1269,
    n521
  );


  buf
  g951
  (
    n932,
    n451
  );


  not
  g952
  (
    n940,
    n463
  );


  not
  g953
  (
    n896,
    n242
  );


  buf
  g954
  (
    n1105,
    n492
  );


  not
  g955
  (
    n933,
    n511
  );


  not
  g956
  (
    n1540,
    n584
  );


  buf
  g957
  (
    n1484,
    n225
  );


  not
  g958
  (
    n1164,
    n636
  );


  not
  g959
  (
    n995,
    n486
  );


  not
  g960
  (
    n1440,
    n164
  );


  buf
  g961
  (
    n758,
    n175
  );


  buf
  g962
  (
    n1009,
    n541
  );


  buf
  g963
  (
    n752,
    n252
  );


  not
  g964
  (
    n1010,
    n483
  );


  not
  g965
  (
    n1607,
    n435
  );


  not
  g966
  (
    n826,
    n512
  );


  not
  g967
  (
    n1444,
    n178
  );


  not
  g968
  (
    n1543,
    n640
  );


  buf
  g969
  (
    n782,
    n340
  );


  buf
  g970
  (
    n753,
    n205
  );


  not
  g971
  (
    n1605,
    n504
  );


  buf
  g972
  (
    n1587,
    n260
  );


  not
  g973
  (
    n691,
    n421
  );


  buf
  g974
  (
    n1434,
    n402
  );


  not
  g975
  (
    n1326,
    n246
  );


  buf
  g976
  (
    n1340,
    n631
  );


  not
  g977
  (
    n908,
    n566
  );


  buf
  g978
  (
    n927,
    n476
  );


  not
  g979
  (
    n1161,
    n418
  );


  not
  g980
  (
    n979,
    n412
  );


  not
  g981
  (
    n1364,
    n548
  );


  not
  g982
  (
    n694,
    n469
  );


  buf
  g983
  (
    n1448,
    n231
  );


  buf
  g984
  (
    n1613,
    n244
  );


  not
  g985
  (
    n1429,
    n600
  );


  buf
  g986
  (
    n1496,
    n524
  );


  buf
  g987
  (
    n1044,
    n502
  );


  buf
  g988
  (
    n1303,
    n210
  );


  buf
  g989
  (
    n737,
    n650
  );


  not
  g990
  (
    n1282,
    n384
  );


  buf
  g991
  (
    n1301,
    n467
  );


  not
  g992
  (
    n840,
    n308
  );


  buf
  g993
  (
    n1139,
    n590
  );


  not
  g994
  (
    n1625,
    n383
  );


  not
  g995
  (
    n982,
    n208
  );


  not
  g996
  (
    n1371,
    n665
  );


  buf
  g997
  (
    n1042,
    n167
  );


  buf
  g998
  (
    n728,
    n268
  );


  not
  g999
  (
    n1329,
    n544
  );


  not
  g1000
  (
    n685,
    n597
  );


  not
  g1001
  (
    n1174,
    n479
  );


  not
  g1002
  (
    n1142,
    n632
  );


  buf
  g1003
  (
    n1133,
    n170
  );


  buf
  g1004
  (
    n1682,
    n189
  );


  not
  g1005
  (
    n1551,
    n556
  );


  not
  g1006
  (
    n1545,
    n370
  );


  buf
  g1007
  (
    n1346,
    n637
  );


  not
  g1008
  (
    n1562,
    n494
  );


  not
  g1009
  (
    n1113,
    n637
  );


  not
  g1010
  (
    n1183,
    n355
  );


  not
  g1011
  (
    n1278,
    n381
  );


  buf
  g1012
  (
    n1669,
    n273
  );


  buf
  g1013
  (
    n798,
    n388
  );


  buf
  g1014
  (
    n1411,
    n561
  );


  not
  g1015
  (
    n1281,
    n365
  );


  buf
  g1016
  (
    n1579,
    n350
  );


  not
  g1017
  (
    n1024,
    n416
  );


  not
  g1018
  (
    n1426,
    n614
  );


  not
  g1019
  (
    n1407,
    n653
  );


  not
  g1020
  (
    n1159,
    n554
  );


  buf
  g1021
  (
    n860,
    n197
  );


  not
  g1022
  (
    n1169,
    n390
  );


  not
  g1023
  (
    n1393,
    n391
  );


  not
  g1024
  (
    n1537,
    n381
  );


  buf
  g1025
  (
    n769,
    n647
  );


  not
  g1026
  (
    n1324,
    n270
  );


  buf
  g1027
  (
    n1136,
    n552
  );


  not
  g1028
  (
    n750,
    n359
  );


  not
  g1029
  (
    n1361,
    n581
  );


  buf
  g1030
  (
    n1115,
    n164
  );


  buf
  g1031
  (
    n808,
    n473
  );


  not
  g1032
  (
    n833,
    n474
  );


  not
  g1033
  (
    n1131,
    n448
  );


  buf
  g1034
  (
    n816,
    n420
  );


  not
  g1035
  (
    n878,
    n254
  );


  buf
  g1036
  (
    n807,
    n433
  );


  not
  g1037
  (
    n1302,
    n369
  );


  not
  g1038
  (
    n1047,
    n623
  );


  buf
  g1039
  (
    n1050,
    n214
  );


  not
  g1040
  (
    n1070,
    n340
  );


  not
  g1041
  (
    n697,
    n351
  );


  not
  g1042
  (
    n1614,
    n423
  );


  buf
  g1043
  (
    n1129,
    n264
  );


  buf
  g1044
  (
    n1059,
    n295
  );


  buf
  g1045
  (
    n733,
    n203
  );


  not
  g1046
  (
    n1580,
    n382
  );


  not
  g1047
  (
    n1257,
    n275
  );


  not
  g1048
  (
    n1538,
    n647
  );


  buf
  g1049
  (
    n1653,
    n398
  );


  not
  g1050
  (
    n1355,
    n275
  );


  buf
  g1051
  (
    n715,
    n573
  );


  buf
  g1052
  (
    n791,
    n393
  );


  buf
  g1053
  (
    n1398,
    n607
  );


  buf
  g1054
  (
    n1581,
    n386
  );


  not
  g1055
  (
    n729,
    n560
  );


  not
  g1056
  (
    n707,
    n388
  );


  buf
  g1057
  (
    n1000,
    n426
  );


  buf
  g1058
  (
    n1185,
    n198
  );


  buf
  g1059
  (
    n937,
    n311
  );


  buf
  g1060
  (
    n1100,
    n247
  );


  buf
  g1061
  (
    n1356,
    n594
  );


  not
  g1062
  (
    n1528,
    n241
  );


  not
  g1063
  (
    n893,
    n282
  );


  not
  g1064
  (
    n1485,
    n302
  );


  not
  g1065
  (
    n1197,
    n611
  );


  buf
  g1066
  (
    n767,
    n377
  );


  buf
  g1067
  (
    n938,
    n654
  );


  not
  g1068
  (
    n1110,
    n599
  );


  buf
  g1069
  (
    n735,
    n404
  );


  not
  g1070
  (
    n1390,
    n580
  );


  buf
  g1071
  (
    n1573,
    n306
  );


  buf
  g1072
  (
    n1242,
    n402
  );


  not
  g1073
  (
    n941,
    n387
  );


  not
  g1074
  (
    n1299,
    n347
  );


  not
  g1075
  (
    n717,
    n499
  );


  buf
  g1076
  (
    n1446,
    n367
  );


  buf
  g1077
  (
    n829,
    n638
  );


  buf
  g1078
  (
    n1162,
    n359
  );


  not
  g1079
  (
    n1524,
    n168
  );


  not
  g1080
  (
    n1655,
    n671
  );


  buf
  g1081
  (
    n901,
    n438
  );


  buf
  g1082
  (
    n747,
    n314
  );


  buf
  g1083
  (
    n1207,
    n405
  );


  not
  g1084
  (
    n848,
    n443
  );


  not
  g1085
  (
    n1181,
    n209
  );


  not
  g1086
  (
    n879,
    n244
  );


  buf
  g1087
  (
    n1212,
    n615
  );


  buf
  g1088
  (
    n1026,
    n295
  );


  not
  g1089
  (
    n690,
    n564
  );


  not
  g1090
  (
    n968,
    n439
  );


  buf
  g1091
  (
    n1408,
    n508
  );


  not
  g1092
  (
    n1449,
    n552
  );


  buf
  g1093
  (
    n1414,
    n189
  );


  not
  g1094
  (
    n776,
    n636
  );


  buf
  g1095
  (
    n1217,
    n205
  );


  not
  g1096
  (
    n1486,
    n655
  );


  not
  g1097
  (
    n1045,
    n535
  );


  not
  g1098
  (
    n1253,
    n161
  );


  buf
  g1099
  (
    n1516,
    n638
  );


  buf
  g1100
  (
    n981,
    n308
  );


  buf
  g1101
  (
    n1560,
    n302
  );


  not
  g1102
  (
    n1167,
    n201
  );


  not
  g1103
  (
    n1227,
    n363
  );


  not
  g1104
  (
    n955,
    n276
  );


  buf
  g1105
  (
    n676,
    n298
  );


  not
  g1106
  (
    n1049,
    n550
  );


  buf
  g1107
  (
    n1287,
    n357
  );


  buf
  g1108
  (
    n689,
    n441
  );


  not
  g1109
  (
    n1402,
    n637
  );


  buf
  g1110
  (
    n705,
    n606
  );


  buf
  g1111
  (
    n1377,
    n662
  );


  not
  g1112
  (
    n1011,
    n257
  );


  not
  g1113
  (
    n731,
    n175
  );


  not
  g1114
  (
    n1673,
    n371
  );


  not
  g1115
  (
    n951,
    n495
  );


  not
  g1116
  (
    n813,
    n428
  );


  not
  g1117
  (
    n1001,
    n263
  );


  buf
  g1118
  (
    n1184,
    n295
  );


  not
  g1119
  (
    n1003,
    n199
  );


  not
  g1120
  (
    n1274,
    n425
  );


  buf
  g1121
  (
    n866,
    n488
  );


  not
  g1122
  (
    n990,
    n667
  );


  buf
  g1123
  (
    n774,
    n455
  );


  buf
  g1124
  (
    n1482,
    n238
  );


  not
  g1125
  (
    n1186,
    n287
  );


  buf
  g1126
  (
    n1622,
    n272
  );


  buf
  g1127
  (
    n845,
    n616
  );


  buf
  g1128
  (
    n762,
    n365
  );


  not
  g1129
  (
    n1022,
    n657
  );


  not
  g1130
  (
    n741,
    n410
  );


  not
  g1131
  (
    n1246,
    n169
  );


  not
  g1132
  (
    n1195,
    n488
  );


  not
  g1133
  (
    n1118,
    n587
  );


  not
  g1134
  (
    n880,
    n469
  );


  not
  g1135
  (
    n925,
    n234
  );


  buf
  g1136
  (
    n1107,
    n348
  );


  buf
  g1137
  (
    n1627,
    n535
  );


  not
  g1138
  (
    n1690,
    n319
  );


  buf
  g1139
  (
    n1569,
    n407
  );


  buf
  g1140
  (
    n926,
    n170
  );


  buf
  g1141
  (
    n1526,
    n229
  );


  not
  g1142
  (
    n881,
    n338
  );


  not
  g1143
  (
    n777,
    n587
  );


  not
  g1144
  (
    n1582,
    n322
  );


  buf
  g1145
  (
    n775,
    n502
  );


  not
  g1146
  (
    n989,
    n514
  );


  buf
  g1147
  (
    n1443,
    n599
  );


  not
  g1148
  (
    n852,
    n164
  );


  buf
  g1149
  (
    n1455,
    n239
  );


  buf
  g1150
  (
    n1168,
    n380
  );


  not
  g1151
  (
    n1660,
    n248
  );


  buf
  g1152
  (
    n1515,
    n366
  );


  not
  g1153
  (
    n1514,
    n168
  );


  buf
  g1154
  (
    n1464,
    n569
  );


  buf
  g1155
  (
    n1205,
    n626
  );


  not
  g1156
  (
    n1387,
    n431
  );


  not
  g1157
  (
    n1630,
    n300
  );


  buf
  g1158
  (
    n1155,
    n389
  );


  buf
  g1159
  (
    n1284,
    n266
  );


  not
  g1160
  (
    n1472,
    n427
  );


  buf
  g1161
  (
    n1376,
    n582
  );


  not
  g1162
  (
    n978,
    n600
  );


  not
  g1163
  (
    n1574,
    n450
  );


  not
  g1164
  (
    n895,
    n626
  );


  buf
  g1165
  (
    n1002,
    n413
  );


  buf
  g1166
  (
    n924,
    n292
  );


  buf
  g1167
  (
    n1178,
    n487
  );


  not
  g1168
  (
    n1564,
    n502
  );


  buf
  g1169
  (
    n1423,
    n536
  );


  not
  g1170
  (
    n1476,
    n595
  );


  buf
  g1171
  (
    n1638,
    n446
  );


  buf
  g1172
  (
    n1215,
    n571
  );


  not
  g1173
  (
    n1016,
    n256
  );


  not
  g1174
  (
    n1293,
    n424
  );


  buf
  g1175
  (
    n745,
    n471
  );


  buf
  g1176
  (
    n1591,
    n383
  );


  not
  g1177
  (
    n815,
    n464
  );


  not
  g1178
  (
    n1202,
    n623
  );


  not
  g1179
  (
    n942,
    n422
  );


  buf
  g1180
  (
    n1193,
    n511
  );


  buf
  g1181
  (
    n1401,
    n635
  );


  buf
  g1182
  (
    n964,
    n216
  );


  not
  g1183
  (
    n1453,
    n413
  );


  buf
  g1184
  (
    n788,
    n305
  );


  buf
  g1185
  (
    n1123,
    n166
  );


  buf
  g1186
  (
    n1436,
    n518
  );


  not
  g1187
  (
    n962,
    n379
  );


  buf
  g1188
  (
    n1478,
    n483
  );


  not
  g1189
  (
    n1040,
    n368
  );


  buf
  g1190
  (
    n1315,
    n551
  );


  not
  g1191
  (
    n743,
    n337
  );


  buf
  g1192
  (
    n1291,
    n172
  );


  buf
  g1193
  (
    n1372,
    n527
  );


  buf
  g1194
  (
    n1276,
    n225
  );


  buf
  g1195
  (
    n1511,
    n443
  );


  buf
  g1196
  (
    n746,
    n315
  );


  not
  g1197
  (
    n1238,
    n584
  );


  not
  g1198
  (
    n1633,
    n458
  );


  buf
  g1199
  (
    n1146,
    n339
  );


  not
  g1200
  (
    n1313,
    n218
  );


  buf
  g1201
  (
    n1432,
    n372
  );


  buf
  g1202
  (
    n1610,
    n475
  );


  buf
  g1203
  (
    n783,
    n249
  );


  not
  g1204
  (
    n1557,
    n183
  );


  buf
  g1205
  (
    n1068,
    n391
  );


  not
  g1206
  (
    n1081,
    n318
  );


  not
  g1207
  (
    n1288,
    n378
  );


  not
  g1208
  (
    n1675,
    n357
  );


  not
  g1209
  (
    n1091,
    n406
  );


  not
  g1210
  (
    n1006,
    n235
  );


  buf
  g1211
  (
    n1684,
    n290
  );


  buf
  g1212
  (
    n725,
    n527
  );


  buf
  g1213
  (
    n993,
    n309
  );


  not
  g1214
  (
    n1025,
    n415
  );


  not
  g1215
  (
    n724,
    n184
  );


  not
  g1216
  (
    n1265,
    n464
  );


  not
  g1217
  (
    n1342,
    n410
  );


  buf
  g1218
  (
    n948,
    n414
  );


  not
  g1219
  (
    n922,
    n299
  );


  not
  g1220
  (
    n1343,
    n456
  );


  buf
  g1221
  (
    n1273,
    n602
  );


  buf
  g1222
  (
    n681,
    n467
  );


  not
  g1223
  (
    n1127,
    n404
  );


  buf
  g1224
  (
    n786,
    n212
  );


  not
  g1225
  (
    n678,
    n547
  );


  buf
  g1226
  (
    n883,
    n211
  );


  not
  g1227
  (
    n830,
    n654
  );


  buf
  g1228
  (
    n1619,
    n353
  );


  not
  g1229
  (
    n1286,
    n391
  );


  buf
  g1230
  (
    n1662,
    n419
  );


  buf
  g1231
  (
    n929,
    n543
  );


  not
  g1232
  (
    n1541,
    n664
  );


  not
  g1233
  (
    n773,
    n227
  );


  not
  g1234
  (
    n900,
    n521
  );


  not
  g1235
  (
    n718,
    n204
  );


  not
  g1236
  (
    n1198,
    n326
  );


  buf
  g1237
  (
    n1416,
    n523
  );


  not
  g1238
  (
    n994,
    n248
  );


  buf
  g1239
  (
    n936,
    n496
  );


  buf
  g1240
  (
    n1465,
    n174
  );


  not
  g1241
  (
    n723,
    n525
  );


  not
  g1242
  (
    n1677,
    n609
  );


  buf
  g1243
  (
    n1663,
    n297
  );


  buf
  g1244
  (
    n1208,
    n318
  );


  not
  g1245
  (
    n1599,
    n662
  );


  not
  g1246
  (
    n686,
    n540
  );


  buf
  g1247
  (
    n749,
    n466
  );


  not
  g1248
  (
    n870,
    n517
  );


  not
  g1249
  (
    n1314,
    n319
  );


  not
  g1250
  (
    n1307,
    n220
  );


  not
  g1251
  (
    n1051,
    n219
  );


  not
  g1252
  (
    n748,
    n457
  );


  buf
  g1253
  (
    n1644,
    n361
  );


  not
  g1254
  (
    n886,
    n437
  );


  not
  g1255
  (
    n1424,
    n324
  );


  not
  g1256
  (
    n1121,
    n262
  );


  not
  g1257
  (
    n931,
    n485
  );


  not
  g1258
  (
    n930,
    n543
  );


  not
  g1259
  (
    n1404,
    n166
  );


  buf
  g1260
  (
    n1567,
    n343
  );


  not
  g1261
  (
    n1311,
    n305
  );


  not
  g1262
  (
    n751,
    n489
  );


  not
  g1263
  (
    n1452,
    n339
  );


  buf
  g1264
  (
    n1076,
    n329
  );


  not
  g1265
  (
    n1616,
    n662
  );


  not
  g1266
  (
    n1338,
    n611
  );


  buf
  g1267
  (
    n1536,
    n670
  );


  not
  g1268
  (
    n1642,
    n166
  );


  buf
  g1269
  (
    n1512,
    n182
  );


  not
  g1270
  (
    n1035,
    n226
  );


  buf
  g1271
  (
    n802,
    n587
  );


  buf
  g1272
  (
    n1532,
    n478
  );


  buf
  g1273
  (
    n1530,
    n505
  );


  buf
  g1274
  (
    n1437,
    n572
  );


  not
  g1275
  (
    n1015,
    n579
  );


  buf
  g1276
  (
    n789,
    n345
  );


  buf
  g1277
  (
    n1392,
    n246
  );


  buf
  g1278
  (
    n712,
    n283
  );


  not
  g1279
  (
    n1219,
    n540
  );


  not
  g1280
  (
    n1572,
    n208
  );


  not
  g1281
  (
    n793,
    n429
  );


  not
  g1282
  (
    n1457,
    n219
  );


  buf
  g1283
  (
    n1189,
    n438
  );


  not
  g1284
  (
    n698,
    n272
  );


  not
  g1285
  (
    n684,
    n245
  );


  buf
  g1286
  (
    n1032,
    n462
  );


  not
  g1287
  (
    n1041,
    n669
  );


  buf
  g1288
  (
    n1544,
    n648
  );


  buf
  g1289
  (
    n905,
    n354
  );


  not
  g1290
  (
    n1691,
    n231
  );


  not
  g1291
  (
    n673,
    n259
  );


  buf
  g1292
  (
    n889,
    n201
  );


  not
  g1293
  (
    n1125,
    n179
  );


  not
  g1294
  (
    n1368,
    n639
  );


  buf
  g1295
  (
    n1137,
    n189
  );


  buf
  g1296
  (
    n899,
    n228
  );


  not
  g1297
  (
    n911,
    n356
  );


  buf
  g1298
  (
    n1108,
    n658
  );


  buf
  g1299
  (
    n1106,
    n444
  );


  not
  g1300
  (
    n1676,
    n492
  );


  not
  g1301
  (
    n1012,
    n493
  );


  buf
  g1302
  (
    n1092,
    n286
  );


  buf
  g1303
  (
    n1054,
    n516
  );


  buf
  g1304
  (
    n1501,
    n522
  );


  not
  g1305
  (
    n1349,
    n527
  );


  not
  g1306
  (
    n1391,
    n288
  );


  buf
  g1307
  (
    n1234,
    n629
  );


  not
  g1308
  (
    n858,
    n500
  );


  not
  g1309
  (
    n956,
    n620
  );


  not
  g1310
  (
    n1323,
    n313
  );


  not
  g1311
  (
    n1645,
    n412
  );


  buf
  g1312
  (
    n1348,
    n581
  );


  not
  g1313
  (
    n706,
    n291
  );


  buf
  g1314
  (
    n1029,
    n381
  );


  not
  g1315
  (
    n1549,
    n194
  );


  not
  g1316
  (
    n847,
    n256
  );


  buf
  g1317
  (
    n755,
    n615
  );


  not
  g1318
  (
    n1369,
    n531
  );


  buf
  g1319
  (
    n1568,
    n389
  );


  and
  g1320
  (
    n742,
    n274,
    n627
  );


  and
  g1321
  (
    n797,
    n218,
    n411,
    n352,
    n178
  );


  xor
  g1322
  (
    n861,
    n546,
    n205,
    n187,
    n279
  );


  or
  g1323
  (
    n1177,
    n325,
    n413,
    n387,
    n658
  );


  or
  g1324
  (
    n1421,
    n236,
    n333,
    n506,
    n417
  );


  and
  g1325
  (
    n823,
    n424,
    n161,
    n196,
    n233
  );


  xnor
  g1326
  (
    n1153,
    n652,
    n378,
    n213,
    n563
  );


  xor
  g1327
  (
    n1308,
    n622,
    n395,
    n562,
    n481
  );


  xor
  g1328
  (
    n1621,
    n189,
    n483,
    n609,
    n263
  );


  xor
  g1329
  (
    n1463,
    n313,
    n265,
    n628,
    n201
  );


  and
  g1330
  (
    n1379,
    n356,
    n283,
    n652,
    n640
  );


  nand
  g1331
  (
    n1097,
    n508,
    n291,
    n281,
    n671
  );


  xor
  g1332
  (
    n1088,
    n418,
    n253,
    n629,
    n307
  );


  xnor
  g1333
  (
    n855,
    n630,
    n309,
    n596,
    n276
  );


  xnor
  g1334
  (
    n872,
    n173,
    n464,
    n557,
    n336
  );


  xnor
  g1335
  (
    n969,
    n544,
    n372,
    n222,
    n192
  );


  nand
  g1336
  (
    n1033,
    n482,
    n421,
    n353,
    n444
  );


  nor
  g1337
  (
    n1008,
    n575,
    n226,
    n206,
    n364
  );


  xor
  g1338
  (
    n859,
    n162,
    n299,
    n267,
    n428
  );


  or
  g1339
  (
    n1553,
    n624,
    n548,
    n386,
    n448
  );


  xnor
  g1340
  (
    n1039,
    n433,
    n412,
    n429,
    n533
  );


  nand
  g1341
  (
    n1061,
    n184,
    n330,
    n498,
    n470
  );


  and
  g1342
  (
    n679,
    n363,
    n233,
    n566,
    n273
  );


  or
  g1343
  (
    n757,
    n661,
    n517,
    n325,
    n468
  );


  and
  g1344
  (
    n1085,
    n237,
    n335,
    n664,
    n263
  );


  nor
  g1345
  (
    n1518,
    n285,
    n611,
    n271,
    n598
  );


  xor
  g1346
  (
    n1611,
    n192,
    n218,
    n302,
    n539
  );


  or
  g1347
  (
    n1428,
    n298,
    n449,
    n459,
    n198
  );


  xnor
  g1348
  (
    n1074,
    n659,
    n293,
    n207,
    n277
  );


  and
  g1349
  (
    n1182,
    n375,
    n563,
    n311,
    n656
  );


  nand
  g1350
  (
    n740,
    n236,
    n522,
    n588,
    n633
  );


  xor
  g1351
  (
    n1320,
    n279,
    n404,
    n342,
    n386
  );


  nand
  g1352
  (
    n1163,
    n536,
    n539,
    n635,
    n494
  );


  xnor
  g1353
  (
    n1353,
    n304,
    n635,
    n286,
    n559
  );


  xnor
  g1354
  (
    n693,
    n660,
    n311,
    n385,
    n225
  );


  or
  g1355
  (
    n846,
    n232,
    n227,
    n394,
    n223
  );


  nand
  g1356
  (
    n909,
    n167,
    n274,
    n214,
    n435
  );


  nand
  g1357
  (
    n1588,
    n408,
    n553,
    n395,
    n406
  );


  or
  g1358
  (
    n1247,
    n603,
    n270,
    n645,
    n644
  );


  nand
  g1359
  (
    n1508,
    n339,
    n444,
    n599,
    n261
  );


  xor
  g1360
  (
    n888,
    n630,
    n437,
    n278,
    n432
  );


  or
  g1361
  (
    n785,
    n566,
    n570,
    n473,
    n393
  );


  nand
  g1362
  (
    n1296,
    n641,
    n163,
    n251,
    n556
  );


  nor
  g1363
  (
    n1231,
    n642,
    n254,
    n331,
    n253
  );


  nor
  g1364
  (
    n760,
    n495,
    n215,
    n329,
    n538
  );


  nand
  g1365
  (
    n1339,
    n289,
    n659,
    n300,
    n587
  );


  nor
  g1366
  (
    n1140,
    n393,
    n593,
    n196,
    n305
  );


  nand
  g1367
  (
    n1629,
    n355,
    n537,
    n212,
    n472
  );


  or
  g1368
  (
    n1199,
    n660,
    n539,
    n528,
    n394
  );


  or
  g1369
  (
    n1654,
    n285,
    n670,
    n570,
    n370
  );


  xnor
  g1370
  (
    n1053,
    n262,
    n396,
    n575,
    n334
  );


  xor
  g1371
  (
    n1067,
    n508,
    n206,
    n241,
    n612
  );


  nand
  g1372
  (
    n1285,
    n375,
    n324,
    n171,
    n377
  );


  xnor
  g1373
  (
    n1664,
    n337,
    n469,
    n441,
    n584
  );


  nor
  g1374
  (
    n1023,
    n235,
    n473,
    n595,
    n352
  );


  and
  g1375
  (
    n1445,
    n612,
    n297,
    n165,
    n313
  );


  and
  g1376
  (
    n1206,
    n491,
    n494,
    n373,
    n442
  );


  xor
  g1377
  (
    n1419,
    n191,
    n563,
    n461,
    n176
  );


  xnor
  g1378
  (
    n1593,
    n424,
    n641,
    n454,
    n271
  );


  xnor
  g1379
  (
    n1672,
    n594,
    n367,
    n385,
    n322
  );


  xor
  g1380
  (
    n1469,
    n600,
    n627,
    n586,
    n239
  );


  nor
  g1381
  (
    n1321,
    n479,
    n330,
    n593,
    n237
  );


  xor
  g1382
  (
    n1534,
    n642,
    n307,
    n200,
    n446
  );


  nor
  g1383
  (
    n915,
    n405,
    n480,
    n320,
    n220
  );


  xnor
  g1384
  (
    n1636,
    n579,
    n177,
    n235,
    n383
  );


  nand
  g1385
  (
    n1565,
    n516,
    n376,
    n553,
    n667
  );


  xnor
  g1386
  (
    n947,
    n274,
    n646,
    n554,
    n529
  );


  and
  g1387
  (
    n1261,
    n413,
    n250,
    n242,
    n183
  );


  nand
  g1388
  (
    n957,
    n628,
    n462,
    n502,
    n450
  );


  xor
  g1389
  (
    n967,
    n493,
    n475,
    n227,
    n321
  );


  nor
  g1390
  (
    n1450,
    n311,
    n312,
    n665,
    n443
  );


  and
  g1391
  (
    n1300,
    n522,
    n230,
    n472,
    n369
  );


  nor
  g1392
  (
    n1451,
    n276,
    n573,
    n643,
    n653
  );


  xnor
  g1393
  (
    n1228,
    n176,
    n207,
    n331,
    n437
  );


  nor
  g1394
  (
    n1080,
    n379,
    n662,
    n625,
    n585
  );


  nand
  g1395
  (
    n1535,
    n449,
    n185,
    n346,
    n303
  );


  xor
  g1396
  (
    n1577,
    n561,
    n374,
    n289,
    n392
  );


  and
  g1397
  (
    n984,
    n509,
    n462,
    n544,
    n475
  );


  and
  g1398
  (
    n1255,
    n664,
    n365,
    n525,
    n571
  );


  xnor
  g1399
  (
    n695,
    n279,
    n426,
    n497,
    n544
  );


  nand
  g1400
  (
    n1134,
    n498,
    n382,
    n163,
    n255
  );


  nor
  g1401
  (
    n975,
    n324,
    n448,
    n208,
    n582
  );


  nor
  g1402
  (
    n1686,
    n398,
    n211,
    n468,
    n280
  );


  xnor
  g1403
  (
    n1667,
    n652,
    n303,
    n324,
    n550
  );


  nand
  g1404
  (
    n1196,
    n583,
    n390,
    n217,
    n483
  );


  nor
  g1405
  (
    n1375,
    n343,
    n532,
    n451,
    n430
  );


  xnor
  g1406
  (
    n997,
    n565,
    n593,
    n271,
    n333
  );


  nand
  g1407
  (
    n1226,
    n172,
    n542,
    n545,
    n485
  );


  xor
  g1408
  (
    n1470,
    n250,
    n590,
    n526,
    n251
  );


  nand
  g1409
  (
    n1641,
    n397,
    n466,
    n341,
    n193
  );


  nor
  g1410
  (
    n1506,
    n513,
    n515,
    n417,
    n387
  );


  or
  g1411
  (
    n1417,
    n461,
    n217,
    n446,
    n654
  );


  and
  g1412
  (
    n1158,
    n503,
    n321,
    n287,
    n579
  );


  xor
  g1413
  (
    n1632,
    n349,
    n171,
    n579,
    n240
  );


  nor
  g1414
  (
    n1150,
    n618,
    n656,
    n399,
    n259
  );


  xnor
  g1415
  (
    n1192,
    n332,
    n268,
    n636,
    n266
  );


  or
  g1416
  (
    n1410,
    n265,
    n478,
    n300,
    n347
  );


  xor
  g1417
  (
    n873,
    n601,
    n209,
    n452,
    n463
  );


  xor
  g1418
  (
    n1646,
    n610,
    n654,
    n511,
    n607
  );


  xor
  g1419
  (
    n863,
    n482,
    n162,
    n604,
    n625
  );


  xnor
  g1420
  (
    n1210,
    n494,
    n212,
    n338,
    n370
  );


  nand
  g1421
  (
    n1649,
    n591,
    n336,
    n620,
    n510
  );


  and
  g1422
  (
    n1256,
    n234,
    n216,
    n598,
    n375
  );


  xor
  g1423
  (
    n1149,
    n656,
    n249,
    n454,
    n503
  );


  and
  g1424
  (
    n1639,
    n241,
    n374,
    n407,
    n356
  );


  nand
  g1425
  (
    n1344,
    n285,
    n447,
    n346,
    n450
  );


  xnor
  g1426
  (
    n831,
    n465,
    n177,
    n519,
    n557
  );


  nor
  g1427
  (
    n832,
    n335,
    n430,
    n190,
    n551
  );


  nand
  g1428
  (
    n1317,
    n433,
    n423,
    n267,
    n188
  );


  nor
  g1429
  (
    n1038,
    n445,
    n275,
    n657,
    n251
  );


  and
  g1430
  (
    n839,
    n171,
    n266,
    n565,
    n457
  );


  nand
  g1431
  (
    n1109,
    n573,
    n368,
    n520,
    n639
  );


  or
  g1432
  (
    n801,
    n234,
    n382,
    n515,
    n294
  );


  or
  g1433
  (
    n1260,
    n420,
    n207,
    n341,
    n343
  );


  xor
  g1434
  (
    n1017,
    n390,
    n580,
    n583,
    n401
  );


  nand
  g1435
  (
    n1529,
    n420,
    n284,
    n466,
    n433
  );


  xor
  g1436
  (
    n756,
    n232,
    n607,
    n486,
    n588
  );


  xnor
  g1437
  (
    n1224,
    n335,
    n210,
    n369,
    n349
  );


  xor
  g1438
  (
    n1688,
    n595,
    n248,
    n247,
    n283
  );


  or
  g1439
  (
    n1351,
    n445,
    n456,
    n485,
    n574
  );


  xnor
  g1440
  (
    n1143,
    n357,
    n247,
    n341,
    n340
  );


  xor
  g1441
  (
    n1648,
    n349,
    n314,
    n323,
    n603
  );


  or
  g1442
  (
    n1280,
    n242,
    n476,
    n431,
    n663
  );


  nor
  g1443
  (
    n884,
    n327,
    n277,
    n524,
    n356
  );


  or
  g1444
  (
    n1020,
    n621,
    n569,
    n319,
    n608
  );


  nor
  g1445
  (
    n910,
    n434,
    n663,
    n612,
    n512
  );


  xnor
  g1446
  (
    n1661,
    n281,
    n485,
    n360,
    n636
  );


  xor
  g1447
  (
    n790,
    n641,
    n423,
    n436,
    n257
  );


  or
  g1448
  (
    n1533,
    n498,
    n322,
    n655,
    n500
  );


  xnor
  g1449
  (
    n1409,
    n237,
    n210,
    n213,
    n484
  );


  or
  g1450
  (
    n1095,
    n173,
    n347,
    n459,
    n548
  );


  xnor
  g1451
  (
    n1063,
    n604,
    n261,
    n235,
    n460
  );


  xor
  g1452
  (
    n1160,
    n328,
    n504,
    n665,
    n581
  );


  nand
  g1453
  (
    n1119,
    n410,
    n252,
    n262,
    n323
  );


  and
  g1454
  (
    n1084,
    n318,
    n627,
    n540,
    n350
  );


  xnor
  g1455
  (
    n836,
    n176,
    n379,
    n585,
    n240
  );


  and
  g1456
  (
    n1165,
    n608,
    n648,
    n611,
    n455
  );


  xor
  g1457
  (
    n976,
    n290,
    n535,
    n309,
    n269
  );


  nor
  g1458
  (
    n1370,
    n283,
    n642,
    n401,
    n287
  );


  nor
  g1459
  (
    n1122,
    n562,
    n614,
    n306,
    n564
  );


  xnor
  g1460
  (
    n963,
    n549,
    n195,
    n325,
    n596
  );


  xnor
  g1461
  (
    n986,
    n422,
    n451,
    n354,
    n480
  );


  nor
  g1462
  (
    n779,
    n396,
    n515,
    n441,
    n516
  );


  or
  g1463
  (
    n1493,
    n170,
    n572,
    n634,
    n501
  );


  nand
  g1464
  (
    n919,
    n417,
    n389,
    n198,
    n294
  );


  xor
  g1465
  (
    n1216,
    n617,
    n519,
    n453,
    n632
  );


  nor
  g1466
  (
    n1268,
    n480,
    n634,
    n439
  );


  nor
  g1467
  (
    n1489,
    n254,
    n173,
    n187,
    n648
  );


  and
  g1468
  (
    n772,
    n567,
    n301,
    n562,
    n299
  );


  or
  g1469
  (
    n1328,
    n353,
    n269,
    n268,
    n303
  );


  and
  g1470
  (
    n1583,
    n293,
    n551,
    n216,
    n374
  );


  or
  g1471
  (
    n1229,
    n361,
    n414,
    n574,
    n644
  );


  or
  g1472
  (
    n1128,
    n444,
    n490,
    n195,
    n492
  );


  or
  g1473
  (
    n851,
    n351,
    n602,
    n632,
    n459
  );


  nor
  g1474
  (
    n1144,
    n180,
    n202,
    n418,
    n251
  );


  or
  g1475
  (
    n771,
    n597,
    n354,
    n270,
    n415
  );


  xnor
  g1476
  (
    n1503,
    n599,
    n233,
    n489,
    n415
  );


  nand
  g1477
  (
    n1225,
    n633,
    n565,
    n456,
    n454
  );


  xor
  g1478
  (
    n1681,
    n622,
    n548,
    n376,
    n445
  );


  xor
  g1479
  (
    n965,
    n194,
    n301,
    n312,
    n180
  );


  xnor
  g1480
  (
    n714,
    n546,
    n610,
    n577,
    n197
  );


  xnor
  g1481
  (
    n1559,
    n668,
    n664,
    n630,
    n594
  );


  nand
  g1482
  (
    n828,
    n360,
    n322,
    n198,
    n464
  );


  or
  g1483
  (
    n1525,
    n161,
    n373,
    n653,
    n491
  );


  and
  g1484
  (
    n780,
    n176,
    n613,
    n523,
    n282
  );


  nor
  g1485
  (
    n1222,
    n349,
    n213,
    n272,
    n488
  );


  or
  g1486
  (
    n1380,
    n358,
    n547,
    n613,
    n344
  );


  nor
  g1487
  (
    n1471,
    n512,
    n576,
    n547,
    n575
  );


  nor
  g1488
  (
    n891,
    n609,
    n499,
    n529,
    n537
  );


  and
  g1489
  (
    n946,
    n624,
    n625,
    n541,
    n571
  );


  xnor
  g1490
  (
    n1065,
    n291,
    n296,
    n447,
    n606
  );


  nand
  g1491
  (
    n952,
    n317,
    n553,
    n597,
    n388
  );


  nor
  g1492
  (
    n914,
    n354,
    n641,
    n368,
    n477
  );


  xor
  g1493
  (
    n885,
    n214,
    n304,
    n278,
    n651
  );


  and
  g1494
  (
    n1606,
    n269,
    n603,
    n649,
    n511
  );


  xor
  g1495
  (
    n1297,
    n530,
    n545,
    n192,
    n240
  );


  or
  g1496
  (
    n1258,
    n514,
    n224,
    n208,
    n358
  );


  xnor
  g1497
  (
    n1187,
    n183,
    n193,
    n392,
    n550
  );


  xor
  g1498
  (
    n1474,
    n391,
    n484,
    n334,
    n367
  );


  nor
  g1499
  (
    n1294,
    n586,
    n282,
    n455,
    n206
  );


  xor
  g1500
  (
    n1399,
    n474,
    n610,
    n576,
    n287
  );


  xor
  g1501
  (
    n778,
    n389,
    n229,
    n245,
    n204
  );


  xnor
  g1502
  (
    n1354,
    n434,
    n416,
    n245,
    n439
  );


  xnor
  g1503
  (
    n1057,
    n308,
    n558,
    n626,
    n630
  );


  and
  g1504
  (
    n1336,
    n365,
    n472,
    n489,
    n525
  );


  nor
  g1505
  (
    n1148,
    n410,
    n327,
    n199,
    n669
  );


  nor
  g1506
  (
    n1027,
    n412,
    n273,
    n529,
    n592
  );


  or
  g1507
  (
    n810,
    n214,
    n539,
    n471,
    n436
  );


  nand
  g1508
  (
    n1030,
    n506,
    n299,
    n187,
    n194
  );


  nand
  g1509
  (
    n1563,
    n570,
    n435,
    n308,
    n246
  );


  xnor
  g1510
  (
    n949,
    n320,
    n207,
    n658,
    n231
  );


  nor
  g1511
  (
    n1418,
    n307,
    n277,
    n427,
    n256
  );


  nand
  g1512
  (
    n721,
    n336,
    n234,
    n637,
    n280
  );


  nand
  g1513
  (
    n1608,
    n352,
    n532,
    n487,
    n622
  );


  or
  g1514
  (
    n1221,
    n576,
    n303,
    n358,
    n531
  );


  nand
  g1515
  (
    n803,
    n279,
    n291,
    n643,
    n260
  );


  xnor
  g1516
  (
    n1438,
    n168,
    n515,
    n650,
    n213
  );


  xnor
  g1517
  (
    n1603,
    n490,
    n264,
    n628,
    n325
  );


  nand
  g1518
  (
    n1094,
    n528,
    n474,
    n168,
    n181
  );


  xor
  g1519
  (
    n1254,
    n370,
    n363,
    n451,
    n278
  );


  xnor
  g1520
  (
    n1270,
    n253,
    n181,
    n543,
    n190
  );


  and
  g1521
  (
    n1360,
    n403,
    n669,
    n561,
    n422
  );


  or
  g1522
  (
    n1262,
    n351,
    n184,
    n362,
    n506
  );


  xor
  g1523
  (
    n1386,
    n342,
    n195,
    n661,
    n463
  );


  or
  g1524
  (
    n1104,
    n334,
    n437,
    n578,
    n331
  );


  nand
  g1525
  (
    n1665,
    n612,
    n655,
    n333,
    n243
  );


  or
  g1526
  (
    n954,
    n640,
    n329,
    n559,
    n194
  );


  nor
  g1527
  (
    n1064,
    n408,
    n645,
    n263,
    n273
  );


  nor
  g1528
  (
    n1201,
    n384,
    n217,
    n505,
    n314
  );


  nor
  g1529
  (
    n1156,
    n589,
    n552,
    n594,
    n542
  );


  or
  g1530
  (
    n1497,
    n616,
    n355,
    n646,
    n272
  );


  and
  g1531
  (
    n945,
    n239,
    n493,
    n614,
    n443
  );


  xnor
  g1532
  (
    n1214,
    n618,
    n533,
    n209
  );


  or
  g1533
  (
    n921,
    n258,
    n345,
    n591,
    n327
  );


  xor
  g1534
  (
    n1180,
    n169,
    n184,
    n285,
    n254
  );


  nor
  g1535
  (
    n1048,
    n310,
    n222,
    n169,
    n218
  );


  or
  g1536
  (
    n700,
    n226,
    n414,
    n407,
    n644
  );


  and
  g1537
  (
    n1425,
    n538,
    n360,
    n200
  );


  xnor
  g1538
  (
    n734,
    n472,
    n372,
    n623,
    n486
  );


  or
  g1539
  (
    n754,
    n428,
    n216,
    n477,
    n385
  );


  xnor
  g1540
  (
    n1687,
    n395,
    n341,
    n436,
    n509
  );


  nand
  g1541
  (
    n1093,
    n403,
    n255,
    n300,
    n210
  );


  xor
  g1542
  (
    n1347,
    n416,
    n634,
    n491,
    n523
  );


  xor
  g1543
  (
    n1643,
    n533,
    n536,
    n369,
    n167
  );


  xor
  g1544
  (
    n768,
    n262,
    n615,
    n442,
    n455
  );


  and
  g1545
  (
    n917,
    n197,
    n429,
    n617,
    n321
  );


  and
  g1546
  (
    n875,
    n638,
    n165,
    n328,
    n588
  );


  or
  g1547
  (
    n971,
    n465,
    n172,
    n639,
    n501
  );


  nand
  g1548
  (
    n1334,
    n401,
    n362,
    n556,
    n223
  );


  and
  g1549
  (
    n720,
    n256,
    n388,
    n447,
    n616
  );


  nor
  g1550
  (
    n1279,
    n596,
    n394,
    n364,
    n187
  );


  xor
  g1551
  (
    n1586,
    n417,
    n411,
    n315,
    n521
  );


  or
  g1552
  (
    n1433,
    n400,
    n380,
    n174,
    n390
  );


  xnor
  g1553
  (
    n894,
    n538,
    n538,
    n224,
    n496
  );


  nor
  g1554
  (
    n1575,
    n230,
    n238,
    n265,
    n512
  );


  or
  g1555
  (
    n850,
    n313,
    n419,
    n224,
    n290
  );


  nor
  g1556
  (
    n953,
    n655,
    n621,
    n259,
    n261
  );


  nand
  g1557
  (
    n1612,
    n426,
    n409,
    n458,
    n568
  );


  nand
  g1558
  (
    n960,
    n191,
    n554,
    n258,
    n228
  );


  xnor
  g1559
  (
    n1266,
    n362,
    n229,
    n530,
    n487
  );


  xor
  g1560
  (
    n1130,
    n644,
    n182,
    n522,
    n568
  );


  nand
  g1561
  (
    n1306,
    n310,
    n220,
    n381,
    n398
  );


  nor
  g1562
  (
    n1634,
    n577,
    n364,
    n447,
    n651
  );


  nand
  g1563
  (
    n944,
    n383,
    n185,
    n608,
    n534
  );


  xnor
  g1564
  (
    n1412,
    n296,
    n531,
    n668,
    n161
  );


  or
  g1565
  (
    n1590,
    n567,
    n167,
    n602,
    n392
  );


  xnor
  g1566
  (
    n1498,
    n596,
    n384,
    n520,
    n540
  );


  nor
  g1567
  (
    n1271,
    n626,
    n309,
    n423,
    n546
  );


  nand
  g1568
  (
    n1468,
    n526,
    n555,
    n660
  );


  nand
  g1569
  (
    n1325,
    n605,
    n557,
    n586,
    n536
  );


  nor
  g1570
  (
    n1087,
    n617,
    n408,
    n517,
    n337
  );


  xor
  g1571
  (
    n1628,
    n628,
    n532,
    n342,
    n290
  );


  xor
  g1572
  (
    n1504,
    n425,
    n278,
    n615,
    n651
  );


  xor
  g1573
  (
    n688,
    n568,
    n490,
    n270,
    n496
  );


  xnor
  g1574
  (
    n1505,
    n342,
    n469,
    n334,
    n606
  );


  or
  g1575
  (
    n1267,
    n201,
    n614,
    n284,
    n301
  );


  or
  g1576
  (
    n759,
    n288,
    n595,
    n344,
    n578
  );


  or
  g1577
  (
    n1241,
    n281,
    n166,
    n534,
    n297
  );


  xnor
  g1578
  (
    n1179,
    n657,
    n510,
    n382,
    n415
  );


  or
  g1579
  (
    n853,
    n320,
    n525,
    n380,
    n267
  );


  xor
  g1580
  (
    n804,
    n316,
    n601,
    n591,
    n222
  );


  or
  g1581
  (
    n1689,
    n228,
    n284,
    n190,
    n280
  );


  and
  g1582
  (
    n1513,
    n361,
    n163,
    n518,
    n326
  );


  or
  g1583
  (
    n825,
    n492,
    n188,
    n521,
    n286
  );


  nor
  g1584
  (
    n849,
    n645,
    n211,
    n238,
    n470
  );


  nand
  g1585
  (
    n1600,
    n209,
    n202,
    n284,
    n567
  );


  xor
  g1586
  (
    n1312,
    n473,
    n245,
    n204,
    n330
  );


  xor
  g1587
  (
    n1077,
    n513,
    n537,
    n489,
    n561
  );


  xnor
  g1588
  (
    n1668,
    n399,
    n609,
    n361,
    n663
  );


  nand
  g1589
  (
    n1232,
    n442,
    n477,
    n445,
    n406
  );


  or
  g1590
  (
    n711,
    n608,
    n405,
    n468,
    n524
  );


  xor
  g1591
  (
    n1079,
    n373,
    n225,
    n202,
    n534
  );


  and
  g1592
  (
    n1335,
    n376,
    n427,
    n179,
    n233
  );


  xnor
  g1593
  (
    n1458,
    n452,
    n516,
    n364,
    n378
  );


  nand
  g1594
  (
    n1640,
    n598,
    n317,
    n617,
    n458
  );


  nor
  g1595
  (
    n1490,
    n535,
    n616,
    n465,
    n501
  );


  and
  g1596
  (
    n1692,
    n457,
    n232,
    n432,
    n255
  );


  xor
  g1597
  (
    n1357,
    n604,
    n478,
    n241,
    n506
  );


  xor
  g1598
  (
    n761,
    n312,
    n564,
    n531,
    n362
  );


  and
  g1599
  (
    n1331,
    n292,
    n219,
    n495,
    n186
  );


  nor
  g1600
  (
    n999,
    n560,
    n440,
    n294,
    n418
  );


  nor
  g1601
  (
    n1243,
    n547,
    n453,
    n440,
    n619
  );


  nand
  g1602
  (
    n950,
    n294,
    n468,
    n583,
    n624
  );


  nand
  g1603
  (
    n1019,
    n321,
    n250,
    n558,
    n429
  );


  nor
  g1604
  (
    n1609,
    n377,
    n523,
    n505,
    n567
  );


  xor
  g1605
  (
    n877,
    n239,
    n642,
    n289,
    n346
  );


  xor
  g1606
  (
    n1086,
    n221,
    n199,
    n405,
    n409
  );


  nand
  g1607
  (
    n1072,
    n202,
    n224,
    n386,
    n520
  );


  xnor
  g1608
  (
    n918,
    n471,
    n320,
    n215,
    n293
  );


  nand
  g1609
  (
    n792,
    n543,
    n221,
    n306,
    n527
  );


  or
  g1610
  (
    n857,
    n573,
    n259,
    n432,
    n479
  );


  xnor
  g1611
  (
    n1657,
    n297,
    n379,
    n380,
    n318
  );


  nor
  g1612
  (
    n1062,
    n428,
    n180,
    n560,
    n638
  );


  xor
  g1613
  (
    n1203,
    n419,
    n499,
    n248,
    n601
  );


  nor
  g1614
  (
    n1461,
    n400,
    n670,
    n244,
    n558
  );


  nor
  g1615
  (
    n1141,
    n230,
    n649,
    n420,
    n571
  );


  or
  g1616
  (
    n1188,
    n338,
    n229,
    n509,
    n293
  );


  and
  g1617
  (
    n1236,
    n243,
    n366,
    n394,
    n669
  );


  and
  g1618
  (
    n1345,
    n474,
    n395,
    n411,
    n371
  );


  or
  g1619
  (
    n763,
    n288,
    n619,
    n427
  );


  xnor
  g1620
  (
    n1373,
    n546,
    n331,
    n572,
    n467
  );


  and
  g1621
  (
    n1058,
    n173,
    n174,
    n238,
    n348
  );


  nand
  g1622
  (
    n1685,
    n659,
    n421,
    n353,
    n606
  );


  and
  g1623
  (
    n1103,
    n460,
    n440,
    n329,
    n518
  );


  or
  g1624
  (
    n1018,
    n408,
    n424,
    n438,
    n572
  );


  xnor
  g1625
  (
    n1083,
    n181,
    n668,
    n514,
    n500
  );


  and
  g1626
  (
    n1298,
    n649,
    n269,
    n590,
    n550
  );


  nor
  g1627
  (
    n1502,
    n648,
    n215,
    n350,
    n532
  );


  or
  g1628
  (
    n1066,
    n661,
    n371,
    n344,
    n426
  );


  nand
  g1629
  (
    n818,
    n352,
    n260,
    n203,
    n236
  );


  or
  g1630
  (
    n817,
    n257,
    n180,
    n591,
    n347
  );


  nand
  g1631
  (
    n1659,
    n605,
    n165,
    n195,
    n575
  );


  and
  g1632
  (
    n874,
    n191,
    n217,
    n657,
    n542
  );


  xnor
  g1633
  (
    n867,
    n666,
    n583,
    n481,
    n373
  );


  nand
  g1634
  (
    n1385,
    n190,
    n647,
    n453,
    n305
  );


  nor
  g1635
  (
    n1384,
    n646,
    n588,
    n651,
    n584
  );


  nand
  g1636
  (
    n1459,
    n162,
    n436,
    n585,
    n497
  );


  xor
  g1637
  (
    n766,
    n440,
    n371,
    n557,
    n530
  );


  nor
  g1638
  (
    n1570,
    n164,
    n328,
    n302,
    n542
  );


  xor
  g1639
  (
    n1495,
    n482,
    n384,
    n319,
    n622
  );


  nand
  g1640
  (
    n680,
    n215,
    n457,
    n179,
    n602
  );


  nor
  g1641
  (
    n1585,
    n403,
    n607,
    n392,
    n524
  );


  xor
  g1642
  (
    n935,
    n507,
    n576,
    n620,
    n541
  );


  xnor
  g1643
  (
    n1462,
    n570,
    n623,
    n564,
    n618
  );


  nor
  g1644
  (
    n1631,
    n670,
    n495,
    n597,
    n497
  );


  nand
  g1645
  (
    n985,
    n363,
    n400,
    n185,
    n569
  );


  xnor
  g1646
  (
    n1175,
    n310,
    n449,
    n459,
    n193
  );


  xnor
  g1647
  (
    n692,
    n643,
    n537,
    n578,
    n223
  );


  nand
  g1648
  (
    n710,
    n586,
    n416,
    n549,
    n432
  );


  xnor
  g1649
  (
    n1295,
    n458,
    n666,
    n624,
    n414
  );


  nor
  g1650
  (
    n1571,
    n507,
    n631,
    n520,
    n378
  );


  and
  g1651
  (
    n827,
    n312,
    n454,
    n268,
    n529
  );


  nor
  g1652
  (
    n784,
    n589,
    n345,
    n605,
    n545
  );


  xnor
  g1653
  (
    n814,
    n304,
    n501,
    n656,
    n237
  );


  nor
  g1654
  (
    n812,
    n430,
    n260,
    n360,
    n265
  );


  xor
  g1655
  (
    n1071,
    n409,
    n267,
    n503,
    n344
  );


  or
  g1656
  (
    n1473,
    n510,
    n348,
    n461,
    n621
  );


  or
  g1657
  (
    n787,
    n186,
    n452,
    n647,
    n338
  );


  xnor
  g1658
  (
    n970,
    n526,
    n377,
    n399,
    n244
  );


  xnor
  g1659
  (
    n1637,
    n314,
    n629,
    n663,
    n317
  );


  or
  g1660
  (
    n902,
    n476,
    n484,
    n503,
    n221
  );


  not
  g1661
  (
    n1713,
    n694
  );


  buf
  g1662
  (
    n1709,
    n674
  );


  not
  g1663
  (
    n1714,
    n698
  );


  buf
  g1664
  (
    n1694,
    n682
  );


  not
  g1665
  (
    n1705,
    n688
  );


  buf
  g1666
  (
    n1707,
    n693
  );


  buf
  g1667
  (
    n1696,
    n683
  );


  not
  g1668
  (
    n1712,
    n697
  );


  not
  g1669
  (
    n1703,
    n692
  );


  buf
  g1670
  (
    n1695,
    n695
  );


  buf
  g1671
  (
    n1704,
    n680
  );


  buf
  g1672
  (
    n1699,
    n678
  );


  not
  g1673
  (
    n1702,
    n689
  );


  buf
  g1674
  (
    n1711,
    n691
  );


  buf
  g1675
  (
    n1701,
    n686
  );


  not
  g1676
  (
    n1708,
    n687
  );


  or
  g1677
  (
    n1698,
    n699,
    n676
  );


  or
  g1678
  (
    n1710,
    n673,
    n690
  );


  nor
  g1679
  (
    n1700,
    n684,
    n685
  );


  nand
  g1680
  (
    n1697,
    n681,
    n677
  );


  nor
  g1681
  (
    n1715,
    n679,
    n700
  );


  nor
  g1682
  (
    n1706,
    n696,
    n675
  );


  not
  g1683
  (
    n1736,
    n721
  );


  not
  g1684
  (
    n1721,
    n1710
  );


  not
  g1685
  (
    n1716,
    n703
  );


  buf
  g1686
  (
    n1728,
    n725
  );


  buf
  g1687
  (
    n1730,
    n1713
  );


  buf
  g1688
  (
    n1723,
    n726
  );


  not
  g1689
  (
    n1732,
    n710
  );


  not
  g1690
  (
    n1718,
    n730
  );


  and
  g1691
  (
    n1717,
    n1705,
    n1715,
    n1708,
    n708
  );


  nand
  g1692
  (
    n1719,
    n1700,
    n711,
    n722,
    n738
  );


  and
  g1693
  (
    n1737,
    n1714,
    n1712,
    n735,
    n740
  );


  nand
  g1694
  (
    n1727,
    n1697,
    n709,
    n1707,
    n712
  );


  xnor
  g1695
  (
    n1720,
    n1698,
    n736,
    n1695,
    n705
  );


  xnor
  g1696
  (
    n1731,
    n1694,
    n723,
    n1704,
    n718
  );


  xor
  g1697
  (
    n1726,
    n1696,
    n1706,
    n720,
    n739
  );


  nand
  g1698
  (
    n1725,
    n715,
    n701,
    n1711,
    n1709
  );


  xnor
  g1699
  (
    n1729,
    n713,
    n732,
    n729,
    n741
  );


  nor
  g1700
  (
    n1734,
    n704,
    n702,
    n1703,
    n714
  );


  nand
  g1701
  (
    n1735,
    n728,
    n1701,
    n719,
    n706
  );


  nor
  g1702
  (
    n1733,
    n727,
    n742,
    n717,
    n734
  );


  xor
  g1703
  (
    n1724,
    n731,
    n716,
    n1702,
    n724
  );


  xnor
  g1704
  (
    n1722,
    n707,
    n1699,
    n737,
    n733
  );


  not
  g1705
  (
    n1739,
    n1717
  );


  buf
  g1706
  (
    n1741,
    n1716
  );


  not
  g1707
  (
    n1750,
    n1719
  );


  buf
  g1708
  (
    n1746,
    n1716
  );


  not
  g1709
  (
    n1748,
    n1719
  );


  not
  g1710
  (
    n1740,
    n1716
  );


  buf
  g1711
  (
    n1751,
    n1717
  );


  not
  g1712
  (
    n1744,
    n1720
  );


  buf
  g1713
  (
    n1738,
    n1717
  );


  buf
  g1714
  (
    n1755,
    n1717
  );


  buf
  g1715
  (
    n1749,
    n1718
  );


  not
  g1716
  (
    n1745,
    n1718
  );


  buf
  g1717
  (
    n1754,
    n1720
  );


  not
  g1718
  (
    n1742,
    n1718
  );


  buf
  g1719
  (
    n1743,
    n1716
  );


  buf
  g1720
  (
    n1753,
    n1719
  );


  not
  g1721
  (
    n1752,
    n1719
  );


  not
  g1722
  (
    n1747,
    n1718
  );


  buf
  g1723
  (
    n1765,
    n1741
  );


  not
  g1724
  (
    n1770,
    n746
  );


  buf
  g1725
  (
    n1760,
    n1743
  );


  not
  g1726
  (
    n1777,
    n763
  );


  not
  g1727
  (
    n1761,
    n1738
  );


  not
  g1728
  (
    n1758,
    n776
  );


  and
  g1729
  (
    n1776,
    n765,
    n1722,
    n1742
  );


  nand
  g1730
  (
    n1757,
    n1740,
    n1739,
    n1738,
    n1741
  );


  xor
  g1731
  (
    n1759,
    n743,
    n774,
    n758,
    n748
  );


  xor
  g1732
  (
    n1774,
    n761,
    n772,
    n1738,
    n1720
  );


  nand
  g1733
  (
    n1773,
    n771,
    n766,
    n745,
    n754
  );


  nor
  g1734
  (
    n1771,
    n768,
    n1723,
    n1721,
    n1740
  );


  xnor
  g1735
  (
    n1769,
    n1742,
    n1743,
    n767,
    n1738
  );


  nand
  g1736
  (
    n1763,
    n753,
    n751,
    n1741,
    n1723
  );


  xnor
  g1737
  (
    n1778,
    n1721,
    n752,
    n1740,
    n1739
  );


  or
  g1738
  (
    n1766,
    n1722,
    n1724,
    n775,
    n749
  );


  nand
  g1739
  (
    n1756,
    n1741,
    n759,
    n747,
    n762
  );


  and
  g1740
  (
    n1772,
    n1721,
    n770,
    n1720,
    n756
  );


  xnor
  g1741
  (
    n1775,
    n764,
    n1742,
    n1721,
    n1723
  );


  xor
  g1742
  (
    n1764,
    n744,
    n755,
    n757,
    n1739
  );


  and
  g1743
  (
    n1768,
    n1723,
    n750,
    n1722,
    n760
  );


  xnor
  g1744
  (
    n1762,
    n1739,
    n1740,
    n1724,
    n777
  );


  and
  g1745
  (
    n1767,
    n1742,
    n769,
    n773,
    n1743
  );


  buf
  g1746
  (
    n1824,
    n1726
  );


  buf
  g1747
  (
    n1840,
    n1770
  );


  not
  g1748
  (
    n1810,
    n1757
  );


  buf
  g1749
  (
    n1818,
    n1773
  );


  buf
  g1750
  (
    n1821,
    n1761
  );


  not
  g1751
  (
    n1839,
    n1762
  );


  not
  g1752
  (
    n1861,
    n1724
  );


  buf
  g1753
  (
    n1827,
    n1733
  );


  buf
  g1754
  (
    n1864,
    n672
  );


  buf
  g1755
  (
    n1831,
    n1772
  );


  not
  g1756
  (
    n1852,
    n1774
  );


  buf
  g1757
  (
    n1847,
    n672
  );


  not
  g1758
  (
    n1826,
    n1753
  );


  not
  g1759
  (
    n1799,
    n1771
  );


  not
  g1760
  (
    n1843,
    n1729
  );


  not
  g1761
  (
    n1855,
    n1756
  );


  not
  g1762
  (
    n1851,
    n1730
  );


  not
  g1763
  (
    n1785,
    n1748
  );


  not
  g1764
  (
    n1804,
    n1772
  );


  not
  g1765
  (
    n1813,
    n1766
  );


  not
  g1766
  (
    n1850,
    n1763
  );


  buf
  g1767
  (
    n1808,
    n785
  );


  buf
  g1768
  (
    n1869,
    n1767
  );


  buf
  g1769
  (
    n1781,
    n1746
  );


  not
  g1770
  (
    n1825,
    n1775
  );


  buf
  g1771
  (
    n1844,
    n1771
  );


  not
  g1772
  (
    n1860,
    n1764
  );


  buf
  g1773
  (
    n1867,
    n1730
  );


  not
  g1774
  (
    n1858,
    n1727
  );


  not
  g1775
  (
    n1868,
    n1762
  );


  buf
  g1776
  (
    n1823,
    n1744
  );


  buf
  g1777
  (
    n1788,
    n1730
  );


  buf
  g1778
  (
    n1820,
    n780
  );


  not
  g1779
  (
    n1801,
    n1760
  );


  buf
  g1780
  (
    n1782,
    n1767
  );


  buf
  g1781
  (
    n1833,
    n1727
  );


  buf
  g1782
  (
    n1836,
    n1749
  );


  buf
  g1783
  (
    n1791,
    n1744
  );


  buf
  g1784
  (
    n1816,
    n1774
  );


  not
  g1785
  (
    n1790,
    n1776
  );


  buf
  g1786
  (
    n1779,
    n1765
  );


  not
  g1787
  (
    n1805,
    n1758
  );


  not
  g1788
  (
    n1800,
    n783
  );


  buf
  g1789
  (
    n1854,
    n1733
  );


  buf
  g1790
  (
    n1786,
    n1750
  );


  buf
  g1791
  (
    n1784,
    n1727
  );


  not
  g1792
  (
    n1837,
    n1759
  );


  not
  g1793
  (
    n1856,
    n1769
  );


  not
  g1794
  (
    n1783,
    n1754
  );


  not
  g1795
  (
    n1819,
    n1745
  );


  not
  g1796
  (
    n1841,
    n1775
  );


  not
  g1797
  (
    n1806,
    n1765
  );


  buf
  g1798
  (
    n1817,
    n1752
  );


  buf
  g1799
  (
    n1842,
    n1763
  );


  not
  g1800
  (
    n1787,
    n1767
  );


  not
  g1801
  (
    n1870,
    n1752
  );


  buf
  g1802
  (
    n1809,
    n1769
  );


  buf
  g1803
  (
    n1792,
    n1766
  );


  not
  g1804
  (
    n1848,
    n1751
  );


  buf
  g1805
  (
    n1853,
    n1726
  );


  or
  g1806
  (
    n1803,
    n1776,
    n1769,
    n1753
  );


  or
  g1807
  (
    n1812,
    n1774,
    n1732,
    n672,
    n1729
  );


  nor
  g1808
  (
    n1846,
    n1727,
    n1725,
    n1770,
    n1728
  );


  and
  g1809
  (
    n1815,
    n1765,
    n1731,
    n1776
  );


  xor
  g1810
  (
    n1795,
    n1751,
    n1778,
    n1769,
    n1759
  );


  or
  g1811
  (
    n1794,
    n778,
    n1768,
    n782,
    n1749
  );


  nor
  g1812
  (
    n1862,
    n1764,
    n1753,
    n1766,
    n1750
  );


  xnor
  g1813
  (
    n1845,
    n671,
    n1725,
    n1759,
    n1767
  );


  or
  g1814
  (
    n1789,
    n1757,
    n671,
    n1772,
    n786
  );


  xor
  g1815
  (
    n1798,
    n1777,
    n779,
    n672,
    n784
  );


  and
  g1816
  (
    n1807,
    n1745,
    n1760,
    n1748,
    n1768
  );


  and
  g1817
  (
    n1780,
    n1746,
    n1777,
    n1749,
    n787
  );


  xnor
  g1818
  (
    n1859,
    n1761,
    n1744,
    n1759,
    n1752
  );


  nand
  g1819
  (
    n1797,
    n1732,
    n1756,
    n1748,
    n1757
  );


  nand
  g1820
  (
    n1857,
    n1748,
    n1777,
    n1771,
    n1760
  );


  xor
  g1821
  (
    n1834,
    n1761,
    n1751,
    n1747,
    n1770
  );


  and
  g1822
  (
    n1802,
    n1744,
    n1758,
    n1762,
    n1753
  );


  and
  g1823
  (
    n1796,
    n1757,
    n1725,
    n1729,
    n1772
  );


  xor
  g1824
  (
    n1793,
    n1751,
    n1768,
    n1745,
    n1731
  );


  xnor
  g1825
  (
    n1866,
    n1758,
    n1746,
    n1774,
    n1766
  );


  xor
  g1826
  (
    n1830,
    n1726,
    n1771,
    n1729,
    n1730
  );


  nand
  g1827
  (
    n1814,
    n1773,
    n1756,
    n1728,
    n1777
  );


  xor
  g1828
  (
    n1832,
    n1764,
    n1732,
    n1758,
    n781
  );


  xor
  g1829
  (
    n1829,
    n1760,
    n1765,
    n1726,
    n1749
  );


  or
  g1830
  (
    n1811,
    n1778,
    n1761,
    n1731,
    n1768
  );


  xor
  g1831
  (
    n1828,
    n1775,
    n1747,
    n1773,
    n1728
  );


  or
  g1832
  (
    n1863,
    n1775,
    n1776,
    n1747,
    n1773
  );


  or
  g1833
  (
    n1838,
    n1764,
    n1733,
    n1762,
    n1752
  );


  xor
  g1834
  (
    n1865,
    n1770,
    n1763,
    n1750
  );


  or
  g1835
  (
    n1835,
    n1745,
    n1725,
    n1724,
    n1756
  );


  and
  g1836
  (
    n1849,
    n1747,
    n1743,
    n1728,
    n1746
  );


  nand
  g1837
  (
    n1822,
    n1778,
    n1778,
    n1750,
    n1732
  );


  and
  g1838
  (
    n2112,
    n838,
    n1001,
    n1530,
    n1267
  );


  and
  g1839
  (
    n2097,
    n1804,
    n1838,
    n1552,
    n932
  );


  nand
  g1840
  (
    n1935,
    n1206,
    n810,
    n1484,
    n1850
  );


  or
  g1841
  (
    n1988,
    n1553,
    n1814,
    n1328,
    n1072
  );


  or
  g1842
  (
    n1987,
    n941,
    n1807,
    n1582,
    n1504
  );


  xor
  g1843
  (
    n1938,
    n1411,
    n1816,
    n1089,
    n1021
  );


  nand
  g1844
  (
    n2223,
    n867,
    n1841,
    n1852,
    n1073
  );


  xnor
  g1845
  (
    n1882,
    n892,
    n1854,
    n1188,
    n855
  );


  nand
  g1846
  (
    n2233,
    n1289,
    n1168,
    n1843,
    n1550
  );


  xnor
  g1847
  (
    n1931,
    n1347,
    n1503,
    n1789,
    n1568
  );


  xnor
  g1848
  (
    n2080,
    n1505,
    n1846,
    n1085,
    n1115
  );


  xnor
  g1849
  (
    n2207,
    n984,
    n1499,
    n1383,
    n1086
  );


  xor
  g1850
  (
    n2237,
    n1562,
    n881,
    n1533,
    n1836
  );


  xor
  g1851
  (
    n2222,
    n1503,
    n1851,
    n1343,
    n1076
  );


  and
  g1852
  (
    n2060,
    n1233,
    n1795,
    n1507,
    n1514
  );


  xnor
  g1853
  (
    n2004,
    n1578,
    n1532,
    n1531,
    n896
  );


  or
  g1854
  (
    n1894,
    n1101,
    n1208,
    n1544,
    n1003
  );


  nor
  g1855
  (
    n1930,
    n1791,
    n1811,
    n1575,
    n1521
  );


  and
  g1856
  (
    n2106,
    n1858,
    n1528,
    n1275,
    n1274
  );


  xor
  g1857
  (
    n2216,
    n1813,
    n1568,
    n1494,
    n1565
  );


  and
  g1858
  (
    n2122,
    n1415,
    n1509,
    n1390,
    n1398
  );


  nor
  g1859
  (
    n2092,
    n1506,
    n1377,
    n1358,
    n1134
  );


  nor
  g1860
  (
    n1985,
    n1801,
    n1791,
    n1488,
    n1822
  );


  nor
  g1861
  (
    n2232,
    n1577,
    n1843,
    n1791,
    n1408
  );


  nand
  g1862
  (
    n2126,
    n1498,
    n1321,
    n1435,
    n1005
  );


  and
  g1863
  (
    n2057,
    n989,
    n1380,
    n1477,
    n1563
  );


  and
  g1864
  (
    n1989,
    n1554,
    n1501,
    n1490,
    n933
  );


  nor
  g1865
  (
    n2046,
    n1230,
    n1551,
    n1848,
    n1829
  );


  or
  g1866
  (
    n2010,
    n1393,
    n1024,
    n1309,
    n1784
  );


  nor
  g1867
  (
    n2059,
    n1792,
    n1186,
    n1229,
    n1580
  );


  and
  g1868
  (
    n1909,
    n1818,
    n1163,
    n1786,
    n1084
  );


  or
  g1869
  (
    n2017,
    n829,
    n1433,
    n1786,
    n1048
  );


  nand
  g1870
  (
    n1918,
    n953,
    n1570,
    n1442,
    n1536
  );


  or
  g1871
  (
    n1976,
    n791,
    n1258,
    n1199,
    n1057
  );


  xnor
  g1872
  (
    n1887,
    n899,
    n1870,
    n1805,
    n1098
  );


  nand
  g1873
  (
    n2054,
    n1251,
    n1535,
    n1547,
    n1810
  );


  nor
  g1874
  (
    n1967,
    n1823,
    n1491,
    n1847,
    n1296
  );


  xnor
  g1875
  (
    n2152,
    n1491,
    n1834,
    n903,
    n1837
  );


  and
  g1876
  (
    n2063,
    n1530,
    n1825,
    n1504,
    n936
  );


  and
  g1877
  (
    n2028,
    n1512,
    n1805,
    n1410,
    n1558
  );


  nor
  g1878
  (
    n1945,
    n1853,
    n1849,
    n1254,
    n1356
  );


  xnor
  g1879
  (
    n2016,
    n1864,
    n1523,
    n821,
    n1449
  );


  nand
  g1880
  (
    n2191,
    n1424,
    n1417,
    n1302,
    n1856
  );


  and
  g1881
  (
    n1982,
    n1409,
    n923,
    n1569,
    n1531
  );


  nor
  g1882
  (
    n2081,
    n1534,
    n1518,
    n1510,
    n1840
  );


  or
  g1883
  (
    n1914,
    n1448,
    n1558,
    n1496,
    n1528
  );


  nand
  g1884
  (
    n1903,
    n1497,
    n859,
    n1787,
    n1493
  );


  nor
  g1885
  (
    n1875,
    n1486,
    n1845,
    n1344,
    n1827
  );


  and
  g1886
  (
    n2133,
    n1524,
    n1470,
    n973,
    n1789
  );


  xnor
  g1887
  (
    n2026,
    n1174,
    n1848,
    n1121,
    n1780
  );


  and
  g1888
  (
    n2173,
    n1158,
    n1521,
    n865,
    n1815
  );


  or
  g1889
  (
    n2039,
    n1118,
    n1821,
    n1378,
    n1571
  );


  xor
  g1890
  (
    n1934,
    n1837,
    n1007,
    n904,
    n1492
  );


  xnor
  g1891
  (
    n1933,
    n1431,
    n1800,
    n866,
    n1831
  );


  or
  g1892
  (
    n2023,
    n1536,
    n1529,
    n1368,
    n1833
  );


  xnor
  g1893
  (
    n1980,
    n1787,
    n1544,
    n1371,
    n1191
  );


  xor
  g1894
  (
    n2238,
    n958,
    n1169,
    n1288,
    n1815
  );


  or
  g1895
  (
    n2182,
    n1574,
    n1861,
    n1799,
    n1227
  );


  xnor
  g1896
  (
    n2022,
    n1846,
    n1543,
    n1555,
    n1303
  );


  nor
  g1897
  (
    n2181,
    n1567,
    n843,
    n956,
    n1561
  );


  nand
  g1898
  (
    n2119,
    n1402,
    n1506,
    n1489,
    n1479
  );


  xor
  g1899
  (
    n2035,
    n841,
    n1498,
    n1542,
    n1562
  );


  and
  g1900
  (
    n2163,
    n1058,
    n1526,
    n1137,
    n1162
  );


  and
  g1901
  (
    n2069,
    n1515,
    n1451,
    n789,
    n1803
  );


  xnor
  g1902
  (
    n2211,
    n979,
    n1459,
    n1160,
    n1326
  );


  nor
  g1903
  (
    n2091,
    n795,
    n988,
    n1485,
    n980
  );


  xnor
  g1904
  (
    n1881,
    n1783,
    n1855,
    n1096,
    n1210
  );


  and
  g1905
  (
    n2187,
    n1833,
    n1310,
    n1348,
    n1499
  );


  xnor
  g1906
  (
    n2066,
    n1099,
    n1552,
    n1109,
    n1520
  );


  or
  g1907
  (
    n2032,
    n1418,
    n1495,
    n1531,
    n1808
  );


  xor
  g1908
  (
    n1908,
    n1242,
    n1868,
    n1232,
    n1523
  );


  and
  g1909
  (
    n2186,
    n1486,
    n1521,
    n868,
    n1011
  );


  or
  g1910
  (
    n2072,
    n1157,
    n1107,
    n1038,
    n1250
  );


  nor
  g1911
  (
    n2014,
    n1811,
    n1804,
    n1009,
    n1809
  );


  or
  g1912
  (
    n2030,
    n1853,
    n1807,
    n1481,
    n1815
  );


  xnor
  g1913
  (
    n1893,
    n1520,
    n1090,
    n1859,
    n1171
  );


  and
  g1914
  (
    n1962,
    n1581,
    n1847,
    n1858,
    n1827
  );


  xnor
  g1915
  (
    n1970,
    n835,
    n946,
    n1503,
    n1216
  );


  xor
  g1916
  (
    n1951,
    n1282,
    n1814,
    n1530,
    n1117
  );


  and
  g1917
  (
    n2145,
    n848,
    n1824,
    n1806,
    n871
  );


  nor
  g1918
  (
    n1927,
    n1554,
    n1848,
    n1558,
    n802
  );


  or
  g1919
  (
    n2228,
    n1285,
    n1796,
    n1133,
    n1533
  );


  xnor
  g1920
  (
    n1975,
    n1823,
    n1565,
    n1394,
    n1782
  );


  xnor
  g1921
  (
    n2204,
    n1537,
    n793,
    n1033,
    n974
  );


  nor
  g1922
  (
    n1889,
    n1862,
    n1802,
    n1549,
    n965
  );


  nor
  g1923
  (
    n1956,
    n827,
    n1395,
    n1054,
    n1487
  );


  xnor
  g1924
  (
    n2224,
    n1083,
    n1575,
    n1502,
    n836
  );


  and
  g1925
  (
    n1977,
    n1419,
    n824,
    n1838,
    n1797
  );


  nand
  g1926
  (
    n1900,
    n1113,
    n1851,
    n889,
    n1287
  );


  nor
  g1927
  (
    n2158,
    n1545,
    n1359,
    n1023,
    n792
  );


  nand
  g1928
  (
    n2079,
    n1403,
    n1064,
    n1124,
    n1032
  );


  or
  g1929
  (
    n2220,
    n1488,
    n1278,
    n1573,
    n1512
  );


  xor
  g1930
  (
    n2073,
    n1824,
    n1580,
    n1859,
    n977
  );


  xnor
  g1931
  (
    n2093,
    n1535,
    n1841,
    n837,
    n1443
  );


  nand
  g1932
  (
    n1963,
    n994,
    n1836,
    n1172
  );


  nand
  g1933
  (
    n2180,
    n885,
    n1517,
    n1780,
    n1379
  );


  xor
  g1934
  (
    n2213,
    n798,
    n1543,
    n1807,
    n1147
  );


  xnor
  g1935
  (
    n1965,
    n1813,
    n1316,
    n1051,
    n1497
  );


  or
  g1936
  (
    n2104,
    n1518,
    n897,
    n931,
    n952
  );


  or
  g1937
  (
    n2212,
    n1492,
    n1006,
    n1519,
    n858
  );


  xnor
  g1938
  (
    n1922,
    n1177,
    n1856,
    n993,
    n1854
  );


  or
  g1939
  (
    n2088,
    n876,
    n1798,
    n982,
    n1401
  );


  xnor
  g1940
  (
    n2047,
    n1346,
    n1796,
    n1566,
    n1543
  );


  nor
  g1941
  (
    n2229,
    n1837,
    n1867,
    n1387,
    n1535
  );


  xnor
  g1942
  (
    n2040,
    n1537,
    n1789,
    n1792,
    n1036
  );


  or
  g1943
  (
    n1901,
    n959,
    n1266,
    n1563,
    n1835
  );


  xor
  g1944
  (
    n2219,
    n1845,
    n1821,
    n1222,
    n1523
  );


  or
  g1945
  (
    n1878,
    n1412,
    n1780,
    n1175,
    n1844
  );


  nor
  g1946
  (
    n2114,
    n887,
    n1010,
    n1803,
    n1399
  );


  xor
  g1947
  (
    n2235,
    n1508,
    n1528,
    n1483,
    n1166
  );


  nand
  g1948
  (
    n2147,
    n1820,
    n1322,
    n1828,
    n1785
  );


  and
  g1949
  (
    n2227,
    n910,
    n1865,
    n1122,
    n794
  );


  xor
  g1950
  (
    n2000,
    n1272,
    n1865,
    n1313,
    n1179
  );


  nor
  g1951
  (
    n2195,
    n1780,
    n1557,
    n1217,
    n1146
  );


  xor
  g1952
  (
    n1883,
    n1853,
    n1165,
    n804,
    n1796
  );


  nor
  g1953
  (
    n1904,
    n1350,
    n1542,
    n1025,
    n1514
  );


  nand
  g1954
  (
    n2027,
    n1159,
    n1464,
    n1803,
    n1560
  );


  or
  g1955
  (
    n2018,
    n1560,
    n926,
    n1838,
    n1794
  );


  nor
  g1956
  (
    n2169,
    n1816,
    n1552,
    n981,
    n1441
  );


  nor
  g1957
  (
    n2124,
    n1375,
    n884,
    n1830,
    n1487
  );


  xnor
  g1958
  (
    n2143,
    n1511,
    n1819,
    n1204,
    n1182
  );


  nand
  g1959
  (
    n2174,
    n1856,
    n1252,
    n1534,
    n1556
  );


  nor
  g1960
  (
    n2151,
    n1542,
    n834,
    n1226,
    n1480
  );


  xor
  g1961
  (
    n2061,
    n1213,
    n1583,
    n1816,
    n970
  );


  nand
  g1962
  (
    n1899,
    n1529,
    n1804,
    n1860,
    n1506
  );


  xor
  g1963
  (
    n2146,
    n1231,
    n1514,
    n1013,
    n949
  );


  or
  g1964
  (
    n1876,
    n1335,
    n1547,
    n1820,
    n1839
  );


  or
  g1965
  (
    n2005,
    n1511,
    n1573,
    n1480,
    n1488
  );


  and
  g1966
  (
    n2154,
    n1325,
    n1869,
    n1525,
    n1787
  );


  nand
  g1967
  (
    n2123,
    n1192,
    n1161,
    n1126,
    n1571
  );


  xor
  g1968
  (
    n2076,
    n1805,
    n1019,
    n1131,
    n1342
  );


  xnor
  g1969
  (
    n2012,
    n1784,
    n1547,
    n944,
    n1546
  );


  nand
  g1970
  (
    n2214,
    n1564,
    n1237,
    n1494,
    n1793
  );


  xnor
  g1971
  (
    n1950,
    n1142,
    n1212,
    n1564,
    n1849
  );


  and
  g1972
  (
    n1926,
    n1841,
    n1510,
    n1817,
    n1565
  );


  or
  g1973
  (
    n2085,
    n924,
    n1822,
    n895,
    n800
  );


  nand
  g1974
  (
    n2140,
    n1830,
    n1262,
    n1513,
    n831
  );


  and
  g1975
  (
    n1952,
    n1014,
    n1869,
    n1203,
    n1835
  );


  xnor
  g1976
  (
    n2206,
    n1576,
    n1050,
    n1857,
    n1863
  );


  xnor
  g1977
  (
    n1979,
    n872,
    n1119,
    n1140,
    n1824
  );


  nand
  g1978
  (
    n2194,
    n1311,
    n1517,
    n1538,
    n1572
  );


  and
  g1979
  (
    n2234,
    n1555,
    n1516,
    n1340,
    n1509
  );


  or
  g1980
  (
    n1954,
    n1522,
    n1503,
    n1385,
    n939
  );


  xnor
  g1981
  (
    n2115,
    n1813,
    n1284,
    n1811,
    n1077
  );


  or
  g1982
  (
    n1913,
    n1246,
    n1129,
    n1800,
    n1215
  );


  xor
  g1983
  (
    n2208,
    n1314,
    n1345,
    n846,
    n1079
  );


  nor
  g1984
  (
    n2162,
    n1432,
    n805,
    n912,
    n893
  );


  nand
  g1985
  (
    n2013,
    n1568,
    n1526,
    n975,
    n1461
  );


  or
  g1986
  (
    n2230,
    n925,
    n1540,
    n890,
    n1502
  );


  xnor
  g1987
  (
    n1949,
    n1423,
    n1053,
    n1496,
    n1855
  );


  and
  g1988
  (
    n2002,
    n1308,
    n1063,
    n1788,
    n1490
  );


  nor
  g1989
  (
    n1948,
    n1810,
    n920,
    n1806,
    n1553
  );


  nand
  g1990
  (
    n2177,
    n1545,
    n1211,
    n1357,
    n1505
  );


  or
  g1991
  (
    n1923,
    n1483,
    n1148,
    n1365,
    n1793
  );


  and
  g1992
  (
    n2164,
    n1529,
    n1551,
    n1082,
    n935
  );


  nor
  g1993
  (
    n2120,
    n1798,
    n1847,
    n1537,
    n1787
  );


  xor
  g1994
  (
    n1873,
    n1551,
    n1840,
    n1544,
    n1286
  );


  xor
  g1995
  (
    n2007,
    n1505,
    n916,
    n1518,
    n797
  );


  nand
  g1996
  (
    n1897,
    n1548,
    n1537,
    n1535,
    n1504
  );


  and
  g1997
  (
    n2130,
    n1806,
    n1790,
    n1180,
    n1527
  );


  xnor
  g1998
  (
    n2189,
    n1482,
    n1225,
    n1151,
    n1139
  );


  nor
  g1999
  (
    n2041,
    n1088,
    n1834,
    n796,
    n1829
  );


  or
  g2000
  (
    n2065,
    n1257,
    n1141,
    n1506,
    n1436
  );


  nor
  g2001
  (
    n2170,
    n1547,
    n1797,
    n1505,
    n1533
  );


  xnor
  g2002
  (
    n1983,
    n898,
    n1297,
    n1261,
    n1801
  );


  and
  g2003
  (
    n2201,
    n1843,
    n1827,
    n1559,
    n1854
  );


  and
  g2004
  (
    n1896,
    n1193,
    n1138,
    n1484,
    n1291
  );


  nor
  g2005
  (
    n2056,
    n819,
    n1809,
    n1015,
    n1145
  );


  nand
  g2006
  (
    n2183,
    n929,
    n880,
    n825,
    n1781
  );


  nor
  g2007
  (
    n2210,
    n1823,
    n987,
    n1507,
    n985
  );


  or
  g2008
  (
    n1929,
    n950,
    n1458,
    n1332,
    n1469
  );


  xnor
  g2009
  (
    n2121,
    n1582,
    n1406,
    n1801,
    n1494
  );


  or
  g2010
  (
    n2083,
    n1388,
    n1339,
    n1559,
    n1018
  );


  nand
  g2011
  (
    n2064,
    n1525,
    n814,
    n911,
    n1052
  );


  nor
  g2012
  (
    n2110,
    n1799,
    n940,
    n1574,
    n1369
  );


  or
  g2013
  (
    n2067,
    n850,
    n1798,
    n1307,
    n1854
  );


  xnor
  g2014
  (
    n2205,
    n1570,
    n1548,
    n1842,
    n1824
  );


  xnor
  g2015
  (
    n2129,
    n1067,
    n1154,
    n1858,
    n1807
  );


  and
  g2016
  (
    n2084,
    n1870,
    n1524,
    n967,
    n969
  );


  nor
  g2017
  (
    n2141,
    n1498,
    n1319,
    n863,
    n1864
  );


  nor
  g2018
  (
    n2175,
    n1794,
    n1489,
    n788,
    n1136
  );


  and
  g2019
  (
    n1978,
    n1802,
    n1153,
    n1831,
    n1569
  );


  or
  g2020
  (
    n1884,
    n1515,
    n1508,
    n955,
    n1334
  );


  nand
  g2021
  (
    n1968,
    n1539,
    n1555,
    n1849,
    n1571
  );


  nand
  g2022
  (
    n2196,
    n1114,
    n801,
    n1573,
    n1370
  );


  nand
  g2023
  (
    n1973,
    n1224,
    n1866,
    n1392,
    n1835
  );


  or
  g2024
  (
    n1888,
    n1508,
    n1527,
    n905,
    n1207
  );


  or
  g2025
  (
    n2165,
    n1463,
    n815,
    n1499,
    n1045
  );


  and
  g2026
  (
    n1961,
    n1366,
    n1198,
    n1579,
    n1475
  );


  and
  g2027
  (
    n1941,
    n1381,
    n1783,
    n1318,
    n1808
  );


  nor
  g2028
  (
    n1991,
    n1788,
    n1452,
    n1020,
    n1799
  );


  xor
  g2029
  (
    n1920,
    n1414,
    n1839,
    n1851,
    n1540
  );


  nand
  g2030
  (
    n2155,
    n1525,
    n1864,
    n1455,
    n938
  );


  xor
  g2031
  (
    n2082,
    n877,
    n1556,
    n1864,
    n883
  );


  nor
  g2032
  (
    n1906,
    n1189,
    n1812,
    n1447,
    n1457
  );


  or
  g2033
  (
    n2144,
    n1839,
    n1277,
    n1517,
    n1548
  );


  or
  g2034
  (
    n2149,
    n1299,
    n1490,
    n1810,
    n1819
  );


  or
  g2035
  (
    n2006,
    n1810,
    n1492,
    n906,
    n960
  );


  or
  g2036
  (
    n2209,
    n1080,
    n1812,
    n1476,
    n927
  );


  xnor
  g2037
  (
    n2025,
    n1523,
    n1298,
    n839,
    n1243
  );


  xor
  g2038
  (
    n2105,
    n806,
    n1304,
    n1330,
    n1108
  );


  and
  g2039
  (
    n1981,
    n1784,
    n1800,
    n1571,
    n1485
  );


  nand
  g2040
  (
    n2095,
    n1790,
    n1561,
    n1554,
    n1529
  );


  and
  g2041
  (
    n1890,
    n1513,
    n1835,
    n1248,
    n1220
  );


  xnor
  g2042
  (
    n2150,
    n1317,
    n1473,
    n1413,
    n828
  );


  and
  g2043
  (
    n2168,
    n1495,
    n997,
    n1558,
    n1800
  );


  nor
  g2044
  (
    n2179,
    n1034,
    n1793,
    n826,
    n922
  );


  nand
  g2045
  (
    n2078,
    n1214,
    n1576,
    n1532
  );


  or
  g2046
  (
    n2068,
    n1561,
    n1430,
    n1047,
    n918
  );


  nand
  g2047
  (
    n1944,
    n1543,
    n1312,
    n1305,
    n860
  );


  nor
  g2048
  (
    n2089,
    n1779,
    n1029,
    n1078,
    n1264
  );


  and
  g2049
  (
    n2117,
    n807,
    n1583,
    n851,
    n1819
  );


  or
  g2050
  (
    n2107,
    n1826,
    n1853,
    n1527,
    n1502
  );


  nand
  g2051
  (
    n2161,
    n1804,
    n1572,
    n1306,
    n1236
  );


  xnor
  g2052
  (
    n2070,
    n1533,
    n1555,
    n1861,
    n1509
  );


  and
  g2053
  (
    n2075,
    n1575,
    n1574,
    n1868,
    n1509
  );


  nor
  g2054
  (
    n2051,
    n1559,
    n1544,
    n1405,
    n934
  );


  nor
  g2055
  (
    n2188,
    n1828,
    n1794,
    n1783,
    n1815
  );


  or
  g2056
  (
    n2218,
    n1487,
    n1796,
    n1241,
    n1511
  );


  nand
  g2057
  (
    n1925,
    n1219,
    n832,
    n1367,
    n818
  );


  nand
  g2058
  (
    n1994,
    n1524,
    n1539,
    n1580,
    n1320
  );


  xor
  g2059
  (
    n2193,
    n1579,
    n1416,
    n1797,
    n1070
  );


  or
  g2060
  (
    n2131,
    n1831,
    n1238,
    n1566,
    n972
  );


  or
  g2061
  (
    n2074,
    n1818,
    n1839,
    n1071,
    n1106
  );


  xor
  g2062
  (
    n2157,
    n1549,
    n1836,
    n817,
    n1454
  );


  xor
  g2063
  (
    n2031,
    n1040,
    n1860,
    n930,
    n1427
  );


  and
  g2064
  (
    n2167,
    n1842,
    n961,
    n882,
    n874
  );


  or
  g2065
  (
    n1960,
    n1870,
    n803,
    n1338,
    n1852
  );


  nand
  g2066
  (
    n1940,
    n921,
    n1061,
    n1293,
    n1549
  );


  nand
  g2067
  (
    n2049,
    n1323,
    n888,
    n1536,
    n1112
  );


  and
  g2068
  (
    n2045,
    n919,
    n957,
    n845,
    n1862
  );


  nor
  g2069
  (
    n1932,
    n1567,
    n1860,
    n1373,
    n1362
  );


  nor
  g2070
  (
    n2148,
    n1046,
    n811,
    n1481,
    n1527
  );


  nand
  g2071
  (
    n1872,
    n1273,
    n1548,
    n1540,
    n1843
  );


  and
  g2072
  (
    n2003,
    n1551,
    n1028,
    n1259,
    n1069
  );


  or
  g2073
  (
    n1943,
    n1363,
    n1382,
    n1528,
    n854
  );


  nand
  g2074
  (
    n2036,
    n1516,
    n1026,
    n1781,
    n1577
  );


  nand
  g2075
  (
    n2055,
    n1143,
    n1562,
    n1235,
    n1164
  );


  nand
  g2076
  (
    n2021,
    n1865,
    n1845,
    n901,
    n1822
  );


  or
  g2077
  (
    n2020,
    n1499,
    n1779,
    n1315,
    n1867
  );


  nor
  g2078
  (
    n1937,
    n844,
    n1579,
    n1031,
    n833
  );


  and
  g2079
  (
    n2171,
    n1861,
    n1167,
    n1290,
    n1786
  );


  nor
  g2080
  (
    n2015,
    n1578,
    n1280,
    n1181,
    n1825
  );


  xor
  g2081
  (
    n2008,
    n1557,
    n1445,
    n1829
  );


  and
  g2082
  (
    n2153,
    n1197,
    n1438,
    n1542,
    n1858
  );


  xnor
  g2083
  (
    n2087,
    n1256,
    n1517,
    n1281,
    n1283
  );


  xor
  g2084
  (
    n1942,
    n1518,
    n1869,
    n1795,
    n1812
  );


  and
  g2085
  (
    n1898,
    n1522,
    n1176,
    n1782,
    n1268
  );


  xor
  g2086
  (
    n2011,
    n1850,
    n1827,
    n1553,
    n978
  );


  xnor
  g2087
  (
    n1924,
    n1486,
    n1105,
    n1271,
    n1825
  );


  and
  g2088
  (
    n1955,
    n1111,
    n1841,
    n1498,
    n1056
  );


  nor
  g2089
  (
    n2100,
    n1516,
    n1552,
    n999,
    n1574
  );


  or
  g2090
  (
    n2058,
    n954,
    n1104,
    n1265,
    n1239
  );


  or
  g2091
  (
    n2048,
    n1301,
    n1802,
    n1779,
    n1863
  );


  or
  g2092
  (
    n2019,
    n1194,
    n1255,
    n1200,
    n908
  );


  xnor
  g2093
  (
    n1995,
    n1324,
    n1128,
    n1855,
    n1538
  );


  and
  g2094
  (
    n1921,
    n1516,
    n820,
    n1566,
    n1546
  );


  nand
  g2095
  (
    n2138,
    n1530,
    n1127,
    n1333,
    n1495
  );


  nand
  g2096
  (
    n1895,
    n1572,
    n1850,
    n1428,
    n1466
  );


  and
  g2097
  (
    n1874,
    n1486,
    n1862,
    n1785,
    n1008
  );


  nor
  g2098
  (
    n2176,
    n1055,
    n1269,
    n1812,
    n1515
  );


  nand
  g2099
  (
    n2009,
    n1514,
    n875,
    n1043,
    n1789
  );


  xor
  g2100
  (
    n2086,
    n900,
    n1279,
    n948,
    n1862
  );


  and
  g2101
  (
    n1959,
    n1538,
    n1563,
    n1474,
    n1802
  );


  nor
  g2102
  (
    n2139,
    n1244,
    n964,
    n1481,
    n1489
  );


  nand
  g2103
  (
    n1915,
    n1512,
    n1779,
    n1068,
    n1818
  );


  xor
  g2104
  (
    n1902,
    n1521,
    n1524,
    n1857,
    n1818
  );


  and
  g2105
  (
    n1958,
    n1444,
    n1788,
    n873,
    n1292
  );


  nor
  g2106
  (
    n2043,
    n1825,
    n1569,
    n1355,
    n1472
  );


  xnor
  g2107
  (
    n2200,
    n1792,
    n1218,
    n894,
    n951
  );


  nand
  g2108
  (
    n2199,
    n1821,
    n1861,
    n1336,
    n1792
  );


  xnor
  g2109
  (
    n2001,
    n1832,
    n1270,
    n1513,
    n1196
  );


  nand
  g2110
  (
    n1916,
    n1519,
    n1581,
    n840,
    n1453
  );


  xor
  g2111
  (
    n1999,
    n1781,
    n1566,
    n861,
    n996
  );


  xor
  g2112
  (
    n2113,
    n1508,
    n1859,
    n991,
    n1519
  );


  xor
  g2113
  (
    n2052,
    n1173,
    n1062,
    n968,
    n1549
  );


  nand
  g2114
  (
    n1911,
    n847,
    n853,
    n1563,
    n1022
  );


  nor
  g2115
  (
    n1936,
    n1795,
    n1178,
    n1183,
    n990
  );


  xnor
  g2116
  (
    n2125,
    n1353,
    n1482,
    n1842,
    n1234
  );


  and
  g2117
  (
    n2142,
    n1867,
    n1545,
    n1569,
    n1095
  );


  xor
  g2118
  (
    n1997,
    n1809,
    n1844,
    n1481,
    n1471
  );


  xor
  g2119
  (
    n1946,
    n1500,
    n1581,
    n790,
    n1116
  );


  nor
  g2120
  (
    n2221,
    n1830,
    n1579,
    n1790,
    n1846
  );


  or
  g2121
  (
    n1990,
    n1352,
    n1500,
    n809,
    n1834
  );


  xnor
  g2122
  (
    n1969,
    n799,
    n1130,
    n1102,
    n902
  );


  and
  g2123
  (
    n2029,
    n1493,
    n1135,
    n1201,
    n1501
  );


  xor
  g2124
  (
    n1953,
    n928,
    n1110,
    n1833,
    n1828
  );


  xor
  g2125
  (
    n2077,
    n1814,
    n1221,
    n1826,
    n1017
  );


  nor
  g2126
  (
    n2202,
    n1391,
    n1863,
    n1832,
    n1866
  );


  xor
  g2127
  (
    n2098,
    n1100,
    n1785,
    n1404,
    n1223
  );


  nand
  g2128
  (
    n2156,
    n1300,
    n1426,
    n1042,
    n1550
  );


  nor
  g2129
  (
    n1966,
    n1846,
    n1337,
    n1519,
    n1568
  );


  or
  g2130
  (
    n1928,
    n1496,
    n852,
    n943,
    n1539
  );


  nand
  g2131
  (
    n1907,
    n1074,
    n1245,
    n891,
    n1247
  );


  nor
  g2132
  (
    n1871,
    n1550,
    n998,
    n1570,
    n1575
  );


  xor
  g2133
  (
    n2109,
    n1540,
    n1425,
    n1170,
    n1794
  );


  or
  g2134
  (
    n1996,
    n1799,
    n1578,
    n1819,
    n1567
  );


  xnor
  g2135
  (
    n1998,
    n1041,
    n1087,
    n1856,
    n1478
  );


  xnor
  g2136
  (
    n2135,
    n1541,
    n1495,
    n1798,
    n1833
  );


  and
  g2137
  (
    n1957,
    n1205,
    n1360,
    n1483,
    n1811
  );


  or
  g2138
  (
    n2116,
    n1538,
    n1791,
    n1823,
    n1507
  );


  or
  g2139
  (
    n2136,
    n1497,
    n1097,
    n1185,
    n1857
  );


  nand
  g2140
  (
    n2044,
    n1828,
    n1795,
    n1550,
    n1565
  );


  and
  g2141
  (
    n2024,
    n1832,
    n1276,
    n1240,
    n1190
  );


  nor
  g2142
  (
    n2197,
    n1361,
    n1817,
    n1782,
    n976
  );


  nor
  g2143
  (
    n1880,
    n813,
    n1572,
    n1081,
    n992
  );


  xnor
  g2144
  (
    n2101,
    n1840,
    n1493,
    n1497,
    n1253
  );


  nand
  g2145
  (
    n1974,
    n1460,
    n1867,
    n1783,
    n1030
  );


  nand
  g2146
  (
    n2160,
    n937,
    n915,
    n1000,
    n1793
  );


  nand
  g2147
  (
    n2128,
    n1816,
    n1092,
    n1567,
    n1557
  );


  xnor
  g2148
  (
    n2111,
    n1577,
    n1546,
    n1786,
    n1560
  );


  xor
  g2149
  (
    n1886,
    n1801,
    n1576,
    n1831,
    n1456
  );


  nor
  g2150
  (
    n2062,
    n1781,
    n1513,
    n1044,
    n857
  );


  xor
  g2151
  (
    n1917,
    n1863,
    n1806,
    n1532,
    n1860
  );


  xnor
  g2152
  (
    n2102,
    n1144,
    n1525,
    n1837,
    n1209
  );


  nand
  g2153
  (
    n2226,
    n1016,
    n1489,
    n1520,
    n1487
  );


  nor
  g2154
  (
    n2185,
    n1556,
    n945,
    n1838,
    n1500
  );


  nand
  g2155
  (
    n2127,
    n1094,
    n1582,
    n1397,
    n1826
  );


  nand
  g2156
  (
    n2042,
    n1329,
    n1429,
    n1035,
    n816
  );


  nand
  g2157
  (
    n2159,
    n1785,
    n947,
    n1866,
    n822
  );


  xnor
  g2158
  (
    n1877,
    n962,
    n1866,
    n1814,
    n1849
  );


  nor
  g2159
  (
    n2094,
    n1485,
    n862,
    n1422,
    n966
  );


  nand
  g2160
  (
    n1939,
    n1294,
    n1808,
    n1522,
    n1840
  );


  nor
  g2161
  (
    n1972,
    n1065,
    n1132,
    n1384,
    n849
  );


  nand
  g2162
  (
    n2172,
    n1844,
    n1364,
    n1485,
    n1446
  );


  nor
  g2163
  (
    n2192,
    n1012,
    n1556,
    n1491
  );


  xor
  g2164
  (
    n2236,
    n1554,
    n1331,
    n1820,
    n1511
  );


  or
  g2165
  (
    n1892,
    n1842,
    n1483,
    n1504,
    n1493
  );


  xor
  g2166
  (
    n1992,
    n1496,
    n1817,
    n1573,
    n1510
  );


  xnor
  g2167
  (
    n1885,
    n909,
    n1507,
    n878,
    n1826
  );


  nand
  g2168
  (
    n1912,
    n971,
    n864,
    n1421,
    n942
  );


  xor
  g2169
  (
    n1971,
    n1374,
    n1541,
    n1376,
    n1465
  );


  xor
  g2170
  (
    n1910,
    n1002,
    n842,
    n1851,
    n870
  );


  xor
  g2171
  (
    n1986,
    n808,
    n1848,
    n1855,
    n1195
  );


  or
  g2172
  (
    n2033,
    n1349,
    n1049,
    n1868,
    n1502
  );


  nor
  g2173
  (
    n2225,
    n913,
    n1437,
    n1484,
    n1372
  );


  xnor
  g2174
  (
    n2037,
    n1536,
    n1557,
    n917,
    n1492
  );


  nand
  g2175
  (
    n2118,
    n1564,
    n1578,
    n1450,
    n1560
  );


  xnor
  g2176
  (
    n1891,
    n1488,
    n1539,
    n1559,
    n1327
  );


  xnor
  g2177
  (
    n2108,
    n1059,
    n1484,
    n1400,
    n1249
  );


  xnor
  g2178
  (
    n2071,
    n1467,
    n983,
    n1821,
    n1870
  );


  and
  g2179
  (
    n2134,
    n1149,
    n1490,
    n1152,
    n1809
  );


  nand
  g2180
  (
    n2231,
    n1060,
    n1817,
    n1832,
    n914
  );


  or
  g2181
  (
    n2217,
    n1562,
    n1027,
    n1570,
    n1790
  );


  xor
  g2182
  (
    n1905,
    n1852,
    n1541,
    n986,
    n1534
  );


  xor
  g2183
  (
    n1879,
    n1420,
    n879,
    n1091,
    n1482
  );


  xor
  g2184
  (
    n2090,
    n1784,
    n1526,
    n1123,
    n1263
  );


  and
  g2185
  (
    n2198,
    n1782,
    n907,
    n1501,
    n1580
  );


  nand
  g2186
  (
    n2103,
    n1813,
    n1093,
    n1500,
    n823
  );


  nor
  g2187
  (
    n2178,
    n1075,
    n1260,
    n1039,
    n1845
  );


  nand
  g2188
  (
    n2132,
    n1847,
    n1541,
    n1859,
    n1351
  );


  xnor
  g2189
  (
    n2034,
    n1797,
    n1577,
    n1805,
    n1857
  );


  xnor
  g2190
  (
    n2215,
    n1576,
    n1407,
    n1295,
    n1534
  );


  and
  g2191
  (
    n2137,
    n1788,
    n1482,
    n1004,
    n1494
  );


  and
  g2192
  (
    n1993,
    n1389,
    n1440,
    n1515,
    n1865
  );


  or
  g2193
  (
    n2050,
    n1522,
    n1520,
    n963,
    n1803
  );


  or
  g2194
  (
    n2203,
    n1510,
    n886,
    n856,
    n1037
  );


  xor
  g2195
  (
    n2099,
    n1852,
    n1808,
    n1120,
    n1354
  );


  nand
  g2196
  (
    n1919,
    n1869,
    n1850,
    n1581,
    n1822
  );


  xnor
  g2197
  (
    n1964,
    n1103,
    n1582,
    n869,
    n1546
  );


  xor
  g2198
  (
    n2166,
    n1526,
    n1564,
    n1844,
    n1184
  );


  nor
  g2199
  (
    n2190,
    n1545,
    n1125,
    n1439,
    n1341
  );


  xor
  g2200
  (
    n1947,
    n1228,
    n1820,
    n1202,
    n1531
  );


  or
  g2201
  (
    n2184,
    n1561,
    n1834,
    n1512,
    n1155
  );


  nor
  g2202
  (
    n2053,
    n1462,
    n995,
    n1553,
    n1396
  );


  or
  g2203
  (
    n1984,
    n1830,
    n1468,
    n812,
    n1434
  );


  xnor
  g2204
  (
    n2096,
    n1150,
    n830,
    n1187,
    n1066
  );


  nor
  g2205
  (
    n2038,
    n1868,
    n1501,
    n1156,
    n1386
  );


  buf
  g2206
  (
    n2704,
    n1914
  );


  not
  g2207
  (
    n2349,
    n1603
  );


  buf
  g2208
  (
    n2461,
    n1934
  );


  not
  g2209
  (
    n2751,
    n1949
  );


  not
  g2210
  (
    n2666,
    n1997
  );


  buf
  g2211
  (
    n2576,
    n1940
  );


  not
  g2212
  (
    n2363,
    n1632
  );


  not
  g2213
  (
    n2332,
    n1992
  );


  buf
  g2214
  (
    n2846,
    n2010
  );


  not
  g2215
  (
    n2488,
    n1978
  );


  buf
  g2216
  (
    n2493,
    n1945
  );


  not
  g2217
  (
    n2469,
    n1597
  );


  not
  g2218
  (
    n2863,
    n1964
  );


  not
  g2219
  (
    n2570,
    n1933
  );


  buf
  g2220
  (
    n2723,
    n2025
  );


  buf
  g2221
  (
    n2647,
    n1969
  );


  not
  g2222
  (
    n2522,
    n1877
  );


  buf
  g2223
  (
    n2333,
    n1951
  );


  not
  g2224
  (
    n2478,
    n1919
  );


  not
  g2225
  (
    n2633,
    n1991
  );


  buf
  g2226
  (
    n2595,
    n1633
  );


  not
  g2227
  (
    n2599,
    n2012
  );


  not
  g2228
  (
    n2643,
    n1905
  );


  buf
  g2229
  (
    n2631,
    n1626
  );


  not
  g2230
  (
    n2555,
    n1635
  );


  not
  g2231
  (
    n2372,
    n1884
  );


  not
  g2232
  (
    n2362,
    n1976
  );


  not
  g2233
  (
    n2521,
    n1872
  );


  buf
  g2234
  (
    n2625,
    n1970
  );


  not
  g2235
  (
    n2515,
    n1938
  );


  not
  g2236
  (
    n2621,
    n1603
  );


  buf
  g2237
  (
    n2826,
    n2003
  );


  buf
  g2238
  (
    n2542,
    n2006
  );


  buf
  g2239
  (
    n2280,
    n1941
  );


  buf
  g2240
  (
    n2698,
    n1612
  );


  buf
  g2241
  (
    n2779,
    n1961
  );


  not
  g2242
  (
    n2414,
    n1618
  );


  not
  g2243
  (
    n2271,
    n2014
  );


  not
  g2244
  (
    n2302,
    n1604
  );


  not
  g2245
  (
    n2530,
    n1872
  );


  not
  g2246
  (
    n2244,
    n1605
  );


  buf
  g2247
  (
    n2771,
    n1949
  );


  not
  g2248
  (
    n2578,
    n1970
  );


  buf
  g2249
  (
    n2240,
    n1987
  );


  not
  g2250
  (
    n2465,
    n1959
  );


  not
  g2251
  (
    n2516,
    n1952
  );


  buf
  g2252
  (
    n2344,
    n1892
  );


  not
  g2253
  (
    n2401,
    n1876
  );


  buf
  g2254
  (
    n2588,
    n1995
  );


  buf
  g2255
  (
    n2550,
    n1918
  );


  buf
  g2256
  (
    n2374,
    n1881
  );


  not
  g2257
  (
    n2498,
    n1920
  );


  not
  g2258
  (
    n2736,
    n1969
  );


  buf
  g2259
  (
    n2691,
    n1928
  );


  buf
  g2260
  (
    n2822,
    n1613
  );


  buf
  g2261
  (
    n2426,
    n1973
  );


  buf
  g2262
  (
    n2632,
    n1878
  );


  buf
  g2263
  (
    n2580,
    n1634
  );


  not
  g2264
  (
    n2501,
    n1925
  );


  buf
  g2265
  (
    n2371,
    n1987
  );


  not
  g2266
  (
    n2430,
    n1635
  );


  not
  g2267
  (
    n2749,
    n1959
  );


  buf
  g2268
  (
    n2834,
    n2003
  );


  not
  g2269
  (
    n2513,
    n1909
  );


  not
  g2270
  (
    n2316,
    n1994
  );


  not
  g2271
  (
    n2671,
    n1956
  );


  buf
  g2272
  (
    n2268,
    n1923
  );


  not
  g2273
  (
    n2353,
    n2018
  );


  buf
  g2274
  (
    n2299,
    n1947
  );


  not
  g2275
  (
    n2340,
    n1612
  );


  buf
  g2276
  (
    n2446,
    n1955
  );


  buf
  g2277
  (
    n2709,
    n1904
  );


  buf
  g2278
  (
    n2778,
    n1879
  );


  buf
  g2279
  (
    n2350,
    n1880
  );


  not
  g2280
  (
    n2806,
    n2018
  );


  not
  g2281
  (
    n2597,
    n1915
  );


  buf
  g2282
  (
    n2334,
    n2014
  );


  not
  g2283
  (
    n2861,
    n2012
  );


  not
  g2284
  (
    n2460,
    n2013
  );


  buf
  g2285
  (
    n2559,
    n1604
  );


  buf
  g2286
  (
    n2812,
    n2015
  );


  not
  g2287
  (
    n2398,
    n1922
  );


  buf
  g2288
  (
    n2719,
    n1904
  );


  buf
  g2289
  (
    n2788,
    n1974
  );


  buf
  g2290
  (
    n2748,
    n1900
  );


  buf
  g2291
  (
    n2512,
    n1590
  );


  buf
  g2292
  (
    n2844,
    n1933
  );


  not
  g2293
  (
    n2352,
    n2000
  );


  buf
  g2294
  (
    n2718,
    n1606
  );


  not
  g2295
  (
    n2531,
    n1931
  );


  not
  g2296
  (
    n2304,
    n1964
  );


  buf
  g2297
  (
    n2517,
    n1610
  );


  buf
  g2298
  (
    n2435,
    n1938
  );


  buf
  g2299
  (
    n2775,
    n1871
  );


  not
  g2300
  (
    n2707,
    n2001
  );


  buf
  g2301
  (
    n2745,
    n1594
  );


  not
  g2302
  (
    n2840,
    n2024
  );


  not
  g2303
  (
    n2303,
    n1587
  );


  buf
  g2304
  (
    n2524,
    n1601
  );


  not
  g2305
  (
    n2477,
    n1584
  );


  buf
  g2306
  (
    n2641,
    n1979
  );


  not
  g2307
  (
    n2475,
    n1629
  );


  buf
  g2308
  (
    n2708,
    n1896
  );


  buf
  g2309
  (
    n2450,
    n1908
  );


  not
  g2310
  (
    n2319,
    n2026
  );


  not
  g2311
  (
    n2637,
    n1900
  );


  buf
  g2312
  (
    n2688,
    n1919
  );


  not
  g2313
  (
    n2623,
    n2019
  );


  buf
  g2314
  (
    n2440,
    n1615
  );


  not
  g2315
  (
    n2308,
    n1939
  );


  buf
  g2316
  (
    n2835,
    n1604
  );


  buf
  g2317
  (
    n2594,
    n1955
  );


  not
  g2318
  (
    n2791,
    n1998
  );


  not
  g2319
  (
    n2821,
    n1897
  );


  not
  g2320
  (
    n2467,
    n1629
  );


  buf
  g2321
  (
    n2654,
    n1910
  );


  not
  g2322
  (
    n2568,
    n1876
  );


  not
  g2323
  (
    n2830,
    n1916
  );


  not
  g2324
  (
    n2620,
    n1947
  );


  buf
  g2325
  (
    n2545,
    n1888
  );


  buf
  g2326
  (
    n2589,
    n1614
  );


  buf
  g2327
  (
    n2658,
    n1924
  );


  buf
  g2328
  (
    n2764,
    n2021
  );


  buf
  g2329
  (
    n2312,
    n1899
  );


  not
  g2330
  (
    n2548,
    n1969
  );


  buf
  g2331
  (
    n2758,
    n1895
  );


  buf
  g2332
  (
    n2697,
    n1975
  );


  buf
  g2333
  (
    n2701,
    n1988
  );


  not
  g2334
  (
    n2714,
    n1915
  );


  not
  g2335
  (
    n2805,
    n1630
  );


  not
  g2336
  (
    n2455,
    n1997
  );


  buf
  g2337
  (
    n2848,
    n1596
  );


  not
  g2338
  (
    n2479,
    n1929
  );


  not
  g2339
  (
    n2413,
    n1599
  );


  not
  g2340
  (
    n2661,
    n1922
  );


  not
  g2341
  (
    n2556,
    n1962
  );


  buf
  g2342
  (
    n2511,
    n1608
  );


  not
  g2343
  (
    n2611,
    n1921
  );


  buf
  g2344
  (
    n2560,
    n1963
  );


  buf
  g2345
  (
    n2575,
    n1929
  );


  buf
  g2346
  (
    n2800,
    n1983
  );


  buf
  g2347
  (
    n2505,
    n1585
  );


  buf
  g2348
  (
    n2403,
    n1618
  );


  not
  g2349
  (
    n2818,
    n1935
  );


  buf
  g2350
  (
    n2711,
    n1996
  );


  not
  g2351
  (
    n2810,
    n1997
  );


  buf
  g2352
  (
    n2616,
    n1948
  );


  not
  g2353
  (
    n2744,
    n1974
  );


  buf
  g2354
  (
    n2321,
    n1925
  );


  buf
  g2355
  (
    n2470,
    n1980
  );


  buf
  g2356
  (
    n2429,
    n1621
  );


  buf
  g2357
  (
    n2689,
    n1999
  );


  not
  g2358
  (
    n2640,
    n1991
  );


  not
  g2359
  (
    n2842,
    n1944
  );


  buf
  g2360
  (
    n2535,
    n1939
  );


  buf
  g2361
  (
    n2665,
    n1591
  );


  buf
  g2362
  (
    n2668,
    n1952
  );


  not
  g2363
  (
    n2253,
    n2005
  );


  not
  g2364
  (
    n2648,
    n1907
  );


  buf
  g2365
  (
    n2504,
    n1902
  );


  not
  g2366
  (
    n2390,
    n2015
  );


  not
  g2367
  (
    n2459,
    n1924
  );


  buf
  g2368
  (
    n2770,
    n1966
  );


  buf
  g2369
  (
    n2416,
    n1586
  );


  not
  g2370
  (
    n2552,
    n1890
  );


  buf
  g2371
  (
    n2410,
    n1893
  );


  not
  g2372
  (
    n2502,
    n1988
  );


  buf
  g2373
  (
    n2254,
    n2013
  );


  not
  g2374
  (
    n2445,
    n1996
  );


  not
  g2375
  (
    n2828,
    n1994
  );


  not
  g2376
  (
    n2617,
    n1601
  );


  buf
  g2377
  (
    n2281,
    n1990
  );


  not
  g2378
  (
    n2419,
    n1935
  );


  not
  g2379
  (
    n2603,
    n1638
  );


  not
  g2380
  (
    n2610,
    n1630
  );


  not
  g2381
  (
    n2600,
    n2016
  );


  not
  g2382
  (
    n2307,
    n1916
  );


  buf
  g2383
  (
    n2762,
    n1929
  );


  buf
  g2384
  (
    n2823,
    n1881
  );


  not
  g2385
  (
    n2629,
    n2000
  );


  buf
  g2386
  (
    n2262,
    n1965
  );


  buf
  g2387
  (
    n2694,
    n1956
  );


  buf
  g2388
  (
    n2767,
    n1910
  );


  not
  g2389
  (
    n2624,
    n2026
  );


  buf
  g2390
  (
    n2251,
    n1995
  );


  not
  g2391
  (
    n2797,
    n1949
  );


  buf
  g2392
  (
    n2782,
    n2008
  );


  not
  g2393
  (
    n2754,
    n1993
  );


  buf
  g2394
  (
    n2412,
    n1903
  );


  buf
  g2395
  (
    n2259,
    n1631
  );


  buf
  g2396
  (
    n2539,
    n1626
  );


  not
  g2397
  (
    n2305,
    n1950
  );


  buf
  g2398
  (
    n2664,
    n1618
  );


  buf
  g2399
  (
    n2265,
    n2007
  );


  buf
  g2400
  (
    n2546,
    n1624
  );


  buf
  g2401
  (
    n2678,
    n1624
  );


  not
  g2402
  (
    n2355,
    n1921
  );


  not
  g2403
  (
    n2759,
    n1971
  );


  not
  g2404
  (
    n2602,
    n1938
  );


  buf
  g2405
  (
    n2402,
    n1627
  );


  not
  g2406
  (
    n2366,
    n2014
  );


  buf
  g2407
  (
    n2761,
    n1925
  );


  buf
  g2408
  (
    n2456,
    n1968
  );


  buf
  g2409
  (
    n2618,
    n1609
  );


  buf
  g2410
  (
    n2804,
    n1882
  );


  not
  g2411
  (
    n2388,
    n1583
  );


  not
  g2412
  (
    n2464,
    n1993
  );


  buf
  g2413
  (
    n2337,
    n1898
  );


  not
  g2414
  (
    n2604,
    n1953
  );


  buf
  g2415
  (
    n2549,
    n1976
  );


  buf
  g2416
  (
    n2418,
    n1880
  );


  not
  g2417
  (
    n2293,
    n1975
  );


  not
  g2418
  (
    n2529,
    n1631
  );


  not
  g2419
  (
    n2572,
    n1908
  );


  not
  g2420
  (
    n2541,
    n2021
  );


  not
  g2421
  (
    n2851,
    n1971
  );


  not
  g2422
  (
    n2301,
    n1932
  );


  not
  g2423
  (
    n2292,
    n1598
  );


  not
  g2424
  (
    n2283,
    n1888
  );


  buf
  g2425
  (
    n2424,
    n1620
  );


  buf
  g2426
  (
    n2533,
    n1912
  );


  not
  g2427
  (
    n2562,
    n1602
  );


  buf
  g2428
  (
    n2590,
    n1974
  );


  buf
  g2429
  (
    n2483,
    n2009
  );


  not
  g2430
  (
    n2267,
    n1967
  );


  buf
  g2431
  (
    n2432,
    n1630
  );


  buf
  g2432
  (
    n2428,
    n1917
  );


  buf
  g2433
  (
    n2650,
    n1611
  );


  not
  g2434
  (
    n2538,
    n1948
  );


  not
  g2435
  (
    n2389,
    n1920
  );


  buf
  g2436
  (
    n2785,
    n1977
  );


  buf
  g2437
  (
    n2655,
    n1616
  );


  not
  g2438
  (
    n2720,
    n1962
  );


  buf
  g2439
  (
    n2392,
    n1883
  );


  buf
  g2440
  (
    n2793,
    n1610
  );


  not
  g2441
  (
    n2296,
    n1606
  );


  buf
  g2442
  (
    n2466,
    n1902
  );


  buf
  g2443
  (
    n2360,
    n1976
  );


  buf
  g2444
  (
    n2703,
    n1586
  );


  buf
  g2445
  (
    n2606,
    n1613
  );


  buf
  g2446
  (
    n2506,
    n1941
  );


  not
  g2447
  (
    n2270,
    n2019
  );


  not
  g2448
  (
    n2309,
    n1632
  );


  buf
  g2449
  (
    n2406,
    n1983
  );


  buf
  g2450
  (
    n2518,
    n1942
  );


  buf
  g2451
  (
    n2690,
    n2016
  );


  not
  g2452
  (
    n2443,
    n1886
  );


  buf
  g2453
  (
    n2747,
    n2000
  );


  not
  g2454
  (
    n2803,
    n1925
  );


  not
  g2455
  (
    n2566,
    n1905
  );


  not
  g2456
  (
    n2476,
    n1975
  );


  buf
  g2457
  (
    n2728,
    n1625
  );


  buf
  g2458
  (
    n2250,
    n1998
  );


  buf
  g2459
  (
    n2628,
    n1946
  );


  buf
  g2460
  (
    n2490,
    n1638
  );


  buf
  g2461
  (
    n2646,
    n1952
  );


  buf
  g2462
  (
    n2645,
    n1904
  );


  buf
  g2463
  (
    n2323,
    n1621
  );


  not
  g2464
  (
    n2756,
    n1946
  );


  buf
  g2465
  (
    n2784,
    n1923
  );


  buf
  g2466
  (
    n2261,
    n1607
  );


  not
  g2467
  (
    n2525,
    n2024
  );


  not
  g2468
  (
    n2528,
    n1619
  );


  buf
  g2469
  (
    n2514,
    n1928
  );


  buf
  g2470
  (
    n2675,
    n2021
  );


  not
  g2471
  (
    n2471,
    n1953
  );


  buf
  g2472
  (
    n2526,
    n2024
  );


  buf
  g2473
  (
    n2373,
    n1983
  );


  not
  g2474
  (
    n2423,
    n1611
  );


  not
  g2475
  (
    n2347,
    n1946
  );


  not
  g2476
  (
    n2480,
    n1635
  );


  buf
  g2477
  (
    n2613,
    n1593
  );


  not
  g2478
  (
    n2384,
    n1939
  );


  not
  g2479
  (
    n2731,
    n1887
  );


  buf
  g2480
  (
    n2790,
    n1978
  );


  buf
  g2481
  (
    n2485,
    n1958
  );


  buf
  g2482
  (
    n2329,
    n1954
  );


  buf
  g2483
  (
    n2626,
    n2023
  );


  buf
  g2484
  (
    n2472,
    n1906
  );


  buf
  g2485
  (
    n2266,
    n1887
  );


  buf
  g2486
  (
    n2750,
    n1937
  );


  not
  g2487
  (
    n2831,
    n1875
  );


  buf
  g2488
  (
    n2378,
    n1975
  );


  buf
  g2489
  (
    n2642,
    n1920
  );


  buf
  g2490
  (
    n2593,
    n1616
  );


  not
  g2491
  (
    n2792,
    n1937
  );


  buf
  g2492
  (
    n2619,
    n1945
  );


  not
  g2493
  (
    n2370,
    n2022
  );


  not
  g2494
  (
    n2382,
    n1626
  );


  not
  g2495
  (
    n2827,
    n1981
  );


  buf
  g2496
  (
    n2581,
    n2017
  );


  buf
  g2497
  (
    n2369,
    n1924
  );


  not
  g2498
  (
    n2462,
    n1896
  );


  buf
  g2499
  (
    n2365,
    n1957
  );


  buf
  g2500
  (
    n2682,
    n1997
  );


  not
  g2501
  (
    n2579,
    n1893
  );


  not
  g2502
  (
    n2781,
    n1979
  );


  buf
  g2503
  (
    n2252,
    n2020
  );


  not
  g2504
  (
    n2313,
    n2003
  );


  not
  g2505
  (
    n2519,
    n1947
  );


  buf
  g2506
  (
    n2853,
    n1901
  );


  not
  g2507
  (
    n2434,
    n1998
  );


  buf
  g2508
  (
    n2447,
    n2016
  );


  buf
  g2509
  (
    n2260,
    n1873
  );


  buf
  g2510
  (
    n2729,
    n1608
  );


  buf
  g2511
  (
    n2284,
    n1631
  );


  not
  g2512
  (
    n2285,
    n2022
  );


  buf
  g2513
  (
    n2439,
    n1589
  );


  buf
  g2514
  (
    n2656,
    n1621
  );


  not
  g2515
  (
    n2702,
    n1973
  );


  not
  g2516
  (
    n2359,
    n1940
  );


  buf
  g2517
  (
    n2786,
    n1619
  );


  not
  g2518
  (
    n2487,
    n1951
  );


  not
  g2519
  (
    n2544,
    n1933
  );


  not
  g2520
  (
    n2441,
    n1877
  );


  not
  g2521
  (
    n2421,
    n1930
  );


  buf
  g2522
  (
    n2492,
    n1589
  );


  buf
  g2523
  (
    n2507,
    n1625
  );


  not
  g2524
  (
    n2614,
    n1609
  );


  buf
  g2525
  (
    n2540,
    n1613
  );


  buf
  g2526
  (
    n2816,
    n1979
  );


  buf
  g2527
  (
    n2553,
    n1992
  );


  buf
  g2528
  (
    n2569,
    n1601
  );


  buf
  g2529
  (
    n2351,
    n1606
  );


  not
  g2530
  (
    n2817,
    n1989
  );


  not
  g2531
  (
    n2862,
    n1999
  );


  buf
  g2532
  (
    n2393,
    n1931
  );


  buf
  g2533
  (
    n2315,
    n1977
  );


  buf
  g2534
  (
    n2753,
    n1880
  );


  not
  g2535
  (
    n2243,
    n1622
  );


  buf
  g2536
  (
    n2564,
    n1969
  );


  buf
  g2537
  (
    n2543,
    n1884
  );


  not
  g2538
  (
    n2328,
    n1926
  );


  buf
  g2539
  (
    n2536,
    n1882
  );


  not
  g2540
  (
    n2290,
    n2016
  );


  not
  g2541
  (
    n2696,
    n1954
  );


  not
  g2542
  (
    n2789,
    n1893
  );


  buf
  g2543
  (
    n2659,
    n1615
  );


  not
  g2544
  (
    n2341,
    n1600
  );


  buf
  g2545
  (
    n2381,
    n1875
  );


  buf
  g2546
  (
    n2241,
    n1595
  );


  buf
  g2547
  (
    n2425,
    n1638
  );


  buf
  g2548
  (
    n2634,
    n1961
  );


  not
  g2549
  (
    n2367,
    n1594
  );


  not
  g2550
  (
    n2699,
    n1616
  );


  not
  g2551
  (
    n2780,
    n1914
  );


  buf
  g2552
  (
    n2852,
    n1902
  );


  buf
  g2553
  (
    n2486,
    n2005
  );


  not
  g2554
  (
    n2760,
    n1873
  );


  not
  g2555
  (
    n2832,
    n1935
  );


  buf
  g2556
  (
    n2380,
    n1943
  );


  buf
  g2557
  (
    n2712,
    n1943
  );


  not
  g2558
  (
    n2433,
    n2008
  );


  buf
  g2559
  (
    n2652,
    n1605
  );


  buf
  g2560
  (
    n2739,
    n2011
  );


  buf
  g2561
  (
    n2755,
    n1945
  );


  buf
  g2562
  (
    n2277,
    n2007
  );


  not
  g2563
  (
    n2345,
    n1933
  );


  buf
  g2564
  (
    n2317,
    n1963
  );


  not
  g2565
  (
    n2571,
    n2004
  );


  not
  g2566
  (
    n2807,
    n1983
  );


  not
  g2567
  (
    n2438,
    n1959
  );


  buf
  g2568
  (
    n2335,
    n1985
  );


  buf
  g2569
  (
    n2422,
    n1626
  );


  not
  g2570
  (
    n2713,
    n1603
  );


  not
  g2571
  (
    n2776,
    n1636
  );


  not
  g2572
  (
    n2407,
    n1934
  );


  not
  g2573
  (
    n2651,
    n1637
  );


  buf
  g2574
  (
    n2310,
    n1951
  );


  not
  g2575
  (
    n2499,
    n1627
  );


  not
  g2576
  (
    n2742,
    n1974
  );


  buf
  g2577
  (
    n2777,
    n2001
  );


  buf
  g2578
  (
    n2692,
    n1600
  );


  not
  g2579
  (
    n2582,
    n1960
  );


  not
  g2580
  (
    n2605,
    n2023
  );


  buf
  g2581
  (
    n2399,
    n1966
  );


  not
  g2582
  (
    n2849,
    n1611
  );


  not
  g2583
  (
    n2554,
    n1980
  );


  buf
  g2584
  (
    n2839,
    n1988
  );


  buf
  g2585
  (
    n2358,
    n1608
  );


  buf
  g2586
  (
    n2583,
    n1589
  );


  not
  g2587
  (
    n2375,
    n1893
  );


  buf
  g2588
  (
    n2385,
    n1957
  );


  buf
  g2589
  (
    n2495,
    n1927
  );


  not
  g2590
  (
    n2444,
    n1937
  );


  buf
  g2591
  (
    n2397,
    n1967
  );


  not
  g2592
  (
    n2452,
    n2002
  );


  buf
  g2593
  (
    n2584,
    n2011
  );


  not
  g2594
  (
    n2395,
    n1907
  );


  not
  g2595
  (
    n2357,
    n1970
  );


  not
  g2596
  (
    n2765,
    n1965
  );


  buf
  g2597
  (
    n2705,
    n1878
  );


  not
  g2598
  (
    n2481,
    n1905
  );


  not
  g2599
  (
    n2473,
    n2010
  );


  not
  g2600
  (
    n2809,
    n1999
  );


  buf
  g2601
  (
    n2567,
    n1919
  );


  not
  g2602
  (
    n2772,
    n1959
  );


  not
  g2603
  (
    n2587,
    n1957
  );


  not
  g2604
  (
    n2306,
    n1973
  );


  buf
  g2605
  (
    n2275,
    n1601
  );


  not
  g2606
  (
    n2561,
    n1604
  );


  not
  g2607
  (
    n2676,
    n1894
  );


  not
  g2608
  (
    n2442,
    n1593
  );


  not
  g2609
  (
    n2769,
    n1986
  );


  not
  g2610
  (
    n2242,
    n2021
  );


  not
  g2611
  (
    n2297,
    n1611
  );


  not
  g2612
  (
    n2746,
    n2022
  );


  buf
  g2613
  (
    n2574,
    n2018
  );


  buf
  g2614
  (
    n2245,
    n1872
  );


  not
  g2615
  (
    n2318,
    n2019
  );


  not
  g2616
  (
    n2819,
    n2007
  );


  not
  g2617
  (
    n2774,
    n1918
  );


  not
  g2618
  (
    n2269,
    n1965
  );


  buf
  g2619
  (
    n2740,
    n1632
  );


  buf
  g2620
  (
    n2300,
    n1956
  );


  buf
  g2621
  (
    n2508,
    n2009
  );


  not
  g2622
  (
    n2649,
    n1980
  );


  buf
  g2623
  (
    n2463,
    n1960
  );


  not
  g2624
  (
    n2282,
    n1588
  );


  not
  g2625
  (
    n2339,
    n1982
  );


  not
  g2626
  (
    n2657,
    n1990
  );


  buf
  g2627
  (
    n2537,
    n1960
  );


  not
  g2628
  (
    n2523,
    n1970
  );


  not
  g2629
  (
    n2420,
    n1990
  );


  buf
  g2630
  (
    n2417,
    n1876
  );


  buf
  g2631
  (
    n2348,
    n1871
  );


  buf
  g2632
  (
    n2732,
    n1943
  );


  buf
  g2633
  (
    n2294,
    n1585
  );


  buf
  g2634
  (
    n2394,
    n2003
  );


  not
  g2635
  (
    n2386,
    n1935
  );


  buf
  g2636
  (
    n2356,
    n1584
  );


  buf
  g2637
  (
    n2725,
    n1883
  );


  not
  g2638
  (
    n2630,
    n1903
  );


  not
  g2639
  (
    n2437,
    n1617
  );


  not
  g2640
  (
    n2336,
    n1932
  );


  buf
  g2641
  (
    n2860,
    n1620
  );


  not
  g2642
  (
    n2276,
    n1627
  );


  buf
  g2643
  (
    n2258,
    n1878
  );


  not
  g2644
  (
    n2474,
    n1887
  );


  not
  g2645
  (
    n2721,
    n1895
  );


  buf
  g2646
  (
    n2563,
    n1620
  );


  not
  g2647
  (
    n2427,
    n1912
  );


  not
  g2648
  (
    n2814,
    n1892
  );


  not
  g2649
  (
    n2601,
    n2001
  );


  buf
  g2650
  (
    n2741,
    n1936
  );


  not
  g2651
  (
    n2609,
    n1885
  );


  buf
  g2652
  (
    n2248,
    n1936
  );


  buf
  g2653
  (
    n2263,
    n1908
  );


  buf
  g2654
  (
    n2660,
    n1913
  );


  buf
  g2655
  (
    n2325,
    n1622
  );


  not
  g2656
  (
    n2457,
    n1913
  );


  not
  g2657
  (
    n2565,
    n1590
  );


  buf
  g2658
  (
    n2551,
    n1599
  );


  not
  g2659
  (
    n2342,
    n1613
  );


  not
  g2660
  (
    n2500,
    n1928
  );


  buf
  g2661
  (
    n2757,
    n1936
  );


  not
  g2662
  (
    n2391,
    n2019
  );


  buf
  g2663
  (
    n2256,
    n1992
  );


  buf
  g2664
  (
    n2272,
    n1939
  );


  buf
  g2665
  (
    n2364,
    n2018
  );


  not
  g2666
  (
    n2679,
    n1637
  );


  not
  g2667
  (
    n2409,
    n1592
  );


  not
  g2668
  (
    n2607,
    n1628
  );


  buf
  g2669
  (
    n2653,
    n1875
  );


  buf
  g2670
  (
    n2615,
    n1895
  );


  not
  g2671
  (
    n2346,
    n1899
  );


  not
  g2672
  (
    n2327,
    n1930
  );


  not
  g2673
  (
    n2458,
    n1919
  );


  buf
  g2674
  (
    n2249,
    n1873
  );


  not
  g2675
  (
    n2838,
    n1948
  );


  buf
  g2676
  (
    n2820,
    n2023
  );


  not
  g2677
  (
    n2598,
    n2006
  );


  not
  g2678
  (
    n2331,
    n1587
  );


  not
  g2679
  (
    n2496,
    n1625
  );


  buf
  g2680
  (
    n2796,
    n1990
  );


  buf
  g2681
  (
    n2833,
    n1633
  );


  buf
  g2682
  (
    n2733,
    n1591
  );


  buf
  g2683
  (
    n2663,
    n1620
  );


  buf
  g2684
  (
    n2255,
    n1602
  );


  buf
  g2685
  (
    n2843,
    n1914
  );


  buf
  g2686
  (
    n2639,
    n2007
  );


  buf
  g2687
  (
    n2815,
    n1986
  );


  not
  g2688
  (
    n2855,
    n1585
  );


  not
  g2689
  (
    n2247,
    n1876
  );


  buf
  g2690
  (
    n2794,
    n1892
  );


  buf
  g2691
  (
    n2787,
    n1871
  );


  not
  g2692
  (
    n2377,
    n1986
  );


  buf
  g2693
  (
    n2257,
    n1874
  );


  not
  g2694
  (
    n2783,
    n1609
  );


  not
  g2695
  (
    n2847,
    n2015
  );


  buf
  g2696
  (
    n2289,
    n1595
  );


  not
  g2697
  (
    n2239,
    n1951
  );


  not
  g2698
  (
    n2726,
    n1900
  );


  buf
  g2699
  (
    n2311,
    n1595
  );


  buf
  g2700
  (
    n2383,
    n1591
  );


  buf
  g2701
  (
    n2730,
    n1938
  );


  buf
  g2702
  (
    n2436,
    n1985
  );


  not
  g2703
  (
    n2738,
    n1889
  );


  buf
  g2704
  (
    n2453,
    n1623
  );


  not
  g2705
  (
    n2693,
    n1596
  );


  not
  g2706
  (
    n2431,
    n1902
  );


  buf
  g2707
  (
    n2813,
    n1940
  );


  buf
  g2708
  (
    n2577,
    n1930
  );


  not
  g2709
  (
    n2534,
    n1884
  );


  buf
  g2710
  (
    n2722,
    n2004
  );


  not
  g2711
  (
    n2558,
    n2008
  );


  buf
  g2712
  (
    n2811,
    n1993
  );


  not
  g2713
  (
    n2387,
    n1946
  );


  buf
  g2714
  (
    n2586,
    n1612
  );


  buf
  g2715
  (
    n2354,
    n1584
  );


  not
  g2716
  (
    n2510,
    n1879
  );


  not
  g2717
  (
    n2801,
    n1597
  );


  not
  g2718
  (
    n2527,
    n1598
  );


  not
  g2719
  (
    n2681,
    n1920
  );


  buf
  g2720
  (
    n2857,
    n1950
  );


  not
  g2721
  (
    n2622,
    n1906
  );


  buf
  g2722
  (
    n2291,
    n1917
  );


  buf
  g2723
  (
    n2677,
    n2000
  );


  not
  g2724
  (
    n2324,
    n1891
  );


  not
  g2725
  (
    n2273,
    n1955
  );


  buf
  g2726
  (
    n2246,
    n2002
  );


  buf
  g2727
  (
    n2338,
    n1624
  );


  buf
  g2728
  (
    n2850,
    n1945
  );


  buf
  g2729
  (
    n2379,
    n1963
  );


  buf
  g2730
  (
    n2824,
    n2005
  );


  buf
  g2731
  (
    n2695,
    n1636
  );


  buf
  g2732
  (
    n2368,
    n1590
  );


  not
  g2733
  (
    n2408,
    n1964
  );


  buf
  g2734
  (
    n2859,
    n1610
  );


  not
  g2735
  (
    n2451,
    n1962
  );


  buf
  g2736
  (
    n2454,
    n1916
  );


  buf
  g2737
  (
    n2735,
    n2017
  );


  buf
  g2738
  (
    n2644,
    n1930
  );


  buf
  g2739
  (
    n2724,
    n1992
  );


  buf
  g2740
  (
    n2638,
    n1630
  );


  buf
  g2741
  (
    n2715,
    n1877
  );


  not
  g2742
  (
    n2320,
    n1619
  );


  not
  g2743
  (
    n2858,
    n1587
  );


  buf
  g2744
  (
    n2669,
    n1583
  );


  buf
  g2745
  (
    n2662,
    n1600
  );


  not
  g2746
  (
    n2808,
    n1996
  );


  buf
  g2747
  (
    n2829,
    n1995
  );


  buf
  g2748
  (
    n2700,
    n1588
  );


  buf
  g2749
  (
    n2264,
    n1998
  );


  buf
  g2750
  (
    n2503,
    n1965
  );


  not
  g2751
  (
    n2573,
    n1608
  );


  buf
  g2752
  (
    n2743,
    n2005
  );


  not
  g2753
  (
    n2547,
    n1917
  );


  buf
  g2754
  (
    n2286,
    n1871
  );


  buf
  g2755
  (
    n2673,
    n2020
  );


  buf
  g2756
  (
    n2376,
    n1596
  );


  not
  g2757
  (
    n2343,
    n1896
  );


  or
  g2758
  (
    n2287,
    n1588,
    n1932,
    n2026,
    n1587
  );


  xor
  g2759
  (
    n2497,
    n1874,
    n1589,
    n1596,
    n1913
  );


  xnor
  g2760
  (
    n2298,
    n2027,
    n1958,
    n1894,
    n1910
  );


  or
  g2761
  (
    n2845,
    n1978,
    n1942,
    n1909,
    n1917
  );


  xnor
  g2762
  (
    n2491,
    n1614,
    n1986,
    n1593,
    n2020
  );


  or
  g2763
  (
    n2415,
    n1982,
    n1628,
    n1584,
    n1906
  );


  or
  g2764
  (
    n2591,
    n1964,
    n1906,
    n1931,
    n1619
  );


  nor
  g2765
  (
    n2295,
    n1995,
    n1981,
    n1922,
    n1609
  );


  or
  g2766
  (
    n2405,
    n1875,
    n1623,
    n1873,
    n1890
  );


  xor
  g2767
  (
    n2279,
    n1980,
    n1976,
    n1918,
    n1602
  );


  or
  g2768
  (
    n2468,
    n2009,
    n1614,
    n1634,
    n1895
  );


  xnor
  g2769
  (
    n2509,
    n1890,
    n1993,
    n1898,
    n2010
  );


  nand
  g2770
  (
    n2684,
    n1926,
    n1889,
    n1996,
    n1949
  );


  xnor
  g2771
  (
    n2687,
    n1908,
    n1897,
    n1606,
    n1900
  );


  or
  g2772
  (
    n2596,
    n2012,
    n1622,
    n1953,
    n1888
  );


  nand
  g2773
  (
    n2635,
    n1961,
    n1924,
    n1944,
    n1928
  );


  nor
  g2774
  (
    n2322,
    n1956,
    n1944,
    n1605,
    n1890
  );


  or
  g2775
  (
    n2449,
    n1940,
    n1989,
    n1614,
    n2008
  );


  xor
  g2776
  (
    n2766,
    n1892,
    n1882,
    n2025,
    n1999
  );


  xor
  g2777
  (
    n2799,
    n1889,
    n1966,
    n1962,
    n1592
  );


  and
  g2778
  (
    n2585,
    n1911,
    n1592,
    n1927,
    n1897
  );


  nor
  g2779
  (
    n2326,
    n1960,
    n1877,
    n1977,
    n1898
  );


  nor
  g2780
  (
    n2864,
    n1961,
    n1981,
    n1634,
    n1879
  );


  nor
  g2781
  (
    n2636,
    n1886,
    n1607,
    n1981,
    n1615
  );


  xor
  g2782
  (
    n2489,
    n1931,
    n1985,
    n1592,
    n1926
  );


  nor
  g2783
  (
    n2557,
    n1958,
    n1979,
    n1904,
    n1891
  );


  nand
  g2784
  (
    n2706,
    n1941,
    n2025,
    n1913,
    n1911
  );


  xor
  g2785
  (
    n2400,
    n1907,
    n1991,
    n1598,
    n1911
  );


  or
  g2786
  (
    n2841,
    n1874,
    n1897,
    n1624,
    n1598
  );


  xnor
  g2787
  (
    n2734,
    n2010,
    n1988,
    n1909,
    n1618
  );


  nor
  g2788
  (
    n2274,
    n1586,
    n1972,
    n2017,
    n1936
  );


  xor
  g2789
  (
    n2717,
    n1954,
    n1909,
    n1991,
    n1586
  );


  nand
  g2790
  (
    n2670,
    n1627,
    n1994,
    n2004,
    n1597
  );


  xor
  g2791
  (
    n2856,
    n1885,
    n1907,
    n1968,
    n1903
  );


  xnor
  g2792
  (
    n2482,
    n1923,
    n1599,
    n1989,
    n1607
  );


  nor
  g2793
  (
    n2773,
    n1953,
    n1987,
    n1985,
    n1887
  );


  xnor
  g2794
  (
    n2763,
    n1941,
    n1602,
    n1880,
    n1600
  );


  xor
  g2795
  (
    n2494,
    n1896,
    n1954,
    n1927,
    n1957
  );


  xor
  g2796
  (
    n2592,
    n1934,
    n1921,
    n1593,
    n2020
  );


  xor
  g2797
  (
    n2532,
    n1591,
    n1881,
    n1966,
    n1889
  );


  xnor
  g2798
  (
    n2795,
    n1881,
    n1994,
    n1915,
    n1916
  );


  nand
  g2799
  (
    n2710,
    n1638,
    n1888,
    n1879,
    n1958
  );


  and
  g2800
  (
    n2330,
    n2012,
    n1914,
    n1634,
    n1912
  );


  and
  g2801
  (
    n2752,
    n1883,
    n1633,
    n1927,
    n1612
  );


  xor
  g2802
  (
    n2836,
    n1594,
    n1891,
    n1982,
    n2002
  );


  nand
  g2803
  (
    n2680,
    n1984,
    n1972,
    n1617,
    n1944
  );


  nand
  g2804
  (
    n2484,
    n1982,
    n1963,
    n1922,
    n2011
  );


  xnor
  g2805
  (
    n2727,
    n1903,
    n1978,
    n2022,
    n1899
  );


  or
  g2806
  (
    n2854,
    n1615,
    n1952,
    n1894,
    n1968
  );


  and
  g2807
  (
    n2686,
    n1894,
    n1597,
    n1899,
    n2013
  );


  xnor
  g2808
  (
    n2404,
    n1972,
    n1637,
    n1915,
    n1617
  );


  or
  g2809
  (
    n2411,
    n1948,
    n1901,
    n1950,
    n1616
  );


  nand
  g2810
  (
    n2768,
    n2002,
    n1623,
    n2006,
    n1911
  );


  nand
  g2811
  (
    n2667,
    n1984,
    n1603,
    n2017,
    n2004
  );


  xor
  g2812
  (
    n2520,
    n1629,
    n1886,
    n1588,
    n1882
  );


  and
  g2813
  (
    n2685,
    n1955,
    n1950,
    n1905,
    n1885
  );


  nand
  g2814
  (
    n2837,
    n1595,
    n2014,
    n1872,
    n1884
  );


  or
  g2815
  (
    n2314,
    n2024,
    n1901,
    n1636,
    n2013
  );


  xnor
  g2816
  (
    n2683,
    n1631,
    n1878,
    n1633,
    n1594
  );


  xnor
  g2817
  (
    n2825,
    n1637,
    n1599,
    n2026,
    n1628
  );


  nand
  g2818
  (
    n2608,
    n2011,
    n1942,
    n2009,
    n1967
  );


  nand
  g2819
  (
    n2448,
    n1901,
    n1898,
    n1628,
    n1971
  );


  nor
  g2820
  (
    n2674,
    n1632,
    n1605,
    n1635,
    n1910
  );


  xor
  g2821
  (
    n2612,
    n1973,
    n1943,
    n1610,
    n1977
  );


  and
  g2822
  (
    n2737,
    n1934,
    n1987,
    n1984,
    n1942
  );


  nand
  g2823
  (
    n2361,
    n2001,
    n1918,
    n1932,
    n1629
  );


  nand
  g2824
  (
    n2802,
    n1912,
    n2015,
    n1921,
    n1984
  );


  xnor
  g2825
  (
    n2672,
    n1923,
    n1585,
    n2006,
    n1937
  );


  nor
  g2826
  (
    n2396,
    n2027,
    n1885,
    n1972,
    n2023
  );


  nand
  g2827
  (
    n2288,
    n1607,
    n1623,
    n1967,
    n1625
  );


  xor
  g2828
  (
    n2798,
    n1989,
    n1617,
    n2025,
    n1621
  );


  nor
  g2829
  (
    n2278,
    n1971,
    n1947,
    n1622,
    n1874
  );


  nor
  g2830
  (
    n2627,
    n1590,
    n1886,
    n1929,
    n1636
  );


  and
  g2831
  (
    n2716,
    n1968,
    n1883,
    n1926,
    n1891
  );


  buf
  g2832
  (
    n2877,
    n2241
  );


  buf
  g2833
  (
    n2879,
    n2248
  );


  buf
  g2834
  (
    n2868,
    n2247
  );


  not
  g2835
  (
    n2867,
    n2249
  );


  not
  g2836
  (
    n2871,
    n2240
  );


  not
  g2837
  (
    n2873,
    n2245
  );


  not
  g2838
  (
    n2865,
    n2239
  );


  not
  g2839
  (
    n2866,
    n2243
  );


  not
  g2840
  (
    n2880,
    n2251
  );


  not
  g2841
  (
    n2872,
    n2242
  );


  buf
  g2842
  (
    n2869,
    n2254
  );


  buf
  g2843
  (
    n2875,
    n2250
  );


  not
  g2844
  (
    n2876,
    n2244
  );


  buf
  g2845
  (
    n2874,
    n2252
  );


  not
  g2846
  (
    n2870,
    n2253
  );


  buf
  g2847
  (
    n2878,
    n2246
  );


  not
  g2848
  (
    n2890,
    n2869
  );


  not
  g2849
  (
    n2891,
    n2875
  );


  not
  g2850
  (
    n2894,
    n2874
  );


  not
  g2851
  (
    n2893,
    n2873
  );


  buf
  g2852
  (
    n2883,
    n2866
  );


  buf
  g2853
  (
    n2884,
    n2875
  );


  not
  g2854
  (
    n2886,
    n2868
  );


  buf
  g2855
  (
    n2888,
    n2871
  );


  buf
  g2856
  (
    n2882,
    n2874
  );


  not
  g2857
  (
    n2889,
    n2870
  );


  not
  g2858
  (
    n2887,
    n2872
  );


  buf
  g2859
  (
    n2885,
    n2865
  );


  buf
  g2860
  (
    n2881,
    n2867
  );


  buf
  g2861
  (
    n2892,
    n2873
  );


  not
  g2862
  (
    n2916,
    n2042
  );


  not
  g2863
  (
    n2908,
    n2032
  );


  buf
  g2864
  (
    n2922,
    n2045
  );


  buf
  g2865
  (
    n2933,
    n2889
  );


  not
  g2866
  (
    n2927,
    n2040
  );


  not
  g2867
  (
    n2913,
    n2027
  );


  not
  g2868
  (
    n2912,
    n2032
  );


  buf
  g2869
  (
    n2940,
    n2881
  );


  not
  g2870
  (
    n2899,
    n2885
  );


  not
  g2871
  (
    n2896,
    n2045
  );


  buf
  g2872
  (
    n2947,
    n2040
  );


  not
  g2873
  (
    n2950,
    n2039
  );


  buf
  g2874
  (
    n2921,
    n2884
  );


  buf
  g2875
  (
    n2932,
    n2886
  );


  buf
  g2876
  (
    n2924,
    n2893
  );


  buf
  g2877
  (
    n2926,
    n2035
  );


  buf
  g2878
  (
    n2902,
    n2043
  );


  not
  g2879
  (
    n2949,
    n2036
  );


  not
  g2880
  (
    n2914,
    n2888
  );


  buf
  g2881
  (
    n2948,
    n2039
  );


  not
  g2882
  (
    n2944,
    n2033
  );


  not
  g2883
  (
    n2943,
    n2882
  );


  buf
  g2884
  (
    n2907,
    n2032
  );


  buf
  g2885
  (
    n2903,
    n2894
  );


  not
  g2886
  (
    n2930,
    n2893
  );


  not
  g2887
  (
    n2920,
    n2883
  );


  not
  g2888
  (
    n2919,
    n2030
  );


  buf
  g2889
  (
    n2904,
    n2034
  );


  nand
  g2890
  (
    n2925,
    n2041,
    n2256
  );


  nand
  g2891
  (
    n2895,
    n2041,
    n2891,
    n2881,
    n2887
  );


  xnor
  g2892
  (
    n2941,
    n2030,
    n2033,
    n2886,
    n2882
  );


  or
  g2893
  (
    n2910,
    n2029,
    n2039,
    n2894,
    n2044
  );


  nor
  g2894
  (
    n2918,
    n2044,
    n2891,
    n2888,
    n2882
  );


  xor
  g2895
  (
    n2901,
    n2890,
    n2028,
    n2034,
    n2881
  );


  nor
  g2896
  (
    n2942,
    n2891,
    n2028,
    n2042,
    n2030
  );


  xor
  g2897
  (
    n2939,
    n2890,
    n2875,
    n2031
  );


  xor
  g2898
  (
    n2936,
    n2890,
    n2255,
    n2028,
    n2892
  );


  or
  g2899
  (
    n2900,
    n2034,
    n2885,
    n2037,
    n2045
  );


  xnor
  g2900
  (
    n2923,
    n2030,
    n2888,
    n2037,
    n2041
  );


  nand
  g2901
  (
    n2898,
    n2038,
    n2889,
    n2890,
    n2036
  );


  xor
  g2902
  (
    n2909,
    n2884,
    n2045,
    n2036,
    n2892
  );


  nor
  g2903
  (
    n2931,
    n2892,
    n2893,
    n2035
  );


  xnor
  g2904
  (
    n2934,
    n2887,
    n2042,
    n2029,
    n2046
  );


  and
  g2905
  (
    n2938,
    n2043,
    n2035,
    n2040,
    n2876
  );


  or
  g2906
  (
    n2937,
    n2027,
    n2893,
    n2038,
    n2044
  );


  xnor
  g2907
  (
    n2935,
    n2044,
    n2891,
    n2028,
    n2038
  );


  xnor
  g2908
  (
    n2946,
    n2036,
    n2040,
    n2887,
    n2876
  );


  nand
  g2909
  (
    n2929,
    n2882,
    n2883,
    n2894,
    n2037
  );


  nor
  g2910
  (
    n2915,
    n2042,
    n2031,
    n2892
  );


  and
  g2911
  (
    n2911,
    n2885,
    n2883,
    n2038
  );


  nand
  g2912
  (
    n2906,
    n2884,
    n2033,
    n2885,
    n2029
  );


  or
  g2913
  (
    n2928,
    n2041,
    n2886,
    n2881
  );


  xnor
  g2914
  (
    n2897,
    n2033,
    n2032,
    n2039,
    n2887
  );


  xor
  g2915
  (
    n2905,
    n2029,
    n2888,
    n2876,
    n2884
  );


  xnor
  g2916
  (
    n2917,
    n2031,
    n2043,
    n2037
  );


  nand
  g2917
  (
    n2945,
    n2894,
    n2889,
    n2034
  );


  nand
  g2918
  (
    n3132,
    n2821,
    n2925,
    n2290,
    n2927
  );


  nand
  g2919
  (
    n3042,
    n2303,
    n2907,
    n2788,
    n2362
  );


  or
  g2920
  (
    n3000,
    n2809,
    n2620,
    n2499,
    n2790
  );


  xor
  g2921
  (
    n3002,
    n2819,
    n2921,
    n2802,
    n2280
  );


  xnor
  g2922
  (
    n2995,
    n2764,
    n2657,
    n2934,
    n2455
  );


  xor
  g2923
  (
    n3039,
    n2947,
    n2724,
    n2429,
    n2744
  );


  or
  g2924
  (
    n3126,
    n2603,
    n2722,
    n2310,
    n2335
  );


  nand
  g2925
  (
    n3019,
    n2918,
    n2318,
    n2590,
    n2440
  );


  xnor
  g2926
  (
    n3057,
    n2917,
    n2918,
    n2287,
    n2766
  );


  xor
  g2927
  (
    n2971,
    n2906,
    n2943,
    n2827,
    n2904
  );


  and
  g2928
  (
    n3112,
    n2598,
    n2946,
    n2941,
    n2388
  );


  xnor
  g2929
  (
    n2984,
    n2288,
    n2810,
    n2820,
    n2930
  );


  xor
  g2930
  (
    n3158,
    n2322,
    n2907,
    n2291,
    n2732
  );


  xor
  g2931
  (
    n3139,
    n2940,
    n2597,
    n2914,
    n2739
  );


  and
  g2932
  (
    n3147,
    n2470,
    n2793,
    n2929,
    n2803
  );


  and
  g2933
  (
    n3053,
    n2917,
    n2822,
    n2258,
    n2825
  );


  xor
  g2934
  (
    n3157,
    n2457,
    n2771,
    n2497,
    n2430
  );


  and
  g2935
  (
    n2981,
    n2344,
    n2824,
    n2905,
    n2391
  );


  nor
  g2936
  (
    n3058,
    n2814,
    n2336,
    n2758,
    n2784
  );


  xor
  g2937
  (
    n3099,
    n2338,
    n2553,
    n2899,
    n2804
  );


  xnor
  g2938
  (
    n3030,
    n2697,
    n2301,
    n2692,
    n2802
  );


  and
  g2939
  (
    n3050,
    n2273,
    n2815,
    n2465,
    n2902
  );


  nor
  g2940
  (
    n3078,
    n2762,
    n2292,
    n2792,
    n2749
  );


  nand
  g2941
  (
    n3172,
    n2320,
    n2816,
    n2809,
    n2921
  );


  nand
  g2942
  (
    n3013,
    n2895,
    n2817,
    n2294,
    n2750
  );


  xor
  g2943
  (
    n3017,
    n2793,
    n2549,
    n2935,
    n2932
  );


  xor
  g2944
  (
    n3137,
    n2913,
    n2263,
    n2488,
    n2786
  );


  xnor
  g2945
  (
    n3026,
    n2542,
    n2915,
    n2912,
    n2560
  );


  xnor
  g2946
  (
    n2998,
    n2752,
    n2803,
    n2467,
    n2348
  );


  and
  g2947
  (
    n3118,
    n2307,
    n2928,
    n2803,
    n2541
  );


  nor
  g2948
  (
    n2954,
    n2368,
    n2920,
    n2821,
    n2330
  );


  nor
  g2949
  (
    n3110,
    n2899,
    n2458,
    n2407,
    n2933
  );


  xor
  g2950
  (
    n3065,
    n2577,
    n2478,
    n2921,
    n2668
  );


  and
  g2951
  (
    n3051,
    n2340,
    n2936,
    n2587,
    n2647
  );


  xnor
  g2952
  (
    n3055,
    n2600,
    n2791,
    n2796,
    n2581
  );


  and
  g2953
  (
    n3084,
    n2919,
    n2398,
    n2944,
    n2820
  );


  nor
  g2954
  (
    n3034,
    n2801,
    n2686,
    n2923,
    n2910
  );


  nand
  g2955
  (
    n3029,
    n2930,
    n2828,
    n2895,
    n2713
  );


  and
  g2956
  (
    n2970,
    n2460,
    n2919,
    n2576,
    n2923
  );


  xor
  g2957
  (
    n3136,
    n2903,
    n2807,
    n2937,
    n2765
  );


  xnor
  g2958
  (
    n3040,
    n2548,
    n2259,
    n2622,
    n2511
  );


  xnor
  g2959
  (
    n3038,
    n2828,
    n2510,
    n2520,
    n2527
  );


  xnor
  g2960
  (
    n3125,
    n2373,
    n2902,
    n2694,
    n2566
  );


  or
  g2961
  (
    n2992,
    n2439,
    n2437,
    n2534,
    n2760
  );


  or
  g2962
  (
    n2976,
    n2350,
    n2289,
    n2804,
    n2803
  );


  nand
  g2963
  (
    n3075,
    n2896,
    n2660,
    n2923,
    n2674
  );


  or
  g2964
  (
    n2969,
    n2742,
    n2611,
    n2905,
    n2798
  );


  and
  g2965
  (
    n3074,
    n2807,
    n2471,
    n2354,
    n2826
  );


  nor
  g2966
  (
    n3062,
    n2926,
    n2821,
    n2333,
    n2450
  );


  or
  g2967
  (
    n2983,
    n2526,
    n2789,
    n2297,
    n2942
  );


  xor
  g2968
  (
    n3047,
    n2516,
    n2494,
    n2818,
    n2403
  );


  nor
  g2969
  (
    n2997,
    n2571,
    n2311,
    n2939,
    n2356
  );


  or
  g2970
  (
    n2991,
    n2706,
    n2945,
    n2802,
    n2613
  );


  and
  g2971
  (
    n3120,
    n2504,
    n2932,
    n2824,
    n2814
  );


  xnor
  g2972
  (
    n3024,
    n2931,
    n2808,
    n2917,
    n2740
  );


  or
  g2973
  (
    n3117,
    n2924,
    n2279,
    n2769,
    n2767
  );


  or
  g2974
  (
    n3077,
    n2777,
    n2423,
    n2591,
    n2296
  );


  or
  g2975
  (
    n3022,
    n2519,
    n2737,
    n2559,
    n2916
  );


  xnor
  g2976
  (
    n2961,
    n2472,
    n2807,
    n2524,
    n2721
  );


  nor
  g2977
  (
    n3079,
    n2912,
    n2770,
    n2808,
    n2947
  );


  nor
  g2978
  (
    n3091,
    n2905,
    n2941,
    n2409,
    n2321
  );


  xnor
  g2979
  (
    n2965,
    n2349,
    n2378,
    n2826,
    n2907
  );


  and
  g2980
  (
    n3031,
    n2772,
    n2924,
    n2480,
    n2512
  );


  and
  g2981
  (
    n3054,
    n2655,
    n2275,
    n2919,
    n2584
  );


  nor
  g2982
  (
    n2975,
    n2284,
    n2334,
    n2332,
    n2546
  );


  nor
  g2983
  (
    n2964,
    n2736,
    n2552,
    n2416,
    n2308
  );


  or
  g2984
  (
    n3119,
    n2323,
    n2897,
    n2756,
    n2693
  );


  xor
  g2985
  (
    n3066,
    n2948,
    n2950,
    n2313,
    n2570
  );


  xor
  g2986
  (
    n3138,
    n2930,
    n2901,
    n2940,
    n2386
  );


  nor
  g2987
  (
    n3086,
    n2650,
    n2822,
    n2942,
    n2343
  );


  xnor
  g2988
  (
    n3169,
    n2493,
    n2895,
    n2918,
    n2666
  );


  nand
  g2989
  (
    n3060,
    n2537,
    n2325,
    n2824,
    n2466
  );


  or
  g2990
  (
    n3015,
    n2902,
    n2896,
    n2446,
    n2353
  );


  nor
  g2991
  (
    n2953,
    n2947,
    n2813,
    n2469,
    n2811
  );


  nand
  g2992
  (
    n3048,
    n2578,
    n2747,
    n2714,
    n2539
  );


  xnor
  g2993
  (
    n3063,
    n2705,
    n2827,
    n2417,
    n2931
  );


  xnor
  g2994
  (
    n3166,
    n2561,
    n2640,
    n2806,
    n2532
  );


  xnor
  g2995
  (
    n2999,
    n2932,
    n2574,
    n2726,
    n2808
  );


  and
  g2996
  (
    n2972,
    n2910,
    n2932,
    n2648,
    n2933
  );


  and
  g2997
  (
    n3127,
    n2729,
    n2509,
    n2925,
    n2798
  );


  or
  g2998
  (
    n3056,
    n2627,
    n2669,
    n2486,
    n2695
  );


  xnor
  g2999
  (
    n3155,
    n2635,
    n2501,
    n2934,
    n2923
  );


  xor
  g3000
  (
    n3011,
    n2445,
    n2656,
    n2634,
    n2496
  );


  or
  g3001
  (
    n3076,
    n2804,
    n2704,
    n2625,
    n2431
  );


  xor
  g3002
  (
    n3100,
    n2911,
    n2420,
    n2805,
    n2929
  );


  or
  g3003
  (
    n3059,
    n2940,
    n2817,
    n2408,
    n2828
  );


  and
  g3004
  (
    n3016,
    n2926,
    n2376,
    n2557,
    n2393
  );


  xor
  g3005
  (
    n3068,
    n2502,
    n2814,
    n2707,
    n2346
  );


  nand
  g3006
  (
    n3144,
    n2565,
    n2616,
    n2468,
    n2367
  );


  xor
  g3007
  (
    n3160,
    n2528,
    n2361,
    n2935,
    n2801
  );


  or
  g3008
  (
    n3089,
    n2505,
    n2819,
    n2283,
    n2271
  );


  xor
  g3009
  (
    n3010,
    n2305,
    n2806,
    n2435,
    n2529
  );


  or
  g3010
  (
    n3090,
    n2944,
    n2691,
    n2612,
    n2643
  );


  nand
  g3011
  (
    n3174,
    n2931,
    n2454,
    n2795,
    n2823
  );


  or
  g3012
  (
    n3148,
    n2298,
    n2916,
    n2461,
    n2898
  );


  nand
  g3013
  (
    n3064,
    n2799,
    n2508,
    n2943,
    n2517
  );


  nor
  g3014
  (
    n3161,
    n2820,
    n2915,
    n2272,
    n2825
  );


  nor
  g3015
  (
    n3122,
    n2751,
    n2935,
    n2823,
    n2599
  );


  and
  g3016
  (
    n2967,
    n2910,
    n2820,
    n2500,
    n2649
  );


  and
  g3017
  (
    n3130,
    n2276,
    n2473,
    n2452,
    n2422
  );


  or
  g3018
  (
    n2958,
    n2937,
    n2658,
    n2914,
    n2268
  );


  nor
  g3019
  (
    n3025,
    n2818,
    n2813,
    n2897,
    n2347
  );


  nand
  g3020
  (
    n3101,
    n2352,
    n2608,
    n2463,
    n2938
  );


  nand
  g3021
  (
    n3008,
    n2802,
    n2383,
    n2942,
    n2829
  );


  xnor
  g3022
  (
    n3097,
    n2806,
    n2949,
    n2776,
    n2646
  );


  and
  g3023
  (
    n3107,
    n2918,
    n2490,
    n2567,
    n2360
  );


  and
  g3024
  (
    n2988,
    n2782,
    n2927,
    n2487,
    n2815
  );


  nor
  g3025
  (
    n3071,
    n2538,
    n2653,
    n2719,
    n2741
  );


  xnor
  g3026
  (
    n2977,
    n2413,
    n2941,
    n2909,
    n2810
  );


  xnor
  g3027
  (
    n3082,
    n2579,
    n2588,
    n2926,
    n2483
  );


  nand
  g3028
  (
    n3044,
    n2518,
    n2485,
    n2949,
    n2916
  );


  or
  g3029
  (
    n2955,
    n2700,
    n2324,
    n2451,
    n2545
  );


  nor
  g3030
  (
    n3020,
    n2796,
    n2896,
    n2807,
    n2339
  );


  xor
  g3031
  (
    n2986,
    n2269,
    n2922,
    n2811,
    n2651
  );


  xnor
  g3032
  (
    n2962,
    n2474,
    n2394,
    n2641,
    n2908
  );


  or
  g3033
  (
    n3141,
    n2441,
    n2787,
    n2319,
    n2639
  );


  xor
  g3034
  (
    n3093,
    n2604,
    n2927,
    n2895,
    n2946
  );


  or
  g3035
  (
    n3168,
    n2937,
    n2621,
    n2723,
    n2819
  );


  or
  g3036
  (
    n3046,
    n2626,
    n2609,
    n2628,
    n2551
  );


  xnor
  g3037
  (
    n3165,
    n2901,
    n2950,
    n2817,
    n2903
  );


  xnor
  g3038
  (
    n3072,
    n2358,
    n2733,
    n2790,
    n2414
  );


  or
  g3039
  (
    n3032,
    n2900,
    n2773,
    n2444,
    n2369
  );


  xnor
  g3040
  (
    n3043,
    n2825,
    n2533,
    n2709,
    n2810
  );


  xor
  g3041
  (
    n3087,
    n2816,
    n2663,
    n2811,
    n2925
  );


  nand
  g3042
  (
    n3061,
    n2531,
    n2816,
    n2933,
    n2428
  );


  and
  g3043
  (
    n3142,
    n2827,
    n2938,
    n2920,
    n2679
  );


  xnor
  g3044
  (
    n2960,
    n2902,
    n2944,
    n2905,
    n2900
  );


  xor
  g3045
  (
    n3096,
    n2822,
    n2899,
    n2406,
    n2400
  );


  and
  g3046
  (
    n2996,
    n2931,
    n2933,
    n2906,
    n2809
  );


  nand
  g3047
  (
    n3083,
    n2690,
    n2909,
    n2285,
    n2915
  );


  and
  g3048
  (
    n3067,
    n2788,
    n2754,
    n2712,
    n2415
  );


  xnor
  g3049
  (
    n3114,
    n2375,
    n2645,
    n2521,
    n2898
  );


  nor
  g3050
  (
    n3081,
    n2900,
    n2665,
    n2728,
    n2464
  );


  and
  g3051
  (
    n3124,
    n2904,
    n2914,
    n2359,
    n2642
  );


  nand
  g3052
  (
    n3146,
    n2936,
    n2947,
    n2513,
    n2912
  );


  xor
  g3053
  (
    n3153,
    n2783,
    n2427,
    n2326,
    n2564
  );


  and
  g3054
  (
    n3092,
    n2506,
    n2936,
    n2572,
    n2731
  );


  nand
  g3055
  (
    n3103,
    n2928,
    n2593,
    n2794,
    n2812
  );


  nand
  g3056
  (
    n3111,
    n2934,
    n2816,
    n2396,
    n2688
  );


  xnor
  g3057
  (
    n3045,
    n2791,
    n2780,
    n2799,
    n2329
  );


  xor
  g3058
  (
    n3121,
    n2921,
    n2805,
    n2677,
    n2372
  );


  xor
  g3059
  (
    n3105,
    n2476,
    n2821,
    n2814,
    n2795
  );


  nand
  g3060
  (
    n3036,
    n2392,
    n2948,
    n2462,
    n2730
  );


  nand
  g3061
  (
    n2987,
    n2312,
    n2805,
    n2675,
    n2926
  );


  nand
  g3062
  (
    n3143,
    n2436,
    n2337,
    n2936,
    n2897
  );


  xor
  g3063
  (
    n3080,
    n2390,
    n2395,
    n2274,
    n2586
  );


  xor
  g3064
  (
    n3085,
    n2607,
    n2257,
    n2922,
    n2550
  );


  or
  g3065
  (
    n3028,
    n2819,
    n2940,
    n2797,
    n2738
  );


  xor
  g3066
  (
    n2980,
    n2699,
    n2810,
    n2569,
    n2759
  );


  xnor
  g3067
  (
    n3129,
    n2778,
    n2911,
    n2498,
    n2535
  );


  or
  g3068
  (
    n3151,
    n2374,
    n2351,
    n2380,
    n2619
  );


  xnor
  g3069
  (
    n3167,
    n2681,
    n2278,
    n2671,
    n2265
  );


  xor
  g3070
  (
    n3171,
    n2734,
    n2379,
    n2629,
    n2727
  );


  xnor
  g3071
  (
    n3149,
    n2913,
    n2903,
    n2503,
    n2575
  );


  xnor
  g3072
  (
    n2978,
    n2815,
    n2410,
    n2633,
    n2904
  );


  and
  g3073
  (
    n2951,
    n2624,
    n2264,
    n2689,
    n2768
  );


  nor
  g3074
  (
    n3006,
    n2680,
    n2293,
    n2585,
    n2781
  );


  nand
  g3075
  (
    n3037,
    n2456,
    n2295,
    n2632,
    n2929
  );


  xor
  g3076
  (
    n3007,
    n2302,
    n2914,
    n2421,
    n2667
  );


  xor
  g3077
  (
    n3021,
    n2748,
    n2755,
    n2939,
    n2397
  );


  or
  g3078
  (
    n3049,
    n2716,
    n2911,
    n2568,
    n2910
  );


  nor
  g3079
  (
    n3052,
    n2725,
    n2774,
    n2753,
    n2507
  );


  and
  g3080
  (
    n3140,
    n2345,
    n2594,
    n2554,
    n2948
  );


  or
  g3081
  (
    n2952,
    n2434,
    n2698,
    n2911,
    n2818
  );


  or
  g3082
  (
    n3163,
    n2826,
    n2939,
    n2491,
    n2827
  );


  and
  g3083
  (
    n3113,
    n2381,
    n2525,
    n2938,
    n2828
  );


  xor
  g3084
  (
    n2959,
    n2443,
    n2662,
    n2328,
    n2806
  );


  xnor
  g3085
  (
    n2982,
    n2479,
    n2913,
    n2946,
    n2556
  );


  nor
  g3086
  (
    n3005,
    n2630,
    n2904,
    n2299,
    n2711
  );


  nand
  g3087
  (
    n3154,
    n2929,
    n2654,
    n2672,
    n2907
  );


  xor
  g3088
  (
    n3162,
    n2897,
    n2419,
    n2637,
    n2946
  );


  nand
  g3089
  (
    n3123,
    n2787,
    n2797,
    n2636,
    n2615
  );


  and
  g3090
  (
    n3027,
    n2823,
    n2934,
    n2514,
    n2364
  );


  xnor
  g3091
  (
    n2985,
    n2614,
    n2922,
    n2924,
    n2573
  );


  nand
  g3092
  (
    n3069,
    n2717,
    n2592,
    n2304,
    n2453
  );


  nor
  g3093
  (
    n3145,
    n2949,
    n2913,
    n2377,
    n2813
  );


  xnor
  g3094
  (
    n3134,
    n2331,
    n2266,
    n2523,
    n2945
  );


  nor
  g3095
  (
    n3088,
    n2327,
    n2558,
    n2306,
    n2363
  );


  or
  g3096
  (
    n3152,
    n2481,
    n2425,
    n2915,
    n2402
  );


  or
  g3097
  (
    n3108,
    n2316,
    n2908,
    n2950,
    n2815
  );


  xor
  g3098
  (
    n2973,
    n2638,
    n2687,
    n2432,
    n2366
  );


  nor
  g3099
  (
    n3115,
    n2938,
    n2644,
    n2900,
    n2829
  );


  and
  g3100
  (
    n2963,
    n2829,
    n2785,
    n2606,
    n2922
  );


  or
  g3101
  (
    n3070,
    n2401,
    n2543,
    n2399,
    n2424
  );


  or
  g3102
  (
    n3001,
    n2605,
    n2903,
    n2261,
    n2670
  );


  xnor
  g3103
  (
    n3133,
    n2365,
    n2286,
    n2300,
    n2384
  );


  or
  g3104
  (
    n3102,
    n2925,
    n2817,
    n2812,
    n2342
  );


  xor
  g3105
  (
    n3170,
    n2919,
    n2314,
    n2530,
    n2805
  );


  or
  g3106
  (
    n2994,
    n2617,
    n2522,
    n2950,
    n2942
  );


  nand
  g3107
  (
    n3164,
    n2735,
    n2899,
    n2448,
    n2580
  );


  xnor
  g3108
  (
    n3135,
    n2673,
    n2928,
    n2482,
    n2909
  );


  nor
  g3109
  (
    n3109,
    n2935,
    n2800,
    n2411,
    n2555
  );


  or
  g3110
  (
    n3159,
    n2812,
    n2659,
    n2610,
    n2405
  );


  nand
  g3111
  (
    n2993,
    n2357,
    n2449,
    n2618,
    n2652
  );


  nor
  g3112
  (
    n3018,
    n2418,
    n2908,
    n2917,
    n2433
  );


  nand
  g3113
  (
    n2957,
    n2924,
    n2949,
    n2825,
    n2582
  );


  xor
  g3114
  (
    n3014,
    n2631,
    n2794,
    n2927,
    n2916
  );


  or
  g3115
  (
    n2966,
    n2945,
    n2941,
    n2901,
    n2315
  );


  nand
  g3116
  (
    n3073,
    n2563,
    n2761,
    n2696,
    n2341
  );


  xor
  g3117
  (
    n3095,
    n2822,
    n2896,
    n2710,
    n2601
  );


  or
  g3118
  (
    n3104,
    n2945,
    n2757,
    n2912,
    n2676
  );


  nand
  g3119
  (
    n3041,
    n2811,
    n2412,
    n2678,
    n2370
  );


  nand
  g3120
  (
    n2956,
    n2715,
    n2743,
    n2824,
    n2426
  );


  nand
  g3121
  (
    n2989,
    n2544,
    n2826,
    n2515,
    n2355
  );


  nand
  g3122
  (
    n3033,
    n2702,
    n2901,
    n2562,
    n2829
  );


  or
  g3123
  (
    n3023,
    n2489,
    n2939,
    n2718,
    n2492
  );


  or
  g3124
  (
    n3173,
    n2906,
    n2685,
    n2746,
    n2909
  );


  nor
  g3125
  (
    n3106,
    n2583,
    n2812,
    n2438,
    n2270
  );


  xnor
  g3126
  (
    n3131,
    n2495,
    n2371,
    n2937,
    n2664
  );


  xor
  g3127
  (
    n2968,
    n2908,
    n2906,
    n2898,
    n2701
  );


  xor
  g3128
  (
    n2979,
    n2720,
    n2683,
    n2404,
    n2944
  );


  and
  g3129
  (
    n3156,
    n2385,
    n2818,
    n2763,
    n2602
  );


  xor
  g3130
  (
    n3004,
    n2317,
    n2930,
    n2948,
    n2898
  );


  and
  g3131
  (
    n3116,
    n2682,
    n2928,
    n2745,
    n2389
  );


  nor
  g3132
  (
    n3009,
    n2459,
    n2475,
    n2789,
    n2920
  );


  nor
  g3133
  (
    n3012,
    n2387,
    n2267,
    n2943,
    n2309
  );


  nor
  g3134
  (
    n3035,
    n2808,
    n2382,
    n2595,
    n2262
  );


  or
  g3135
  (
    n3094,
    n2282,
    n2804,
    n2661,
    n2800
  );


  xnor
  g3136
  (
    n3003,
    n2943,
    n2442,
    n2540,
    n2596
  );


  xor
  g3137
  (
    n3128,
    n2809,
    n2920,
    n2779,
    n2623
  );


  xnor
  g3138
  (
    n3098,
    n2447,
    n2708,
    n2823,
    n2684
  );


  nor
  g3139
  (
    n3150,
    n2589,
    n2484,
    n2703,
    n2260
  );


  xor
  g3140
  (
    n2974,
    n2477,
    n2775,
    n2792,
    n2547
  );


  nand
  g3141
  (
    n2990,
    n2277,
    n2281,
    n2536,
    n2813
  );


  buf
  g3142
  (
    n3285,
    n3083
  );


  not
  g3143
  (
    n3242,
    n2100
  );


  buf
  g3144
  (
    n3478,
    n2217
  );


  buf
  g3145
  (
    n3504,
    n2050
  );


  not
  g3146
  (
    n3331,
    n2118
  );


  not
  g3147
  (
    n3458,
    n3031
  );


  buf
  g3148
  (
    n3464,
    n2999
  );


  buf
  g3149
  (
    n3404,
    n3056
  );


  not
  g3150
  (
    n3309,
    n2066
  );


  not
  g3151
  (
    n3320,
    n2996
  );


  not
  g3152
  (
    n3395,
    n2140
  );


  not
  g3153
  (
    n3381,
    n2108
  );


  not
  g3154
  (
    n3586,
    n3010
  );


  buf
  g3155
  (
    n3451,
    n3020
  );


  buf
  g3156
  (
    n3313,
    n3015
  );


  buf
  g3157
  (
    n3317,
    n2976
  );


  buf
  g3158
  (
    n3352,
    n2230
  );


  buf
  g3159
  (
    n3449,
    n3134
  );


  buf
  g3160
  (
    n3348,
    n2061
  );


  not
  g3161
  (
    n3343,
    n2173
  );


  not
  g3162
  (
    n3355,
    n3031
  );


  buf
  g3163
  (
    n3253,
    n2169
  );


  not
  g3164
  (
    n3578,
    n3157
  );


  buf
  g3165
  (
    n3558,
    n3131
  );


  buf
  g3166
  (
    n3333,
    n3062
  );


  buf
  g3167
  (
    n3608,
    n2105
  );


  buf
  g3168
  (
    n3514,
    n3058
  );


  not
  g3169
  (
    n3367,
    n3125
  );


  buf
  g3170
  (
    n3209,
    n2222
  );


  buf
  g3171
  (
    n3374,
    n2053
  );


  buf
  g3172
  (
    n3393,
    n3139
  );


  buf
  g3173
  (
    n3548,
    n2053
  );


  buf
  g3174
  (
    n3216,
    n2128
  );


  not
  g3175
  (
    n3254,
    n3148
  );


  not
  g3176
  (
    n3516,
    n3068
  );


  buf
  g3177
  (
    n3403,
    n2981
  );


  buf
  g3178
  (
    n3314,
    n3050
  );


  not
  g3179
  (
    n3480,
    n3071
  );


  buf
  g3180
  (
    n3214,
    n2059
  );


  buf
  g3181
  (
    n3509,
    n2195
  );


  not
  g3182
  (
    n3197,
    n2166
  );


  not
  g3183
  (
    n3294,
    n2064
  );


  not
  g3184
  (
    n3524,
    n3109
  );


  buf
  g3185
  (
    n3231,
    n3041
  );


  not
  g3186
  (
    n3570,
    n2974
  );


  not
  g3187
  (
    n3398,
    n2091
  );


  not
  g3188
  (
    n3501,
    n2103
  );


  not
  g3189
  (
    n3500,
    n3030
  );


  not
  g3190
  (
    n3202,
    n2225
  );


  buf
  g3191
  (
    n3421,
    n2065
  );


  buf
  g3192
  (
    n3468,
    n2086
  );


  buf
  g3193
  (
    n3407,
    n2082
  );


  not
  g3194
  (
    n3566,
    n2114
  );


  not
  g3195
  (
    n3511,
    n2998
  );


  buf
  g3196
  (
    n3342,
    n3129
  );


  and
  g3197
  (
    n3510,
    n2049,
    n3151,
    n2972,
    n3032
  );


  xnor
  g3198
  (
    n3267,
    n2086,
    n2174,
    n3159,
    n2101
  );


  and
  g3199
  (
    n3584,
    n2142,
    n3143,
    n2055,
    n2219
  );


  and
  g3200
  (
    n3463,
    n2076,
    n2997,
    n3113,
    n3068
  );


  or
  g3201
  (
    n3571,
    n2973,
    n3007,
    n2102,
    n3063
  );


  or
  g3202
  (
    n3327,
    n2149,
    n3013,
    n2173,
    n3116
  );


  nor
  g3203
  (
    n3349,
    n2183,
    n3065,
    n3083,
    n3073
  );


  nor
  g3204
  (
    n3498,
    n3014,
    n2076,
    n2077,
    n3141
  );


  nand
  g3205
  (
    n3459,
    n2160,
    n2111,
    n3092,
    n2994
  );


  or
  g3206
  (
    n3567,
    n2143,
    n2124,
    n2995,
    n2993
  );


  nor
  g3207
  (
    n3465,
    n3093,
    n3160,
    n2071,
    n3051
  );


  or
  g3208
  (
    n3235,
    n3087,
    n3152,
    n3124,
    n2160
  );


  xor
  g3209
  (
    n3519,
    n2977,
    n2163,
    n2068,
    n2137
  );


  nand
  g3210
  (
    n3603,
    n2150,
    n2092,
    n3096,
    n2078
  );


  nand
  g3211
  (
    n3472,
    n3139,
    n3035,
    n2063,
    n3089
  );


  or
  g3212
  (
    n3225,
    n2193,
    n2107,
    n3140,
    n3129
  );


  nand
  g3213
  (
    n3453,
    n3144,
    n3100,
    n2212,
    n2119
  );


  nor
  g3214
  (
    n3534,
    n2062,
    n3117,
    n3151,
    n3167
  );


  xnor
  g3215
  (
    n3298,
    n3069,
    n3023,
    n2194,
    n2170
  );


  and
  g3216
  (
    n3536,
    n3099,
    n2145,
    n2154,
    n2210
  );


  or
  g3217
  (
    n3264,
    n3132,
    n3035,
    n2989,
    n3028
  );


  xnor
  g3218
  (
    n3321,
    n3033,
    n2093,
    n2191,
    n2184
  );


  xnor
  g3219
  (
    n3185,
    n3074,
    n3128,
    n3019,
    n2101
  );


  xor
  g3220
  (
    n3555,
    n3047,
    n3129,
    n2070,
    n2175
  );


  nor
  g3221
  (
    n3375,
    n2154,
    n2069,
    n2231,
    n3159
  );


  xnor
  g3222
  (
    n3268,
    n2205,
    n2089,
    n3144,
    n2153
  );


  xor
  g3223
  (
    n3383,
    n2083,
    n3102,
    n3060,
    n2214
  );


  xor
  g3224
  (
    n3433,
    n2228,
    n2952,
    n2951,
    n2134
  );


  xnor
  g3225
  (
    n3290,
    n2066,
    n2971,
    n2151,
    n2122
  );


  nor
  g3226
  (
    n3420,
    n2048,
    n2206,
    n2200,
    n2150
  );


  nand
  g3227
  (
    n3310,
    n2157,
    n2219,
    n3040,
    n3052
  );


  xnor
  g3228
  (
    n3585,
    n3134,
    n3146,
    n3097,
    n3057
  );


  or
  g3229
  (
    n3488,
    n2052,
    n3114,
    n2146,
    n3005
  );


  nor
  g3230
  (
    n3605,
    n2234,
    n3110,
    n2192,
    n2227
  );


  xor
  g3231
  (
    n3543,
    n2057,
    n3010,
    n2088,
    n2062
  );


  or
  g3232
  (
    n3508,
    n2072,
    n3149,
    n3087,
    n3074
  );


  xnor
  g3233
  (
    n3426,
    n3137,
    n3153,
    n2982,
    n2231
  );


  xor
  g3234
  (
    n3416,
    n2057,
    n2157,
    n3018,
    n2201
  );


  nor
  g3235
  (
    n3410,
    n3000,
    n2059,
    n3070,
    n3038
  );


  and
  g3236
  (
    n3588,
    n2223,
    n2124,
    n3127,
    n3082
  );


  nand
  g3237
  (
    n3184,
    n3155,
    n2983,
    n2170,
    n2076
  );


  xor
  g3238
  (
    n3366,
    n3155,
    n2118,
    n3004,
    n3092
  );


  nand
  g3239
  (
    n3556,
    n3011,
    n3093,
    n2073,
    n3136
  );


  or
  g3240
  (
    n3182,
    n2112,
    n2147,
    n3044,
    n2218
  );


  and
  g3241
  (
    n3391,
    n2155,
    n2131,
    n2215,
    n2085
  );


  nor
  g3242
  (
    n3428,
    n2055,
    n2156,
    n3041,
    n3037
  );


  xor
  g3243
  (
    n3476,
    n3114,
    n2183,
    n2961,
    n2139
  );


  nand
  g3244
  (
    n3210,
    n3131,
    n3150,
    n3066,
    n3142
  );


  and
  g3245
  (
    n3568,
    n3063,
    n2989,
    n3137,
    n2990
  );


  nor
  g3246
  (
    n3271,
    n2992,
    n3084,
    n3153,
    n2154
  );


  xnor
  g3247
  (
    n3292,
    n2067,
    n3130,
    n2164,
    n3137
  );


  nor
  g3248
  (
    n3221,
    n2086,
    n3105,
    n2211,
    n2116
  );


  nand
  g3249
  (
    n3546,
    n2120,
    n2133,
    n2106,
    n2997
  );


  xor
  g3250
  (
    n3579,
    n2064,
    n2097,
    n2963,
    n2115
  );


  or
  g3251
  (
    n3191,
    n2229,
    n2213,
    n3032,
    n3099
  );


  xnor
  g3252
  (
    n3339,
    n2134,
    n2067,
    n3058,
    n3138
  );


  and
  g3253
  (
    n3582,
    n2121,
    n2096,
    n2063,
    n3058
  );


  xnor
  g3254
  (
    n3441,
    n3045,
    n2972,
    n2159,
    n2046
  );


  xnor
  g3255
  (
    n3477,
    n2173,
    n3101,
    n3116,
    n2147
  );


  nor
  g3256
  (
    n3539,
    n2204,
    n3073,
    n3143,
    n3095
  );


  xor
  g3257
  (
    n3545,
    n2206,
    n2954,
    n3022,
    n2995
  );


  xnor
  g3258
  (
    n3380,
    n3011,
    n3052,
    n2968,
    n2127
  );


  xnor
  g3259
  (
    n3286,
    n2127,
    n2162,
    n2192,
    n3072
  );


  xnor
  g3260
  (
    n3295,
    n2117,
    n3122,
    n2217,
    n2228
  );


  or
  g3261
  (
    n3212,
    n3030,
    n2203,
    n2122,
    n3098
  );


  and
  g3262
  (
    n3576,
    n2992,
    n2970,
    n2096,
    n2224
  );


  xor
  g3263
  (
    n3345,
    n2234,
    n3059,
    n3045,
    n3096
  );


  nand
  g3264
  (
    n3564,
    n2083,
    n2211,
    n3000,
    n3018
  );


  and
  g3265
  (
    n3373,
    n3050,
    n3081,
    n3114,
    n3147
  );


  or
  g3266
  (
    n3200,
    n2190,
    n2127,
    n3006,
    n2233
  );


  xnor
  g3267
  (
    n3434,
    n3008,
    n2092,
    n2141,
    n2121
  );


  and
  g3268
  (
    n3276,
    n2978,
    n3076,
    n3001,
    n3094
  );


  xor
  g3269
  (
    n3293,
    n2067,
    n3036,
    n2128,
    n2980
  );


  and
  g3270
  (
    n3474,
    n2988,
    n3123,
    n2061,
    n2126
  );


  xor
  g3271
  (
    n3283,
    n2082,
    n2078,
    n2096,
    n2181
  );


  or
  g3272
  (
    n3418,
    n2211,
    n3163,
    n2187,
    n3025
  );


  nor
  g3273
  (
    n3540,
    n2097,
    n3029,
    n2185,
    n2224
  );


  or
  g3274
  (
    n3394,
    n2991,
    n2985,
    n2965,
    n2975
  );


  xor
  g3275
  (
    n3354,
    n2047,
    n2991,
    n2146,
    n3143
  );


  xnor
  g3276
  (
    n3178,
    n3013,
    n3104,
    n3043,
    n3091
  );


  nor
  g3277
  (
    n3388,
    n2087,
    n3152,
    n2984,
    n2977
  );


  nor
  g3278
  (
    n3204,
    n2109,
    n3127,
    n2989,
    n2999
  );


  nand
  g3279
  (
    n3487,
    n2157,
    n3154,
    n2226,
    n2050
  );


  xor
  g3280
  (
    n3466,
    n3157,
    n2075,
    n2109,
    n3088
  );


  nand
  g3281
  (
    n3311,
    n3122,
    n2189,
    n3014,
    n2979
  );


  nand
  g3282
  (
    n3413,
    n2075,
    n2181,
    n3027,
    n3166
  );


  or
  g3283
  (
    n3213,
    n2103,
    n2174,
    n2048,
    n2168
  );


  xor
  g3284
  (
    n3219,
    n3122,
    n3001,
    n2981,
    n3050
  );


  xnor
  g3285
  (
    n3587,
    n3015,
    n3078,
    n3034,
    n2069
  );


  nand
  g3286
  (
    n3520,
    n2137,
    n2218,
    n2101,
    n2070
  );


  xor
  g3287
  (
    n3201,
    n3135,
    n2091,
    n2202,
    n2189
  );


  nand
  g3288
  (
    n3440,
    n3087,
    n3087,
    n3061,
    n3053
  );


  xnor
  g3289
  (
    n3217,
    n2975,
    n2162,
    n2177,
    n3022
  );


  and
  g3290
  (
    n3246,
    n3015,
    n2115,
    n2120,
    n3065
  );


  nor
  g3291
  (
    n3351,
    n2121,
    n2205,
    n3045,
    n2235
  );


  and
  g3292
  (
    n3319,
    n2136,
    n2957,
    n2196,
    n2087
  );


  nand
  g3293
  (
    n3256,
    n3091,
    n2113,
    n3025
  );


  nand
  g3294
  (
    n3456,
    n2208,
    n3048,
    n2197,
    n2155
  );


  or
  g3295
  (
    n3505,
    n2074,
    n2102,
    n3100,
    n3156
  );


  or
  g3296
  (
    n3419,
    n3090,
    n2074,
    n2156,
    n3077
  );


  and
  g3297
  (
    n3553,
    n2221,
    n2195,
    n2087,
    n2107
  );


  xor
  g3298
  (
    n3390,
    n2092,
    n2171,
    n3090,
    n2164
  );


  xor
  g3299
  (
    n3565,
    n2094,
    n3040,
    n2206,
    n3032
  );


  or
  g3300
  (
    n3377,
    n2153,
    n3100,
    n2985,
    n2194
  );


  nand
  g3301
  (
    n3360,
    n2144,
    n3043,
    n2133,
    n3103
  );


  nand
  g3302
  (
    n3289,
    n2983,
    n3018,
    n2188,
    n3009
  );


  or
  g3303
  (
    n3382,
    n2233,
    n2126,
    n3049,
    n2079
  );


  xor
  g3304
  (
    n3356,
    n2201,
    n2232,
    n2969,
    n3070
  );


  nor
  g3305
  (
    n3412,
    n2055,
    n2078,
    n2995,
    n2227
  );


  nand
  g3306
  (
    n3535,
    n3030,
    n2233,
    n2145,
    n2985
  );


  nor
  g3307
  (
    n3439,
    n3142,
    n2220,
    n3105,
    n3101
  );


  nand
  g3308
  (
    n3262,
    n2110,
    n3146,
    n2058,
    n2198
  );


  xnor
  g3309
  (
    n3411,
    n2132,
    n3066,
    n2175,
    n3091
  );


  nor
  g3310
  (
    n3423,
    n3121,
    n2100,
    n2132,
    n3060
  );


  xor
  g3311
  (
    n3340,
    n2111,
    n2118,
    n2190,
    n2081
  );


  or
  g3312
  (
    n3469,
    n3110,
    n2106,
    n3074,
    n3014
  );


  xnor
  g3313
  (
    n3260,
    n2052,
    n2047,
    n2178,
    n3048
  );


  nand
  g3314
  (
    n3591,
    n3152,
    n2058,
    n2199,
    n2966
  );


  xnor
  g3315
  (
    n3338,
    n3130,
    n2175,
    n2988,
    n2181
  );


  or
  g3316
  (
    n3503,
    n2179,
    n3047,
    n2202,
    n3080
  );


  and
  g3317
  (
    n3482,
    n3049,
    n3126,
    n3047,
    n2061
  );


  and
  g3318
  (
    n3518,
    n3142,
    n3075,
    n2143,
    n2960
  );


  nand
  g3319
  (
    n3180,
    n2131,
    n3024,
    n2142,
    n3079
  );


  nor
  g3320
  (
    n3496,
    n3119,
    n2083,
    n3024,
    n3167
  );


  nand
  g3321
  (
    n3357,
    n2049,
    n2127,
    n2073,
    n3107
  );


  or
  g3322
  (
    n3497,
    n2143,
    n3000,
    n2065,
    n2082
  );


  nor
  g3323
  (
    n3492,
    n2192,
    n2968,
    n3006,
    n2174
  );


  xor
  g3324
  (
    n3606,
    n3147,
    n3086,
    n3163,
    n2135
  );


  or
  g3325
  (
    n3563,
    n2169,
    n2225,
    n2083,
    n2182
  );


  xnor
  g3326
  (
    n3248,
    n2141,
    n3076,
    n2106,
    n3068
  );


  xor
  g3327
  (
    n3288,
    n3150,
    n2991,
    n3155,
    n3120
  );


  nor
  g3328
  (
    n3430,
    n2052,
    n3084,
    n3062,
    n3146
  );


  nand
  g3329
  (
    n3601,
    n3048,
    n3095,
    n2228,
    n2152
  );


  xor
  g3330
  (
    n3247,
    n2955,
    n2176,
    n2123,
    n3102
  );


  xor
  g3331
  (
    n3208,
    n3016,
    n2985,
    n2224,
    n2144
  );


  xnor
  g3332
  (
    n3562,
    n3140,
    n2225,
    n2074,
    n3061
  );


  or
  g3333
  (
    n3572,
    n2203,
    n3156,
    n2071,
    n3165
  );


  and
  g3334
  (
    n3250,
    n2184,
    n2984,
    n2065,
    n2123
  );


  xnor
  g3335
  (
    n3192,
    n3085,
    n3020,
    n2090,
    n2110
  );


  nor
  g3336
  (
    n3551,
    n2225,
    n3055,
    n2986,
    n3025
  );


  or
  g3337
  (
    n3303,
    n2106,
    n2967,
    n3067,
    n3160
  );


  xor
  g3338
  (
    n3280,
    n2198,
    n2216,
    n3003,
    n2223
  );


  nor
  g3339
  (
    n3527,
    n3102,
    n2184,
    n2197,
    n3144
  );


  xor
  g3340
  (
    n3595,
    n2053,
    n2974,
    n3064,
    n3148
  );


  xnor
  g3341
  (
    n3532,
    n3094,
    n3158,
    n2168,
    n3128
  );


  nor
  g3342
  (
    n3341,
    n2219,
    n2195,
    n2175,
    n2126
  );


  or
  g3343
  (
    n3218,
    n3054,
    n2969,
    n3091,
    n2216
  );


  xnor
  g3344
  (
    n3387,
    n3168,
    n2211,
    n3122,
    n3123
  );


  nand
  g3345
  (
    n3424,
    n2124,
    n2120,
    n3057,
    n2046
  );


  nand
  g3346
  (
    n3350,
    n3063,
    n3121,
    n3152,
    n2095
  );


  and
  g3347
  (
    n3446,
    n2129,
    n2208,
    n2105,
    n3116
  );


  and
  g3348
  (
    n3232,
    n3140,
    n2205,
    n3028,
    n2125
  );


  xor
  g3349
  (
    n3245,
    n3160,
    n2161,
    n3054,
    n3097
  );


  nor
  g3350
  (
    n3187,
    n3039,
    n2987,
    n3053,
    n3017
  );


  xor
  g3351
  (
    n3305,
    n2179,
    n2980,
    n3019,
    n2999
  );


  and
  g3352
  (
    n3526,
    n2084,
    n3106,
    n3163,
    n3125
  );


  and
  g3353
  (
    n3176,
    n2198,
    n3119,
    n2976,
    n2135
  );


  and
  g3354
  (
    n3244,
    n2222,
    n2984,
    n2052,
    n3082
  );


  xor
  g3355
  (
    n3226,
    n2986,
    n2060,
    n2123,
    n2071
  );


  xor
  g3356
  (
    n3330,
    n2071,
    n2148,
    n3075,
    n2080
  );


  xor
  g3357
  (
    n3175,
    n2159,
    n2222,
    n3023,
    n2080
  );


  xnor
  g3358
  (
    n3442,
    n2196,
    n2975,
    n3141,
    n2079
  );


  nand
  g3359
  (
    n3598,
    n2084,
    n2200,
    n2994,
    n3071
  );


  nor
  g3360
  (
    n3344,
    n2172,
    n2236,
    n3051,
    n3028
  );


  xor
  g3361
  (
    n3379,
    n2122,
    n3127,
    n2997,
    n2063
  );


  xor
  g3362
  (
    n3353,
    n3037,
    n3107,
    n2176,
    n3079
  );


  xnor
  g3363
  (
    n3542,
    n3106,
    n2097,
    n2234,
    n2994
  );


  xor
  g3364
  (
    n3486,
    n3150,
    n2188,
    n2172,
    n2140
  );


  xnor
  g3365
  (
    n3177,
    n2190,
    n2226,
    n2177,
    n2092
  );


  and
  g3366
  (
    n3241,
    n2167,
    n2134,
    n2215,
    n3096
  );


  xnor
  g3367
  (
    n3389,
    n2098,
    n2190,
    n3158,
    n2069
  );


  nor
  g3368
  (
    n3277,
    n2226,
    n2137,
    n2142
  );


  xor
  g3369
  (
    n3236,
    n2059,
    n3133,
    n3108,
    n2133
  );


  nand
  g3370
  (
    n3365,
    n2172,
    n2157,
    n2093,
    n2967
  );


  xor
  g3371
  (
    n3189,
    n2191,
    n3058,
    n3027,
    n2216
  );


  nor
  g3372
  (
    n3223,
    n3060,
    n2163,
    n3034,
    n3043
  );


  or
  g3373
  (
    n3179,
    n2076,
    n3102,
    n3112,
    n3166
  );


  and
  g3374
  (
    n3452,
    n2170,
    n2077,
    n2200,
    n3052
  );


  and
  g3375
  (
    n3194,
    n3029,
    n2978,
    n2141,
    n2072
  );


  xor
  g3376
  (
    n3266,
    n2996,
    n2981,
    n2113,
    n3072
  );


  nor
  g3377
  (
    n3368,
    n3110,
    n2144,
    n3004,
    n2065
  );


  xor
  g3378
  (
    n3450,
    n2174,
    n2200,
    n3151,
    n3005
  );


  xor
  g3379
  (
    n3425,
    n3031,
    n3109,
    n2213,
    n2178
  );


  xnor
  g3380
  (
    n3228,
    n2085,
    n2104,
    n3090,
    n3138
  );


  xnor
  g3381
  (
    n3550,
    n2210,
    n2213,
    n3035,
    n2165
  );


  or
  g3382
  (
    n3485,
    n2139,
    n2199,
    n2118,
    n3028
  );


  nand
  g3383
  (
    n3279,
    n2159,
    n2981,
    n3008,
    n3121
  );


  xor
  g3384
  (
    n3322,
    n2197,
    n3084,
    n3080,
    n2993
  );


  nor
  g3385
  (
    n3399,
    n3056,
    n2100,
    n3013,
    n2197
  );


  nand
  g3386
  (
    n3346,
    n2993,
    n2144,
    n3016,
    n2992
  );


  nand
  g3387
  (
    n3602,
    n2172,
    n3044,
    n2067,
    n3051
  );


  xor
  g3388
  (
    n3318,
    n3158,
    n3071,
    n3023,
    n3106
  );


  nor
  g3389
  (
    n3337,
    n3060,
    n2123,
    n3017,
    n2980
  );


  or
  g3390
  (
    n3538,
    n2980,
    n3062,
    n3111,
    n2231
  );


  or
  g3391
  (
    n3335,
    n2109,
    n2196,
    n2084,
    n2166
  );


  xor
  g3392
  (
    n3363,
    n3120,
    n2204,
    n2163,
    n2990
  );


  nand
  g3393
  (
    n3610,
    n3162,
    n3005,
    n2081,
    n3016
  );


  xor
  g3394
  (
    n3237,
    n2089,
    n3097,
    n2215,
    n2060
  );


  or
  g3395
  (
    n3265,
    n2102,
    n2073,
    n3092,
    n2066
  );


  xnor
  g3396
  (
    n3336,
    n3118,
    n2227,
    n2058,
    n3109
  );


  xor
  g3397
  (
    n3592,
    n3126,
    n3123,
    n3148,
    n2176
  );


  nand
  g3398
  (
    n3401,
    n2132,
    n2971,
    n3003,
    n2164
  );


  nor
  g3399
  (
    n3196,
    n3041,
    n2136,
    n2130,
    n2114
  );


  xnor
  g3400
  (
    n3300,
    n2090,
    n3017,
    n2148,
    n2158
  );


  nand
  g3401
  (
    n3299,
    n2191,
    n3069,
    n3057,
    n3036
  );


  and
  g3402
  (
    n3502,
    n3053,
    n3115,
    n2138,
    n3066
  );


  nand
  g3403
  (
    n3443,
    n2974,
    n3147,
    n2107,
    n3159
  );


  xnor
  g3404
  (
    n3415,
    n2992,
    n3089,
    n3149,
    n3073
  );


  or
  g3405
  (
    n3541,
    n3128,
    n3065,
    n3115,
    n3079
  );


  xor
  g3406
  (
    n3255,
    n2166,
    n3154,
    n3002,
    n2051
  );


  nor
  g3407
  (
    n3275,
    n2103,
    n2224,
    n2117,
    n2047
  );


  xnor
  g3408
  (
    n3359,
    n3097,
    n2977,
    n2132,
    n3165
  );


  xor
  g3409
  (
    n3481,
    n3138,
    n2964,
    n3133,
    n2986
  );


  nor
  g3410
  (
    n3557,
    n2150,
    n3044,
    n2097,
    n3103
  );


  xnor
  g3411
  (
    n3229,
    n3070,
    n3117,
    n2070,
    n2056
  );


  xnor
  g3412
  (
    n3522,
    n2959,
    n3064,
    n3132,
    n2230
  );


  or
  g3413
  (
    n3205,
    n2122,
    n3099,
    n3100,
    n3001
  );


  and
  g3414
  (
    n3521,
    n2998,
    n2119,
    n2178,
    n2997
  );


  nand
  g3415
  (
    n3364,
    n3082,
    n3039,
    n2093,
    n3010
  );


  xnor
  g3416
  (
    n3243,
    n2969,
    n3101,
    n3080,
    n2956
  );


  nor
  g3417
  (
    n3549,
    n3042,
    n2232,
    n2153,
    n2183
  );


  and
  g3418
  (
    n3561,
    n2088,
    n2085,
    n3106,
    n3047
  );


  nor
  g3419
  (
    n3405,
    n3151,
    n3124,
    n3002,
    n2166
  );


  and
  g3420
  (
    n3460,
    n2094,
    n3105,
    n3046,
    n2223
  );


  and
  g3421
  (
    n3188,
    n2064,
    n3042,
    n3024,
    n2147
  );


  or
  g3422
  (
    n3222,
    n3162,
    n3155,
    n2962,
    n2151
  );


  and
  g3423
  (
    n3435,
    n3027,
    n3008,
    n2223,
    n3135
  );


  xnor
  g3424
  (
    n3239,
    n3090,
    n3063,
    n2195,
    n3117
  );


  and
  g3425
  (
    n3537,
    n2193,
    n3078,
    n2049,
    n2116
  );


  nor
  g3426
  (
    n3581,
    n2978,
    n3020,
    n3010,
    n3165
  );


  xor
  g3427
  (
    n3457,
    n2054,
    n2152,
    n3088,
    n3011
  );


  nand
  g3428
  (
    n3569,
    n2165,
    n3089,
    n2979,
    n3072
  );


  and
  g3429
  (
    n3307,
    n2209,
    n2161,
    n2140,
    n3069
  );


  and
  g3430
  (
    n3291,
    n2108,
    n2168,
    n2114,
    n2161
  );


  or
  g3431
  (
    n3369,
    n3067,
    n2048,
    n2169,
    n3164
  );


  nor
  g3432
  (
    n3238,
    n2189,
    n2072,
    n3128,
    n3154
  );


  or
  g3433
  (
    n3328,
    n2991,
    n3120,
    n2094,
    n2987
  );


  nand
  g3434
  (
    n3583,
    n2176,
    n3038,
    n3160,
    n2114
  );


  xnor
  g3435
  (
    n3429,
    n2972,
    n3018,
    n3129,
    n3017
  );


  nand
  g3436
  (
    n3575,
    n2219,
    n2098,
    n2177,
    n2142
  );


  nor
  g3437
  (
    n3507,
    n3084,
    n2119,
    n2203,
    n3026
  );


  nor
  g3438
  (
    n3371,
    n3103,
    n2160,
    n3022,
    n2103
  );


  xor
  g3439
  (
    n3580,
    n3036,
    n3158,
    n3086,
    n3042
  );


  and
  g3440
  (
    n3400,
    n3033,
    n2180,
    n3059,
    n2979
  );


  or
  g3441
  (
    n3397,
    n3139,
    n3074,
    n3049,
    n3110
  );


  nor
  g3442
  (
    n3259,
    n3093,
    n3067,
    n3124,
    n2136
  );


  nand
  g3443
  (
    n3198,
    n2229,
    n3085,
    n3029,
    n2233
  );


  xor
  g3444
  (
    n3489,
    n3055,
    n3125,
    n2171,
    n2220
  );


  nor
  g3445
  (
    n3529,
    n2188,
    n2209,
    n2218,
    n3002
  );


  nor
  g3446
  (
    n3523,
    n3007,
    n2138,
    n3139,
    n2171
  );


  nand
  g3447
  (
    n3384,
    n2095,
    n3117,
    n3118,
    n2982
  );


  or
  g3448
  (
    n3408,
    n3111,
    n3009,
    n2051,
    n2165
  );


  or
  g3449
  (
    n3325,
    n2072,
    n2131,
    n2138,
    n2968
  );


  xor
  g3450
  (
    n3361,
    n2152,
    n2117,
    n2120,
    n3166
  );


  nand
  g3451
  (
    n3252,
    n2113,
    n3118,
    n2159,
    n2180
  );


  or
  g3452
  (
    n3554,
    n3095,
    n2107,
    n2170,
    n3044
  );


  nor
  g3453
  (
    n3274,
    n3112,
    n2201,
    n2050,
    n2193
  );


  nor
  g3454
  (
    n3517,
    n2080,
    n2970,
    n2094,
    n2126
  );


  nand
  g3455
  (
    n3491,
    n3161,
    n3133,
    n3046,
    n3041
  );


  nand
  g3456
  (
    n3406,
    n2102,
    n3154,
    n3056,
    n3126
  );


  xor
  g3457
  (
    n3594,
    n3118,
    n2158,
    n2125,
    n2994
  );


  and
  g3458
  (
    n3417,
    n2202,
    n2046,
    n3051,
    n3161
  );


  or
  g3459
  (
    n3372,
    n2167,
    n2060,
    n2080,
    n3071
  );


  or
  g3460
  (
    n3467,
    n2212,
    n3104,
    n3159,
    n2973
  );


  or
  g3461
  (
    n3461,
    n2192,
    n2073,
    n2152,
    n2130
  );


  nor
  g3462
  (
    n3479,
    n2145,
    n2112,
    n3040,
    n2217
  );


  or
  g3463
  (
    n3302,
    n2079,
    n3083,
    n2148,
    n3114
  );


  xnor
  g3464
  (
    n3533,
    n3157,
    n2953,
    n2139,
    n2207
  );


  and
  g3465
  (
    n3181,
    n2212,
    n2112,
    n2062,
    n2183
  );


  nor
  g3466
  (
    n3560,
    n2974,
    n2105,
    n2158,
    n3078
  );


  nand
  g3467
  (
    n3251,
    n2151,
    n2968,
    n2131,
    n3002
  );


  xnor
  g3468
  (
    n3211,
    n3061,
    n3111,
    n2216,
    n2199
  );


  xor
  g3469
  (
    n3577,
    n2165,
    n2138,
    n2978,
    n2054
  );


  nor
  g3470
  (
    n3438,
    n2182,
    n3141,
    n2099,
    n3023
  );


  or
  g3471
  (
    n3547,
    n2983,
    n2050,
    n3046,
    n2990
  );


  or
  g3472
  (
    n3597,
    n2220,
    n3068,
    n3040,
    n3056
  );


  xnor
  g3473
  (
    n3263,
    n3045,
    n2112,
    n3113,
    n2104
  );


  nand
  g3474
  (
    n3455,
    n3161,
    n3081,
    n2207,
    n3012
  );


  nor
  g3475
  (
    n3206,
    n2056,
    n3101,
    n2221,
    n3116
  );


  and
  g3476
  (
    n3432,
    n2088,
    n2104,
    n3148,
    n2109
  );


  xnor
  g3477
  (
    n3427,
    n2156,
    n2089,
    n2093,
    n3076
  );


  nand
  g3478
  (
    n3278,
    n3093,
    n2125,
    n3003,
    n2210
  );


  and
  g3479
  (
    n3600,
    n2180,
    n3111,
    n3004,
    n2229
  );


  nor
  g3480
  (
    n3490,
    n3024,
    n3112,
    n2116,
    n3133
  );


  nor
  g3481
  (
    n3552,
    n2226,
    n2181,
    n2186,
    n3161
  );


  or
  g3482
  (
    n3448,
    n2099,
    n2207,
    n2973,
    n3107
  );


  or
  g3483
  (
    n3593,
    n3013,
    n3108,
    n3126,
    n3012
  );


  or
  g3484
  (
    n3234,
    n2088,
    n3135,
    n2177,
    n2058
  );


  nor
  g3485
  (
    n3386,
    n3104,
    n2182,
    n2049,
    n2188
  );


  and
  g3486
  (
    n3282,
    n2998,
    n2098,
    n3033,
    n3038
  );


  or
  g3487
  (
    n3195,
    n2151,
    n2104,
    n3088,
    n2231
  );


  and
  g3488
  (
    n3445,
    n2185,
    n2193,
    n2982,
    n2206
  );


  xnor
  g3489
  (
    n3190,
    n2075,
    n3066,
    n3004,
    n3166
  );


  nand
  g3490
  (
    n3301,
    n2199,
    n2084,
    n2984,
    n2971
  );


  xor
  g3491
  (
    n3270,
    n3149,
    n3059,
    n2998,
    n3033
  );


  xor
  g3492
  (
    n3437,
    n2986,
    n2075,
    n2077,
    n2134
  );


  xor
  g3493
  (
    n3392,
    n3108,
    n2105,
    n2221,
    n3153
  );


  or
  g3494
  (
    n3199,
    n2095,
    n2160,
    n3135,
    n2970
  );


  nor
  g3495
  (
    n3329,
    n2155,
    n3031,
    n3164,
    n2230
  );


  and
  g3496
  (
    n3525,
    n2218,
    n3147,
    n2214,
    n2082
  );


  xnor
  g3497
  (
    n3495,
    n3039,
    n2230,
    n2069,
    n2079
  );


  nor
  g3498
  (
    n3249,
    n3137,
    n3080,
    n2091,
    n2051
  );


  or
  g3499
  (
    n3370,
    n2115,
    n2204,
    n2077,
    n2198
  );


  and
  g3500
  (
    n3306,
    n2227,
    n2204,
    n3156,
    n2988
  );


  nand
  g3501
  (
    n3528,
    n2185,
    n3089,
    n3061,
    n3131
  );


  xnor
  g3502
  (
    n3186,
    n3048,
    n3014,
    n3145,
    n3105
  );


  and
  g3503
  (
    n3347,
    n2228,
    n2987,
    n3011,
    n3113
  );


  nand
  g3504
  (
    n3258,
    n2057,
    n2212,
    n3115,
    n2087
  );


  and
  g3505
  (
    n3499,
    n3083,
    n3162,
    n3130,
    n3050
  );


  or
  g3506
  (
    n3447,
    n2208,
    n3006,
    n2207,
    n2090
  );


  nand
  g3507
  (
    n3494,
    n2971,
    n2220,
    n3153,
    n2163
  );


  or
  g3508
  (
    n3281,
    n3143,
    n3104,
    n2161,
    n3008
  );


  xnor
  g3509
  (
    n3573,
    n3131,
    n2054,
    n2056,
    n3134
  );


  nor
  g3510
  (
    n3444,
    n2085,
    n2149,
    n3021,
    n2164
  );


  xor
  g3511
  (
    n3269,
    n3078,
    n3094,
    n3022,
    n3142
  );


  or
  g3512
  (
    n3431,
    n2130,
    n2061,
    n3073,
    n2222
  );


  or
  g3513
  (
    n3297,
    n3064,
    n2089,
    n2987,
    n3127
  );


  and
  g3514
  (
    n3604,
    n2184,
    n2235,
    n3079,
    n2078
  );


  and
  g3515
  (
    n3559,
    n2068,
    n2191,
    n3121,
    n2113
  );


  xor
  g3516
  (
    n3227,
    n3015,
    n2053,
    n2993,
    n2205
  );


  xor
  g3517
  (
    n3462,
    n3070,
    n2140,
    n3085,
    n3019
  );


  nand
  g3518
  (
    n3183,
    n3115,
    n2182,
    n3009,
    n3108
  );


  nand
  g3519
  (
    n3436,
    n2047,
    n2110,
    n3007,
    n2136
  );


  nand
  g3520
  (
    n3471,
    n3145,
    n3000,
    n2187,
    n2995
  );


  nor
  g3521
  (
    n3193,
    n2973,
    n3054,
    n2110,
    n2187
  );


  xnor
  g3522
  (
    n3531,
    n2235,
    n3163,
    n2209,
    n2150
  );


  xnor
  g3523
  (
    n3484,
    n3125,
    n3082,
    n3032,
    n2121
  );


  xnor
  g3524
  (
    n3513,
    n3026,
    n3055,
    n2194,
    n2169
  );


  or
  g3525
  (
    n3590,
    n3026,
    n2119,
    n2128,
    n2976
  );


  or
  g3526
  (
    n3257,
    n2162,
    n2124,
    n3130,
    n2999
  );


  xor
  g3527
  (
    n3589,
    n2095,
    n3146,
    n2066,
    n3059
  );


  and
  g3528
  (
    n3273,
    n3132,
    n2064,
    n2086,
    n3098
  );


  nand
  g3529
  (
    n3402,
    n3164,
    n2108,
    n2229,
    n2099
  );


  and
  g3530
  (
    n3470,
    n3096,
    n3026,
    n3123,
    n2186
  );


  nand
  g3531
  (
    n3530,
    n2158,
    n2975,
    n2057,
    n3006
  );


  xnor
  g3532
  (
    n3220,
    n2969,
    n2117,
    n2129,
    n3020
  );


  xnor
  g3533
  (
    n3287,
    n3036,
    n2171,
    n3088,
    n3112
  );


  nor
  g3534
  (
    n3385,
    n3167,
    n3145,
    n3077,
    n2081
  );


  and
  g3535
  (
    n3312,
    n2185,
    n2187,
    n2146,
    n2180
  );


  xnor
  g3536
  (
    n3272,
    n2130,
    n2111,
    n3167,
    n3150
  );


  nand
  g3537
  (
    n3506,
    n2111,
    n3092,
    n3039,
    n2133
  );


  and
  g3538
  (
    n3396,
    n3049,
    n3136,
    n3107,
    n2983
  );


  xnor
  g3539
  (
    n3454,
    n3095,
    n3038,
    n2149,
    n2179
  );


  nand
  g3540
  (
    n3326,
    n3046,
    n3075,
    n3098,
    n2148
  );


  xnor
  g3541
  (
    n3316,
    n3054,
    n3098,
    n3037,
    n2996
  );


  nor
  g3542
  (
    n3574,
    n2068,
    n2162,
    n2101,
    n2154
  );


  xnor
  g3543
  (
    n3596,
    n2988,
    n2156,
    n2145,
    n3144
  );


  nor
  g3544
  (
    n3308,
    n3012,
    n2070,
    n2234,
    n3029
  );


  xnor
  g3545
  (
    n3240,
    n2108,
    n2056,
    n2129,
    n2143
  );


  and
  g3546
  (
    n3609,
    n3062,
    n3030,
    n2173,
    n3136
  );


  or
  g3547
  (
    n3378,
    n2202,
    n2054,
    n2189,
    n2155
  );


  and
  g3548
  (
    n3233,
    n2167,
    n2982,
    n2059,
    n3003
  );


  and
  g3549
  (
    n3544,
    n2958,
    n3113,
    n3007,
    n2972
  );


  xnor
  g3550
  (
    n3473,
    n2168,
    n2970,
    n2051,
    n2221
  );


  and
  g3551
  (
    n3224,
    n2210,
    n2068,
    n3120,
    n2186
  );


  and
  g3552
  (
    n3324,
    n2055,
    n2186,
    n3077
  );


  xor
  g3553
  (
    n3483,
    n3109,
    n3019,
    n3124,
    n3075
  );


  or
  g3554
  (
    n3414,
    n2979,
    n2178,
    n2139,
    n3069
  );


  nand
  g3555
  (
    n3409,
    n3042,
    n2196,
    n3081,
    n2996
  );


  nor
  g3556
  (
    n3599,
    n2217,
    n2090,
    n3064,
    n3012
  );


  nor
  g3557
  (
    n3332,
    n3157,
    n2100,
    n2135,
    n3085
  );


  or
  g3558
  (
    n3512,
    n2213,
    n2208,
    n2167,
    n3052
  );


  nand
  g3559
  (
    n3422,
    n2179,
    n3136,
    n2128,
    n2125
  );


  nor
  g3560
  (
    n3207,
    n2215,
    n2203,
    n3067,
    n2149
  );


  or
  g3561
  (
    n3334,
    n2990,
    n2201,
    n3034,
    n3164
  );


  nand
  g3562
  (
    n3362,
    n3021,
    n3086,
    n2129,
    n3076
  );


  xor
  g3563
  (
    n3323,
    n3099,
    n3035,
    n3065,
    n2235
  );


  and
  g3564
  (
    n3607,
    n2147,
    n2146,
    n2232,
    n3001
  );


  nand
  g3565
  (
    n3215,
    n3057,
    n3086,
    n2081,
    n3072
  );


  xnor
  g3566
  (
    n3304,
    n2209,
    n3103,
    n2063,
    n2135
  );


  nand
  g3567
  (
    n3315,
    n2062,
    n3141,
    n2060,
    n2099
  );


  nor
  g3568
  (
    n3284,
    n3034,
    n3138,
    n3016,
    n3021
  );


  xor
  g3569
  (
    n3515,
    n3134,
    n3156,
    n2232,
    n2096
  );


  nand
  g3570
  (
    n3296,
    n2048,
    n3094,
    n3140,
    n2989
  );


  xnor
  g3571
  (
    n3261,
    n2153,
    n2214,
    n3162,
    n3119
  );


  or
  g3572
  (
    n3358,
    n2091,
    n3037,
    n3043,
    n2116
  );


  nor
  g3573
  (
    n3230,
    n2074,
    n3165,
    n3009,
    n2194
  );


  and
  g3574
  (
    n3376,
    n2141,
    n2098,
    n2214,
    n3081
  );


  xnor
  g3575
  (
    n3493,
    n3055,
    n3005,
    n3149,
    n3021
  );


  xnor
  g3576
  (
    n3475,
    n2977,
    n3145,
    n3027,
    n2115
  );


  nor
  g3577
  (
    n3203,
    n3132,
    n3119,
    n2976,
    n3053
  );


  and
  g3578
  (
    n3625,
    n3210,
    n3208,
    n3268,
    n3195
  );


  nor
  g3579
  (
    n3622,
    n3206,
    n3272,
    n3191,
    n3277
  );


  xnor
  g3580
  (
    n3611,
    n3179,
    n3278,
    n3248,
    n3258
  );


  and
  g3581
  (
    n3633,
    n3184,
    n3225,
    n3261,
    n3181
  );


  xnor
  g3582
  (
    n3635,
    n3224,
    n3246,
    n3219,
    n3223
  );


  nor
  g3583
  (
    n3613,
    n3244,
    n3249,
    n3259,
    n3215
  );


  nor
  g3584
  (
    n3636,
    n3205,
    n3271,
    n3204,
    n3265
  );


  xnor
  g3585
  (
    n3614,
    n3243,
    n3188,
    n3187,
    n3274
  );


  nand
  g3586
  (
    n3632,
    n3209,
    n3239,
    n3254,
    n3228
  );


  xor
  g3587
  (
    n3612,
    n3260,
    n3229,
    n3202,
    n3226
  );


  xor
  g3588
  (
    n3615,
    n3197,
    n3214,
    n3250,
    n3183
  );


  nand
  g3589
  (
    n3616,
    n3247,
    n3212,
    n3270,
    n3236
  );


  xor
  g3590
  (
    n3627,
    n3255,
    n3192,
    n3177,
    n3234
  );


  or
  g3591
  (
    n3628,
    n3233,
    n3207,
    n3232,
    n3252
  );


  or
  g3592
  (
    n3634,
    n3266,
    n3273,
    n3227,
    n3267
  );


  nor
  g3593
  (
    n3617,
    n3180,
    n3237,
    n3218,
    n3264
  );


  and
  g3594
  (
    n3618,
    n3256,
    n3201,
    n3251,
    n3222
  );


  or
  g3595
  (
    n3629,
    n3245,
    n3213,
    n3230,
    n3221
  );


  or
  g3596
  (
    n3626,
    n3231,
    n3257,
    n3193,
    n3275
  );


  or
  g3597
  (
    n3621,
    n3276,
    n3211,
    n3203,
    n3240
  );


  or
  g3598
  (
    n3631,
    n3238,
    n3200,
    n3253,
    n3175
  );


  xnor
  g3599
  (
    n3620,
    n3189,
    n3241,
    n3190,
    n3196
  );


  nand
  g3600
  (
    n3623,
    n3235,
    n3176,
    n3185,
    n3269
  );


  xor
  g3601
  (
    n3624,
    n3217,
    n3220,
    n3216,
    n3182
  );


  nand
  g3602
  (
    n3630,
    n3178,
    n3186,
    n3194,
    n3198
  );


  and
  g3603
  (
    n3619,
    n3262,
    n3199,
    n3263,
    n3242
  );


  and
  g3604
  (
    n3646,
    n3614,
    n3619,
    n2836,
    n3289
  );


  nor
  g3605
  (
    n3641,
    n3622,
    n3280,
    n3625,
    n2836
  );


  and
  g3606
  (
    n3648,
    n3292,
    n3611,
    n3620,
    n2831
  );


  and
  g3607
  (
    n3647,
    n3281,
    n3287,
    n3293,
    n2830
  );


  xnor
  g3608
  (
    n3638,
    n2832,
    n2832,
    n3615,
    n2830
  );


  xor
  g3609
  (
    n3645,
    n3290,
    n2834,
    n2830,
    n3621
  );


  nand
  g3610
  (
    n3640,
    n3283,
    n3291,
    n2830,
    n3285
  );


  and
  g3611
  (
    n3651,
    n3296,
    n3618,
    n2833,
    n3616
  );


  xor
  g3612
  (
    n3642,
    n3282,
    n2834,
    n3623,
    n3612
  );


  xor
  g3613
  (
    n3643,
    n3624,
    n3294,
    n3613,
    n2833
  );


  nand
  g3614
  (
    n3639,
    n3295,
    n2832,
    n3617,
    n2835
  );


  xnor
  g3615
  (
    n3649,
    n2834,
    n2831
  );


  nand
  g3616
  (
    n3650,
    n3279,
    n2833,
    n3284
  );


  nand
  g3617
  (
    n3637,
    n3286,
    n3288,
    n2835
  );


  and
  g3618
  (
    n3644,
    n2836,
    n2834,
    n2832,
    n2835
  );


  or
  g3619
  (
    n3661,
    n3646,
    n3169,
    n2876,
    n3637
  );


  xnor
  g3620
  (
    n3657,
    n2877,
    n3650,
    n2878,
    n3169
  );


  or
  g3621
  (
    n3655,
    n2838,
    n2878,
    n2879,
    n3634
  );


  or
  g3622
  (
    n3653,
    n2838,
    n2880,
    n3645,
    n3639
  );


  and
  g3623
  (
    n3663,
    n2879,
    n3641,
    n3628,
    n3635
  );


  xnor
  g3624
  (
    n3667,
    n2877,
    n3629,
    n2837,
    n2878
  );


  and
  g3625
  (
    n3666,
    n3649,
    n3627,
    n3636,
    n3632
  );


  xor
  g3626
  (
    n3664,
    n3648,
    n3169,
    n3626,
    n3633
  );


  nor
  g3627
  (
    n3654,
    n2880,
    n2879,
    n3651,
    n3643
  );


  xnor
  g3628
  (
    n3662,
    n3168,
    n3638,
    n3630,
    n2880
  );


  and
  g3629
  (
    n3659,
    n2839,
    n3651,
    n2838,
    n2877
  );


  nor
  g3630
  (
    n3658,
    n3168,
    n2837,
    n3169
  );


  xnor
  g3631
  (
    n3656,
    n3640,
    n3170,
    n2839,
    n2880
  );


  and
  g3632
  (
    n3665,
    n2839,
    n2838,
    n3644,
    n2836
  );


  xor
  g3633
  (
    n3660,
    n2837,
    n3647,
    n2879,
    n2878
  );


  xnor
  g3634
  (
    n3652,
    n3631,
    n2877,
    n3168,
    n3642
  );


  buf
  g3635
  (
    n3671,
    n3653
  );


  not
  g3636
  (
    n3668,
    n3654
  );


  not
  g3637
  (
    n3669,
    n3655
  );


  buf
  g3638
  (
    n3670,
    n3652
  );


  and
  g3639
  (
    n3680,
    n3670,
    n3174
  );


  xnor
  g3640
  (
    n3681,
    n3173,
    n3671
  );


  nor
  g3641
  (
    n3683,
    n3670,
    n3658
  );


  xnor
  g3642
  (
    n3684,
    n3172,
    n3173
  );


  xnor
  g3643
  (
    n3678,
    n3174,
    n3661
  );


  nand
  g3644
  (
    n3674,
    n3670,
    n3662
  );


  or
  g3645
  (
    n3675,
    n3656,
    n3671,
    n3670
  );


  or
  g3646
  (
    n3672,
    n3669,
    n3668,
    n3170
  );


  nor
  g3647
  (
    n3677,
    n3171,
    n3174
  );


  buf
  g3648
  (
    n3682,
    n3171
  );


  nand
  g3649
  (
    n3685,
    n3173,
    n3172,
    n3671
  );


  nor
  g3650
  (
    n3679,
    n3669,
    n3170,
    n3657
  );


  xnor
  g3651
  (
    n3673,
    n3671,
    n3173,
    n3669
  );


  xor
  g3652
  (
    n3676,
    n3660,
    n3659,
    n3172,
    n3668
  );


  nor
  g3653
  (
    n3735,
    n3304,
    n3307,
    n3329,
    n3315
  );


  or
  g3654
  (
    n3719,
    n3357,
    n3399,
    n3402,
    n3396
  );


  xnor
  g3655
  (
    n3695,
    n3346,
    n3675,
    n3310
  );


  nor
  g3656
  (
    n3689,
    n3351,
    n3323,
    n3460,
    n3348
  );


  xnor
  g3657
  (
    n3711,
    n3672,
    n3347,
    n3445,
    n3433
  );


  xnor
  g3658
  (
    n3705,
    n3672,
    n3450,
    n3452,
    n3684
  );


  and
  g3659
  (
    n3729,
    n3308,
    n3684,
    n3377,
    n3311
  );


  or
  g3660
  (
    n3693,
    n3675,
    n3375,
    n3677,
    n3446
  );


  xnor
  g3661
  (
    n3698,
    n3674,
    n3390,
    n3327,
    n3451
  );


  and
  g3662
  (
    n3696,
    n3298,
    n3678,
    n3384,
    n3403
  );


  xnor
  g3663
  (
    n3717,
    n3673,
    n3676,
    n3313,
    n3424
  );


  nand
  g3664
  (
    n3737,
    n3317,
    n3385,
    n3414,
    n3674
  );


  or
  g3665
  (
    n3687,
    n3339,
    n3345,
    n3681,
    n3382
  );


  xor
  g3666
  (
    n3713,
    n3412,
    n3361,
    n3386,
    n3401
  );


  nand
  g3667
  (
    n3715,
    n3378,
    n3343,
    n3428,
    n3355
  );


  or
  g3668
  (
    n3726,
    n3673,
    n3359,
    n3415,
    n3417
  );


  nand
  g3669
  (
    n3736,
    n3332,
    n3350,
    n3408,
    n3391
  );


  xnor
  g3670
  (
    n3728,
    n3392,
    n3437,
    n3443,
    n3677
  );


  nand
  g3671
  (
    n3718,
    n3685,
    n3341,
    n3316,
    n3366
  );


  xor
  g3672
  (
    n3733,
    n3322,
    n3365,
    n3301,
    n3349
  );


  nand
  g3673
  (
    n3694,
    n3336,
    n3342,
    n3369,
    n3681
  );


  nor
  g3674
  (
    n3710,
    n3679,
    n3680,
    n3397,
    n3303
  );


  nor
  g3675
  (
    n3688,
    n3464,
    n3438,
    n3458,
    n3371
  );


  or
  g3676
  (
    n3707,
    n3675,
    n3679,
    n3684,
    n3368
  );


  and
  g3677
  (
    n3701,
    n3672,
    n3676,
    n3326,
    n3325
  );


  xnor
  g3678
  (
    n3716,
    n3374,
    n3425,
    n3320,
    n3448
  );


  nor
  g3679
  (
    n3691,
    n3309,
    n3683,
    n3682,
    n3459
  );


  nor
  g3680
  (
    n3731,
    n3456,
    n3362,
    n3373,
    n3440
  );


  nand
  g3681
  (
    n3708,
    n3398,
    n3422,
    n3455,
    n3370
  );


  nand
  g3682
  (
    n3686,
    n3682,
    n3683,
    n3319
  );


  or
  g3683
  (
    n3739,
    n3673,
    n3685,
    n3334,
    n3331
  );


  nand
  g3684
  (
    n3700,
    n3404,
    n3434,
    n3432,
    n3674
  );


  xor
  g3685
  (
    n3703,
    n3353,
    n3411,
    n3389,
    n3461
  );


  and
  g3686
  (
    n3723,
    n3676,
    n3676,
    n3305,
    n3388
  );


  or
  g3687
  (
    n3712,
    n3685,
    n3435,
    n3410,
    n3297
  );


  nand
  g3688
  (
    n3721,
    n3406,
    n3372,
    n3300,
    n3684
  );


  xnor
  g3689
  (
    n3738,
    n3678,
    n3354,
    n3356,
    n3430
  );


  xnor
  g3690
  (
    n3741,
    n3306,
    n3318,
    n3680,
    n3454
  );


  or
  g3691
  (
    n3702,
    n3681,
    n3395,
    n3299,
    n3427
  );


  nor
  g3692
  (
    n3725,
    n3367,
    n3441,
    n3418,
    n3423
  );


  xnor
  g3693
  (
    n3704,
    n3447,
    n3338,
    n3421,
    n3419
  );


  nand
  g3694
  (
    n3740,
    n3314,
    n3673,
    n3679,
    n3405
  );


  xor
  g3695
  (
    n3706,
    n3439,
    n3444,
    n3680,
    n3674
  );


  nor
  g3696
  (
    n3722,
    n3678,
    n3449,
    n3302,
    n3426
  );


  or
  g3697
  (
    n3709,
    n3463,
    n3364,
    n3429,
    n3677
  );


  or
  g3698
  (
    n3697,
    n3678,
    n3681,
    n3321,
    n3312
  );


  xor
  g3699
  (
    n3692,
    n3409,
    n3453,
    n3400,
    n3381
  );


  and
  g3700
  (
    n3727,
    n3407,
    n3335,
    n3376,
    n3352
  );


  nor
  g3701
  (
    n3724,
    n3677,
    n3340,
    n3683,
    n3380
  );


  nor
  g3702
  (
    n3720,
    n3379,
    n3457,
    n3363,
    n3682
  );


  or
  g3703
  (
    n3690,
    n3394,
    n3442,
    n3462,
    n3337
  );


  nor
  g3704
  (
    n3730,
    n3328,
    n3333,
    n3344,
    n3416
  );


  or
  g3705
  (
    n3714,
    n3420,
    n3358,
    n3680,
    n3393
  );


  xnor
  g3706
  (
    n3699,
    n3682,
    n3330,
    n3436,
    n3679
  );


  or
  g3707
  (
    n3734,
    n3387,
    n3431,
    n3413,
    n3383
  );


  nor
  g3708
  (
    n3732,
    n3360,
    n3672,
    n3324,
    n3685
  );


  nor
  g3709
  (
    n3762,
    n3467,
    n3692
  );


  or
  g3710
  (
    n3770,
    n3480,
    n3701
  );


  and
  g3711
  (
    n3752,
    n3486,
    n3481
  );


  or
  g3712
  (
    n3753,
    n3706,
    n3478
  );


  and
  g3713
  (
    n3745,
    n3484,
    n3713
  );


  and
  g3714
  (
    n3749,
    n3475,
    n3700
  );


  xor
  g3715
  (
    n3767,
    n3711,
    n3689
  );


  xor
  g3716
  (
    n3742,
    n3488,
    n3492
  );


  and
  g3717
  (
    n3746,
    n3482,
    n3490
  );


  or
  g3718
  (
    n3765,
    n3479,
    n3468
  );


  nand
  g3719
  (
    n3750,
    n3697,
    n3473
  );


  and
  g3720
  (
    n3764,
    n3698,
    n3710
  );


  xnor
  g3721
  (
    n3766,
    n3466,
    n3693
  );


  xor
  g3722
  (
    n3759,
    n3483,
    n3474
  );


  nor
  g3723
  (
    n3758,
    n3485,
    n3487
  );


  or
  g3724
  (
    n3744,
    n3690,
    n3703
  );


  or
  g3725
  (
    n3760,
    n3469,
    n3476
  );


  xnor
  g3726
  (
    n3755,
    n3477,
    n3687
  );


  nand
  g3727
  (
    n3761,
    n3493,
    n3707
  );


  nand
  g3728
  (
    n3748,
    n3708,
    n3704
  );


  or
  g3729
  (
    n3743,
    n3465,
    n3696
  );


  and
  g3730
  (
    n3768,
    n3705,
    n3491
  );


  or
  g3731
  (
    n3756,
    n3472,
    n3695
  );


  or
  g3732
  (
    n3769,
    n3694,
    n3699
  );


  or
  g3733
  (
    n3763,
    n3714,
    n3709
  );


  or
  g3734
  (
    n3751,
    n3688,
    n3691
  );


  xnor
  g3735
  (
    n3747,
    n3489,
    n3712
  );


  xor
  g3736
  (
    n3754,
    n3702,
    n3470
  );


  and
  g3737
  (
    n3757,
    n3686,
    n3471
  );


  not
  g3738
  (
    n3771,
    n3749
  );


  not
  g3739
  (
    n3788,
    n3750
  );


  buf
  g3740
  (
    n3782,
    n3751
  );


  buf
  g3741
  (
    n3776,
    n3746
  );


  buf
  g3742
  (
    n3785,
    n3754
  );


  buf
  g3743
  (
    n3789,
    n3752
  );


  buf
  g3744
  (
    n3775,
    n3755
  );


  not
  g3745
  (
    n3777,
    n3743
  );


  not
  g3746
  (
    n3780,
    n3715
  );


  buf
  g3747
  (
    n3772,
    n3745
  );


  not
  g3748
  (
    n3773,
    n3748
  );


  buf
  g3749
  (
    n3783,
    n3753
  );


  not
  g3750
  (
    n3779,
    n3744
  );


  not
  g3751
  (
    n3781,
    n3762
  );


  buf
  g3752
  (
    n3784,
    n3716
  );


  buf
  g3753
  (
    n3774,
    n3747
  );


  buf
  g3754
  (
    n3787,
    n3760
  );


  not
  g3755
  (
    n3786,
    n3718
  );


  nand
  g3756
  (
    n3790,
    n3717,
    n3757
  );


  and
  g3757
  (
    n3778,
    n3756,
    n3761,
    n3759,
    n3758
  );


  xnor
  g3758
  (
    n3798,
    n1639,
    n3500,
    n3775,
    n3495
  );


  nor
  g3759
  (
    n3791,
    n3775,
    n3775,
    n3510,
    n2839
  );


  or
  g3760
  (
    n3793,
    n3503,
    n3494,
    n3512,
    n3502
  );


  and
  g3761
  (
    n3795,
    n3513,
    n3501,
    n3509,
    n3498
  );


  and
  g3762
  (
    n3796,
    n3771,
    n3506,
    n3507,
    n3497
  );


  xnor
  g3763
  (
    n3794,
    n3511,
    n3772,
    n3496,
    n3508
  );


  nand
  g3764
  (
    n3792,
    n3774,
    n3499,
    n3504,
    n3773
  );


  nand
  g3765
  (
    n3797,
    n1639,
    n3505,
    n2840,
    n3775
  );


  xor
  g3766
  (
    n3809,
    n3664,
    n3798,
    n3667,
    n3721
  );


  and
  g3767
  (
    n3800,
    n3517,
    n3794,
    n3662,
    n3798
  );


  nor
  g3768
  (
    n3810,
    n3519,
    n3663,
    n3665,
    n3667
  );


  nand
  g3769
  (
    n3803,
    n3522,
    n3662,
    n3793,
    n3663
  );


  or
  g3770
  (
    n3804,
    n3666,
    n3665,
    n3514,
    n3797
  );


  xnor
  g3771
  (
    n3805,
    n3791,
    n3515,
    n3664,
    n3663
  );


  or
  g3772
  (
    n3802,
    n3798,
    n3516,
    n3664,
    n3665
  );


  xnor
  g3773
  (
    n3806,
    n3667,
    n3796,
    n3719,
    n3521
  );


  or
  g3774
  (
    n3808,
    n3664,
    n3662,
    n3663,
    n3520
  );


  xor
  g3775
  (
    n3799,
    n3797,
    n3798,
    n3792,
    n3795
  );


  or
  g3776
  (
    n3807,
    n3720,
    n3666,
    n3665,
    n3518
  );


  or
  g3777
  (
    n3801,
    n3667,
    n3523,
    n3666
  );


  nor
  g3778
  (
    n3844,
    n3524,
    n1649,
    n3808,
    n1648
  );


  nor
  g3779
  (
    n3840,
    n2236,
    n1661,
    n1659,
    n1654
  );


  nor
  g3780
  (
    n3824,
    n3803,
    n1651,
    n1648,
    n3801
  );


  nand
  g3781
  (
    n3839,
    n1651,
    n1663,
    n3810,
    n3800
  );


  or
  g3782
  (
    n3812,
    n3804,
    n1643,
    n3799,
    n3802
  );


  or
  g3783
  (
    n3832,
    n3807,
    n3799,
    n3805,
    n1668
  );


  nand
  g3784
  (
    n3841,
    n1641,
    n1639,
    n1670,
    n1644
  );


  xnor
  g3785
  (
    n3820,
    n1642,
    n1657,
    n1643,
    n1667
  );


  and
  g3786
  (
    n3850,
    n1661,
    n1645,
    n1660,
    n1664
  );


  or
  g3787
  (
    n3822,
    n1666,
    n3809,
    n3801
  );


  nor
  g3788
  (
    n3843,
    n3809,
    n1654,
    n1658,
    n1646
  );


  and
  g3789
  (
    n3811,
    n1644,
    n3806,
    n1668,
    n2238
  );


  nor
  g3790
  (
    n3854,
    n3799,
    n3800,
    n3805,
    n1642
  );


  nand
  g3791
  (
    n3846,
    n3804,
    n1651,
    n2237,
    n3805
  );


  xor
  g3792
  (
    n3817,
    n3806,
    n1655,
    n3809,
    n3802
  );


  xor
  g3793
  (
    n3842,
    n1665,
    n1665,
    n1653,
    n1649
  );


  nor
  g3794
  (
    n3829,
    n1642,
    n1661,
    n1659,
    n1652
  );


  or
  g3795
  (
    n3836,
    n2238,
    n1650,
    n1640,
    n1647
  );


  xor
  g3796
  (
    n3821,
    n3802,
    n1666,
    n1667,
    n3799
  );


  and
  g3797
  (
    n3818,
    n1662,
    n1733,
    n3800,
    n1648
  );


  or
  g3798
  (
    n3813,
    n1657,
    n1662,
    n2238,
    n1653
  );


  and
  g3799
  (
    n3849,
    n1658,
    n1664,
    n1640,
    n2237
  );


  and
  g3800
  (
    n3823,
    n1647,
    n1671,
    n1645,
    n1667
  );


  nor
  g3801
  (
    n3847,
    n1652,
    n1653,
    n1656,
    n1644
  );


  or
  g3802
  (
    n3833,
    n1646,
    n1668,
    n1652,
    n1650
  );


  and
  g3803
  (
    n3856,
    n3809,
    n1651,
    n1646,
    n1642
  );


  and
  g3804
  (
    n3845,
    n3810,
    n2238,
    n1668,
    n1649
  );


  nand
  g3805
  (
    n3857,
    n1662,
    n1659,
    n1661,
    n3808
  );


  nand
  g3806
  (
    n3826,
    n3526,
    n3804,
    n1670,
    n3807
  );


  xor
  g3807
  (
    n3830,
    n1660,
    n3801,
    n1654,
    n1647
  );


  nand
  g3808
  (
    n3816,
    n3806,
    n3808,
    n1656,
    n1660
  );


  nand
  g3809
  (
    n3825,
    n1666,
    n1645,
    n3802,
    n1663
  );


  xnor
  g3810
  (
    n3814,
    n3803,
    n3808,
    n1666,
    n2237
  );


  xnor
  g3811
  (
    n3828,
    n1640,
    n2237,
    n3805,
    n1656
  );


  xnor
  g3812
  (
    n3852,
    n3803,
    n3807,
    n1650,
    n1646
  );


  and
  g3813
  (
    n3853,
    n1660,
    n3527,
    n1640,
    n3804
  );


  xnor
  g3814
  (
    n3848,
    n1648,
    n3807,
    n3810,
    n1653
  );


  and
  g3815
  (
    n3855,
    n1670,
    n1663,
    n1641,
    n1667
  );


  or
  g3816
  (
    n3834,
    n1665,
    n1643,
    n1639,
    n1671
  );


  and
  g3817
  (
    n3831,
    n1669,
    n1657,
    n1643,
    n1656
  );


  or
  g3818
  (
    n3819,
    n1670,
    n1647,
    n1664,
    n3525
  );


  nand
  g3819
  (
    n3815,
    n1658,
    n1652,
    n1669,
    n1659
  );


  xor
  g3820
  (
    n3851,
    n1663,
    n1641,
    n1655,
    n1658
  );


  nor
  g3821
  (
    n3838,
    n1655,
    n3806,
    n1654,
    n2236
  );


  xnor
  g3822
  (
    n3858,
    n1641,
    n1644,
    n3810,
    n1665
  );


  xnor
  g3823
  (
    n3827,
    n1662,
    n1649,
    n2236,
    n1664
  );


  xnor
  g3824
  (
    n3837,
    n3800,
    n1657,
    n1669,
    n1645
  );


  nand
  g3825
  (
    n3835,
    n1655,
    n1650,
    n3803,
    n1669
  );


  and
  g3826
  (
    n3871,
    n3779,
    n3820,
    n2841,
    n3781
  );


  and
  g3827
  (
    n3863,
    n3534,
    n3780,
    n3779
  );


  xor
  g3828
  (
    n3869,
    n3811,
    n3776,
    n2841,
    n3530
  );


  and
  g3829
  (
    n3870,
    n3777,
    n3782,
    n3813,
    n3536
  );


  nand
  g3830
  (
    n3872,
    n2842,
    n3779,
    n2840
  );


  xnor
  g3831
  (
    n3861,
    n3781,
    n3777,
    n3532,
    n3528
  );


  nor
  g3832
  (
    n3867,
    n3535,
    n3780,
    n2841
  );


  xnor
  g3833
  (
    n3860,
    n3824,
    n3817,
    n3781,
    n3822
  );


  nor
  g3834
  (
    n3859,
    n3812,
    n3529,
    n3816,
    n3825
  );


  or
  g3835
  (
    n3865,
    n3778,
    n3776,
    n3823,
    n3531
  );


  xnor
  g3836
  (
    n3868,
    n2842,
    n3777,
    n3782,
    n2840
  );


  or
  g3837
  (
    n3864,
    n3818,
    n3819,
    n3778,
    n3777
  );


  nand
  g3838
  (
    n3873,
    n3781,
    n3776,
    n3778,
    n3780
  );


  xnor
  g3839
  (
    n3866,
    n3778,
    n3533,
    n3782,
    n3821
  );


  or
  g3840
  (
    n3862,
    n3776,
    n3779,
    n3814,
    n3815
  );


  and
  g3841
  (
    n3880,
    n3725,
    n3540,
    n3736,
    n3723
  );


  or
  g3842
  (
    n3877,
    n3859,
    n3733,
    n3863,
    n3537
  );


  nor
  g3843
  (
    n3882,
    n3538,
    n3866,
    n3735,
    n3868
  );


  nor
  g3844
  (
    n3879,
    n3539,
    n3542,
    n3869,
    n2842
  );


  and
  g3845
  (
    n3883,
    n3541,
    n3737,
    n3726,
    n2843
  );


  nor
  g3846
  (
    n3884,
    n3862,
    n3724,
    n2844,
    n3730
  );


  or
  g3847
  (
    n3874,
    n3729,
    n3860,
    n2844
  );


  nand
  g3848
  (
    n3878,
    n3727,
    n3865,
    n3861,
    n3722
  );


  nand
  g3849
  (
    n3881,
    n3864,
    n3734,
    n3731,
    n3728
  );


  nand
  g3850
  (
    n3876,
    n3867,
    n2843,
    n3738,
    n2842
  );


  xnor
  g3851
  (
    n3875,
    n3732,
    n2843,
    n2844
  );


  xnor
  g3852
  (
    n3886,
    n3768,
    n3551,
    n3544,
    n3884
  );


  or
  g3853
  (
    n3888,
    n3877,
    n3763,
    n3880,
    n3784
  );


  xor
  g3854
  (
    n3885,
    n3765,
    n3878,
    n3764,
    n3547
  );


  xnor
  g3855
  (
    n3893,
    n3784,
    n3770,
    n3883,
    n3783
  );


  xor
  g3856
  (
    n3889,
    n3876,
    n3769,
    n3543,
    n3783
  );


  xor
  g3857
  (
    n3891,
    n3881,
    n3549,
    n1671,
    n3879
  );


  nor
  g3858
  (
    n3890,
    n3548,
    n3784,
    n3783,
    n3882
  );


  xor
  g3859
  (
    n3892,
    n3782,
    n3550,
    n3783,
    n3545
  );


  nand
  g3860
  (
    n3887,
    n3767,
    n3546,
    n3784,
    n3766
  );


  nor
  g3861
  (
    n3903,
    n3886,
    n3891,
    n3828,
    n3892
  );


  nor
  g3862
  (
    n3900,
    n3836,
    n3786,
    n3893,
    n3891
  );


  or
  g3863
  (
    n3907,
    n3787,
    n3893,
    n3832,
    n3790
  );


  nand
  g3864
  (
    n3905,
    n3785,
    n3790,
    n3786,
    n3787
  );


  xnor
  g3865
  (
    n3894,
    n3893,
    n2845,
    n3787,
    n3786
  );


  xor
  g3866
  (
    n3896,
    n3891,
    n3554,
    n3785,
    n3889
  );


  xor
  g3867
  (
    n3895,
    n3845,
    n3839,
    n3833,
    n3838
  );


  nor
  g3868
  (
    n3908,
    n3785,
    n3835,
    n3826,
    n3885
  );


  nand
  g3869
  (
    n3904,
    n3829,
    n3790,
    n3888
  );


  or
  g3870
  (
    n3911,
    n3555,
    n3892,
    n3831,
    n3841
  );


  or
  g3871
  (
    n3899,
    n3890,
    n3558,
    n3893,
    n3552
  );


  nand
  g3872
  (
    n3898,
    n3840,
    n3556,
    n3844,
    n3789
  );


  or
  g3873
  (
    n3906,
    n3846,
    n3842,
    n3789,
    n3892
  );


  nor
  g3874
  (
    n3910,
    n3786,
    n3557,
    n3787,
    n3559
  );


  xnor
  g3875
  (
    n3901,
    n3837,
    n3843,
    n3788,
    n3789
  );


  and
  g3876
  (
    n3897,
    n3892,
    n3834,
    n3788,
    n3827
  );


  nand
  g3877
  (
    n3909,
    n3830,
    n3891,
    n3887,
    n3789
  );


  nor
  g3878
  (
    n3902,
    n3785,
    n3553,
    n3788
  );


  and
  g3879
  (
    n3926,
    n1675,
    n1677,
    n1674,
    n1673
  );


  or
  g3880
  (
    n3916,
    n3898,
    n1679,
    n1682,
    n1675
  );


  nor
  g3881
  (
    n3915,
    n1680,
    n1673,
    n1674
  );


  nand
  g3882
  (
    n3918,
    n1672,
    n1680,
    n3895,
    n1677
  );


  xnor
  g3883
  (
    n3922,
    n1682,
    n1681,
    n1672
  );


  nand
  g3884
  (
    n3921,
    n1678,
    n3898,
    n1671,
    n1676
  );


  and
  g3885
  (
    n3917,
    n1673,
    n3901,
    n1675,
    n1674
  );


  xor
  g3886
  (
    n3913,
    n2845,
    n1679,
    n1672,
    n1681
  );


  xnor
  g3887
  (
    n3912,
    n1676,
    n1681,
    n3900,
    n1679
  );


  xnor
  g3888
  (
    n3925,
    n3894,
    n1680,
    n3900,
    n1678
  );


  xnor
  g3889
  (
    n3923,
    n1679,
    n3897,
    n1680,
    n1677
  );


  nand
  g3890
  (
    n3920,
    n1676,
    n3896,
    n3895
  );


  xnor
  g3891
  (
    n3924,
    n3899,
    n1672,
    n3901,
    n1678
  );


  nor
  g3892
  (
    n3919,
    n1677,
    n3899,
    n3897,
    n1682
  );


  xnor
  g3893
  (
    n3914,
    n1675,
    n1674,
    n1676,
    n1678
  );


  xor
  g3894
  (
    n3930,
    n3571,
    n3569,
    n3561,
    n3562
  );


  and
  g3895
  (
    n3927,
    n3564,
    n3924,
    n3923,
    n3567
  );


  nor
  g3896
  (
    n3929,
    n3563,
    n3568,
    n3926,
    n3570
  );


  or
  g3897
  (
    n3928,
    n3925,
    n3560,
    n3566,
    n3565
  );


  nor
  g3898
  (
    n3934,
    n3929,
    n3855,
    n3930,
    n3574
  );


  and
  g3899
  (
    n3938,
    n1734,
    n3930,
    n1736
  );


  and
  g3900
  (
    n3941,
    n3927,
    n1737,
    n2845,
    n3851
  );


  nor
  g3901
  (
    n3933,
    n1735,
    n3929,
    n1734,
    n3850
  );


  nor
  g3902
  (
    n3939,
    n3572,
    n3929,
    n1734,
    n3857
  );


  nor
  g3903
  (
    n3937,
    n3852,
    n3856,
    n1736,
    n3576
  );


  or
  g3904
  (
    n3932,
    n1735,
    n3849,
    n3930,
    n3928
  );


  nor
  g3905
  (
    n3940,
    n1735,
    n3928,
    n3858,
    n3854
  );


  nor
  g3906
  (
    n3936,
    n3848,
    n3575,
    n1734,
    n1683
  );


  or
  g3907
  (
    n3935,
    n3927,
    n1737,
    n3573,
    n3847
  );


  nand
  g3908
  (
    n3942,
    n1737,
    n1737,
    n1682,
    n3853
  );


  nand
  g3909
  (
    n3931,
    n1736,
    n1735,
    n3930,
    n3929
  );


  or
  g3910
  (
    n3962,
    n3590,
    n3739,
    n3942,
    n3911
  );


  nor
  g3911
  (
    n3953,
    n3589,
    n3931,
    n2849,
    n3583
  );


  xor
  g3912
  (
    n3948,
    n2849,
    n3939,
    n2846,
    n3906
  );


  or
  g3913
  (
    n3979,
    n1690,
    n3940,
    n3935,
    n1754
  );


  and
  g3914
  (
    n3946,
    n3939,
    n3938,
    n1687,
    n3902
  );


  and
  g3915
  (
    n3947,
    n3939,
    n3592,
    n3579,
    n3938
  );


  and
  g3916
  (
    n3958,
    n3935,
    n1684,
    n3580,
    n3933
  );


  and
  g3917
  (
    n3961,
    n3942,
    n3910,
    n3933,
    n3907
  );


  nor
  g3918
  (
    n3955,
    n1683,
    n1690,
    n3938,
    n1754
  );


  or
  g3919
  (
    n3974,
    n1690,
    n3908,
    n2845,
    n3942
  );


  and
  g3920
  (
    n3951,
    n1754,
    n3907,
    n2846,
    n3937
  );


  nor
  g3921
  (
    n3954,
    n3911,
    n3941,
    n2847,
    n3910
  );


  nor
  g3922
  (
    n3960,
    n3908,
    n3741,
    n3584,
    n3935
  );


  nor
  g3923
  (
    n3943,
    n3872,
    n3909,
    n3936,
    n3585
  );


  or
  g3924
  (
    n3977,
    n3905,
    n2848,
    n1686,
    n1755
  );


  and
  g3925
  (
    n3978,
    n1683,
    n3904,
    n2848,
    n1686
  );


  nor
  g3926
  (
    n3963,
    n1690,
    n3905,
    n3740,
    n1686
  );


  xor
  g3927
  (
    n3957,
    n3910,
    n3588,
    n3870,
    n3941
  );


  xor
  g3928
  (
    n3949,
    n2847,
    n3909,
    n3940,
    n1688
  );


  or
  g3929
  (
    n3950,
    n3904,
    n3932,
    n3578,
    n1683
  );


  or
  g3930
  (
    n3952,
    n1689,
    n1689,
    n1684,
    n2847
  );


  and
  g3931
  (
    n3980,
    n3586,
    n3873,
    n3906,
    n1685
  );


  and
  g3932
  (
    n3973,
    n1755,
    n3906,
    n3909,
    n3908
  );


  xnor
  g3933
  (
    n3976,
    n3871,
    n1685,
    n3593,
    n3940
  );


  or
  g3934
  (
    n3971,
    n3908,
    n1684,
    n3903,
    n3911
  );


  or
  g3935
  (
    n3956,
    n1688,
    n3907,
    n2848,
    n1687
  );


  xor
  g3936
  (
    n3965,
    n3591,
    n3941,
    n3910,
    n1691
  );


  nor
  g3937
  (
    n3975,
    n1687,
    n3873,
    n3936,
    n3937
  );


  and
  g3938
  (
    n3966,
    n1755,
    n3936,
    n3937,
    n2847
  );


  and
  g3939
  (
    n3944,
    n2848,
    n3581,
    n3934,
    n3577
  );


  or
  g3940
  (
    n3970,
    n1688,
    n3936,
    n3582,
    n3942
  );


  nand
  g3941
  (
    n3945,
    n3906,
    n3902,
    n1684,
    n1689
  );


  xnor
  g3942
  (
    n3964,
    n1691,
    n1688,
    n2849,
    n1689
  );


  and
  g3943
  (
    n3959,
    n3939,
    n1685,
    n3937
  );


  xor
  g3944
  (
    n3969,
    n1687,
    n2846,
    n1686,
    n1755
  );


  nand
  g3945
  (
    n3968,
    n3935,
    n2846,
    n3909,
    n3903
  );


  nor
  g3946
  (
    n3972,
    n3911,
    n3940,
    n1691,
    n3587
  );


  nand
  g3947
  (
    n3967,
    n3941,
    n3907,
    n3934,
    n3938
  );


  nand
  g3948
  (
    n3992,
    n3957,
    n3966,
    n3594,
    n3959
  );


  nand
  g3949
  (
    n3983,
    n2850,
    n2849,
    n1692,
    n3955
  );


  and
  g3950
  (
    n3986,
    n3974,
    n3956,
    n3965,
    n3977
  );


  nor
  g3951
  (
    n3993,
    n3980,
    n3950,
    n3958,
    n3979
  );


  and
  g3952
  (
    n3994,
    n3977,
    n3600,
    n3970,
    n3961
  );


  and
  g3953
  (
    n3982,
    n3976,
    n3972,
    n3979,
    n3971
  );


  nor
  g3954
  (
    n3981,
    n3945,
    n3954,
    n3980,
    n3979
  );


  or
  g3955
  (
    n3987,
    n3978,
    n3969,
    n3963,
    n3952
  );


  xor
  g3956
  (
    n3989,
    n3962,
    n1692,
    n3596,
    n3980
  );


  xor
  g3957
  (
    n3985,
    n3979,
    n2850,
    n3598,
    n3967
  );


  xnor
  g3958
  (
    AntiSAT_key_wire,
    n3964,
    n3978,
    n3599,
    n3968
  );


  nand
  g3959
  (
    n3984,
    n1692,
    n3946,
    n3975,
    n3978
  );


  nand
  g3960
  (
    n3995,
    n3973,
    n1692,
    n3595,
    n3953
  );


  xor
  g3961
  (
    n3990,
    n3943,
    n1693,
    n2850,
    n1691
  );


  nand
  g3962
  (
    n3991,
    n3949,
    n3597,
    n3947,
    n3978
  );


  nor
  g3963
  (
    n3988,
    n3944,
    n3960,
    n3951,
    n3948
  );


  nor
  g3964
  (
    n3997,
    n3996,
    n1693,
    n3980
  );


  and
  g3965
  (
    n3998,
    n3609,
    n3606,
    n3608,
    n3602
  );


  or
  g3966
  (
    n4000,
    n3603,
    n3997,
    n3605
  );


  and
  g3967
  (
    n4001,
    n3604,
    n3997,
    n3610
  );


  nor
  g3968
  (
    n3999,
    n2851,
    n2850,
    n3607,
    n3601
  );


  and
  g3969
  (
    n4011,
    n2852,
    n2859,
    n3998,
    n3999
  );


  or
  g3970
  (
    n4007,
    n2856,
    n2862,
    n2852,
    n3999
  );


  and
  g3971
  (
    n4016,
    n2853,
    n2862,
    n1693
  );


  or
  g3972
  (
    n4004,
    n2861,
    n2854,
    n2857,
    n2858
  );


  and
  g3973
  (
    n4017,
    n2859,
    n2861,
    n4001,
    n2857
  );


  xor
  g3974
  (
    n4014,
    n2855,
    n2854,
    n2857,
    n2853
  );


  or
  g3975
  (
    n4010,
    n2853,
    n2851,
    n3998,
    n2852
  );


  or
  g3976
  (
    n4006,
    n4001,
    n2858,
    n2859,
    n2853
  );


  nor
  g3977
  (
    n4009,
    n2858,
    n4000,
    n3999,
    n4001
  );


  nand
  g3978
  (
    n4012,
    n2860,
    n2856,
    n4000,
    n2857
  );


  nand
  g3979
  (
    n4003,
    n2855,
    n2856,
    n3998,
    n2862
  );


  and
  g3980
  (
    n4015,
    n2856,
    n2861,
    n3999,
    n4000
  );


  nand
  g3981
  (
    n4002,
    n4000,
    n4001,
    n2855,
    n2860
  );


  xor
  g3982
  (
    n4013,
    n2860,
    n2851,
    n2854,
    n3998
  );


  or
  g3983
  (
    n4005,
    n2858,
    n2851,
    n2852,
    n2859
  );


  xor
  g3984
  (
    n4008,
    n2855,
    n2861,
    n2854,
    n2860
  );


  and
  g3985
  (
    n4025,
    n4003,
    n4013,
    n4014,
    n4015
  );


  xor
  g3986
  (
    n4021,
    n4015,
    n4017,
    n4012
  );


  nand
  g3987
  (
    n4018,
    n4006,
    n2863,
    n4005,
    n2864
  );


  xnor
  g3988
  (
    n4020,
    n2862,
    n4017,
    n4014,
    n4010
  );


  or
  g3989
  (
    n4026,
    n4015,
    n4013,
    n2864,
    n4011
  );


  and
  g3990
  (
    n4022,
    n4008,
    n4013,
    n2864,
    n2863
  );


  xor
  g3991
  (
    n4019,
    n4011,
    n4016,
    n4007,
    n4012
  );


  and
  g3992
  (
    n4027,
    n4015,
    n4017,
    n4013
  );


  xnor
  g3993
  (
    n4024,
    n4016,
    n4016,
    n4014,
    n2863
  );


  xnor
  g3994
  (
    n4029,
    n2863,
    n4002,
    n4004,
    n4012
  );


  xor
  g3995
  (
    n4028,
    n4009,
    n4011
  );


  and
  g3996
  (
    n4023,
    n2864,
    n4016,
    n4010,
    n4014
  );


  nand
  g3997
  (
    n4030,
    n4020,
    n4029,
    n4022,
    n4021
  );


  nand
  g3998
  (
    n4032,
    n4027,
    n4023,
    n4019,
    n4026
  );


  xor
  g3999
  (
    n4031,
    n4024,
    n4025,
    n4018,
    n4028
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n3996,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

