// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_42 written by SynthGen on 2021/04/05 11:08:36
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_42 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n116, n115, n114, n107, n101, n125, n119, n103,
 n112, n111, n117, n129, n113, n126, n109, n110,
 n132, n120, n104, n102, n122, n131, n105, n128,
 n123, n108, n130, n124, n118, n121, n127, n106);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n116, n115, n114, n107, n101, n125, n119, n103,
 n112, n111, n117, n129, n113, n126, n109, n110,
 n132, n120, n104, n102, n122, n131, n105, n128,
 n123, n108, n130, n124, n118, n121, n127, n106;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

not  g0 (n41, n8);
buf  g1 (n38, n6);
buf  g2 (n55, n2);
not  g3 (n51, n11);
not  g4 (n52, n9);
buf  g5 (n56, n8);
buf  g6 (n49, n9);
not  g7 (n36, n10);
buf  g8 (n42, n10);
not  g9 (n37, n8);
not  g10 (n60, n3);
not  g11 (n50, n6);
buf  g12 (n33, n7);
buf  g13 (n58, n7);
buf  g14 (n40, n10);
buf  g15 (n48, n8);
buf  g16 (n54, n9);
buf  g17 (n46, n9);
not  g18 (n34, n1);
not  g19 (n59, n11);
buf  g20 (n57, n7);
buf  g21 (n45, n5);
not  g22 (n39, n10);
not  g23 (n47, n6);
not  g24 (n35, n11);
buf  g25 (n61, n4);
not  g26 (n53, n6);
not  g27 (n43, n7);
not  g28 (n44, n11);
buf  g29 (n68, n33);
not  g30 (n66, n37);
not  g31 (n69, n35);
not  g32 (n67, n37);
buf  g33 (n64, n37);
not  g34 (n63, n36);
not  g35 (n65, n37);
not  g36 (n62, n34);
nand g37 (n79, n20, n29, n67, n17);
or   g38 (n98, n21, n23, n69);
and  g39 (n76, n30, n68, n25, n15);
or   g40 (n87, n39, n65, n66, n14);
or   g41 (n86, n38, n38, n23, n39);
nor  g42 (n73, n68, n12, n21);
xnor g43 (n95, n19, n29, n28);
nor  g44 (n94, n62, n25, n38, n16);
and  g45 (n72, n26, n24, n68, n65);
nor  g46 (n91, n63, n28, n40, n22);
or   g47 (n77, n39, n30, n66, n15);
nand g48 (n96, n32, n64, n14, n63);
nand g49 (n83, n67, n62, n23, n69);
nand g50 (n70, n27, n67, n22);
or   g51 (n97, n27, n31, n30, n17);
or   g52 (n89, n28, n24, n12, n13);
xnor g53 (n82, n22, n14, n27, n68);
and  g54 (n93, n16, n22, n31, n62);
nor  g55 (n100, n64, n23, n13);
nand g56 (n88, n18, n63, n65);
xor  g57 (n78, n40, n19, n64, n30);
and  g58 (n75, n28, n40, n29, n26);
and  g59 (n85, n19, n15, n17, n62);
xnor g60 (n84, n14, n19, n64, n27);
or   g61 (n80, n66, n65, n24, n25);
nand g62 (n99, n18, n16, n31, n20);
xnor g63 (n74, n20, n26, n39, n21);
xnor g64 (n81, n25, n66, n16, n32);
xnor g65 (n92, n18, n38, n24, n15);
xnor g66 (n71, n18, n12, n13, n20);
nor  g67 (n90, n21, n31, n26, n17);
nand g68 (n118, n95, n94, n57, n43);
xnor g69 (n126, n48, n61, n93, n59);
xnor g70 (n132, n47, n99, n100, n56);
nand g71 (n129, n54, n42, n71, n48);
xnor g72 (n110, n45, n47, n98, n44);
xor  g73 (n109, n96, n85, n86, n88);
and  g74 (n125, n55, n60, n80, n41);
xnor g75 (n127, n41, n44, n53, n90);
nor  g76 (n114, n73, n60, n91, n54);
and  g77 (n120, n81, n43, n48, n41);
nand g78 (n111, n99, n51, n74, n40);
and  g79 (n113, n57, n82, n100, n41);
xnor g80 (n128, n51, n46, n45, n56);
nor  g81 (n105, n51, n99, n49);
or   g82 (n121, n98, n54, n57, n60);
nor  g83 (n103, n92, n58, n79, n76);
xnor g84 (n131, n54, n46, n59, n50);
xnor g85 (n106, n97, n56, n99, n58);
nand g86 (n116, n47, n53, n77, n46);
xor  g87 (n115, n78, n44, n100, n98);
and  g88 (n124, n98, n89, n43, n48);
or   g89 (n104, n55, n50, n53, n61);
xnor g90 (n102, n42, n70, n50, n49);
nand g91 (n101, n45, n60, n59, n69);
and  g92 (n107, n42, n44, n52, n58);
xor  g93 (n122, n58, n32, n53, n59);
xnor g94 (n130, n83, n100, n61, n55);
and  g95 (n123, n84, n45, n57, n51);
xnor g96 (n108, n87, n47, n42, n43);
or   g97 (n117, n50, n46, n52, n61);
nand g98 (n119, n72, n49, n52);
and  g99 (n112, n75, n55, n32, n56);
endmodule
