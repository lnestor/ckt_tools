// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_541_1114 written by SynthGen on 2021/05/24 19:47:35
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_541_1114 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31,
 n555, n546, n564, n552, n572, n544, n571, n557,
 n545, n560, n543, n568, n562, n570, n558, n567,
 n550, n551, n556, n554, n547, n565, n549, n559,
 n569, n548, n561, n563, n566, n553);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31;

output n555, n546, n564, n552, n572, n544, n571, n557,
 n545, n560, n543, n568, n562, n570, n558, n567,
 n550, n551, n556, n554, n547, n565, n549, n559,
 n569, n548, n561, n563, n566, n553;

wire n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n402, n403, n404, n405, n406, n407,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n425, n426, n427, n428, n429, n430, n431,
 n432, n433, n434, n435, n436, n437, n438, n439,
 n440, n441, n442, n443, n444, n445, n446, n447,
 n448, n449, n450, n451, n452, n453, n454, n455,
 n456, n457, n458, n459, n460, n461, n462, n463,
 n464, n465, n466, n467, n468, n469, n470, n471,
 n472, n473, n474, n475, n476, n477, n478, n479,
 n480, n481, n482, n483, n484, n485, n486, n487,
 n488, n489, n490, n491, n492, n493, n494, n495,
 n496, n497, n498, n499, n500, n501, n502, n503,
 n504, n505, n506, n507, n508, n509, n510, n511,
 n512, n513, n514, n515, n516, n517, n518, n519,
 n520, n521, n522, n523, n524, n525, n526, n527,
 n528, n529, n530, n531, n532, n533, n534, n535,
 n536, n537, n538, n539, n540, n541, n542;

buf  g0 (n102, n20);
not  g1 (n63, n11);
buf  g2 (n36, n2);
buf  g3 (n97, n9);
buf  g4 (n62, n7);
buf  g5 (n91, n12);
buf  g6 (n41, n1);
buf  g7 (n112, n19);
not  g8 (n106, n14);
not  g9 (n81, n5);
not  g10 (n98, n13);
buf  g11 (n32, n11);
buf  g12 (n118, n7);
not  g13 (n33, n5);
not  g14 (n95, n20);
buf  g15 (n69, n21);
not  g16 (n66, n10);
not  g17 (n61, n12);
buf  g18 (n47, n4);
not  g19 (n84, n16);
buf  g20 (n117, n12);
not  g21 (n50, n18);
buf  g22 (n38, n11);
not  g23 (n67, n6);
buf  g24 (n59, n22);
buf  g25 (n74, n6);
not  g26 (n52, n1);
buf  g27 (n73, n3);
buf  g28 (n44, n1);
buf  g29 (n114, n11);
not  g30 (n88, n5);
buf  g31 (n35, n23);
not  g32 (n49, n18);
not  g33 (n46, n6);
buf  g34 (n54, n17);
buf  g35 (n87, n10);
not  g36 (n104, n14);
buf  g37 (n86, n19);
buf  g38 (n57, n13);
not  g39 (n110, n3);
buf  g40 (n77, n2);
not  g41 (n82, n8);
buf  g42 (n119, n22);
buf  g43 (n72, n5);
buf  g44 (n70, n14);
not  g45 (n83, n15);
not  g46 (n39, n4);
buf  g47 (n96, n14);
not  g48 (n53, n22);
not  g49 (n85, n20);
not  g50 (n56, n21);
buf  g51 (n64, n13);
buf  g52 (n93, n9);
not  g53 (n79, n17);
not  g54 (n55, n21);
buf  g55 (n43, n19);
not  g56 (n45, n2);
buf  g57 (n90, n17);
not  g58 (n71, n9);
not  g59 (n99, n19);
not  g60 (n107, n17);
not  g61 (n58, n6);
buf  g62 (n113, n7);
buf  g63 (n42, n8);
buf  g64 (n48, n10);
not  g65 (n92, n18);
not  g66 (n65, n21);
not  g67 (n109, n7);
buf  g68 (n76, n8);
not  g69 (n34, n16);
buf  g70 (n111, n9);
not  g71 (n89, n16);
not  g72 (n116, n16);
buf  g73 (n101, n15);
buf  g74 (n94, n15);
not  g75 (n37, n1);
not  g76 (n115, n13);
buf  g77 (n108, n18);
buf  g78 (n75, n15);
not  g79 (n103, n3);
not  g80 (n80, n8);
not  g81 (n60, n3);
not  g82 (n78, n20);
buf  g83 (n105, n12);
not  g84 (n120, n4);
buf  g85 (n40, n22);
buf  g86 (n100, n4);
not  g87 (n68, n2);
not  g88 (n51, n10);
not  g89 (n166, n57);
buf  g90 (n197, n91);
not  g91 (n180, n60);
not  g92 (n163, n63);
buf  g93 (n123, n49);
buf  g94 (n243, n32);
not  g95 (n228, n26);
not  g96 (n154, n76);
buf  g97 (n231, n65);
not  g98 (n158, n38);
buf  g99 (n138, n39);
not  g100 (n156, n40);
not  g101 (n160, n54);
not  g102 (n169, n90);
buf  g103 (n238, n27);
buf  g104 (n208, n28);
not  g105 (n130, n61);
not  g106 (n227, n87);
buf  g107 (n142, n30);
buf  g108 (n225, n32);
not  g109 (n239, n95);
buf  g110 (n128, n84);
not  g111 (n162, n46);
buf  g112 (n240, n77);
buf  g113 (n132, n51);
buf  g114 (n233, n48);
buf  g115 (n189, n97);
not  g116 (n146, n61);
not  g117 (n175, n96);
not  g118 (n144, n48);
not  g119 (n215, n74);
not  g120 (n134, n36);
buf  g121 (n224, n62);
buf  g122 (n176, n46);
not  g123 (n196, n79);
not  g124 (n183, n74);
buf  g125 (n192, n33);
not  g126 (n137, n45);
buf  g127 (n125, n26);
buf  g128 (n205, n83);
buf  g129 (n184, n34);
not  g130 (n172, n40);
not  g131 (n157, n88);
buf  g132 (n122, n95);
buf  g133 (n143, n59);
not  g134 (n203, n81);
not  g135 (n164, n53);
not  g136 (n181, n83);
buf  g137 (n139, n23);
not  g138 (n217, n36);
not  g139 (n135, n77);
not  g140 (n234, n65);
not  g141 (n141, n38);
buf  g142 (n165, n77);
buf  g143 (n190, n74);
not  g144 (n121, n69);
not  g145 (n167, n44);
buf  g146 (n178, n48);
buf  g147 (n133, n36);
buf  g148 (n213, n38);
not  g149 (n230, n92);
buf  g150 (n245, n53);
not  g151 (n147, n35);
buf  g152 (n179, n41);
not  g153 (n202, n24);
xor  g154 (n219, n87, n57);
nand g155 (n177, n80, n93, n45, n92);
xnor g156 (n204, n79, n29, n43, n42);
or   g157 (n232, n68, n24, n73, n37);
xnor g158 (n200, n56, n94, n31, n71);
and  g159 (n223, n83, n55, n93, n85);
xor  g160 (n124, n26, n58, n62, n56);
nand g161 (n187, n97, n38, n33);
or   g162 (n155, n75, n52, n96);
nand g163 (n218, n45, n25, n28, n80);
and  g164 (n201, n82, n39, n42, n89);
xor  g165 (n148, n70, n73, n85, n56);
xnor g166 (n131, n76, n72, n53);
nor  g167 (n150, n95, n66, n42, n88);
and  g168 (n193, n56, n72, n62, n68);
xor  g169 (n152, n75, n37, n43, n93);
nor  g170 (n199, n66, n31, n82, n68);
xnor g171 (n216, n43, n65, n74, n58);
and  g172 (n185, n59, n52, n90, n30);
xnor g173 (n171, n25, n57, n46, n31);
or   g174 (n168, n29, n78, n86, n44);
and  g175 (n195, n30, n70, n41, n81);
xnor g176 (n126, n94, n98, n71, n93);
nor  g177 (n236, n90, n34, n94, n76);
nand g178 (n237, n73, n43, n90, n47);
nand g179 (n188, n44, n42, n71, n54);
xnor g180 (n214, n58, n28, n89, n88);
xor  g181 (n226, n86, n73, n41, n25);
or   g182 (n159, n44, n34, n59, n88);
xor  g183 (n229, n81, n39, n64, n34);
nand g184 (n186, n61, n37, n67, n72);
xor  g185 (n174, n67, n52, n69, n92);
xor  g186 (n210, n29, n96, n86, n87);
nand g187 (n222, n32, n54, n23, n31);
nor  g188 (n211, n50, n84);
nor  g189 (n173, n67, n64, n27);
and  g190 (n191, n61, n78, n45, n59);
or   g191 (n149, n63, n50, n79, n55);
nand g192 (n244, n35, n39, n75, n64);
nor  g193 (n207, n77, n47, n70, n85);
nor  g194 (n206, n33, n83, n60, n78);
or   g195 (n136, n27, n35, n55, n89);
or   g196 (n198, n96, n51, n55, n60);
nand g197 (n220, n67, n36, n66, n49);
or   g198 (n194, n76, n98, n80, n62);
xnor g199 (n145, n82, n91, n24);
or   g200 (n140, n32, n47, n58, n80);
xor  g201 (n212, n70, n81, n48, n50);
nor  g202 (n127, n94, n49, n57, n47);
and  g203 (n129, n51, n41, n79, n91);
xnor g204 (n151, n86, n84, n46, n60);
xnor g205 (n182, n75, n85, n68, n66);
xor  g206 (n221, n25, n27, n23, n69);
or   g207 (n241, n35, n63, n78, n71);
or   g208 (n235, n63, n30, n95, n24);
xor  g209 (n209, n28, n54, n26, n97);
nor  g210 (n161, n89, n69, n92, n49);
nor  g211 (n153, n87, n51, n40, n98);
nor  g212 (n242, n97, n98, n40, n65);
or   g213 (n170, n37, n72, n29, n82);
nor  g214 (n251, n134, n127);
xor  g215 (n246, n122, n129);
nand g216 (n250, n126, n133);
not  g217 (n257, n100);
not  g218 (n247, n99);
xor  g219 (n255, n101, n124);
nand g220 (n252, n102, n130);
nand g221 (n260, n121, n131);
or   g222 (n259, n128, n132);
nand g223 (n256, n100, n102);
xor  g224 (n249, n123, n101);
nor  g225 (n253, n125, n135);
nor  g226 (n258, n100, n102);
buf  g227 (n248, n101);
nand g228 (n254, n102, n136);
buf  g229 (n261, n99);
or   g230 (n306, n204, n247, n174, n213);
xnor g231 (n308, n178, n140, n202, n256);
nor  g232 (n302, n164, n154, n179, n210);
xor  g233 (n297, n247, n236, n212, n224);
nor  g234 (n324, n218, n217, n260, n257);
nor  g235 (n307, n236, n208, n249, n220);
or   g236 (n304, n219, n251, n137, n159);
or   g237 (n263, n258, n250, n215, n261);
nor  g238 (n274, n168, n162, n248, n255);
nand g239 (n321, n185, n230, n223, n236);
or   g240 (n270, n251, n225, n214, n221);
and  g241 (n286, n246, n225, n250, n251);
and  g242 (n313, n209, n222, n230, n249);
and  g243 (n294, n246, n252, n233, n220);
and  g244 (n271, n231, n171, n170, n206);
xnor g245 (n293, n250, n227, n226, n201);
or   g246 (n301, n235, n213, n210, n211);
and  g247 (n300, n200, n209, n227, n145);
xnor g248 (n305, n215, n219, n225, n196);
nand g249 (n288, n223, n219, n195, n258);
and  g250 (n280, n218, n235, n225, n252);
nor  g251 (n318, n208, n209, n229, n251);
nor  g252 (n315, n254, n219, n253, n236);
xor  g253 (n285, n214, n249, n246, n216);
and  g254 (n296, n155, n211, n253, n175);
nor  g255 (n299, n138, n217, n218, n246);
and  g256 (n277, n221, n215, n223, n189);
nand g257 (n323, n203, n221, n214, n259);
nand g258 (n264, n161, n226, n228, n180);
or   g259 (n319, n255, n261, n205, n259);
nand g260 (n276, n254, n199, n158, n198);
or   g261 (n303, n222, n231, n253, n252);
nand g262 (n298, n257, n232, n228);
nand g263 (n275, n247, n217, n233, n193);
or   g264 (n278, n207, n226, n248, n234);
xor  g265 (n325, n172, n153, n258, n210);
xnor g266 (n281, n234, n261, n260, n259);
or   g267 (n279, n224, n223, n212, n143);
xor  g268 (n287, n165, n213, n212, n248);
nor  g269 (n322, n257, n247, n206, n148);
nor  g270 (n289, n211, n149, n190, n212);
or   g271 (n290, n235, n142, n257, n144);
nor  g272 (n292, n146, n222, n256, n216);
xnor g273 (n273, n261, n218, n249, n228);
xor  g274 (n311, n228, n255, n224, n151);
nand g275 (n283, n250, n256, n232, n222);
or   g276 (n314, n204, n182, n226, n169);
nor  g277 (n267, n220, n197, n157, n211);
xor  g278 (n272, n207, n254, n230, n233);
and  g279 (n269, n253, n229, n184, n216);
nand g280 (n284, n183, n177, n230, n194);
and  g281 (n310, n156, n208, n207, n206);
xnor g282 (n282, n187, n213, n221, n231);
nor  g283 (n312, n173, n216, n260);
nand g284 (n320, n139, n220, n252, n229);
or   g285 (n266, n248, n235, n166, n191);
nand g286 (n317, n167, n234, n215, n217);
or   g287 (n295, n229, n231, n192, n255);
nand g288 (n268, n254, n186, n227, n188);
and  g289 (n316, n205, n204, n256, n258);
and  g290 (n262, n227, n234, n232, n214);
nor  g291 (n309, n259, n152, n181, n205);
or   g292 (n265, n224, n176, n141, n147);
or   g293 (n291, n160, n150, n233, n163);
xnor g294 (n342, n301, n301, n271, n105);
nor  g295 (n372, n111, n287, n271, n285);
or   g296 (n404, n280, n104, n265, n306);
nand g297 (n379, n108, n239, n286, n273);
xnor g298 (n351, n308, n116, n316, n240);
and  g299 (n341, n320, n290, n322, n112);
xor  g300 (n347, n311, n117, n111, n106);
nand g301 (n326, n264, n280, n313, n274);
xnor g302 (n371, n274, n291, n278, n302);
nand g303 (n334, n310, n109, n299, n117);
and  g304 (n405, n110, n115, n114, n314);
or   g305 (n383, n270, n268, n289, n294);
and  g306 (n346, n299, n317, n312, n320);
nand g307 (n353, n306, n107, n103, n276);
and  g308 (n363, n287, n116, n267, n314);
xnor g309 (n390, n320, n237, n272, n290);
xnor g310 (n381, n314, n104, n283, n313);
and  g311 (n375, n238, n275, n276, n277);
xnor g312 (n344, n272, n110, n268, n310);
and  g313 (n400, n239, n315, n298, n106);
or   g314 (n343, n282, n242, n263, n304);
xor  g315 (n335, n319, n281, n276, n303);
nand g316 (n359, n322, n300, n296, n265);
xor  g317 (n395, n269, n108, n271, n293);
nand g318 (n355, n268, n318, n115, n264);
nand g319 (n370, n299, n296, n111, n276);
xnor g320 (n403, n297, n104, n107, n106);
nand g321 (n399, n115, n238, n289, n273);
and  g322 (n408, n110, n308, n312, n293);
or   g323 (n366, n267, n284, n263, n290);
xnor g324 (n349, n280, n298, n109, n292);
and  g325 (n358, n268, n294, n239, n295);
and  g326 (n350, n300, n310, n262, n114);
nor  g327 (n389, n315, n110, n303, n286);
or   g328 (n402, n273, n314, n319, n270);
or   g329 (n336, n267, n312, n109, n293);
nor  g330 (n388, n322, n275, n283, n115);
xnor g331 (n382, n315, n116, n286, n243);
or   g332 (n329, n309, n305, n311, n244);
nor  g333 (n373, n298, n302, n282, n283);
nor  g334 (n333, n285, n309, n113, n283);
or   g335 (n393, n307, n240, n321, n267);
and  g336 (n376, n114, n288, n291, n295);
or   g337 (n396, n317, n103, n239, n265);
and  g338 (n364, n241, n108, n305, n304);
xor  g339 (n340, n272, n311, n103, n307);
xnor g340 (n332, n303, n262, n318, n294);
xnor g341 (n369, n311, n237, n304, n242);
xnor g342 (n384, n266, n288, n241, n106);
nor  g343 (n338, n238, n306, n322, n278);
nand g344 (n330, n307, n113, n109, n295);
and  g345 (n401, n300, n105, n241, n315);
nand g346 (n394, n305, n275, n320, n107);
nand g347 (n337, n117, n296, n108, n284);
nor  g348 (n368, n321, n321, n105, n297);
xnor g349 (n328, n301, n313, n264, n295);
xor  g350 (n352, n284, n243, n292);
nand g351 (n361, n285, n281, n262, n288);
xnor g352 (n365, n262, n282, n287, n301);
xor  g353 (n345, n302, n242, n277, n285);
and  g354 (n357, n240, n317, n279, n291);
or   g355 (n397, n298, n107, n270, n308);
or   g356 (n360, n237, n305, n242, n277);
xor  g357 (n348, n297, n272, n292, n112);
and  g358 (n354, n313, n280, n303, n266);
xor  g359 (n339, n271, n238, n318, n279);
or   g360 (n385, n296, n273, n240, n241);
or   g361 (n378, n288, n281, n112, n279);
nor  g362 (n356, n297, n266, n243, n308);
xor  g363 (n380, n321, n265, n292, n316);
nor  g364 (n374, n291, n114, n116, n317);
and  g365 (n367, n270, n263, n289, n281);
xor  g366 (n386, n104, n286, n113, n274);
or   g367 (n392, n113, n284, n300, n237);
nor  g368 (n387, n299, n289, n293, n319);
or   g369 (n362, n275, n307, n279, n302);
nand g370 (n398, n269, n309, n318, n310);
or   g371 (n407, n282, n316, n269, n111);
xor  g372 (n327, n278, n312, n319, n264);
xor  g373 (n377, n278, n103, n274, n266);
xor  g374 (n406, n290, n263, n277, n306);
and  g375 (n331, n269, n294, n105, n316);
nor  g376 (n391, n304, n112, n287, n309);
or   g377 (n409, n326, n324);
xor  g378 (n410, n327, n323, n324);
or   g379 (n411, n328, n323);
nor  g380 (n418, n358, n333, n411, n334);
or   g381 (n415, n336, n357, n335, n410);
xnor g382 (n420, n346, n343, n338, n352);
nor  g383 (n416, n410, n411, n354);
and  g384 (n414, n344, n337, n349, n409);
nand g385 (n417, n341, n351, n350, n331);
nor  g386 (n412, n411, n332, n348, n409);
nor  g387 (n419, n353, n339, n410, n330);
and  g388 (n421, n356, n345, n347, n342);
nand g389 (n413, n340, n355, n329, n409);
not  g390 (n451, n118);
not  g391 (n426, n362);
not  g392 (n461, n364);
buf  g393 (n454, n420);
buf  g394 (n450, n368);
buf  g395 (n455, n415);
buf  g396 (n457, n359);
buf  g397 (n438, n412);
buf  g398 (n423, n412);
not  g399 (n428, n420);
not  g400 (n452, n415);
not  g401 (n447, n417);
not  g402 (n425, n417);
buf  g403 (n442, n416);
buf  g404 (n441, n415);
buf  g405 (n435, n418);
buf  g406 (n449, n366);
buf  g407 (n458, n414);
buf  g408 (n431, n416);
not  g409 (n460, n360);
buf  g410 (n433, n420);
buf  g411 (n439, n413);
buf  g412 (n445, n363);
buf  g413 (n448, n361);
buf  g414 (n429, n421);
not  g415 (n440, n118);
not  g416 (n446, n421);
buf  g417 (n436, n415);
not  g418 (n456, n417);
not  g419 (n430, n416);
not  g420 (n424, n412);
buf  g421 (n459, n419);
not  g422 (n434, n419);
not  g423 (n443, n413);
xor  g424 (n437, n370, n117, n417);
nor  g425 (n432, n413, n421);
or   g426 (n444, n414, n413, n418);
xnor g427 (n422, n414, n369, n367, n419);
or   g428 (n453, n365, n420, n414, n418);
and  g429 (n427, n419, n412, n416, n118);
not  g430 (n482, n426);
not  g431 (n479, n424);
buf  g432 (n480, n427);
not  g433 (n465, n424);
not  g434 (n472, n427);
buf  g435 (n462, n426);
not  g436 (n467, n423);
buf  g437 (n474, n427);
not  g438 (n468, n425);
buf  g439 (n483, n424);
buf  g440 (n485, n423);
buf  g441 (n471, n427);
not  g442 (n477, n422);
buf  g443 (n466, n422);
buf  g444 (n484, n425);
not  g445 (n473, n424);
not  g446 (n463, n426);
buf  g447 (n470, n426);
not  g448 (n476, n425);
not  g449 (n481, n423);
buf  g450 (n464, n422);
buf  g451 (n475, n423);
not  g452 (n469, n425);
not  g453 (n478, n422);
nor  g454 (n517, n372, n456, n463, n383);
xnor g455 (n516, n120, n379, n444, n442);
or   g456 (n522, n471, n452, n120, n465);
nor  g457 (n500, n429, n450, n431, n458);
xnor g458 (n529, n119, n391, n440, n459);
or   g459 (n537, n371, n452, n471, n430);
nor  g460 (n526, n458, n463, n438, n472);
or   g461 (n515, n373, n429, n437, n441);
xor  g462 (n520, n437, n431, n438, n119);
xnor g463 (n533, n463, n432, n445, n394);
xnor g464 (n542, n460, n464, n440, n392);
or   g465 (n532, n471, n456, n451, n462);
and  g466 (n541, n444, n433, n387);
and  g467 (n519, n462, n454, n439, n375);
and  g468 (n534, n474, n434, n454, n447);
nand g469 (n499, n437, n435, n432, n445);
nand g470 (n492, n444, n451, n443, n462);
xnor g471 (n502, n469, n461, n457, n433);
xor  g472 (n525, n442, n446, n385, n471);
or   g473 (n535, n448, n468, n453, n475);
and  g474 (n498, n436, n461, n469, n435);
or   g475 (n496, n452, n456, n454, n474);
xor  g476 (n524, n458, n439, n459, n447);
xor  g477 (n528, n475, n470, n389, n458);
and  g478 (n494, n468, n460, n473, n469);
xnor g479 (n491, n462, n442, n120, n445);
nor  g480 (n490, n466, n434, n465, n470);
and  g481 (n527, n453, n118, n465, n436);
and  g482 (n536, n473, n441, n430, n461);
xor  g483 (n501, n448, n430, n457, n396);
nand g484 (n493, n455, n448, n435, n467);
nor  g485 (n503, n438, n437, n382, n429);
or   g486 (n518, n476, n475, n469, n441);
nor  g487 (n514, n464, n457, n460, n442);
xnor g488 (n509, n440, n460, n475, n393);
xnor g489 (n540, n434, n432, n376, n453);
and  g490 (n523, n465, n440, n461, n449);
or   g491 (n497, n466, n377, n431);
and  g492 (n538, n450, n443, n466, n428);
and  g493 (n513, n447, n451, n470);
and  g494 (n495, n464, n473, n450);
or   g495 (n488, n459, n464, n467, n428);
nand g496 (n531, n452, n378, n443, n455);
xnor g497 (n530, n439, n447, n468, n388);
and  g498 (n506, n120, n438, n435, n433);
or   g499 (n510, n472, n446, n470, n381);
nand g500 (n505, n474, n455, n467, n428);
xnor g501 (n539, n446, n443, n455, n474);
nand g502 (n486, n449, n450, n119, n467);
xor  g503 (n487, n446, n463, n457, n374);
xor  g504 (n507, n441, n384, n448, n436);
xnor g505 (n521, n456, n445, n449, n429);
and  g506 (n508, n472, n472, n436, n395);
or   g507 (n489, n466, n386, n439, n449);
xor  g508 (n512, n454, n390, n434, n432);
xnor g509 (n504, n444, n453, n430, n380);
or   g510 (n511, n428, n468, n459, n119);
xnor g511 (n561, n520, n506, n526, n512);
xnor g512 (n548, n325, n477, n503, n497);
nor  g513 (n568, n485, n400, n479, n499);
xor  g514 (n554, n489, n398, n245, n480);
nand g515 (n544, n477, n478, n245, n487);
nor  g516 (n551, n407, n529, n501, n325);
nor  g517 (n550, n524, n324, n522, n538);
or   g518 (n569, n480, n502, n483, n478);
nor  g519 (n555, n495, n397, n401, n521);
nand g520 (n545, n496, n530, n531, n483);
nand g521 (n559, n482, n532, n476, n533);
or   g522 (n547, n244, n518, n483, n481);
xor  g523 (n563, n402, n477, n478, n541);
xnor g524 (n562, n483, n325, n525);
xnor g525 (n560, n484, n482, n504, n244);
nor  g526 (n564, n498, n245, n514, n493);
or   g527 (n570, n540, n527, n399, n488);
nand g528 (n556, n508, n519, n403, n490);
nand g529 (n549, n486, n511, n479, n536);
and  g530 (n572, n523, n404, n484, n479);
and  g531 (n571, n482, n484, n405, n539);
or   g532 (n543, n542, n476, n481);
or   g533 (n546, n510, n478, n477, n482);
xnor g534 (n567, n408, n480, n509, n507);
nor  g535 (n552, n480, n485, n244, n484);
xor  g536 (n553, n535, n505, n515, n500);
nand g537 (n565, n485, n537, n492, n494);
and  g538 (n566, n516, n528, n491, n534);
nand g539 (n557, n485, n245, n406, n479);
or   g540 (n558, n517, n481, n513, n476);
endmodule
