// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_221_421 written by SynthGen on 2021/05/24 19:47:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_221_421 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17,
 n231, n212, n208, n238, n207, n226, n218, n214,
 n220, n227, n234, n235, n228, n222, n223, n209,
 n230, n224, n221, n210, n233, n216, n219, n237,
 n236, n232, n217, n213, n229, n215, n211, n225);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17;

output n231, n212, n208, n238, n207, n226, n218, n214,
 n220, n227, n234, n235, n228, n222, n223, n209,
 n230, n224, n221, n210, n233, n216, n219, n237,
 n236, n232, n217, n213, n229, n215, n211, n225;

wire n18, n19, n20, n21, n22, n23, n24, n25,
 n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206;

not  g0 (n28, n2);
buf  g1 (n18, n3);
not  g2 (n26, n3);
not  g3 (n32, n1);
buf  g4 (n22, n5);
buf  g5 (n30, n1);
buf  g6 (n23, n3);
not  g7 (n25, n5);
buf  g8 (n19, n2);
not  g9 (n21, n5);
not  g10 (n20, n1);
buf  g11 (n29, n4);
buf  g12 (n31, n2);
buf  g13 (n27, n4);
not  g14 (n24, n4);
buf  g15 (n78, n23);
not  g16 (n58, n21);
not  g17 (n53, n22);
not  g18 (n62, n32);
not  g19 (n69, n22);
buf  g20 (n59, n24);
buf  g21 (n48, n21);
buf  g22 (n61, n20);
not  g23 (n67, n26);
not  g24 (n65, n18);
not  g25 (n52, n30);
buf  g26 (n57, n32);
not  g27 (n73, n28);
not  g28 (n40, n31);
not  g29 (n50, n20);
buf  g30 (n43, n23);
not  g31 (n44, n19);
not  g32 (n34, n18);
buf  g33 (n37, n29);
buf  g34 (n42, n25);
not  g35 (n74, n28);
not  g36 (n70, n18);
not  g37 (n41, n27);
not  g38 (n47, n29);
not  g39 (n49, n24);
buf  g40 (n55, n30);
not  g41 (n68, n22);
buf  g42 (n38, n20);
buf  g43 (n64, n28);
buf  g44 (n72, n24);
not  g45 (n33, n27);
buf  g46 (n39, n26);
buf  g47 (n51, n19);
buf  g48 (n54, n30);
not  g49 (n63, n26);
not  g50 (n45, n21);
buf  g51 (n60, n27);
buf  g52 (n75, n32);
buf  g53 (n36, n19);
buf  g54 (n71, n25);
buf  g55 (n77, n31);
buf  g56 (n35, n23);
not  g57 (n66, n32);
not  g58 (n46, n29);
not  g59 (n76, n31);
buf  g60 (n56, n25);
buf  g61 (n174, n33);
buf  g62 (n101, n60);
not  g63 (n94, n45);
buf  g64 (n181, n77);
buf  g65 (n104, n48);
not  g66 (n155, n52);
not  g67 (n201, n9);
buf  g68 (n143, n76);
not  g69 (n91, n71);
buf  g70 (n165, n34);
buf  g71 (n99, n35);
not  g72 (n199, n65);
not  g73 (n106, n77);
not  g74 (n98, n57);
buf  g75 (n176, n53);
buf  g76 (n178, n75);
not  g77 (n108, n17);
not  g78 (n141, n59);
buf  g79 (n150, n45);
not  g80 (n124, n41);
buf  g81 (n203, n77);
not  g82 (n128, n69);
not  g83 (n196, n39);
not  g84 (n102, n67);
buf  g85 (n156, n46);
buf  g86 (n139, n41);
buf  g87 (n205, n78);
buf  g88 (n132, n47);
not  g89 (n127, n50);
not  g90 (n133, n61);
buf  g91 (n197, n60);
buf  g92 (n84, n69);
not  g93 (n136, n78);
buf  g94 (n80, n65);
buf  g95 (n125, n38);
not  g96 (n182, n14);
buf  g97 (n81, n41);
buf  g98 (n112, n7);
buf  g99 (n123, n66);
not  g100 (n160, n14);
buf  g101 (n87, n65);
buf  g102 (n118, n55);
buf  g103 (n138, n36);
not  g104 (n170, n8);
not  g105 (n154, n72);
not  g106 (n188, n70);
not  g107 (n145, n54);
buf  g108 (n137, n44);
not  g109 (n130, n76);
buf  g110 (n206, n73);
buf  g111 (n149, n52);
buf  g112 (n90, n35);
not  g113 (n120, n42);
not  g114 (n192, n8);
not  g115 (n111, n74);
buf  g116 (n117, n74);
buf  g117 (n129, n7);
not  g118 (n202, n15);
not  g119 (n166, n49);
buf  g120 (n114, n6);
buf  g121 (n126, n47);
not  g122 (n142, n59);
not  g123 (n96, n33);
buf  g124 (n147, n15);
buf  g125 (n157, n53);
not  g126 (n97, n34);
buf  g127 (n151, n58);
not  g128 (n183, n10);
not  g129 (n185, n66);
buf  g130 (n169, n64);
buf  g131 (n161, n45);
not  g132 (n92, n73);
not  g133 (n109, n40);
not  g134 (n93, n59);
buf  g135 (n85, n9);
buf  g136 (n131, n74);
not  g137 (n122, n71);
not  g138 (n163, n51);
buf  g139 (n88, n62);
not  g140 (n82, n43);
buf  g141 (n146, n75);
buf  g142 (n193, n40);
buf  g143 (n158, n37);
not  g144 (n152, n50);
buf  g145 (n100, n49);
not  g146 (n140, n71);
buf  g147 (n110, n49);
buf  g148 (n186, n38);
buf  g149 (n191, n57);
not  g150 (n119, n43);
not  g151 (n198, n37);
not  g152 (n194, n37);
not  g153 (n180, n46);
buf  g154 (n162, n48);
buf  g155 (n83, n48);
not  g156 (n148, n66);
buf  g157 (n195, n13);
not  g158 (n95, n54);
not  g159 (n204, n10);
buf  g160 (n86, n14);
buf  g161 (n189, n75);
buf  g162 (n175, n55);
not  g163 (n187, n39);
buf  g164 (n200, n35);
buf  g165 (n168, n73);
not  g166 (n172, n34);
not  g167 (n190, n53);
buf  g168 (n171, n72);
not  g169 (n115, n68);
not  g170 (n79, n61);
buf  g171 (n177, n15);
not  g172 (n153, n33);
nor  g173 (n144, n16, n17);
xor  g174 (n105, n57, n6, n38, n36);
or   g175 (n164, n70, n56, n11, n50);
xor  g176 (n107, n70, n9, n12, n56);
and  g177 (n103, n17, n55, n68, n46);
nand g178 (n179, n10, n78, n6, n16);
nand g179 (n116, n13, n44, n64, n42);
and  g180 (n121, n7, n51, n64, n72);
and  g181 (n184, n39, n44, n8, n47);
and  g182 (n159, n68, n67, n54, n61);
xor  g183 (n173, n60, n16, n58, n52);
xor  g184 (n167, n76, n12, n63, n67);
or   g185 (n134, n62, n63, n69);
xor  g186 (n113, n56, n36, n12, n51);
nor  g187 (n135, n43, n11, n62, n58);
xnor g188 (n89, n13, n40, n11, n42);
xnor g189 (n220, n121, n135, n101, n184);
and  g190 (n222, n204, n199, n196, n119);
nand g191 (n213, n87, n126, n206, n194);
or   g192 (n208, n139, n120, n92, n183);
and  g193 (n219, n154, n198, n202, n163);
and  g194 (n232, n109, n107, n96, n146);
and  g195 (n225, n178, n158, n160, n102);
xnor g196 (n227, n179, n157, n145, n192);
nand g197 (n210, n83, n85, n193, n190);
and  g198 (n218, n86, n182, n156, n148);
xnor g199 (n231, n99, n162, n128, n147);
xor  g200 (n214, n169, n116, n88, n165);
and  g201 (n224, n98, n79, n123, n143);
and  g202 (n238, n104, n134, n132, n108);
nand g203 (n237, n136, n131, n176, n172);
or   g204 (n223, n170, n175, n106, n140);
or   g205 (n216, n186, n166, n168, n82);
and  g206 (n209, n110, n94, n173, n124);
and  g207 (n211, n115, n138, n153, n149);
and  g208 (n215, n195, n111, n137, n100);
nand g209 (n229, n129, n197, n114, n95);
xnor g210 (n234, n151, n122, n91, n81);
nand g211 (n212, n167, n150, n185, n171);
xnor g212 (n217, n187, n103, n152, n203);
and  g213 (n235, n177, n105, n181, n113);
and  g214 (n221, n84, n130, n191, n141);
and  g215 (n230, n188, n161, n200, n180);
or   g216 (n236, n144, n89, n118, n142);
xnor g217 (n226, n112, n125, n97, n164);
nor  g218 (n233, n90, n127, n189, n93);
xor  g219 (n207, n159, n117, n80, n174);
and  g220 (n228, n201, n133, n155, n205);
endmodule
