

module Stat_1162_33_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n805,
  n830,
  n820,
  n809,
  n799,
  n821,
  n831,
  n829,
  n816,
  n832,
  n817,
  n801,
  n813,
  n827,
  n806,
  n804,
  n828,
  n800,
  n798,
  n796,
  n797,
  n1018,
  n1029,
  n1019,
  n1025,
  n1024,
  n1030,
  n1028,
  n1042,
  n1180,
  n1181,
  n1169,
  n1178,
  n1175,
  n1183,
  n1166,
  n1171,
  n1167,
  n1174,
  n1170,
  n1179,
  n1173,
  n1168,
  n1172,
  n1177,
  n1182,
  n1176,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n805;
  output n830;
  output n820;
  output n809;
  output n799;
  output n821;
  output n831;
  output n829;
  output n816;
  output n832;
  output n817;
  output n801;
  output n813;
  output n827;
  output n806;
  output n804;
  output n828;
  output n800;
  output n798;
  output n796;
  output n797;
  output n1018;
  output n1029;
  output n1019;
  output n1025;
  output n1024;
  output n1030;
  output n1028;
  output n1042;
  output n1180;
  output n1181;
  output n1169;
  output n1178;
  output n1175;
  output n1183;
  output n1166;
  output n1171;
  output n1167;
  output n1174;
  output n1170;
  output n1179;
  output n1173;
  output n1168;
  output n1172;
  output n1177;
  output n1182;
  output n1176;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n802;
  wire n803;
  wire n807;
  wire n808;
  wire n810;
  wire n811;
  wire n812;
  wire n814;
  wire n815;
  wire n818;
  wire n819;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1026;
  wire n1027;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n92,
    n13
  );


  buf
  g1
  (
    n71,
    n12
  );


  buf
  g2
  (
    n24,
    n10
  );


  buf
  g3
  (
    n42,
    n15
  );


  not
  g4
  (
    n101,
    n17
  );


  buf
  g5
  (
    n25,
    n17
  );


  buf
  g6
  (
    n45,
    n21
  );


  not
  g7
  (
    n93,
    n17
  );


  buf
  g8
  (
    n54,
    n13
  );


  buf
  g9
  (
    n39,
    n19
  );


  not
  g10
  (
    n38,
    n4
  );


  not
  g11
  (
    n63,
    n4
  );


  not
  g12
  (
    n84,
    n7
  );


  not
  g13
  (
    n105,
    n2
  );


  buf
  g14
  (
    n88,
    n14
  );


  buf
  g15
  (
    n58,
    n19
  );


  not
  g16
  (
    n95,
    n5
  );


  not
  g17
  (
    n40,
    n9
  );


  not
  g18
  (
    n23,
    n3
  );


  buf
  g19
  (
    n64,
    n1
  );


  buf
  g20
  (
    n81,
    n2
  );


  not
  g21
  (
    n57,
    n6
  );


  buf
  g22
  (
    n73,
    n8
  );


  not
  g23
  (
    n37,
    n12
  );


  buf
  g24
  (
    n79,
    n19
  );


  buf
  g25
  (
    n48,
    n14
  );


  not
  g26
  (
    n30,
    n9
  );


  buf
  g27
  (
    n27,
    n9
  );


  buf
  g28
  (
    n99,
    n10
  );


  buf
  g29
  (
    n46,
    n3
  );


  not
  g30
  (
    n98,
    n11
  );


  not
  g31
  (
    n80,
    n11
  );


  not
  g32
  (
    n62,
    n8
  );


  not
  g33
  (
    n86,
    n14
  );


  not
  g34
  (
    n26,
    n16
  );


  not
  g35
  (
    n100,
    n21
  );


  not
  g36
  (
    n60,
    n20
  );


  buf
  g37
  (
    n31,
    n7
  );


  not
  g38
  (
    n65,
    n8
  );


  buf
  g39
  (
    n75,
    n10
  );


  buf
  g40
  (
    n102,
    n11
  );


  buf
  g41
  (
    n41,
    n16
  );


  buf
  g42
  (
    n90,
    n1
  );


  not
  g43
  (
    n52,
    n5
  );


  not
  g44
  (
    n103,
    n4
  );


  not
  g45
  (
    n50,
    n6
  );


  not
  g46
  (
    n28,
    n14
  );


  not
  g47
  (
    n94,
    n18
  );


  buf
  g48
  (
    n44,
    n7
  );


  buf
  g49
  (
    n59,
    n20
  );


  buf
  g50
  (
    n83,
    n15
  );


  buf
  g51
  (
    n89,
    n2
  );


  not
  g52
  (
    n72,
    n4
  );


  not
  g53
  (
    n69,
    n11
  );


  buf
  g54
  (
    n33,
    n19
  );


  not
  g55
  (
    n87,
    n17
  );


  not
  g56
  (
    n70,
    n1
  );


  not
  g57
  (
    n34,
    n18
  );


  buf
  g58
  (
    n76,
    n16
  );


  buf
  g59
  (
    n47,
    n20
  );


  not
  g60
  (
    n67,
    n9
  );


  buf
  g61
  (
    n91,
    n1
  );


  not
  g62
  (
    n66,
    n15
  );


  buf
  g63
  (
    n43,
    n12
  );


  buf
  g64
  (
    n35,
    n18
  );


  buf
  g65
  (
    n55,
    n5
  );


  buf
  g66
  (
    n96,
    n7
  );


  buf
  g67
  (
    n77,
    n10
  );


  buf
  g68
  (
    n74,
    n5
  );


  buf
  g69
  (
    n68,
    n21
  );


  not
  g70
  (
    n36,
    n2
  );


  buf
  g71
  (
    n32,
    n20
  );


  buf
  g72
  (
    n82,
    n6
  );


  buf
  g73
  (
    n56,
    n8
  );


  not
  g74
  (
    n85,
    n18
  );


  buf
  g75
  (
    n97,
    n6
  );


  not
  g76
  (
    n78,
    n12
  );


  not
  g77
  (
    n22,
    n13
  );


  buf
  g78
  (
    KeyWire_0_3,
    n3
  );


  buf
  g79
  (
    n53,
    n21
  );


  not
  g80
  (
    n51,
    n16
  );


  not
  g81
  (
    n29,
    n15
  );


  not
  g82
  (
    n104,
    n13
  );


  buf
  g83
  (
    n49,
    n3
  );


  buf
  g84
  (
    n161,
    n74
  );


  buf
  g85
  (
    n199,
    n36
  );


  buf
  g86
  (
    n379,
    n88
  );


  buf
  g87
  (
    n256,
    n54
  );


  not
  g88
  (
    n343,
    n35
  );


  buf
  g89
  (
    n310,
    n56
  );


  not
  g90
  (
    n368,
    n31
  );


  not
  g91
  (
    n254,
    n89
  );


  buf
  g92
  (
    n266,
    n90
  );


  not
  g93
  (
    n311,
    n52
  );


  not
  g94
  (
    n260,
    n51
  );


  buf
  g95
  (
    n295,
    n72
  );


  buf
  g96
  (
    n158,
    n69
  );


  buf
  g97
  (
    n120,
    n28
  );


  buf
  g98
  (
    n276,
    n74
  );


  not
  g99
  (
    n187,
    n55
  );


  buf
  g100
  (
    n306,
    n72
  );


  not
  g101
  (
    n319,
    n67
  );


  buf
  g102
  (
    n148,
    n82
  );


  not
  g103
  (
    n348,
    n71
  );


  buf
  g104
  (
    n272,
    n62
  );


  not
  g105
  (
    n395,
    n93
  );


  buf
  g106
  (
    n173,
    n37
  );


  not
  g107
  (
    n229,
    n93
  );


  not
  g108
  (
    n278,
    n80
  );


  not
  g109
  (
    n134,
    n52
  );


  buf
  g110
  (
    n154,
    n51
  );


  not
  g111
  (
    n322,
    n84
  );


  not
  g112
  (
    n303,
    n86
  );


  not
  g113
  (
    n338,
    n42
  );


  buf
  g114
  (
    n108,
    n89
  );


  not
  g115
  (
    n224,
    n22
  );


  not
  g116
  (
    n414,
    n37
  );


  buf
  g117
  (
    n222,
    n41
  );


  not
  g118
  (
    n235,
    n74
  );


  buf
  g119
  (
    n172,
    n98
  );


  buf
  g120
  (
    n298,
    n34
  );


  buf
  g121
  (
    n160,
    n65
  );


  buf
  g122
  (
    n234,
    n56
  );


  buf
  g123
  (
    n225,
    n80
  );


  not
  g124
  (
    n334,
    n26
  );


  not
  g125
  (
    n205,
    n33
  );


  buf
  g126
  (
    n244,
    n55
  );


  not
  g127
  (
    n230,
    n94
  );


  not
  g128
  (
    n221,
    n94
  );


  not
  g129
  (
    n378,
    n86
  );


  buf
  g130
  (
    n359,
    n67
  );


  not
  g131
  (
    n410,
    n57
  );


  not
  g132
  (
    n141,
    n27
  );


  not
  g133
  (
    n189,
    n77
  );


  buf
  g134
  (
    n243,
    n70
  );


  not
  g135
  (
    n128,
    n77
  );


  buf
  g136
  (
    n372,
    n62
  );


  not
  g137
  (
    n227,
    n26
  );


  buf
  g138
  (
    n137,
    n45
  );


  not
  g139
  (
    n363,
    n44
  );


  not
  g140
  (
    n146,
    n54
  );


  not
  g141
  (
    n320,
    n81
  );


  buf
  g142
  (
    n316,
    n42
  );


  not
  g143
  (
    n389,
    n79
  );


  buf
  g144
  (
    n210,
    n62
  );


  buf
  g145
  (
    n331,
    n60
  );


  buf
  g146
  (
    n294,
    n25
  );


  buf
  g147
  (
    n408,
    n90
  );


  not
  g148
  (
    n127,
    n41
  );


  not
  g149
  (
    n309,
    n44
  );


  not
  g150
  (
    n250,
    n31
  );


  buf
  g151
  (
    n117,
    n87
  );


  not
  g152
  (
    n124,
    n60
  );


  buf
  g153
  (
    n197,
    n54
  );


  buf
  g154
  (
    n107,
    n95
  );


  buf
  g155
  (
    n126,
    n87
  );


  buf
  g156
  (
    n238,
    n38
  );


  buf
  g157
  (
    n366,
    n82
  );


  not
  g158
  (
    n125,
    n70
  );


  not
  g159
  (
    n269,
    n34
  );


  buf
  g160
  (
    n390,
    n40
  );


  not
  g161
  (
    n214,
    n23
  );


  buf
  g162
  (
    n301,
    n50
  );


  not
  g163
  (
    n209,
    n28
  );


  not
  g164
  (
    n293,
    n67
  );


  not
  g165
  (
    KeyWire_0_11,
    n47
  );


  buf
  g166
  (
    n394,
    n75
  );


  not
  g167
  (
    n195,
    n32
  );


  not
  g168
  (
    n178,
    n79
  );


  not
  g169
  (
    n371,
    n56
  );


  buf
  g170
  (
    n190,
    n32
  );


  not
  g171
  (
    n259,
    n54
  );


  not
  g172
  (
    n242,
    n48
  );


  not
  g173
  (
    n155,
    n84
  );


  buf
  g174
  (
    n404,
    n57
  );


  buf
  g175
  (
    n347,
    n30
  );


  buf
  g176
  (
    n282,
    n78
  );


  not
  g177
  (
    n418,
    n76
  );


  buf
  g178
  (
    n198,
    n47
  );


  not
  g179
  (
    n168,
    n75
  );


  buf
  g180
  (
    n383,
    n70
  );


  not
  g181
  (
    n204,
    n72
  );


  not
  g182
  (
    n240,
    n40
  );


  not
  g183
  (
    KeyWire_0_14,
    n100
  );


  buf
  g184
  (
    n289,
    n85
  );


  buf
  g185
  (
    n133,
    n39
  );


  buf
  g186
  (
    n201,
    n75
  );


  buf
  g187
  (
    n219,
    n46
  );


  not
  g188
  (
    n362,
    n23
  );


  buf
  g189
  (
    n113,
    n79
  );


  buf
  g190
  (
    n318,
    n82
  );


  buf
  g191
  (
    n270,
    n40
  );


  not
  g192
  (
    n370,
    n40
  );


  buf
  g193
  (
    n119,
    n46
  );


  not
  g194
  (
    n220,
    n99
  );


  not
  g195
  (
    n218,
    n52
  );


  not
  g196
  (
    n236,
    n68
  );


  not
  g197
  (
    n180,
    n28
  );


  buf
  g198
  (
    n246,
    n42
  );


  buf
  g199
  (
    n162,
    n83
  );


  not
  g200
  (
    n118,
    n98
  );


  buf
  g201
  (
    n203,
    n61
  );


  buf
  g202
  (
    n279,
    n64
  );


  not
  g203
  (
    n336,
    n99
  );


  not
  g204
  (
    n349,
    n59
  );


  buf
  g205
  (
    n267,
    n23
  );


  not
  g206
  (
    n231,
    n92
  );


  buf
  g207
  (
    n140,
    n89
  );


  not
  g208
  (
    n407,
    n89
  );


  not
  g209
  (
    n129,
    n33
  );


  not
  g210
  (
    n405,
    n22
  );


  not
  g211
  (
    n163,
    n25
  );


  not
  g212
  (
    n340,
    n57
  );


  not
  g213
  (
    n263,
    n66
  );


  buf
  g214
  (
    n109,
    n34
  );


  not
  g215
  (
    n253,
    n47
  );


  not
  g216
  (
    n346,
    n32
  );


  buf
  g217
  (
    n355,
    n92
  );


  buf
  g218
  (
    n403,
    n76
  );


  buf
  g219
  (
    n249,
    n59
  );


  buf
  g220
  (
    n142,
    n97
  );


  not
  g221
  (
    n398,
    n45
  );


  buf
  g222
  (
    n314,
    n86
  );


  not
  g223
  (
    KeyWire_0_10,
    n68
  );


  not
  g224
  (
    n122,
    n49
  );


  not
  g225
  (
    n106,
    n92
  );


  not
  g226
  (
    n159,
    n95
  );


  not
  g227
  (
    n361,
    n29
  );


  not
  g228
  (
    n406,
    n43
  );


  not
  g229
  (
    n115,
    n71
  );


  not
  g230
  (
    n382,
    n84
  );


  buf
  g231
  (
    n354,
    n77
  );


  buf
  g232
  (
    n182,
    n64
  );


  buf
  g233
  (
    n111,
    n30
  );


  buf
  g234
  (
    n364,
    n35
  );


  buf
  g235
  (
    n143,
    n27
  );


  not
  g236
  (
    n174,
    n80
  );


  buf
  g237
  (
    n200,
    n98
  );


  buf
  g238
  (
    n232,
    n48
  );


  buf
  g239
  (
    n123,
    n53
  );


  not
  g240
  (
    n145,
    n97
  );


  not
  g241
  (
    n393,
    n57
  );


  not
  g242
  (
    n144,
    n78
  );


  not
  g243
  (
    n356,
    n66
  );


  buf
  g244
  (
    n164,
    n24
  );


  buf
  g245
  (
    n329,
    n65
  );


  buf
  g246
  (
    n283,
    n76
  );


  buf
  g247
  (
    n265,
    n95
  );


  not
  g248
  (
    n186,
    n69
  );


  not
  g249
  (
    n341,
    n100
  );


  not
  g250
  (
    n376,
    n74
  );


  buf
  g251
  (
    n400,
    n55
  );


  not
  g252
  (
    n284,
    n76
  );


  not
  g253
  (
    n239,
    n81
  );


  not
  g254
  (
    n360,
    n27
  );


  buf
  g255
  (
    n373,
    n87
  );


  buf
  g256
  (
    n112,
    n34
  );


  not
  g257
  (
    n352,
    n49
  );


  buf
  g258
  (
    n365,
    n66
  );


  buf
  g259
  (
    n288,
    n61
  );


  not
  g260
  (
    n328,
    n37
  );


  buf
  g261
  (
    n110,
    n48
  );


  buf
  g262
  (
    n251,
    n36
  );


  buf
  g263
  (
    n402,
    n64
  );


  buf
  g264
  (
    n374,
    n90
  );


  buf
  g265
  (
    n217,
    n50
  );


  not
  g266
  (
    n177,
    n87
  );


  not
  g267
  (
    n228,
    n53
  );


  not
  g268
  (
    n417,
    n96
  );


  not
  g269
  (
    n317,
    n53
  );


  buf
  g270
  (
    n419,
    n33
  );


  buf
  g271
  (
    n255,
    n99
  );


  not
  g272
  (
    n170,
    n73
  );


  not
  g273
  (
    n138,
    n41
  );


  not
  g274
  (
    n175,
    n67
  );


  buf
  g275
  (
    n335,
    n51
  );


  not
  g276
  (
    n321,
    n60
  );


  buf
  g277
  (
    n252,
    n55
  );


  buf
  g278
  (
    n194,
    n82
  );


  not
  g279
  (
    n241,
    n97
  );


  not
  g280
  (
    n131,
    n69
  );


  not
  g281
  (
    n287,
    n47
  );


  not
  g282
  (
    n152,
    n24
  );


  buf
  g283
  (
    n399,
    n98
  );


  not
  g284
  (
    n233,
    n52
  );


  not
  g285
  (
    n193,
    n48
  );


  not
  g286
  (
    n292,
    n50
  );


  buf
  g287
  (
    n345,
    n73
  );


  buf
  g288
  (
    n299,
    n42
  );


  not
  g289
  (
    n271,
    n31
  );


  buf
  g290
  (
    n313,
    n65
  );


  buf
  g291
  (
    n325,
    n83
  );


  not
  g292
  (
    n377,
    n63
  );


  buf
  g293
  (
    n304,
    n96
  );


  buf
  g294
  (
    n327,
    n49
  );


  not
  g295
  (
    n184,
    n83
  );


  not
  g296
  (
    n291,
    n24
  );


  buf
  g297
  (
    n409,
    n43
  );


  buf
  g298
  (
    n237,
    n85
  );


  buf
  g299
  (
    n185,
    n91
  );


  buf
  g300
  (
    n333,
    n51
  );


  not
  g301
  (
    n273,
    n92
  );


  not
  g302
  (
    n135,
    n45
  );


  not
  g303
  (
    n324,
    n32
  );


  buf
  g304
  (
    KeyWire_0_12,
    n65
  );


  not
  g305
  (
    n387,
    n90
  );


  buf
  g306
  (
    n312,
    n99
  );


  not
  g307
  (
    n416,
    n73
  );


  buf
  g308
  (
    n380,
    n94
  );


  buf
  g309
  (
    n188,
    n44
  );


  not
  g310
  (
    n392,
    n39
  );


  buf
  g311
  (
    n257,
    n64
  );


  not
  g312
  (
    n281,
    n78
  );


  not
  g313
  (
    n192,
    n56
  );


  not
  g314
  (
    n176,
    n71
  );


  not
  g315
  (
    n297,
    n50
  );


  not
  g316
  (
    n196,
    n49
  );


  buf
  g317
  (
    n171,
    n43
  );


  buf
  g318
  (
    n339,
    n46
  );


  buf
  g319
  (
    n290,
    n63
  );


  not
  g320
  (
    n315,
    n58
  );


  buf
  g321
  (
    n344,
    n37
  );


  buf
  g322
  (
    n330,
    n85
  );


  buf
  g323
  (
    n121,
    n85
  );


  buf
  g324
  (
    n413,
    n94
  );


  buf
  g325
  (
    KeyWire_0_2,
    n91
  );


  not
  g326
  (
    n147,
    n24
  );


  buf
  g327
  (
    n226,
    n26
  );


  not
  g328
  (
    n307,
    n80
  );


  not
  g329
  (
    n275,
    n68
  );


  buf
  g330
  (
    n114,
    n78
  );


  not
  g331
  (
    n156,
    n26
  );


  not
  g332
  (
    n277,
    n77
  );


  not
  g333
  (
    n150,
    n33
  );


  not
  g334
  (
    n167,
    n22
  );


  not
  g335
  (
    n342,
    n39
  );


  buf
  g336
  (
    n216,
    n35
  );


  buf
  g337
  (
    n211,
    n29
  );


  not
  g338
  (
    n386,
    n58
  );


  buf
  g339
  (
    n262,
    n88
  );


  not
  g340
  (
    n261,
    n81
  );


  buf
  g341
  (
    n358,
    n38
  );


  not
  g342
  (
    n337,
    n83
  );


  buf
  g343
  (
    n367,
    n75
  );


  not
  g344
  (
    n353,
    n41
  );


  not
  g345
  (
    n212,
    n59
  );


  not
  g346
  (
    n308,
    n36
  );


  not
  g347
  (
    n130,
    n22
  );


  not
  g348
  (
    n351,
    n35
  );


  not
  g349
  (
    n165,
    n62
  );


  buf
  g350
  (
    KeyWire_0_8,
    n46
  );


  buf
  g351
  (
    n202,
    n70
  );


  not
  g352
  (
    n396,
    n59
  );


  not
  g353
  (
    n248,
    n29
  );


  not
  g354
  (
    n215,
    n66
  );


  not
  g355
  (
    n397,
    n84
  );


  not
  g356
  (
    n350,
    n81
  );


  buf
  g357
  (
    n132,
    n38
  );


  buf
  g358
  (
    n305,
    n63
  );


  not
  g359
  (
    n116,
    n44
  );


  not
  g360
  (
    n285,
    n88
  );


  not
  g361
  (
    n153,
    n29
  );


  buf
  g362
  (
    n191,
    n73
  );


  not
  g363
  (
    n206,
    n63
  );


  buf
  g364
  (
    n391,
    n86
  );


  not
  g365
  (
    n179,
    n27
  );


  not
  g366
  (
    n384,
    n30
  );


  buf
  g367
  (
    n385,
    n96
  );


  not
  g368
  (
    n332,
    n58
  );


  not
  g369
  (
    n401,
    n93
  );


  not
  g370
  (
    n286,
    n58
  );


  buf
  g371
  (
    n136,
    n91
  );


  not
  g372
  (
    n245,
    n61
  );


  buf
  g373
  (
    n166,
    n25
  );


  not
  g374
  (
    n223,
    n91
  );


  not
  g375
  (
    n149,
    n93
  );


  buf
  g376
  (
    n412,
    n53
  );


  not
  g377
  (
    n169,
    n23
  );


  buf
  g378
  (
    n264,
    n97
  );


  buf
  g379
  (
    n388,
    n96
  );


  not
  g380
  (
    n213,
    n72
  );


  buf
  g381
  (
    n181,
    n61
  );


  not
  g382
  (
    n381,
    n43
  );


  not
  g383
  (
    n207,
    n39
  );


  not
  g384
  (
    n151,
    n25
  );


  buf
  g385
  (
    n208,
    n71
  );


  not
  g386
  (
    n326,
    n36
  );


  buf
  g387
  (
    n296,
    n88
  );


  not
  g388
  (
    n247,
    n38
  );


  buf
  g389
  (
    n274,
    n95
  );


  buf
  g390
  (
    n302,
    n79
  );


  buf
  g391
  (
    n357,
    n68
  );


  not
  g392
  (
    n268,
    n69
  );


  not
  g393
  (
    n157,
    n30
  );


  not
  g394
  (
    n411,
    n60
  );


  not
  g395
  (
    n139,
    n45
  );


  buf
  g396
  (
    n300,
    n31
  );


  not
  g397
  (
    n415,
    n28
  );


  buf
  g398
  (
    n432,
    n113
  );


  not
  g399
  (
    n467,
    n232
  );


  buf
  g400
  (
    n663,
    n231
  );


  not
  g401
  (
    n566,
    n111
  );


  not
  g402
  (
    n607,
    n239
  );


  not
  g403
  (
    n537,
    n178
  );


  not
  g404
  (
    n481,
    n321
  );


  not
  g405
  (
    n435,
    n261
  );


  buf
  g406
  (
    n454,
    n305
  );


  buf
  g407
  (
    n611,
    n349
  );


  buf
  g408
  (
    n501,
    n142
  );


  buf
  g409
  (
    n606,
    n133
  );


  xor
  g410
  (
    n655,
    n348,
    n255,
    n276,
    n134
  );


  nor
  g411
  (
    n688,
    n263,
    n337,
    n277,
    n351
  );


  and
  g412
  (
    n686,
    n249,
    n223,
    n246,
    n354
  );


  and
  g413
  (
    n536,
    n146,
    n111,
    n368,
    n230
  );


  xor
  g414
  (
    n547,
    n192,
    n160,
    n300,
    n190
  );


  xnor
  g415
  (
    n565,
    n298,
    n157,
    n297,
    n204
  );


  xnor
  g416
  (
    n461,
    n256,
    n360,
    n191,
    n335
  );


  or
  g417
  (
    n570,
    n233,
    n307,
    n337,
    n278
  );


  or
  g418
  (
    n690,
    n348,
    n179,
    n308,
    n299
  );


  and
  g419
  (
    n557,
    n181,
    n240,
    n329,
    n323
  );


  nor
  g420
  (
    n603,
    n258,
    n198,
    n359,
    n313
  );


  xor
  g421
  (
    n499,
    n235,
    n290,
    n205,
    n316
  );


  nand
  g422
  (
    n476,
    n216,
    n265,
    n318,
    n243
  );


  xnor
  g423
  (
    n605,
    n346,
    n337,
    n214,
    n223
  );


  nor
  g424
  (
    n666,
    n279,
    n156,
    n344,
    n153
  );


  and
  g425
  (
    n586,
    n315,
    n106,
    n254,
    n212
  );


  xor
  g426
  (
    n575,
    n249,
    n315,
    n127,
    n322
  );


  and
  g427
  (
    n609,
    n352,
    n279,
    n201,
    n145
  );


  and
  g428
  (
    n520,
    n249,
    n106,
    n210,
    n358
  );


  xnor
  g429
  (
    n629,
    n131,
    n347,
    n294,
    n278
  );


  nor
  g430
  (
    n583,
    n253,
    n352,
    n344,
    n203
  );


  nand
  g431
  (
    n525,
    n270,
    n281,
    n228,
    n157
  );


  nor
  g432
  (
    n524,
    n231,
    n125,
    n322,
    n325
  );


  xor
  g433
  (
    n431,
    n341,
    n264,
    n118,
    n190
  );


  xor
  g434
  (
    n612,
    n272,
    n171,
    n319,
    n139
  );


  xnor
  g435
  (
    n594,
    n253,
    n239,
    n233,
    n310
  );


  xnor
  g436
  (
    n692,
    n285,
    n330,
    n226,
    n224
  );


  nor
  g437
  (
    n523,
    n326,
    n286,
    n291,
    n312
  );


  xor
  g438
  (
    n533,
    n364,
    n340,
    n288,
    n363
  );


  nor
  g439
  (
    n452,
    n184,
    n214,
    n205,
    n260
  );


  or
  g440
  (
    n545,
    n364,
    n212,
    n227,
    n243
  );


  xor
  g441
  (
    n538,
    n193,
    n342,
    n119,
    n267
  );


  xor
  g442
  (
    n555,
    n226,
    n279,
    n347,
    n266
  );


  nand
  g443
  (
    n643,
    n158,
    n272,
    n112,
    n171
  );


  or
  g444
  (
    n477,
    n303,
    n340,
    n270,
    n108
  );


  nor
  g445
  (
    n447,
    n345,
    n134,
    n174,
    n236
  );


  xor
  g446
  (
    n656,
    n369,
    n273,
    n190,
    n276
  );


  or
  g447
  (
    n683,
    n237,
    n286,
    n123,
    n269
  );


  xor
  g448
  (
    n622,
    n139,
    n229,
    n133,
    n221
  );


  and
  g449
  (
    n597,
    n154,
    n361,
    n290,
    n282
  );


  or
  g450
  (
    n680,
    n117,
    n210,
    n129,
    n339
  );


  xnor
  g451
  (
    n549,
    n296,
    n269,
    n229,
    n262
  );


  and
  g452
  (
    n584,
    n223,
    n145,
    n149,
    n332
  );


  nor
  g453
  (
    n436,
    n126,
    n367,
    n331,
    n362
  );


  and
  g454
  (
    n540,
    n341,
    n262,
    n177,
    n235
  );


  or
  g455
  (
    n556,
    n222,
    n356,
    n237,
    n315
  );


  or
  g456
  (
    n496,
    n111,
    n186,
    n132,
    n295
  );


  nor
  g457
  (
    n571,
    n325,
    n199,
    n178,
    n212
  );


  or
  g458
  (
    n430,
    n328,
    n343,
    n175,
    n280
  );


  and
  g459
  (
    n553,
    n351,
    n179,
    n152,
    n313
  );


  and
  g460
  (
    n681,
    n242,
    n302,
    n328,
    n179
  );


  nand
  g461
  (
    n649,
    n132,
    n340,
    n220,
    n224
  );


  xor
  g462
  (
    n652,
    n313,
    n300,
    n200,
    n196
  );


  nand
  g463
  (
    n478,
    n302,
    n168,
    n352,
    n272
  );


  xor
  g464
  (
    n591,
    n281,
    n326,
    n300,
    n368
  );


  or
  g465
  (
    n685,
    n219,
    n210,
    n136,
    n339
  );


  or
  g466
  (
    n624,
    n291,
    n327,
    n161,
    n345
  );


  and
  g467
  (
    n492,
    n219,
    n301,
    n262,
    n195
  );


  xor
  g468
  (
    n574,
    n321,
    n363,
    n355,
    n311
  );


  nor
  g469
  (
    n626,
    n186,
    n261,
    n116,
    n231
  );


  xnor
  g470
  (
    n665,
    n352,
    n153,
    n362,
    n175
  );


  xor
  g471
  (
    n651,
    n242,
    n131,
    n261,
    n130
  );


  and
  g472
  (
    n422,
    n266,
    n277,
    n159,
    n129
  );


  or
  g473
  (
    n516,
    n314,
    n256,
    n275,
    n147
  );


  or
  g474
  (
    n608,
    n333,
    n249,
    n309,
    n263
  );


  nor
  g475
  (
    n588,
    n197,
    n296,
    n305,
    n198
  );


  xnor
  g476
  (
    n669,
    n236,
    n362,
    n167,
    n324
  );


  and
  g477
  (
    n635,
    n283,
    n167,
    n181,
    n164
  );


  xnor
  g478
  (
    n488,
    n338,
    n245,
    n154,
    n295
  );


  or
  g479
  (
    n582,
    n127,
    n229,
    n194,
    n224
  );


  or
  g480
  (
    n564,
    n322,
    n298,
    n204,
    n144
  );


  nand
  g481
  (
    n682,
    n120,
    n143,
    n246,
    n187
  );


  nor
  g482
  (
    n676,
    n182,
    n239,
    n167,
    n355
  );


  xnor
  g483
  (
    n433,
    n365,
    n168,
    n216,
    n180
  );


  and
  g484
  (
    n456,
    n271,
    n264,
    n228,
    n293
  );


  nand
  g485
  (
    n465,
    n304,
    n228,
    n199,
    n298
  );


  nor
  g486
  (
    n577,
    n363,
    n252,
    n343,
    n204
  );


  nor
  g487
  (
    n562,
    n345,
    n235,
    n244,
    n361
  );


  xor
  g488
  (
    n617,
    n367,
    n113,
    n271,
    n366
  );


  or
  g489
  (
    n560,
    n250,
    n227,
    n177,
    n137
  );


  nor
  g490
  (
    n552,
    n184,
    n176,
    n146,
    n234
  );


  or
  g491
  (
    n463,
    n230,
    n217,
    n283,
    n247
  );


  nor
  g492
  (
    n502,
    n236,
    n335,
    n189,
    n248
  );


  xor
  g493
  (
    n627,
    n213,
    n111,
    n152,
    n215
  );


  nand
  g494
  (
    n595,
    n302,
    n164,
    n242,
    n174
  );


  and
  g495
  (
    n468,
    n355,
    n360,
    n198,
    n250
  );


  or
  g496
  (
    n678,
    n234,
    n287,
    n230,
    n118
  );


  or
  g497
  (
    n535,
    n368,
    n334,
    n257,
    n156
  );


  nand
  g498
  (
    n512,
    n143,
    n323,
    n135,
    n349
  );


  xor
  g499
  (
    n675,
    n247,
    n107,
    n333,
    n141
  );


  and
  g500
  (
    n539,
    n238,
    n337,
    n360,
    n308
  );


  nand
  g501
  (
    n646,
    n248,
    n217,
    n290,
    n209
  );


  xor
  g502
  (
    n542,
    n339,
    n244,
    n260,
    n209
  );


  nor
  g503
  (
    n509,
    n165,
    n113,
    n319,
    n360
  );


  xnor
  g504
  (
    n519,
    n273,
    n329,
    n288,
    n196
  );


  nand
  g505
  (
    n424,
    n345,
    n299,
    n281,
    n338
  );


  nand
  g506
  (
    n510,
    n247,
    n366,
    n262,
    n127
  );


  nand
  g507
  (
    n670,
    n128,
    n112,
    n286,
    n246
  );


  nand
  g508
  (
    n650,
    n122,
    n126,
    n201,
    n169
  );


  and
  g509
  (
    n647,
    n251,
    n346,
    n168,
    n283
  );


  or
  g510
  (
    n471,
    n347,
    n336,
    n122,
    n178
  );


  xnor
  g511
  (
    n563,
    n124,
    n109,
    n335,
    n126
  );


  nor
  g512
  (
    n448,
    n187,
    n244,
    n342,
    n142
  );


  nand
  g513
  (
    n644,
    n137,
    n221,
    n218,
    n288
  );


  nand
  g514
  (
    n590,
    n133,
    n336,
    n137,
    n146
  );


  nand
  g515
  (
    n440,
    n331,
    n149,
    n260,
    n190
  );


  or
  g516
  (
    n473,
    n172,
    n324,
    n341,
    n204
  );


  xnor
  g517
  (
    n559,
    n181,
    n207,
    n158,
    n164
  );


  nor
  g518
  (
    n446,
    n327,
    n210,
    n160,
    n271
  );


  nand
  g519
  (
    n598,
    n257,
    n303,
    n115,
    n338
  );


  xnor
  g520
  (
    n443,
    n278,
    n150,
    n168,
    n205
  );


  and
  g521
  (
    n439,
    n141,
    n151,
    n273,
    n191
  );


  xnor
  g522
  (
    n593,
    n367,
    n201,
    n208,
    n155
  );


  nand
  g523
  (
    n600,
    n206,
    n233,
    n311,
    n368
  );


  or
  g524
  (
    n687,
    n330,
    n280,
    n174,
    n317
  );


  xor
  g525
  (
    n518,
    n183,
    n267,
    n159,
    n255
  );


  or
  g526
  (
    n462,
    n114,
    n268,
    n251,
    n257
  );


  or
  g527
  (
    n489,
    n207,
    n236,
    n254,
    n211
  );


  or
  g528
  (
    n618,
    n333,
    n177,
    n182,
    n340
  );


  nand
  g529
  (
    n475,
    n240,
    n261,
    n317,
    n125
  );


  xor
  g530
  (
    n581,
    n280,
    n116,
    n163,
    n294
  );


  xor
  g531
  (
    n569,
    n154,
    n175,
    n167,
    n172
  );


  nor
  g532
  (
    n585,
    n180,
    n330,
    n183,
    n306
  );


  and
  g533
  (
    n455,
    n161,
    n275,
    n215,
    n292
  );


  nor
  g534
  (
    n427,
    n274,
    n108,
    n346,
    n211
  );


  xor
  g535
  (
    n548,
    n225,
    n171,
    n234,
    n117
  );


  xor
  g536
  (
    n561,
    n118,
    n356,
    n221,
    n309
  );


  xnor
  g537
  (
    n576,
    n330,
    n335,
    n138,
    n240
  );


  or
  g538
  (
    n531,
    n365,
    n243,
    n323,
    n142
  );


  nor
  g539
  (
    n671,
    n192,
    n124,
    n306,
    n284
  );


  xor
  g540
  (
    n628,
    n241,
    n119,
    n285,
    n320
  );


  nor
  g541
  (
    n495,
    n171,
    n282,
    n197,
    n267
  );


  nor
  g542
  (
    n483,
    n198,
    n271,
    n258,
    n159
  );


  nor
  g543
  (
    n469,
    n234,
    n281,
    n333,
    n274
  );


  xor
  g544
  (
    n485,
    n275,
    n121,
    n276,
    n129
  );


  xor
  g545
  (
    n658,
    n115,
    n341,
    n110,
    n208
  );


  xor
  g546
  (
    n444,
    n191,
    n127,
    n299,
    n259
  );


  xor
  g547
  (
    n638,
    n334,
    n131,
    n216,
    n367
  );


  or
  g548
  (
    n558,
    n359,
    n169,
    n138,
    n346
  );


  xnor
  g549
  (
    n551,
    n233,
    n128,
    n219,
    n134
  );


  xnor
  g550
  (
    n480,
    n219,
    n229,
    n230,
    n123
  );


  and
  g551
  (
    n526,
    n254,
    n301,
    n165,
    n296
  );


  or
  g552
  (
    n550,
    n318,
    n324,
    n290,
    n277
  );


  or
  g553
  (
    n679,
    n185,
    n359,
    n194,
    n269
  );


  nor
  g554
  (
    n451,
    n303,
    n295,
    n354,
    n292
  );


  nor
  g555
  (
    n640,
    n310,
    n228,
    n119,
    n156
  );


  or
  g556
  (
    n623,
    n263,
    n302,
    n196,
    n301
  );


  xor
  g557
  (
    n653,
    n300,
    n170,
    n121,
    n265
  );


  nand
  g558
  (
    n580,
    n176,
    n158,
    n321,
    n180
  );


  and
  g559
  (
    n657,
    n358,
    n304,
    n148,
    n110
  );


  and
  g560
  (
    n472,
    n259,
    n209,
    n369,
    n162
  );


  and
  g561
  (
    n677,
    n213,
    n189,
    n114,
    n157
  );


  xnor
  g562
  (
    n592,
    n160,
    n312,
    n237,
    n307
  );


  nand
  g563
  (
    n601,
    n112,
    n160,
    n313,
    n140
  );


  nand
  g564
  (
    n482,
    n291,
    n117,
    n215,
    n151
  );


  nor
  g565
  (
    n610,
    n169,
    n231,
    n332,
    n156
  );


  nor
  g566
  (
    n641,
    n214,
    n144,
    n199,
    n310
  );


  or
  g567
  (
    n507,
    n116,
    n151,
    n128,
    n140
  );


  and
  g568
  (
    n554,
    n175,
    n196,
    n143,
    n165
  );


  nor
  g569
  (
    n494,
    n289,
    n320,
    n114,
    n152
  );


  xor
  g570
  (
    n498,
    n188,
    n115,
    n317,
    n357
  );


  xnor
  g571
  (
    n514,
    n213,
    n132,
    n323,
    n259
  );


  xor
  g572
  (
    n645,
    n255,
    n252,
    n182,
    n344
  );


  nor
  g573
  (
    n515,
    n170,
    n241,
    n284,
    n220
  );


  xnor
  g574
  (
    n602,
    n314,
    n130,
    n113,
    n324
  );


  and
  g575
  (
    n506,
    n213,
    n173,
    n320,
    n260
  );


  nand
  g576
  (
    n479,
    n207,
    n194,
    n304,
    n144
  );


  xor
  g577
  (
    n659,
    n241,
    n209,
    n134,
    n221
  );


  nor
  g578
  (
    n460,
    n166,
    n208,
    n278,
    n124
  );


  xnor
  g579
  (
    n428,
    n165,
    n159,
    n148
  );


  nand
  g580
  (
    n613,
    n252,
    n206,
    n135,
    n149
  );


  nand
  g581
  (
    n445,
    n166,
    n270,
    n147,
    n253
  );


  xor
  g582
  (
    n529,
    n218,
    n232,
    n235,
    n179
  );


  nor
  g583
  (
    n505,
    n202,
    n307,
    n157,
    n369
  );


  nand
  g584
  (
    n587,
    n294,
    n266,
    n150,
    n153
  );


  nand
  g585
  (
    n648,
    n268,
    n309,
    n297,
    n336
  );


  nor
  g586
  (
    n426,
    n328,
    n255,
    n125,
    n186
  );


  or
  g587
  (
    n425,
    n288,
    n155,
    n366,
    n166
  );


  xnor
  g588
  (
    n497,
    n354,
    n285,
    n172,
    n222
  );


  xor
  g589
  (
    n484,
    n287,
    n327,
    n269,
    n264
  );


  or
  g590
  (
    n672,
    n344,
    n321,
    n297,
    n258
  );


  or
  g591
  (
    n691,
    n350,
    n152,
    n163,
    n169
  );


  and
  g592
  (
    n474,
    n294,
    n325,
    n147,
    n153
  );


  xnor
  g593
  (
    n621,
    n218,
    n308,
    n365,
    n350
  );


  nor
  g594
  (
    n614,
    n329,
    n164,
    n250,
    n146
  );


  nand
  g595
  (
    n573,
    n136,
    n287,
    n238,
    n161
  );


  xnor
  g596
  (
    n620,
    n224,
    n193,
    n121,
    n155
  );


  xor
  g597
  (
    n636,
    n225,
    n185,
    n108,
    n358
  );


  or
  g598
  (
    n654,
    n317,
    n223,
    n145,
    n245
  );


  and
  g599
  (
    n491,
    n256,
    n336,
    n188,
    n142
  );


  and
  g600
  (
    n500,
    n289,
    n353,
    n128,
    n312
  );


  nand
  g601
  (
    n543,
    n274,
    n149,
    n119,
    n232
  );


  nor
  g602
  (
    n578,
    n200,
    n150,
    n272,
    n222
  );


  and
  g603
  (
    n604,
    n215,
    n172,
    n248,
    n122
  );


  and
  g604
  (
    n637,
    n245,
    n109,
    n217,
    n202
  );


  nand
  g605
  (
    n527,
    n206,
    n240,
    n158,
    n348
  );


  nor
  g606
  (
    n464,
    n220,
    n225,
    n200,
    n147
  );


  xor
  g607
  (
    n511,
    n205,
    n273,
    n264,
    n329
  );


  xnor
  g608
  (
    n616,
    n189,
    n203,
    n339,
    n316
  );


  nor
  g609
  (
    n453,
    n285,
    n293,
    n284,
    n226
  );


  xnor
  g610
  (
    n534,
    n174,
    n189,
    n184,
    n141
  );


  nor
  g611
  (
    n508,
    n162,
    n357,
    n350,
    n187
  );


  nor
  g612
  (
    n667,
    n292,
    n114,
    n181,
    n325
  );


  and
  g613
  (
    n450,
    n202,
    n140,
    n143,
    n115
  );


  or
  g614
  (
    n522,
    n299,
    n349,
    n173,
    n123
  );


  nor
  g615
  (
    n684,
    n348,
    n144,
    n328,
    n136
  );


  nand
  g616
  (
    n458,
    n283,
    n130,
    n138,
    n106
  );


  nor
  g617
  (
    n546,
    n185,
    n188,
    n201,
    n180
  );


  nor
  g618
  (
    n486,
    n246,
    n292,
    n133,
    n351
  );


  xnor
  g619
  (
    n532,
    n139,
    n222,
    n310,
    n135
  );


  nor
  g620
  (
    n420,
    n270,
    n298,
    n268,
    n287
  );


  xnor
  g621
  (
    n503,
    n364,
    n122,
    n151,
    n220
  );


  nor
  g622
  (
    n599,
    n326,
    n163,
    n116,
    n291
  );


  or
  g623
  (
    n504,
    n361,
    n206,
    n289,
    n268
  );


  and
  g624
  (
    n596,
    n191,
    n364,
    n301,
    n245
  );


  xor
  g625
  (
    n457,
    n183,
    n173,
    n320,
    n326
  );


  and
  g626
  (
    n673,
    n289,
    n354,
    n319,
    n106
  );


  nor
  g627
  (
    n625,
    n356,
    n279,
    n194,
    n123
  );


  nand
  g628
  (
    n568,
    n186,
    n331,
    n257,
    n248
  );


  or
  g629
  (
    n634,
    n356,
    n107,
    n243,
    n318
  );


  nand
  g630
  (
    n441,
    n109,
    n120,
    n173,
    n311
  );


  or
  g631
  (
    n674,
    n120,
    n358,
    n365,
    n253
  );


  xor
  g632
  (
    n437,
    n132,
    n218,
    n195,
    n211
  );


  xnor
  g633
  (
    n633,
    n314,
    n139,
    n266,
    n251
  );


  nand
  g634
  (
    n459,
    n316,
    n342,
    n343,
    n314
  );


  and
  g635
  (
    n487,
    n347,
    n296,
    n327,
    n124
  );


  and
  g636
  (
    n429,
    n188,
    n342,
    n305,
    n363
  );


  xnor
  g637
  (
    n572,
    n239,
    n284,
    n161,
    n200
  );


  nor
  g638
  (
    n615,
    n162,
    n125,
    n265,
    n332
  );


  xnor
  g639
  (
    n662,
    n238,
    n267,
    n117,
    n112
  );


  xnor
  g640
  (
    n631,
    n254,
    n286,
    n275,
    n237
  );


  or
  g641
  (
    n642,
    n178,
    n227,
    n357
  );


  and
  g642
  (
    n528,
    n241,
    n322,
    n318,
    n357
  );


  or
  g643
  (
    n661,
    n108,
    n118,
    n334,
    n207
  );


  xor
  g644
  (
    n490,
    n244,
    n148,
    n350,
    n110
  );


  xnor
  g645
  (
    n668,
    n195,
    n110,
    n307,
    n331
  );


  nand
  g646
  (
    n664,
    n135,
    n304,
    n353,
    n176
  );


  nand
  g647
  (
    n423,
    n176,
    n225,
    n319,
    n126
  );


  nand
  g648
  (
    n421,
    n141,
    n192,
    n359,
    n131
  );


  xnor
  g649
  (
    n530,
    n184,
    n250,
    n187,
    n195
  );


  xor
  g650
  (
    n567,
    n129,
    n192,
    n137,
    n155
  );


  xor
  g651
  (
    n517,
    n263,
    n232,
    n136,
    n183
  );


  xnor
  g652
  (
    n541,
    n138,
    n217,
    n305,
    n177
  );


  xnor
  g653
  (
    n521,
    n316,
    n362,
    n280,
    n366
  );


  nand
  g654
  (
    n466,
    n369,
    n277,
    n150,
    n203
  );


  xnor
  g655
  (
    n438,
    n211,
    n226,
    n282,
    n121
  );


  nand
  g656
  (
    n493,
    n353,
    n130,
    n265,
    n256
  );


  or
  g657
  (
    n579,
    n162,
    n259,
    n193,
    n197
  );


  xor
  g658
  (
    n689,
    n274,
    n170,
    n251,
    n349
  );


  nor
  g659
  (
    n589,
    n202,
    n306,
    n242
  );


  xnor
  g660
  (
    n470,
    n107,
    n252,
    n214,
    n120
  );


  xor
  g661
  (
    n619,
    n293,
    n312,
    n309,
    n208
  );


  and
  g662
  (
    n639,
    n163,
    n343,
    n303,
    n193
  );


  or
  g663
  (
    n449,
    n203,
    n351,
    n197,
    n293
  );


  nand
  g664
  (
    KeyWire_0_13,
    n276,
    n140,
    n185,
    n258
  );


  xor
  g665
  (
    n544,
    n166,
    n315,
    n247,
    n308
  );


  and
  g666
  (
    n442,
    n216,
    n154,
    n355,
    n282
  );


  or
  g667
  (
    n513,
    n361,
    n297,
    n170,
    n199
  );


  and
  g668
  (
    n660,
    n145,
    n107,
    n295,
    n238
  );


  xor
  g669
  (
    n630,
    n334,
    n338,
    n311,
    n182
  );


  xor
  g670
  (
    n434,
    n332,
    n109,
    n212,
    n353
  );


  buf
  g671
  (
    n730,
    n446
  );


  buf
  g672
  (
    n708,
    n454
  );


  buf
  g673
  (
    n707,
    n448
  );


  buf
  g674
  (
    n717,
    n458
  );


  buf
  g675
  (
    n732,
    n435
  );


  buf
  g676
  (
    n725,
    n461
  );


  buf
  g677
  (
    n701,
    n452
  );


  not
  g678
  (
    n694,
    n424
  );


  not
  g679
  (
    n711,
    n433
  );


  buf
  g680
  (
    n698,
    n428
  );


  buf
  g681
  (
    n713,
    n423
  );


  not
  g682
  (
    n706,
    n456
  );


  buf
  g683
  (
    n727,
    n450
  );


  not
  g684
  (
    n704,
    n444
  );


  buf
  g685
  (
    n729,
    n431
  );


  not
  g686
  (
    n718,
    n451
  );


  not
  g687
  (
    n709,
    n459
  );


  buf
  g688
  (
    n722,
    n427
  );


  not
  g689
  (
    n719,
    n420
  );


  not
  g690
  (
    n715,
    n460
  );


  not
  g691
  (
    n695,
    n425
  );


  buf
  g692
  (
    n703,
    n426
  );


  buf
  g693
  (
    n723,
    n436
  );


  not
  g694
  (
    n712,
    n437
  );


  buf
  g695
  (
    n720,
    n443
  );


  buf
  g696
  (
    n733,
    n447
  );


  not
  g697
  (
    n734,
    n434
  );


  not
  g698
  (
    n724,
    n442
  );


  buf
  g699
  (
    n714,
    n445
  );


  not
  g700
  (
    n726,
    n421
  );


  not
  g701
  (
    KeyWire_0_5,
    n455
  );


  buf
  g702
  (
    n728,
    n422
  );


  not
  g703
  (
    n697,
    n439
  );


  not
  g704
  (
    n716,
    n457
  );


  buf
  g705
  (
    n702,
    n432
  );


  buf
  g706
  (
    n699,
    n440
  );


  buf
  g707
  (
    n721,
    n453
  );


  not
  g708
  (
    n705,
    n430
  );


  not
  g709
  (
    n696,
    n449
  );


  buf
  g710
  (
    n710,
    n429
  );


  buf
  g711
  (
    n693,
    n438
  );


  not
  g712
  (
    n700,
    n441
  );


  buf
  g713
  (
    n747,
    n695
  );


  not
  g714
  (
    KeyWire_0_1,
    n370
  );


  not
  g715
  (
    n742,
    n473
  );


  not
  g716
  (
    n751,
    n708
  );


  buf
  g717
  (
    n746,
    n699
  );


  not
  g718
  (
    n758,
    n463
  );


  buf
  g719
  (
    n739,
    n712
  );


  buf
  g720
  (
    n755,
    n372
  );


  not
  g721
  (
    n745,
    n468
  );


  not
  g722
  (
    n748,
    n462
  );


  not
  g723
  (
    n752,
    n464
  );


  not
  g724
  (
    n756,
    n693
  );


  not
  g725
  (
    n754,
    n696
  );


  buf
  g726
  (
    n749,
    n370
  );


  buf
  g727
  (
    n750,
    n713
  );


  buf
  g728
  (
    n753,
    n702
  );


  and
  g729
  (
    n735,
    n466,
    n707,
    n714,
    n472
  );


  or
  g730
  (
    n744,
    n465,
    n474,
    n371,
    n705
  );


  and
  g731
  (
    n757,
    n698,
    n370,
    n371,
    n469
  );


  nand
  g732
  (
    n740,
    n475,
    n703,
    n715,
    n710
  );


  nor
  g733
  (
    n738,
    n709,
    n697,
    n371,
    n467
  );


  nor
  g734
  (
    n743,
    n470,
    n476,
    n701,
    n716
  );


  nand
  g735
  (
    n741,
    n694,
    n704,
    n700,
    n706
  );


  xnor
  g736
  (
    n736,
    n471,
    n370,
    n371,
    n711
  );


  buf
  g737
  (
    n760,
    n743
  );


  not
  g738
  (
    n762,
    n737
  );


  buf
  g739
  (
    n764,
    n745
  );


  not
  g740
  (
    n768,
    n735
  );


  not
  g741
  (
    n763,
    n741
  );


  not
  g742
  (
    n769,
    n740
  );


  not
  g743
  (
    n766,
    n478
  );


  buf
  g744
  (
    n765,
    n738
  );


  and
  g745
  (
    n767,
    n482,
    n739
  );


  and
  g746
  (
    n761,
    n736,
    n480,
    n742,
    n481
  );


  or
  g747
  (
    n759,
    n477,
    n744,
    n479,
    n483
  );


  not
  g748
  (
    n776,
    n721
  );


  buf
  g749
  (
    n775,
    n760
  );


  not
  g750
  (
    n770,
    n720
  );


  buf
  g751
  (
    n779,
    n717
  );


  not
  g752
  (
    n773,
    n722
  );


  not
  g753
  (
    n772,
    n759
  );


  not
  g754
  (
    n777,
    n760
  );


  or
  g755
  (
    n778,
    n759,
    n760,
    n761,
    n723
  );


  nor
  g756
  (
    n774,
    n719,
    n718,
    n484,
    n725
  );


  and
  g757
  (
    n771,
    n724,
    n759,
    n761
  );


  buf
  g758
  (
    n788,
    n771
  );


  buf
  g759
  (
    n781,
    n775
  );


  nand
  g760
  (
    n794,
    n772,
    n773
  );


  xor
  g761
  (
    n789,
    n776,
    n747,
    n103,
    n754
  );


  nand
  g762
  (
    n780,
    n487,
    n778,
    n779,
    n746
  );


  or
  g763
  (
    n795,
    n105,
    n101,
    n770,
    n774
  );


  xor
  g764
  (
    n792,
    n104,
    n104,
    n778,
    n486
  );


  and
  g765
  (
    n783,
    n776,
    n751,
    n485,
    n105
  );


  and
  g766
  (
    n790,
    n756,
    n755,
    n748,
    n777
  );


  xor
  g767
  (
    n793,
    n757,
    n102,
    n758,
    n753
  );


  nor
  g768
  (
    n785,
    n750,
    n758,
    n103,
    n101
  );


  nor
  g769
  (
    n787,
    n101,
    n102,
    n100,
    n105
  );


  or
  g770
  (
    n791,
    n749,
    n777,
    n752,
    n775
  );


  nor
  g771
  (
    n782,
    n101,
    n104,
    n105,
    n757
  );


  nor
  g772
  (
    n786,
    n104,
    n103,
    n102
  );


  nand
  g773
  (
    n784,
    n774,
    n103,
    n779,
    n100
  );


  xnor
  g774
  (
    n804,
    n767,
    n783,
    n496
  );


  nand
  g775
  (
    n812,
    n780,
    n503,
    n521
  );


  nor
  g776
  (
    n808,
    n789,
    n786,
    n375,
    n764
  );


  or
  g777
  (
    n810,
    n379,
    n490,
    n781,
    n375
  );


  nand
  g778
  (
    n800,
    n382,
    n489,
    n765,
    n374
  );


  xnor
  g779
  (
    n825,
    n780,
    n762,
    n511,
    n512
  );


  nor
  g780
  (
    n797,
    n500,
    n763,
    n510,
    n377
  );


  xor
  g781
  (
    n813,
    n761,
    n381,
    n488,
    n374
  );


  and
  g782
  (
    n824,
    n494,
    n501,
    n516,
    n787
  );


  and
  g783
  (
    n807,
    n373,
    n762,
    n784,
    n492
  );


  xor
  g784
  (
    n805,
    n508,
    n788,
    n375,
    n784
  );


  nand
  g785
  (
    n815,
    n786,
    n520,
    n504,
    n381
  );


  and
  g786
  (
    n811,
    n782,
    n499,
    n383,
    n498
  );


  nand
  g787
  (
    n827,
    n783,
    n382,
    n380,
    n505
  );


  xor
  g788
  (
    n818,
    n764,
    n507,
    n379,
    n373
  );


  and
  g789
  (
    n799,
    n784,
    n372,
    n768,
    n491
  );


  nand
  g790
  (
    n809,
    n376,
    n787,
    n762,
    n514
  );


  nand
  g791
  (
    n816,
    n788,
    n378,
    n764,
    n783
  );


  or
  g792
  (
    n828,
    n509,
    n376,
    n378
  );


  or
  g793
  (
    n817,
    n785,
    n381,
    n766,
    n379
  );


  nand
  g794
  (
    n822,
    n780,
    n765,
    n788,
    n781
  );


  nand
  g795
  (
    n803,
    n383,
    n786,
    n785,
    n765
  );


  and
  g796
  (
    n830,
    n376,
    n762,
    n782,
    n764
  );


  and
  g797
  (
    n826,
    n380,
    n493,
    n787,
    n767
  );


  and
  g798
  (
    n831,
    n765,
    n378,
    n377
  );


  nor
  g799
  (
    n806,
    n381,
    n372,
    n766,
    n784
  );


  and
  g800
  (
    n801,
    n377,
    n767,
    n376,
    n517
  );


  nand
  g801
  (
    n829,
    n782,
    n519,
    n763,
    n781
  );


  xor
  g802
  (
    n820,
    n767,
    n785,
    n515,
    n766
  );


  or
  g803
  (
    n819,
    n785,
    n506,
    n786,
    n781
  );


  and
  g804
  (
    n832,
    n766,
    n783,
    n379,
    n380
  );


  xnor
  g805
  (
    n814,
    n375,
    n763,
    n497,
    n780
  );


  or
  g806
  (
    n796,
    n383,
    n513,
    n495,
    n768
  );


  nand
  g807
  (
    n821,
    n788,
    n374,
    n502,
    n382
  );


  nor
  g808
  (
    n798,
    n518,
    n372,
    n380,
    n374
  );


  xnor
  g809
  (
    n802,
    n782,
    n373,
    n383,
    n763
  );


  or
  g810
  (
    n823,
    n787,
    n761,
    n373,
    n382
  );


  buf
  g811
  (
    KeyWire_0_6,
    n819
  );


  not
  g812
  (
    n833,
    n818
  );


  buf
  g813
  (
    n836,
    n817
  );


  not
  g814
  (
    n834,
    n820
  );


  buf
  g815
  (
    n850,
    n795
  );


  xnor
  g816
  (
    n848,
    n792,
    n836,
    n529
  );


  or
  g817
  (
    n847,
    n792,
    n834,
    n526,
    n833
  );


  xnor
  g818
  (
    n837,
    n522,
    n530,
    n835,
    n525
  );


  nand
  g819
  (
    n841,
    n789,
    n835,
    n792,
    n791
  );


  nand
  g820
  (
    KeyWire_0_4,
    n532,
    n791,
    n728,
    n835
  );


  nor
  g821
  (
    n846,
    n789,
    n794,
    n793,
    n531
  );


  nand
  g822
  (
    n849,
    n523,
    n836,
    n727
  );


  nor
  g823
  (
    n840,
    n833,
    n834
  );


  nor
  g824
  (
    n842,
    n793,
    n795,
    n728,
    n790
  );


  nor
  g825
  (
    n845,
    n794,
    n836,
    n524,
    n790
  );


  nor
  g826
  (
    n851,
    n790,
    n795,
    n794,
    n527
  );


  xnor
  g827
  (
    n838,
    n533,
    n789,
    n793,
    n528
  );


  nand
  g828
  (
    n844,
    n835,
    n791,
    n729,
    n793
  );


  xnor
  g829
  (
    n852,
    n794,
    n836,
    n726,
    n792
  );


  xor
  g830
  (
    n839,
    n791,
    n833,
    n790,
    n834
  );


  not
  g831
  (
    n878,
    n850
  );


  not
  g832
  (
    n857,
    n535
  );


  not
  g833
  (
    n870,
    n840
  );


  not
  g834
  (
    n879,
    n843
  );


  buf
  g835
  (
    n887,
    n845
  );


  buf
  g836
  (
    n905,
    n852
  );


  buf
  g837
  (
    n880,
    n851
  );


  buf
  g838
  (
    n904,
    n845
  );


  buf
  g839
  (
    n858,
    n848
  );


  not
  g840
  (
    n862,
    n840
  );


  not
  g841
  (
    n900,
    n841
  );


  buf
  g842
  (
    n896,
    n837
  );


  buf
  g843
  (
    n884,
    n851
  );


  not
  g844
  (
    n856,
    n839
  );


  buf
  g845
  (
    n910,
    n842
  );


  not
  g846
  (
    n912,
    n841
  );


  not
  g847
  (
    n913,
    n839
  );


  not
  g848
  (
    n875,
    n838
  );


  not
  g849
  (
    n906,
    n850
  );


  buf
  g850
  (
    n891,
    n846
  );


  not
  g851
  (
    n914,
    n845
  );


  buf
  g852
  (
    n898,
    n844
  );


  not
  g853
  (
    n866,
    n845
  );


  not
  g854
  (
    n895,
    n842
  );


  buf
  g855
  (
    n893,
    n837
  );


  not
  g856
  (
    n889,
    n825
  );


  buf
  g857
  (
    n909,
    n844
  );


  buf
  g858
  (
    n864,
    n826
  );


  buf
  g859
  (
    n859,
    n852
  );


  buf
  g860
  (
    n863,
    n838
  );


  not
  g861
  (
    n894,
    n840
  );


  not
  g862
  (
    n888,
    n851
  );


  not
  g863
  (
    n886,
    n842
  );


  buf
  g864
  (
    n868,
    n841
  );


  buf
  g865
  (
    n853,
    n848
  );


  buf
  g866
  (
    n855,
    n841
  );


  not
  g867
  (
    n872,
    n848
  );


  not
  g868
  (
    n883,
    n840
  );


  buf
  g869
  (
    n903,
    n850
  );


  buf
  g870
  (
    n876,
    n839
  );


  not
  g871
  (
    n885,
    n847
  );


  buf
  g872
  (
    n865,
    n827
  );


  not
  g873
  (
    n860,
    n852
  );


  not
  g874
  (
    n890,
    n848
  );


  buf
  g875
  (
    n907,
    n839
  );


  buf
  g876
  (
    n892,
    n846
  );


  buf
  g877
  (
    n867,
    n843
  );


  not
  g878
  (
    n915,
    n852
  );


  buf
  g879
  (
    n861,
    n844
  );


  buf
  g880
  (
    n901,
    n844
  );


  buf
  g881
  (
    n911,
    n822
  );


  not
  g882
  (
    n916,
    n847
  );


  buf
  g883
  (
    n873,
    n821
  );


  buf
  g884
  (
    n897,
    n849
  );


  not
  g885
  (
    n871,
    n824
  );


  not
  g886
  (
    n899,
    n846
  );


  not
  g887
  (
    n854,
    n846
  );


  buf
  g888
  (
    n881,
    n837
  );


  not
  g889
  (
    n877,
    n837
  );


  not
  g890
  (
    n908,
    n847
  );


  not
  g891
  (
    n902,
    n534
  );


  and
  g892
  (
    KeyWire_0_0,
    n838,
    n850,
    n849,
    n823
  );


  or
  g893
  (
    n874,
    n849,
    n843,
    n847
  );


  and
  g894
  (
    n882,
    n849,
    n838,
    n851,
    n842
  );


  buf
  g895
  (
    n917,
    n863
  );


  not
  g896
  (
    n924,
    n857
  );


  not
  g897
  (
    n919,
    n854
  );


  buf
  g898
  (
    n920,
    n862
  );


  buf
  g899
  (
    n925,
    n853
  );


  not
  g900
  (
    n928,
    n855
  );


  buf
  g901
  (
    n923,
    n860
  );


  not
  g902
  (
    n921,
    n858
  );


  not
  g903
  (
    n922,
    n859
  );


  not
  g904
  (
    n927,
    n861
  );


  not
  g905
  (
    n918,
    n856
  );


  not
  g906
  (
    n926,
    n864
  );


  nor
  g907
  (
    n929,
    n924,
    n416,
    n394,
    n400
  );


  xnor
  g908
  (
    n949,
    n409,
    n928,
    n411,
    n921
  );


  or
  g909
  (
    n953,
    n922,
    n404,
    n917,
    n395
  );


  and
  g910
  (
    KeyWire_0_7,
    n925,
    n404,
    n396,
    n400
  );


  and
  g911
  (
    n954,
    n919,
    n925,
    n922,
    n390
  );


  xor
  g912
  (
    n947,
    n400,
    n385,
    n388
  );


  and
  g913
  (
    n946,
    n923,
    n389,
    n920,
    n396
  );


  and
  g914
  (
    n974,
    n918,
    n396,
    n919,
    n920
  );


  xor
  g915
  (
    n971,
    n417,
    n418,
    n391,
    n920
  );


  nor
  g916
  (
    n935,
    n419,
    n410,
    n920,
    n918
  );


  or
  g917
  (
    n951,
    n415,
    n918,
    n917,
    n403
  );


  or
  g918
  (
    n976,
    n413,
    n917,
    n925
  );


  nand
  g919
  (
    n966,
    n408,
    n393,
    n928,
    n412
  );


  xnor
  g920
  (
    n960,
    n386,
    n406,
    n417
  );


  nor
  g921
  (
    n932,
    n412,
    n413,
    n408,
    n407
  );


  nand
  g922
  (
    n965,
    n926,
    n393,
    n917,
    n384
  );


  or
  g923
  (
    n959,
    n399,
    n416,
    n412,
    n921
  );


  nor
  g924
  (
    n938,
    n407,
    n410,
    n416,
    n401
  );


  or
  g925
  (
    n975,
    n385,
    n386,
    n392,
    n403
  );


  xor
  g926
  (
    n943,
    n924,
    n406,
    n395,
    n387
  );


  nand
  g927
  (
    n942,
    n393,
    n387,
    n410,
    n394
  );


  xor
  g928
  (
    n962,
    n397,
    n398,
    n399
  );


  and
  g929
  (
    n958,
    n391,
    n389,
    n919,
    n392
  );


  nor
  g930
  (
    n963,
    n402,
    n412,
    n419,
    n384
  );


  xnor
  g931
  (
    n945,
    n926,
    n402,
    n389,
    n398
  );


  nor
  g932
  (
    n967,
    n402,
    n391,
    n401,
    n385
  );


  nand
  g933
  (
    n930,
    n408,
    n413,
    n926,
    n410
  );


  nor
  g934
  (
    n950,
    n395,
    n388,
    n413,
    n409
  );


  xnor
  g935
  (
    n944,
    n408,
    n395,
    n923,
    n409
  );


  xnor
  g936
  (
    n948,
    n416,
    n923,
    n403,
    n386
  );


  xor
  g937
  (
    n939,
    n418,
    n407,
    n400,
    n397
  );


  xor
  g938
  (
    n955,
    n401,
    n414,
    n918,
    n403
  );


  nand
  g939
  (
    n973,
    n390,
    n396,
    n405,
    n414
  );


  and
  g940
  (
    n933,
    n418,
    n405,
    n402
  );


  xor
  g941
  (
    n957,
    n414,
    n384,
    n388,
    n394
  );


  xnor
  g942
  (
    n934,
    n921,
    n390,
    n922,
    n386
  );


  nor
  g943
  (
    n937,
    n928,
    n404,
    n417,
    n399
  );


  xnor
  g944
  (
    n961,
    n418,
    n407,
    n384,
    n923
  );


  xor
  g945
  (
    n964,
    n406,
    n392,
    n409,
    n387
  );


  xnor
  g946
  (
    n956,
    n419,
    n928,
    n417,
    n415
  );


  and
  g947
  (
    n952,
    n401,
    n387,
    n390,
    n919
  );


  nand
  g948
  (
    n931,
    n397,
    n385,
    n393,
    n391
  );


  nand
  g949
  (
    n970,
    n921,
    n394,
    n411,
    n414
  );


  and
  g950
  (
    n968,
    n927,
    n924,
    n404,
    n926
  );


  xnor
  g951
  (
    n941,
    n924,
    n927,
    n419,
    n415
  );


  nand
  g952
  (
    n940,
    n398,
    n411,
    n392,
    n927
  );


  nor
  g953
  (
    n972,
    n389,
    n922,
    n398,
    n411
  );


  or
  g954
  (
    n969,
    n397,
    n927,
    n405,
    n415
  );


  xnor
  g955
  (
    n977,
    n567,
    n944,
    n576,
    n578
  );


  xor
  g956
  (
    n986,
    n559,
    n557,
    n560,
    n936
  );


  xor
  g957
  (
    n988,
    n577,
    n932,
    n574,
    n569
  );


  xnor
  g958
  (
    n983,
    n550,
    n572,
    n556,
    n939
  );


  nor
  g959
  (
    n989,
    n554,
    n561,
    n582,
    n573
  );


  xnor
  g960
  (
    n984,
    n935,
    n568,
    n934,
    n580
  );


  xnor
  g961
  (
    n981,
    n566,
    n938,
    n549,
    n551
  );


  and
  g962
  (
    n991,
    n544,
    n552,
    n564,
    n545
  );


  xor
  g963
  (
    n987,
    n941,
    n942,
    n553,
    n541
  );


  nor
  g964
  (
    n978,
    n571,
    n536,
    n575,
    n583
  );


  xnor
  g965
  (
    n992,
    n943,
    n562,
    n930,
    n542
  );


  and
  g966
  (
    n982,
    n546,
    n929,
    n548,
    n931
  );


  and
  g967
  (
    n980,
    n563,
    n537,
    n933,
    n579
  );


  nand
  g968
  (
    n979,
    n570,
    n937,
    n555,
    n539
  );


  or
  g969
  (
    n985,
    n565,
    n538,
    n940,
    n547
  );


  and
  g970
  (
    n990,
    n540,
    n558,
    n581,
    n543
  );


  buf
  g971
  (
    KeyWire_0_15,
    n978
  );


  not
  g972
  (
    n996,
    n977
  );


  or
  g973
  (
    n993,
    n587,
    n584
  );


  xnor
  g974
  (
    n995,
    n586,
    n585,
    n978,
    n977
  );


  and
  g975
  (
    n999,
    n967,
    n945,
    n954
  );


  nor
  g976
  (
    n1001,
    n960,
    n994,
    n966
  );


  xnor
  g977
  (
    n1007,
    n970,
    n952,
    n994,
    n964
  );


  and
  g978
  (
    n1003,
    n959,
    n968,
    n953,
    n971
  );


  xnor
  g979
  (
    n998,
    n995,
    n994,
    n950,
    n972
  );


  xnor
  g980
  (
    n1005,
    n955,
    n970,
    n994,
    n958
  );


  nand
  g981
  (
    n1000,
    n957,
    n947,
    n949,
    n993
  );


  and
  g982
  (
    n1004,
    n961,
    n969,
    n951,
    n956
  );


  xor
  g983
  (
    n1006,
    n948,
    n993,
    n968,
    n995
  );


  or
  g984
  (
    n1008,
    n946,
    n971,
    n993,
    n962
  );


  or
  g985
  (
    n1002,
    n967,
    n995,
    n993,
    n969
  );


  xor
  g986
  (
    n997,
    n966,
    n995,
    n963,
    n965
  );


  nor
  g987
  (
    n1015,
    n982,
    n989,
    n997,
    n980
  );


  xor
  g988
  (
    n1011,
    n985,
    n989,
    n983,
    n988
  );


  nand
  g989
  (
    n1017,
    n984,
    n998,
    n988
  );


  nand
  g990
  (
    n1013,
    n983,
    n980,
    n981,
    n999
  );


  and
  g991
  (
    n1012,
    n998,
    n987,
    n984,
    n979
  );


  xor
  g992
  (
    n1014,
    n998,
    n987,
    n997,
    n986
  );


  nor
  g993
  (
    n1009,
    n979,
    n987,
    n985,
    n984
  );


  nand
  g994
  (
    n1010,
    n998,
    n986,
    n985
  );


  nor
  g995
  (
    n1016,
    n981,
    n997,
    n982,
    n999
  );


  xnor
  g996
  (
    n1029,
    n896,
    n886,
    n1011,
    n867
  );


  and
  g997
  (
    n1022,
    n1010,
    n866,
    n878,
    n996
  );


  or
  g998
  (
    n1026,
    n1012,
    n869,
    n996,
    n873
  );


  xnor
  g999
  (
    n1018,
    n888,
    n1014,
    n897,
    n1013
  );


  nand
  g1000
  (
    n1023,
    n996,
    n868,
    n876,
    n882
  );


  xnor
  g1001
  (
    n1025,
    n881,
    n1011,
    n1009,
    n1010
  );


  nand
  g1002
  (
    n1027,
    n870,
    n1009,
    n1014,
    n871
  );


  nor
  g1003
  (
    n1031,
    n891,
    n1012,
    n879
  );


  xnor
  g1004
  (
    n1028,
    n884,
    n1013,
    n889,
    n877
  );


  or
  g1005
  (
    n1024,
    n1012,
    n872,
    n898,
    n1011
  );


  nor
  g1006
  (
    n1019,
    n588,
    n875,
    n890,
    n883
  );


  or
  g1007
  (
    n1030,
    n887,
    n865,
    n892,
    n885
  );


  nor
  g1008
  (
    n1032,
    n1014,
    n1010,
    n996,
    n1013
  );


  xnor
  g1009
  (
    n1020,
    n1011,
    n895,
    n874,
    n1013
  );


  xnor
  g1010
  (
    n1021,
    n1014,
    n894,
    n880,
    n893
  );


  and
  g1011
  (
    n1036,
    n593,
    n1032,
    n1003,
    n1002
  );


  xor
  g1012
  (
    n1038,
    n1027,
    n1002,
    n1029,
    n592
  );


  nor
  g1013
  (
    n1035,
    n1031,
    n596,
    n1000
  );


  xor
  g1014
  (
    n1037,
    n1028,
    n1001,
    n594,
    n1003
  );


  or
  g1015
  (
    n1040,
    n1002,
    n1000,
    n589,
    n1030
  );


  nand
  g1016
  (
    n1039,
    n999,
    n1001,
    n1000
  );


  or
  g1017
  (
    n1034,
    n1026,
    n591,
    n999,
    n1025
  );


  xnor
  g1018
  (
    n1033,
    n595,
    n1002,
    n1001,
    n590
  );


  nand
  g1019
  (
    n1041,
    n1034,
    n598,
    n599,
    n600
  );


  xor
  g1020
  (
    n1042,
    n1033,
    n601,
    n597,
    n602
  );


  xor
  g1021
  (
    n1043,
    n603,
    n604,
    n605,
    n1042
  );


  buf
  g1022
  (
    n1044,
    n1043
  );


  nor
  g1023
  (
    n1045,
    n606,
    n1043,
    n607
  );


  nor
  g1024
  (
    n1046,
    n610,
    n608,
    n1044,
    n609
  );


  buf
  g1025
  (
    n1049,
    n1046
  );


  not
  g1026
  (
    n1048,
    n611
  );


  buf
  g1027
  (
    n1047,
    n1046
  );


  not
  g1028
  (
    n1050,
    n1048
  );


  not
  g1029
  (
    n1051,
    n1048
  );


  buf
  g1030
  (
    n1053,
    n1048
  );


  nor
  g1031
  (
    n1052,
    n612,
    n1045,
    n1047
  );


  and
  g1032
  (
    n1055,
    n1050,
    n972
  );


  nand
  g1033
  (
    n1058,
    n990,
    n992,
    n1036
  );


  xor
  g1034
  (
    n1056,
    n990,
    n1035,
    n991,
    n1050
  );


  or
  g1035
  (
    n1054,
    n1050,
    n991,
    n1051
  );


  xnor
  g1036
  (
    n1057,
    n990,
    n1050,
    n992,
    n989
  );


  not
  g1037
  (
    n1062,
    n1055
  );


  buf
  g1038
  (
    KeyWire_0_9,
    n1054
  );


  buf
  g1039
  (
    n1061,
    n1054
  );


  buf
  g1040
  (
    n1059,
    n1054
  );


  xnor
  g1041
  (
    n1070,
    n734,
    n1061,
    n1008,
    n1059
  );


  or
  g1042
  (
    n1075,
    n1003,
    n1004,
    n831
  );


  nor
  g1043
  (
    n1066,
    n1006,
    n1003,
    n1053,
    n729
  );


  nand
  g1044
  (
    n1073,
    n733,
    n1006,
    n1052,
    n1060
  );


  and
  g1045
  (
    n1069,
    n1061,
    n1062,
    n1007,
    n731
  );


  and
  g1046
  (
    n1074,
    n1059,
    n1006,
    n1053
  );


  or
  g1047
  (
    n1064,
    n829,
    n732,
    n1051,
    n1004
  );


  xor
  g1048
  (
    n1063,
    n830,
    n828,
    n731,
    n1061
  );


  xnor
  g1049
  (
    n1076,
    n1005,
    n1007,
    n730
  );


  xnor
  g1050
  (
    n1071,
    n730,
    n1059,
    n1060,
    n795
  );


  nor
  g1051
  (
    n1065,
    n1061,
    n1060,
    n1006,
    n1059
  );


  and
  g1052
  (
    n1067,
    n1008,
    n1008,
    n1051,
    n1052
  );


  and
  g1053
  (
    n1068,
    n1007,
    n1005,
    n1062
  );


  nor
  g1054
  (
    n1077,
    n1008,
    n1005,
    n733
  );


  and
  g1055
  (
    n1078,
    n1060,
    n1062,
    n732,
    n1053
  );


  xnor
  g1056
  (
    n1072,
    n1004,
    n1052,
    n1051
  );


  xnor
  g1057
  (
    n1091,
    n1066,
    n626,
    n639,
    n1063
  );


  xnor
  g1058
  (
    n1080,
    n1064,
    n616,
    n1058,
    n1066
  );


  xor
  g1059
  (
    n1090,
    n628,
    n621,
    n641,
    n1067
  );


  nor
  g1060
  (
    n1079,
    n1058,
    n635,
    n1067,
    n1056
  );


  or
  g1061
  (
    n1089,
    n1058,
    n624,
    n1055,
    n629
  );


  or
  g1062
  (
    n1085,
    n1064,
    n1058,
    n1065,
    n627
  );


  xnor
  g1063
  (
    n1087,
    n1056,
    n1056,
    n1055,
    n1067
  );


  xor
  g1064
  (
    n1086,
    n642,
    n632,
    n620,
    n614
  );


  nand
  g1065
  (
    n1092,
    n613,
    n618,
    n619,
    n630
  );


  nand
  g1066
  (
    n1088,
    n1057,
    n640,
    n1064,
    n615
  );


  or
  g1067
  (
    n1082,
    n1065,
    n1066,
    n1063,
    n622
  );


  or
  g1068
  (
    n1093,
    n625,
    n623,
    n636,
    n1057
  );


  or
  g1069
  (
    n1081,
    n633,
    n637,
    n638,
    n1057
  );


  nand
  g1070
  (
    n1084,
    n631,
    n1056,
    n617,
    n1057
  );


  nor
  g1071
  (
    n1083,
    n1055,
    n634,
    n1065,
    n1068
  );


  buf
  g1072
  (
    n1105,
    n1080
  );


  buf
  g1073
  (
    n1131,
    n906
  );


  buf
  g1074
  (
    n1126,
    n1093
  );


  buf
  g1075
  (
    n1127,
    n913
  );


  not
  g1076
  (
    n1133,
    n1085
  );


  not
  g1077
  (
    n1116,
    n908
  );


  buf
  g1078
  (
    n1102,
    n1015
  );


  buf
  g1079
  (
    n1118,
    n1087
  );


  buf
  g1080
  (
    n1115,
    n1090
  );


  not
  g1081
  (
    n1106,
    n1082
  );


  buf
  g1082
  (
    n1108,
    n1091
  );


  buf
  g1083
  (
    n1099,
    n912
  );


  not
  g1084
  (
    n1135,
    n1091
  );


  not
  g1085
  (
    n1111,
    n1015
  );


  buf
  g1086
  (
    n1123,
    n899
  );


  not
  g1087
  (
    n1100,
    n1016
  );


  buf
  g1088
  (
    n1129,
    n1093
  );


  not
  g1089
  (
    n1120,
    n1080
  );


  buf
  g1090
  (
    n1096,
    n1090
  );


  buf
  g1091
  (
    n1119,
    n1080
  );


  buf
  g1092
  (
    n1113,
    n1091
  );


  buf
  g1093
  (
    n1112,
    n912
  );


  not
  g1094
  (
    n1132,
    n1084
  );


  not
  g1095
  (
    n1122,
    n1084
  );


  buf
  g1096
  (
    n1117,
    n915
  );


  buf
  g1097
  (
    n1125,
    n910
  );


  not
  g1098
  (
    n1114,
    n1085
  );


  not
  g1099
  (
    n1121,
    n904
  );


  buf
  g1100
  (
    n1109,
    n1017
  );


  or
  g1101
  (
    n1110,
    n769,
    n911,
    n1082
  );


  xnor
  g1102
  (
    n1128,
    n1085,
    n1016,
    n910,
    n1082
  );


  xnor
  g1103
  (
    n1107,
    n1081,
    n914,
    n832,
    n906
  );


  xor
  g1104
  (
    n1137,
    n1017,
    n1088,
    n1081,
    n1092
  );


  nand
  g1105
  (
    n1095,
    n1084,
    n914,
    n769,
    n1016
  );


  and
  g1106
  (
    n1097,
    n1015,
    n1087,
    n907,
    n913
  );


  xor
  g1107
  (
    n1124,
    n1083,
    n643,
    n1088
  );


  nor
  g1108
  (
    n1103,
    n1092,
    n1017,
    n1083,
    n901
  );


  nor
  g1109
  (
    n1140,
    n1081,
    n905,
    n1089,
    n1079
  );


  or
  g1110
  (
    n1139,
    n1086,
    n1046,
    n1089
  );


  xor
  g1111
  (
    n1098,
    n645,
    n1015,
    n902,
    n1079
  );


  nor
  g1112
  (
    n1134,
    n1090,
    n644,
    n1091,
    n769
  );


  xor
  g1113
  (
    n1104,
    n904,
    n903,
    n1017,
    n1087
  );


  or
  g1114
  (
    n1101,
    n769,
    n1092,
    n734,
    n1016
  );


  or
  g1115
  (
    n1094,
    n905,
    n909,
    n908,
    n907
  );


  xnor
  g1116
  (
    n1136,
    n915,
    n1086,
    n1093
  );


  and
  g1117
  (
    n1138,
    n768,
    n1092,
    n1083,
    n900
  );


  nand
  g1118
  (
    n1130,
    n768,
    n1093,
    n911,
    n909
  );


  or
  g1119
  (
    n1146,
    n1116,
    n1049,
    n1114,
    n1038
  );


  xor
  g1120
  (
    n1141,
    n1039,
    n1048,
    n1075,
    n1100
  );


  or
  g1121
  (
    n1164,
    n1108,
    n1132,
    n1128,
    n1074
  );


  nand
  g1122
  (
    n1162,
    n1120,
    n1037,
    n1133,
    n1071
  );


  or
  g1123
  (
    n1142,
    n1075,
    n1073,
    n1077,
    n1127
  );


  or
  g1124
  (
    n1156,
    n1077,
    n1126,
    n1068
  );


  and
  g1125
  (
    n1159,
    n1118,
    n974,
    n1075,
    n973
  );


  xor
  g1126
  (
    n1144,
    n1102,
    n1140,
    n1136,
    n1072
  );


  xor
  g1127
  (
    n1152,
    n1112,
    n1099,
    n1139,
    n1131
  );


  or
  g1128
  (
    n1153,
    n1106,
    n1130,
    n1077,
    n916
  );


  xnor
  g1129
  (
    n1161,
    n1069,
    n1076,
    n1049,
    n1095
  );


  nor
  g1130
  (
    n1154,
    n1078,
    n1123,
    n1071,
    n1138
  );


  and
  g1131
  (
    n1148,
    n1129,
    n1073,
    n1049,
    n1097
  );


  nand
  g1132
  (
    n1165,
    n976,
    n975,
    n1074,
    n1110
  );


  and
  g1133
  (
    n1143,
    n1137,
    n1072,
    n1122,
    n1070
  );


  or
  g1134
  (
    n1145,
    n1040,
    n1096,
    n1094,
    n1078
  );


  nor
  g1135
  (
    n1157,
    n1078,
    n1078,
    n1073,
    n1121
  );


  nand
  g1136
  (
    n1150,
    n1076,
    n1098,
    n1072,
    n1107
  );


  and
  g1137
  (
    n1155,
    n1109,
    n976,
    n1135,
    n1074
  );


  nand
  g1138
  (
    n1147,
    n1115,
    n1069,
    n1101
  );


  nand
  g1139
  (
    n1158,
    n1049,
    n1124,
    n1104,
    n1071
  );


  xor
  g1140
  (
    n1149,
    n1103,
    n916,
    n1119,
    n1117
  );


  nand
  g1141
  (
    n1163,
    n1105,
    n973,
    n976,
    n974
  );


  nand
  g1142
  (
    n1151,
    n1070,
    n1125,
    n1076,
    n1111
  );


  or
  g1143
  (
    n1160,
    n1070,
    n1113,
    n975,
    n1134
  );


  xor
  g1144
  (
    n1177,
    n1150,
    n669,
    n649,
    n668
  );


  and
  g1145
  (
    n1172,
    n680,
    n1157,
    n674,
    n1164
  );


  nor
  g1146
  (
    n1166,
    n1142,
    n653,
    n651,
    n1151
  );


  nand
  g1147
  (
    n1167,
    n661,
    n1165,
    n1162,
    n1161
  );


  xnor
  g1148
  (
    n1171,
    n656,
    n1152,
    n663,
    n1156
  );


  nor
  g1149
  (
    n1178,
    n658,
    n676,
    n662,
    n648
  );


  xor
  g1150
  (
    n1182,
    n652,
    n1147,
    n1146,
    n1153
  );


  xnor
  g1151
  (
    n1183,
    n685,
    n1155,
    n1143,
    n1145
  );


  xnor
  g1152
  (
    n1170,
    n660,
    n1159,
    n1141,
    n684
  );


  and
  g1153
  (
    n1179,
    n675,
    n650,
    n681,
    n678
  );


  and
  g1154
  (
    n1169,
    n682,
    n1148,
    n690,
    n677
  );


  xnor
  g1155
  (
    n1174,
    n692,
    n671,
    n672,
    n683
  );


  nor
  g1156
  (
    n1175,
    n688,
    n689,
    n1149,
    n657
  );


  nor
  g1157
  (
    n1173,
    n659,
    n666,
    n1154,
    n673
  );


  and
  g1158
  (
    n1181,
    n647,
    n664,
    n1160,
    n646
  );


  nand
  g1159
  (
    n1176,
    n655,
    n1144,
    n1158,
    n654
  );


  and
  g1160
  (
    n1168,
    n670,
    n665,
    n686,
    n1163
  );


  xnor
  g1161
  (
    n1180,
    n679,
    n687,
    n691,
    n667
  );


  xnor
  KeyGate_0_0
  (
    n869,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n737,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n183,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n61,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n843,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n731,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n835,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n936,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n369,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1060,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n258,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n323,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n280,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n632,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n375,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n994,
    KeyNOTWire_0_15
  );


endmodule

