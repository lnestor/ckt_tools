

module Stat_1153_20_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n792,
  n798,
  n959,
  n961,
  n1163,
  n1162,
  n1174,
  n1157,
  n1156,
  n1159,
  n1172,
  n1169,
  n1171,
  n1158,
  n1164,
  n1161,
  n1165,
  n1173,
  n1166,
  n1154,
  n1175,
  n1167,
  n1168,
  n1155,
  n1160,
  n1170,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n792;
  output n798;
  output n959;
  output n961;
  output n1163;
  output n1162;
  output n1174;
  output n1157;
  output n1156;
  output n1159;
  output n1172;
  output n1169;
  output n1171;
  output n1158;
  output n1164;
  output n1161;
  output n1165;
  output n1173;
  output n1166;
  output n1154;
  output n1175;
  output n1167;
  output n1168;
  output n1155;
  output n1160;
  output n1170;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n960;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n107,
    n11
  );


  not
  g1
  (
    n53,
    n10
  );


  not
  g2
  (
    n98,
    n20
  );


  buf
  g3
  (
    n84,
    n13
  );


  not
  g4
  (
    n30,
    n4
  );


  not
  g5
  (
    n93,
    n16
  );


  buf
  g6
  (
    n102,
    n1
  );


  not
  g7
  (
    n50,
    n17
  );


  not
  g8
  (
    n96,
    n11
  );


  buf
  g9
  (
    n54,
    n7
  );


  buf
  g10
  (
    n68,
    n15
  );


  buf
  g11
  (
    n88,
    n22
  );


  not
  g12
  (
    n110,
    n1
  );


  not
  g13
  (
    n82,
    n12
  );


  not
  g14
  (
    n73,
    n5
  );


  not
  g15
  (
    n33,
    n15
  );


  not
  g16
  (
    KeyWire_0_48,
    n19
  );


  buf
  g17
  (
    n62,
    n11
  );


  not
  g18
  (
    n46,
    n16
  );


  not
  g19
  (
    KeyWire_0_10,
    n12
  );


  not
  g20
  (
    n61,
    n7
  );


  buf
  g21
  (
    n70,
    n13
  );


  not
  g22
  (
    n76,
    n10
  );


  buf
  g23
  (
    n25,
    n4
  );


  buf
  g24
  (
    n74,
    n4
  );


  buf
  g25
  (
    n32,
    n3
  );


  not
  g26
  (
    n80,
    n19
  );


  not
  g27
  (
    n37,
    n4
  );


  buf
  g28
  (
    n78,
    n8
  );


  not
  g29
  (
    n75,
    n14
  );


  buf
  g30
  (
    n35,
    n8
  );


  buf
  g31
  (
    n44,
    n21
  );


  not
  g32
  (
    n104,
    n13
  );


  not
  g33
  (
    n55,
    n18
  );


  buf
  g34
  (
    n72,
    n13
  );


  not
  g35
  (
    n51,
    n19
  );


  not
  g36
  (
    n95,
    n16
  );


  buf
  g37
  (
    n42,
    n6
  );


  not
  g38
  (
    KeyWire_0_23,
    n10
  );


  not
  g39
  (
    KeyWire_0_55,
    n9
  );


  not
  g40
  (
    n47,
    n21
  );


  not
  g41
  (
    n87,
    n19
  );


  buf
  g42
  (
    n45,
    n16
  );


  buf
  g43
  (
    n86,
    n22
  );


  not
  g44
  (
    n103,
    n17
  );


  not
  g45
  (
    n100,
    n3
  );


  buf
  g46
  (
    n34,
    n14
  );


  buf
  g47
  (
    n79,
    n8
  );


  buf
  g48
  (
    n31,
    n6
  );


  buf
  g49
  (
    n94,
    n10
  );


  not
  g50
  (
    n49,
    n2
  );


  not
  g51
  (
    n43,
    n3
  );


  buf
  g52
  (
    n83,
    n9
  );


  not
  g53
  (
    n41,
    n15
  );


  buf
  g54
  (
    n105,
    n12
  );


  not
  g55
  (
    n90,
    n2
  );


  buf
  g56
  (
    n92,
    n14
  );


  not
  g57
  (
    n65,
    n3
  );


  buf
  g58
  (
    n64,
    n21
  );


  not
  g59
  (
    n27,
    n5
  );


  not
  g60
  (
    KeyWire_0_30,
    n5
  );


  buf
  g61
  (
    n48,
    n18
  );


  not
  g62
  (
    n77,
    n9
  );


  buf
  g63
  (
    n85,
    n6
  );


  not
  g64
  (
    n29,
    n17
  );


  buf
  g65
  (
    n56,
    n7
  );


  buf
  g66
  (
    n63,
    n5
  );


  not
  g67
  (
    n24,
    n1
  );


  not
  g68
  (
    n23,
    n18
  );


  not
  g69
  (
    n60,
    n17
  );


  not
  g70
  (
    n67,
    n20
  );


  buf
  g71
  (
    n108,
    n22
  );


  buf
  g72
  (
    n81,
    n7
  );


  not
  g73
  (
    n69,
    n21
  );


  buf
  g74
  (
    n97,
    n2
  );


  buf
  g75
  (
    n99,
    n20
  );


  buf
  g76
  (
    n106,
    n1
  );


  buf
  g77
  (
    n57,
    n18
  );


  not
  g78
  (
    n59,
    n20
  );


  not
  g79
  (
    n91,
    n9
  );


  buf
  g80
  (
    n66,
    n15
  );


  not
  g81
  (
    n109,
    n22
  );


  buf
  g82
  (
    n89,
    n8
  );


  buf
  g83
  (
    n101,
    n12
  );


  buf
  g84
  (
    n58,
    n11
  );


  buf
  g85
  (
    n71,
    n6
  );


  not
  g86
  (
    n28,
    n14
  );


  buf
  g87
  (
    n39,
    n2
  );


  not
  g88
  (
    n390,
    n88
  );


  not
  g89
  (
    n241,
    n28
  );


  buf
  g90
  (
    n113,
    n26
  );


  not
  g91
  (
    n146,
    n44
  );


  not
  g92
  (
    n298,
    n96
  );


  buf
  g93
  (
    n315,
    n62
  );


  buf
  g94
  (
    n358,
    n88
  );


  not
  g95
  (
    KeyWire_0_63,
    n67
  );


  buf
  g96
  (
    n306,
    n97
  );


  buf
  g97
  (
    n222,
    n87
  );


  not
  g98
  (
    n258,
    n73
  );


  buf
  g99
  (
    n225,
    n63
  );


  not
  g100
  (
    KeyWire_0_49,
    n98
  );


  not
  g101
  (
    n294,
    n64
  );


  not
  g102
  (
    n310,
    n99
  );


  not
  g103
  (
    n169,
    n43
  );


  buf
  g104
  (
    n190,
    n108
  );


  not
  g105
  (
    n453,
    n65
  );


  not
  g106
  (
    n249,
    n46
  );


  buf
  g107
  (
    n205,
    n52
  );


  not
  g108
  (
    n313,
    n40
  );


  buf
  g109
  (
    n280,
    n67
  );


  buf
  g110
  (
    n250,
    n36
  );


  buf
  g111
  (
    n409,
    n88
  );


  buf
  g112
  (
    n174,
    n60
  );


  buf
  g113
  (
    n179,
    n92
  );


  not
  g114
  (
    KeyWire_0_21,
    n106
  );


  not
  g115
  (
    n340,
    n92
  );


  buf
  g116
  (
    n213,
    n32
  );


  not
  g117
  (
    n426,
    n86
  );


  buf
  g118
  (
    n286,
    n36
  );


  not
  g119
  (
    n263,
    n27
  );


  buf
  g120
  (
    n439,
    n58
  );


  not
  g121
  (
    n383,
    n48
  );


  not
  g122
  (
    n418,
    n75
  );


  buf
  g123
  (
    n337,
    n82
  );


  not
  g124
  (
    n207,
    n56
  );


  not
  g125
  (
    n406,
    n81
  );


  not
  g126
  (
    n323,
    n81
  );


  buf
  g127
  (
    n212,
    n47
  );


  buf
  g128
  (
    n376,
    n39
  );


  buf
  g129
  (
    n299,
    n32
  );


  buf
  g130
  (
    n118,
    n92
  );


  not
  g131
  (
    n303,
    n81
  );


  buf
  g132
  (
    n317,
    n68
  );


  not
  g133
  (
    n292,
    n42
  );


  not
  g134
  (
    n233,
    n70
  );


  not
  g135
  (
    n437,
    n90
  );


  not
  g136
  (
    n265,
    n105
  );


  not
  g137
  (
    n279,
    n73
  );


  not
  g138
  (
    n391,
    n24
  );


  not
  g139
  (
    n287,
    n47
  );


  not
  g140
  (
    n132,
    n24
  );


  buf
  g141
  (
    n382,
    n48
  );


  not
  g142
  (
    n341,
    n86
  );


  buf
  g143
  (
    n304,
    n102
  );


  buf
  g144
  (
    n434,
    n94
  );


  not
  g145
  (
    n199,
    n66
  );


  not
  g146
  (
    n264,
    n26
  );


  buf
  g147
  (
    n202,
    n77
  );


  buf
  g148
  (
    n324,
    n50
  );


  not
  g149
  (
    n343,
    n78
  );


  buf
  g150
  (
    n136,
    n28
  );


  buf
  g151
  (
    n380,
    n103
  );


  buf
  g152
  (
    n175,
    n61
  );


  not
  g153
  (
    n411,
    n33
  );


  buf
  g154
  (
    n447,
    n104
  );


  buf
  g155
  (
    n442,
    n85
  );


  buf
  g156
  (
    n262,
    n71
  );


  buf
  g157
  (
    n374,
    n43
  );


  buf
  g158
  (
    n339,
    n100
  );


  buf
  g159
  (
    n452,
    n34
  );


  buf
  g160
  (
    n415,
    n50
  );


  buf
  g161
  (
    n256,
    n42
  );


  buf
  g162
  (
    n166,
    n30
  );


  buf
  g163
  (
    n230,
    n108
  );


  buf
  g164
  (
    n328,
    n53
  );


  not
  g165
  (
    n122,
    n80
  );


  buf
  g166
  (
    n234,
    n32
  );


  buf
  g167
  (
    n261,
    n80
  );


  not
  g168
  (
    n384,
    n99
  );


  buf
  g169
  (
    n318,
    n60
  );


  buf
  g170
  (
    KeyWire_0_4,
    n64
  );


  not
  g171
  (
    n277,
    n66
  );


  not
  g172
  (
    n274,
    n27
  );


  buf
  g173
  (
    n289,
    n68
  );


  not
  g174
  (
    n117,
    n88
  );


  buf
  g175
  (
    n111,
    n57
  );


  not
  g176
  (
    n236,
    n45
  );


  buf
  g177
  (
    n240,
    n104
  );


  not
  g178
  (
    n217,
    n83
  );


  not
  g179
  (
    n346,
    n102
  );


  not
  g180
  (
    n273,
    n74
  );


  buf
  g181
  (
    n229,
    n67
  );


  not
  g182
  (
    n260,
    n97
  );


  not
  g183
  (
    n291,
    n51
  );


  not
  g184
  (
    n319,
    n45
  );


  not
  g185
  (
    KeyWire_0_41,
    n40
  );


  not
  g186
  (
    KeyWire_0_14,
    n49
  );


  not
  g187
  (
    n422,
    n108
  );


  not
  g188
  (
    n177,
    n79
  );


  buf
  g189
  (
    n367,
    n28
  );


  buf
  g190
  (
    n401,
    n48
  );


  buf
  g191
  (
    n393,
    n72
  );


  buf
  g192
  (
    n191,
    n61
  );


  not
  g193
  (
    n445,
    n97
  );


  buf
  g194
  (
    n345,
    n41
  );


  buf
  g195
  (
    n235,
    n71
  );


  not
  g196
  (
    n246,
    n65
  );


  buf
  g197
  (
    n115,
    n35
  );


  not
  g198
  (
    n395,
    n44
  );


  not
  g199
  (
    n369,
    n95
  );


  buf
  g200
  (
    n278,
    n41
  );


  not
  g201
  (
    n377,
    n107
  );


  buf
  g202
  (
    n413,
    n55
  );


  buf
  g203
  (
    n128,
    n35
  );


  buf
  g204
  (
    n251,
    n80
  );


  buf
  g205
  (
    n275,
    n83
  );


  not
  g206
  (
    KeyWire_0_40,
    n106
  );


  buf
  g207
  (
    n360,
    n101
  );


  not
  g208
  (
    n402,
    n84
  );


  buf
  g209
  (
    n145,
    n75
  );


  not
  g210
  (
    n446,
    n77
  );


  buf
  g211
  (
    n267,
    n69
  );


  buf
  g212
  (
    n160,
    n37
  );


  buf
  g213
  (
    n331,
    n49
  );


  not
  g214
  (
    n206,
    n64
  );


  buf
  g215
  (
    n405,
    n23
  );


  not
  g216
  (
    n435,
    n93
  );


  not
  g217
  (
    KeyWire_0_33,
    n37
  );


  not
  g218
  (
    n394,
    n25
  );


  buf
  g219
  (
    n255,
    n59
  );


  buf
  g220
  (
    KeyWire_0_36,
    n45
  );


  not
  g221
  (
    n125,
    n53
  );


  not
  g222
  (
    n215,
    n89
  );


  buf
  g223
  (
    n312,
    n69
  );


  buf
  g224
  (
    n432,
    n62
  );


  buf
  g225
  (
    n444,
    n75
  );


  buf
  g226
  (
    n149,
    n31
  );


  not
  g227
  (
    n144,
    n89
  );


  buf
  g228
  (
    n398,
    n78
  );


  buf
  g229
  (
    n150,
    n96
  );


  buf
  g230
  (
    n158,
    n23
  );


  buf
  g231
  (
    n112,
    n37
  );


  not
  g232
  (
    n335,
    n38
  );


  buf
  g233
  (
    n300,
    n101
  );


  not
  g234
  (
    n427,
    n41
  );


  buf
  g235
  (
    n410,
    n47
  );


  not
  g236
  (
    n269,
    n69
  );


  buf
  g237
  (
    KeyWire_0_43,
    n57
  );


  not
  g238
  (
    n407,
    n37
  );


  not
  g239
  (
    n314,
    n98
  );


  not
  g240
  (
    n363,
    n57
  );


  not
  g241
  (
    n139,
    n96
  );


  not
  g242
  (
    n424,
    n56
  );


  buf
  g243
  (
    n354,
    n99
  );


  not
  g244
  (
    n387,
    n79
  );


  buf
  g245
  (
    n211,
    n87
  );


  not
  g246
  (
    n309,
    n67
  );


  not
  g247
  (
    n326,
    n42
  );


  buf
  g248
  (
    n414,
    n84
  );


  buf
  g249
  (
    n214,
    n28
  );


  buf
  g250
  (
    n428,
    n27
  );


  buf
  g251
  (
    n378,
    n91
  );


  buf
  g252
  (
    n172,
    n51
  );


  not
  g253
  (
    n259,
    n39
  );


  not
  g254
  (
    n334,
    n52
  );


  not
  g255
  (
    n403,
    n93
  );


  buf
  g256
  (
    n436,
    n43
  );


  buf
  g257
  (
    n220,
    n96
  );


  buf
  g258
  (
    n219,
    n71
  );


  not
  g259
  (
    n283,
    n84
  );


  buf
  g260
  (
    n288,
    n70
  );


  buf
  g261
  (
    KeyWire_0_38,
    n95
  );


  not
  g262
  (
    n189,
    n77
  );


  not
  g263
  (
    n182,
    n59
  );


  buf
  g264
  (
    n336,
    n86
  );


  buf
  g265
  (
    n124,
    n108
  );


  buf
  g266
  (
    n218,
    n59
  );


  not
  g267
  (
    n114,
    n102
  );


  buf
  g268
  (
    n448,
    n68
  );


  buf
  g269
  (
    n252,
    n92
  );


  not
  g270
  (
    n186,
    n107
  );


  buf
  g271
  (
    n173,
    n30
  );


  buf
  g272
  (
    n420,
    n103
  );


  buf
  g273
  (
    n359,
    n80
  );


  not
  g274
  (
    n171,
    n70
  );


  buf
  g275
  (
    n194,
    n90
  );


  not
  g276
  (
    n440,
    n40
  );


  buf
  g277
  (
    n301,
    n107
  );


  buf
  g278
  (
    n221,
    n40
  );


  buf
  g279
  (
    n148,
    n86
  );


  not
  g280
  (
    n272,
    n24
  );


  buf
  g281
  (
    n242,
    n29
  );


  buf
  g282
  (
    n399,
    n34
  );


  buf
  g283
  (
    n170,
    n23
  );


  buf
  g284
  (
    n181,
    n41
  );


  buf
  g285
  (
    n308,
    n79
  );


  not
  g286
  (
    n167,
    n51
  );


  not
  g287
  (
    n133,
    n106
  );


  buf
  g288
  (
    n322,
    n61
  );


  not
  g289
  (
    n438,
    n56
  );


  buf
  g290
  (
    n404,
    n104
  );


  buf
  g291
  (
    n227,
    n25
  );


  not
  g292
  (
    n385,
    n87
  );


  buf
  g293
  (
    n356,
    n25
  );


  buf
  g294
  (
    n134,
    n91
  );


  not
  g295
  (
    n184,
    n85
  );


  buf
  g296
  (
    n126,
    n61
  );


  buf
  g297
  (
    n327,
    n39
  );


  not
  g298
  (
    n163,
    n72
  );


  buf
  g299
  (
    n130,
    n105
  );


  not
  g300
  (
    n187,
    n33
  );


  buf
  g301
  (
    n325,
    n34
  );


  not
  g302
  (
    n129,
    n101
  );


  buf
  g303
  (
    n281,
    n58
  );


  buf
  g304
  (
    n381,
    n83
  );


  buf
  g305
  (
    n348,
    n82
  );


  not
  g306
  (
    n153,
    n53
  );


  not
  g307
  (
    n450,
    n45
  );


  not
  g308
  (
    n154,
    n100
  );


  buf
  g309
  (
    n231,
    n55
  );


  buf
  g310
  (
    n425,
    n62
  );


  not
  g311
  (
    n349,
    n47
  );


  buf
  g312
  (
    n423,
    n50
  );


  not
  g313
  (
    n197,
    n94
  );


  buf
  g314
  (
    n185,
    n49
  );


  not
  g315
  (
    n350,
    n33
  );


  buf
  g316
  (
    n237,
    n75
  );


  buf
  g317
  (
    n151,
    n69
  );


  buf
  g318
  (
    n178,
    n81
  );


  not
  g319
  (
    n243,
    n78
  );


  not
  g320
  (
    n386,
    n43
  );


  not
  g321
  (
    n198,
    n105
  );


  buf
  g322
  (
    KeyWire_0_1,
    n85
  );


  not
  g323
  (
    n296,
    n72
  );


  not
  g324
  (
    n152,
    n103
  );


  not
  g325
  (
    n375,
    n55
  );


  buf
  g326
  (
    n372,
    n104
  );


  buf
  g327
  (
    n364,
    n63
  );


  not
  g328
  (
    n142,
    n46
  );


  buf
  g329
  (
    n119,
    n58
  );


  buf
  g330
  (
    n270,
    n91
  );


  not
  g331
  (
    n311,
    n36
  );


  buf
  g332
  (
    n183,
    n97
  );


  buf
  g333
  (
    n266,
    n68
  );


  not
  g334
  (
    n138,
    n73
  );


  not
  g335
  (
    n431,
    n66
  );


  buf
  g336
  (
    n379,
    n54
  );


  not
  g337
  (
    n305,
    n31
  );


  buf
  g338
  (
    n164,
    n38
  );


  buf
  g339
  (
    n408,
    n30
  );


  not
  g340
  (
    n362,
    n93
  );


  buf
  g341
  (
    KeyWire_0_7,
    n106
  );


  not
  g342
  (
    n451,
    n100
  );


  not
  g343
  (
    n247,
    n38
  );


  not
  g344
  (
    n200,
    n53
  );


  not
  g345
  (
    n392,
    n89
  );


  buf
  g346
  (
    n429,
    n63
  );


  buf
  g347
  (
    n188,
    n77
  );


  not
  g348
  (
    n176,
    n27
  );


  buf
  g349
  (
    n293,
    n101
  );


  not
  g350
  (
    KeyWire_0_57,
    n55
  );


  not
  g351
  (
    n123,
    n38
  );


  not
  g352
  (
    n141,
    n52
  );


  buf
  g353
  (
    n344,
    n46
  );


  buf
  g354
  (
    n120,
    n54
  );


  not
  g355
  (
    n290,
    n70
  );


  not
  g356
  (
    n239,
    n62
  );


  not
  g357
  (
    n333,
    n29
  );


  not
  g358
  (
    n271,
    n78
  );


  not
  g359
  (
    n155,
    n36
  );


  not
  g360
  (
    n297,
    n71
  );


  buf
  g361
  (
    n371,
    n74
  );


  not
  g362
  (
    n357,
    n44
  );


  not
  g363
  (
    n370,
    n79
  );


  buf
  g364
  (
    n159,
    n94
  );


  buf
  g365
  (
    n208,
    n76
  );


  not
  g366
  (
    n400,
    n34
  );


  not
  g367
  (
    n162,
    n103
  );


  buf
  g368
  (
    n116,
    n31
  );


  not
  g369
  (
    KeyWire_0_27,
    n59
  );


  not
  g370
  (
    n389,
    n99
  );


  buf
  g371
  (
    n285,
    n54
  );


  buf
  g372
  (
    KeyWire_0_44,
    n85
  );


  not
  g373
  (
    n366,
    n48
  );


  buf
  g374
  (
    n449,
    n52
  );


  buf
  g375
  (
    n302,
    n60
  );


  buf
  g376
  (
    n210,
    n90
  );


  not
  g377
  (
    n223,
    n63
  );


  buf
  g378
  (
    n421,
    n107
  );


  not
  g379
  (
    n396,
    n29
  );


  buf
  g380
  (
    n388,
    n51
  );


  not
  g381
  (
    KeyWire_0_0,
    n74
  );


  not
  g382
  (
    n216,
    n42
  );


  not
  g383
  (
    n203,
    n105
  );


  not
  g384
  (
    n127,
    n26
  );


  buf
  g385
  (
    n196,
    n87
  );


  buf
  g386
  (
    n137,
    n58
  );


  buf
  g387
  (
    KeyWire_0_19,
    n102
  );


  buf
  g388
  (
    n321,
    n94
  );


  buf
  g389
  (
    n180,
    n72
  );


  not
  g390
  (
    n254,
    n60
  );


  not
  g391
  (
    n168,
    n76
  );


  buf
  g392
  (
    n228,
    n24
  );


  not
  g393
  (
    n245,
    n25
  );


  not
  g394
  (
    n238,
    n100
  );


  not
  g395
  (
    n192,
    n44
  );


  not
  g396
  (
    n143,
    n56
  );


  buf
  g397
  (
    n351,
    n91
  );


  not
  g398
  (
    n419,
    n54
  );


  not
  g399
  (
    n365,
    n49
  );


  buf
  g400
  (
    n248,
    n26
  );


  buf
  g401
  (
    n209,
    n30
  );


  not
  g402
  (
    n330,
    n23
  );


  not
  g403
  (
    n268,
    n76
  );


  buf
  g404
  (
    n454,
    n82
  );


  buf
  g405
  (
    n441,
    n29
  );


  buf
  g406
  (
    n433,
    n50
  );


  not
  g407
  (
    n443,
    n98
  );


  buf
  g408
  (
    n347,
    n98
  );


  not
  g409
  (
    KeyWire_0_16,
    n82
  );


  not
  g410
  (
    n131,
    n31
  );


  buf
  g411
  (
    n430,
    n90
  );


  not
  g412
  (
    n353,
    n32
  );


  not
  g413
  (
    n412,
    n46
  );


  not
  g414
  (
    n361,
    n66
  );


  not
  g415
  (
    n224,
    n95
  );


  buf
  g416
  (
    n193,
    n35
  );


  not
  g417
  (
    n135,
    n95
  );


  buf
  g418
  (
    n416,
    n84
  );


  buf
  g419
  (
    n156,
    n73
  );


  not
  g420
  (
    n161,
    n83
  );


  not
  g421
  (
    KeyWire_0_50,
    n64
  );


  not
  g422
  (
    n232,
    n39
  );


  buf
  g423
  (
    n332,
    n74
  );


  not
  g424
  (
    n320,
    n65
  );


  buf
  g425
  (
    n157,
    n33
  );


  not
  g426
  (
    n417,
    n93
  );


  not
  g427
  (
    n226,
    n76
  );


  not
  g428
  (
    KeyWire_0_61,
    n89
  );


  buf
  g429
  (
    KeyWire_0_45,
    n57
  );


  buf
  g430
  (
    n355,
    n65
  );


  not
  g431
  (
    n352,
    n35
  );


  buf
  g432
  (
    n628,
    n234
  );


  buf
  g433
  (
    n587,
    n122
  );


  buf
  g434
  (
    n675,
    n373
  );


  buf
  g435
  (
    n667,
    n315
  );


  buf
  g436
  (
    n676,
    n238
  );


  buf
  g437
  (
    n589,
    n254
  );


  not
  g438
  (
    n478,
    n236
  );


  buf
  g439
  (
    n653,
    n211
  );


  not
  g440
  (
    n641,
    n216
  );


  not
  g441
  (
    n548,
    n282
  );


  buf
  g442
  (
    n522,
    n165
  );


  not
  g443
  (
    n688,
    n155
  );


  buf
  g444
  (
    n605,
    n276
  );


  not
  g445
  (
    n476,
    n219
  );


  buf
  g446
  (
    KeyWire_0_35,
    n372
  );


  not
  g447
  (
    n582,
    n330
  );


  buf
  g448
  (
    n669,
    n308
  );


  buf
  g449
  (
    n594,
    n240
  );


  not
  g450
  (
    n515,
    n239
  );


  buf
  g451
  (
    n520,
    n264
  );


  buf
  g452
  (
    n693,
    n167
  );


  not
  g453
  (
    KeyWire_0_13,
    n251
  );


  not
  g454
  (
    n531,
    n337
  );


  not
  g455
  (
    n483,
    n280
  );


  buf
  g456
  (
    n664,
    n255
  );


  buf
  g457
  (
    n597,
    n363
  );


  not
  g458
  (
    n622,
    n192
  );


  not
  g459
  (
    n464,
    n183
  );


  not
  g460
  (
    n658,
    n268
  );


  buf
  g461
  (
    n497,
    n299
  );


  not
  g462
  (
    n636,
    n375
  );


  not
  g463
  (
    n460,
    n259
  );


  not
  g464
  (
    n543,
    n289
  );


  buf
  g465
  (
    n540,
    n343
  );


  not
  g466
  (
    KeyWire_0_53,
    n179
  );


  not
  g467
  (
    n640,
    n228
  );


  not
  g468
  (
    n561,
    n168
  );


  buf
  g469
  (
    n519,
    n116
  );


  not
  g470
  (
    KeyWire_0_20,
    n333
  );


  buf
  g471
  (
    n612,
    n172
  );


  not
  g472
  (
    KeyWire_0_42,
    n244
  );


  buf
  g473
  (
    n484,
    n344
  );


  buf
  g474
  (
    n506,
    n233
  );


  buf
  g475
  (
    n526,
    n341
  );


  not
  g476
  (
    n695,
    n279
  );


  not
  g477
  (
    n678,
    n128
  );


  buf
  g478
  (
    n595,
    n366
  );


  buf
  g479
  (
    n538,
    n371
  );


  buf
  g480
  (
    n643,
    n326
  );


  buf
  g481
  (
    n705,
    n121
  );


  not
  g482
  (
    n498,
    n209
  );


  buf
  g483
  (
    n701,
    n364
  );


  not
  g484
  (
    n647,
    n367
  );


  not
  g485
  (
    n603,
    n360
  );


  buf
  g486
  (
    n635,
    n295
  );


  buf
  g487
  (
    n652,
    n294
  );


  not
  g488
  (
    n475,
    n150
  );


  not
  g489
  (
    n558,
    n374
  );


  not
  g490
  (
    n691,
    n277
  );


  not
  g491
  (
    n720,
    n114
  );


  not
  g492
  (
    n521,
    n199
  );


  not
  g493
  (
    n474,
    n307
  );


  not
  g494
  (
    n586,
    n328
  );


  buf
  g495
  (
    n591,
    n217
  );


  buf
  g496
  (
    n549,
    n313
  );


  not
  g497
  (
    n513,
    n296
  );


  not
  g498
  (
    n662,
    n317
  );


  buf
  g499
  (
    n651,
    n169
  );


  buf
  g500
  (
    n655,
    n229
  );


  not
  g501
  (
    n683,
    n113
  );


  buf
  g502
  (
    n562,
    n298
  );


  buf
  g503
  (
    n629,
    n250
  );


  buf
  g504
  (
    n479,
    n325
  );


  buf
  g505
  (
    n552,
    n272
  );


  buf
  g506
  (
    n539,
    n306
  );


  buf
  g507
  (
    n670,
    n186
  );


  buf
  g508
  (
    n523,
    n348
  );


  buf
  g509
  (
    n510,
    n257
  );


  buf
  g510
  (
    n639,
    n245
  );


  buf
  g511
  (
    n455,
    n370
  );


  not
  g512
  (
    n596,
    n133
  );


  buf
  g513
  (
    n686,
    n349
  );


  buf
  g514
  (
    KeyWire_0_5,
    n119
  );


  not
  g515
  (
    n576,
    n120
  );


  not
  g516
  (
    n575,
    n231
  );


  not
  g517
  (
    n713,
    n152
  );


  buf
  g518
  (
    n637,
    n124
  );


  not
  g519
  (
    n490,
    n287
  );


  buf
  g520
  (
    n516,
    n300
  );


  not
  g521
  (
    n661,
    n178
  );


  not
  g522
  (
    n602,
    n158
  );


  buf
  g523
  (
    n660,
    n314
  );


  not
  g524
  (
    KeyWire_0_60,
    n278
  );


  buf
  g525
  (
    n709,
    n241
  );


  buf
  g526
  (
    n710,
    n196
  );


  buf
  g527
  (
    n617,
    n310
  );


  buf
  g528
  (
    n625,
    n157
  );


  not
  g529
  (
    n524,
    n204
  );


  buf
  g530
  (
    n545,
    n146
  );


  not
  g531
  (
    n489,
    n225
  );


  not
  g532
  (
    n493,
    n297
  );


  buf
  g533
  (
    n703,
    n227
  );


  not
  g534
  (
    n467,
    n352
  );


  buf
  g535
  (
    n465,
    n160
  );


  buf
  g536
  (
    n624,
    n362
  );


  buf
  g537
  (
    n495,
    n164
  );


  not
  g538
  (
    n699,
    n135
  );


  not
  g539
  (
    n459,
    n347
  );


  buf
  g540
  (
    n588,
    n291
  );


  buf
  g541
  (
    n638,
    n117
  );


  buf
  g542
  (
    n657,
    n329
  );


  not
  g543
  (
    n674,
    n324
  );


  buf
  g544
  (
    KeyWire_0_39,
    n214
  );


  buf
  g545
  (
    n557,
    n187
  );


  not
  g546
  (
    KeyWire_0_32,
    n208
  );


  not
  g547
  (
    n700,
    n321
  );


  not
  g548
  (
    n466,
    n185
  );


  not
  g549
  (
    n572,
    n207
  );


  not
  g550
  (
    n458,
    n200
  );


  not
  g551
  (
    n611,
    n222
  );


  not
  g552
  (
    n554,
    n191
  );


  buf
  g553
  (
    n537,
    n145
  );


  buf
  g554
  (
    n716,
    n248
  );


  not
  g555
  (
    n619,
    n267
  );


  not
  g556
  (
    KeyWire_0_2,
    n170
  );


  not
  g557
  (
    KeyWire_0_54,
    n127
  );


  not
  g558
  (
    n491,
    n198
  );


  buf
  g559
  (
    n461,
    n184
  );


  not
  g560
  (
    KeyWire_0_37,
    n258
  );


  buf
  g561
  (
    n579,
    n355
  );


  not
  g562
  (
    n599,
    n223
  );


  buf
  g563
  (
    n604,
    n327
  );


  not
  g564
  (
    KeyWire_0_25,
    n309
  );


  buf
  g565
  (
    n573,
    n288
  );


  not
  g566
  (
    n477,
    n115
  );


  buf
  g567
  (
    n518,
    n320
  );


  not
  g568
  (
    n634,
    n260
  );


  buf
  g569
  (
    n690,
    n205
  );


  buf
  g570
  (
    n616,
    n273
  );


  not
  g571
  (
    n481,
    n190
  );


  not
  g572
  (
    n566,
    n256
  );


  buf
  g573
  (
    n470,
    n351
  );


  buf
  g574
  (
    n463,
    n141
  );


  not
  g575
  (
    n544,
    n318
  );


  not
  g576
  (
    n711,
    n226
  );


  buf
  g577
  (
    n666,
    n266
  );


  not
  g578
  (
    n528,
    n206
  );


  buf
  g579
  (
    n584,
    n131
  );


  not
  g580
  (
    n712,
    n215
  );


  not
  g581
  (
    n564,
    n130
  );


  not
  g582
  (
    n512,
    n358
  );


  buf
  g583
  (
    n677,
    n175
  );


  buf
  g584
  (
    n646,
    n147
  );


  buf
  g585
  (
    n472,
    n247
  );


  not
  g586
  (
    n671,
    n177
  );


  buf
  g587
  (
    n719,
    n243
  );


  not
  g588
  (
    n456,
    n202
  );


  not
  g589
  (
    n650,
    n357
  );


  buf
  g590
  (
    n680,
    n249
  );


  buf
  g591
  (
    n697,
    n305
  );


  buf
  g592
  (
    n621,
    n335
  );


  buf
  g593
  (
    n536,
    n189
  );


  buf
  g594
  (
    n718,
    n353
  );


  buf
  g595
  (
    n694,
    n293
  );


  not
  g596
  (
    n644,
    n144
  );


  buf
  g597
  (
    n482,
    n230
  );


  buf
  g598
  (
    n567,
    n292
  );


  not
  g599
  (
    KeyWire_0_24,
    n159
  );


  not
  g600
  (
    KeyWire_0_6,
    n336
  );


  not
  g601
  (
    n684,
    n220
  );


  not
  g602
  (
    n468,
    n193
  );


  not
  g603
  (
    n620,
    n376
  );


  buf
  g604
  (
    n606,
    n261
  );


  not
  g605
  (
    n608,
    n224
  );


  not
  g606
  (
    n668,
    n125
  );


  not
  g607
  (
    n626,
    n232
  );


  not
  g608
  (
    n714,
    n302
  );


  buf
  g609
  (
    n601,
    n195
  );


  buf
  g610
  (
    n457,
    n162
  );


  buf
  g611
  (
    n574,
    n253
  );


  buf
  g612
  (
    n535,
    n369
  );


  not
  g613
  (
    n673,
    n180
  );


  buf
  g614
  (
    KeyWire_0_8,
    n161
  );


  not
  g615
  (
    n532,
    n118
  );


  buf
  g616
  (
    n631,
    n286
  );


  not
  g617
  (
    n698,
    n213
  );


  buf
  g618
  (
    n559,
    n263
  );


  not
  g619
  (
    n501,
    n181
  );


  buf
  g620
  (
    n663,
    n111
  );


  buf
  g621
  (
    KeyWire_0_29,
    n359
  );


  not
  g622
  (
    n496,
    n346
  );


  not
  g623
  (
    n530,
    n342
  );


  buf
  g624
  (
    n534,
    n163
  );


  buf
  g625
  (
    n682,
    n140
  );


  not
  g626
  (
    n615,
    n143
  );


  not
  g627
  (
    n648,
    n194
  );


  buf
  g628
  (
    n485,
    n262
  );


  not
  g629
  (
    n642,
    n174
  );


  buf
  g630
  (
    n614,
    n156
  );


  not
  g631
  (
    n565,
    n271
  );


  not
  g632
  (
    n715,
    n284
  );


  not
  g633
  (
    n585,
    n301
  );


  buf
  g634
  (
    n627,
    n126
  );


  buf
  g635
  (
    n581,
    n138
  );


  not
  g636
  (
    n488,
    n149
  );


  not
  g637
  (
    n471,
    n123
  );


  buf
  g638
  (
    n480,
    n265
  );


  not
  g639
  (
    n609,
    n203
  );


  not
  g640
  (
    n499,
    n171
  );


  buf
  g641
  (
    n578,
    n212
  );


  buf
  g642
  (
    n577,
    n303
  );


  not
  g643
  (
    n509,
    n345
  );


  not
  g644
  (
    n473,
    n323
  );


  buf
  g645
  (
    KeyWire_0_52,
    n142
  );


  buf
  g646
  (
    n503,
    n129
  );


  not
  g647
  (
    KeyWire_0_46,
    n350
  );


  not
  g648
  (
    n681,
    n356
  );


  not
  g649
  (
    KeyWire_0_12,
    n237
  );


  buf
  g650
  (
    n462,
    n270
  );


  not
  g651
  (
    n659,
    n153
  );


  not
  g652
  (
    n689,
    n112
  );


  buf
  g653
  (
    n555,
    n197
  );


  not
  g654
  (
    n560,
    n368
  );


  buf
  g655
  (
    n704,
    n331
  );


  not
  g656
  (
    n533,
    n274
  );


  buf
  g657
  (
    n486,
    n173
  );


  buf
  g658
  (
    n563,
    n201
  );


  buf
  g659
  (
    n656,
    n188
  );


  not
  g660
  (
    n571,
    n285
  );


  buf
  g661
  (
    n502,
    n242
  );


  buf
  g662
  (
    n525,
    n269
  );


  not
  g663
  (
    n580,
    n275
  );


  buf
  g664
  (
    n529,
    n137
  );


  not
  g665
  (
    n547,
    n339
  );


  buf
  g666
  (
    KeyWire_0_59,
    n136
  );


  not
  g667
  (
    n504,
    n134
  );


  buf
  g668
  (
    n672,
    n154
  );


  not
  g669
  (
    n665,
    n361
  );


  not
  g670
  (
    n550,
    n332
  );


  buf
  g671
  (
    n632,
    n304
  );


  not
  g672
  (
    n487,
    n252
  );


  buf
  g673
  (
    n592,
    n132
  );


  buf
  g674
  (
    n553,
    n166
  );


  not
  g675
  (
    n654,
    n139
  );


  not
  g676
  (
    n568,
    n311
  );


  buf
  g677
  (
    n607,
    n218
  );


  buf
  g678
  (
    n593,
    n354
  );


  not
  g679
  (
    n556,
    n221
  );


  buf
  g680
  (
    n623,
    n338
  );


  not
  g681
  (
    n570,
    n148
  );


  buf
  g682
  (
    n692,
    n246
  );


  not
  g683
  (
    n687,
    n151
  );


  not
  g684
  (
    n590,
    n283
  );


  buf
  g685
  (
    n551,
    n334
  );


  buf
  g686
  (
    n508,
    n319
  );


  buf
  g687
  (
    n542,
    n235
  );


  not
  g688
  (
    n569,
    n290
  );


  buf
  g689
  (
    n598,
    n322
  );


  buf
  g690
  (
    n505,
    n182
  );


  not
  g691
  (
    n685,
    n176
  );


  buf
  g692
  (
    n600,
    n316
  );


  not
  g693
  (
    n469,
    n340
  );


  not
  g694
  (
    n633,
    n365
  );


  buf
  g695
  (
    n527,
    n210
  );


  not
  g696
  (
    n645,
    n281
  );


  buf
  g697
  (
    n649,
    n312
  );


  not
  g698
  (
    n732,
    n456
  );


  not
  g699
  (
    n724,
    n474
  );


  buf
  g700
  (
    n740,
    n109
  );


  buf
  g701
  (
    n731,
    n465
  );


  not
  g702
  (
    n738,
    n458
  );


  not
  g703
  (
    n726,
    n470
  );


  not
  g704
  (
    n734,
    n467
  );


  not
  g705
  (
    n727,
    n110
  );


  buf
  g706
  (
    n736,
    n469
  );


  not
  g707
  (
    n741,
    n110
  );


  buf
  g708
  (
    n737,
    n461
  );


  not
  g709
  (
    n739,
    n462
  );


  not
  g710
  (
    n728,
    n463
  );


  buf
  g711
  (
    n723,
    n475
  );


  not
  g712
  (
    n729,
    n455
  );


  buf
  g713
  (
    n722,
    n459
  );


  not
  g714
  (
    n725,
    n457
  );


  buf
  g715
  (
    n735,
    n110
  );


  xor
  g716
  (
    n733,
    n468,
    n109
  );


  xnor
  g717
  (
    n721,
    n466,
    n109,
    n471,
    n472
  );


  xor
  g718
  (
    n730,
    n460,
    n464,
    n473,
    n109
  );


  nor
  g719
  (
    n744,
    n387,
    n388,
    n390,
    n381
  );


  and
  g720
  (
    n743,
    n378,
    n385,
    n386,
    n721
  );


  xnor
  g721
  (
    n742,
    n391,
    n379,
    n722,
    n389
  );


  nor
  g722
  (
    n745,
    n721,
    n721,
    n382,
    n377
  );


  xor
  g723
  (
    n746,
    n383,
    n384,
    n380,
    n721
  );


  buf
  g724
  (
    n756,
    n744
  );


  buf
  g725
  (
    n754,
    n745
  );


  buf
  g726
  (
    n752,
    n743
  );


  not
  g727
  (
    n750,
    n746
  );


  buf
  g728
  (
    n755,
    n745
  );


  buf
  g729
  (
    n753,
    n744
  );


  not
  g730
  (
    n748,
    n746
  );


  not
  g731
  (
    n751,
    n746
  );


  not
  g732
  (
    n749,
    n742
  );


  not
  g733
  (
    n747,
    n746
  );


  or
  g734
  (
    n757,
    n570,
    n555,
    n724,
    n565
  );


  xnor
  g735
  (
    n769,
    n756,
    n573,
    n753,
    n748
  );


  and
  g736
  (
    n767,
    n509,
    n723,
    n722,
    n559
  );


  or
  g737
  (
    n796,
    n581,
    n748,
    n750,
    n499
  );


  nor
  g738
  (
    n766,
    n569,
    n537,
    n545,
    n747
  );


  and
  g739
  (
    n764,
    n492,
    n749,
    n723,
    n479
  );


  nand
  g740
  (
    n792,
    n562,
    n481,
    n755,
    n513
  );


  and
  g741
  (
    n794,
    n501,
    n483,
    n477,
    n753
  );


  xnor
  g742
  (
    n784,
    n533,
    n502,
    n564,
    n482
  );


  xnor
  g743
  (
    n773,
    n560,
    n529,
    n514,
    n568
  );


  nor
  g744
  (
    KeyWire_0_28,
    n519,
    n500,
    n556,
    n749
  );


  xor
  g745
  (
    n776,
    n486,
    n756,
    n579,
    n722
  );


  nor
  g746
  (
    n775,
    n561,
    n751,
    n574,
    n554
  );


  or
  g747
  (
    n786,
    n520,
    n724,
    n539,
    n522
  );


  and
  g748
  (
    n785,
    n582,
    n532,
    n535,
    n753
  );


  nand
  g749
  (
    n770,
    n542,
    n480,
    n505,
    n750
  );


  or
  g750
  (
    n774,
    n498,
    n507,
    n755
  );


  xor
  g751
  (
    n779,
    n752,
    n495,
    n546,
    n563
  );


  xor
  g752
  (
    n758,
    n572,
    n516,
    n724,
    n547
  );


  and
  g753
  (
    n790,
    n530,
    n577,
    n724,
    n747
  );


  nor
  g754
  (
    n793,
    n750,
    n749,
    n752,
    n511
  );


  or
  g755
  (
    n795,
    n755,
    n557,
    n576,
    n578
  );


  xnor
  g756
  (
    n781,
    n536,
    n566,
    n749,
    n747
  );


  and
  g757
  (
    KeyWire_0_11,
    n506,
    n508,
    n521,
    n484
  );


  nand
  g758
  (
    n762,
    n752,
    n754,
    n751,
    n515
  );


  xor
  g759
  (
    n780,
    n723,
    n490,
    n534,
    n524
  );


  xor
  g760
  (
    n760,
    n494,
    n722,
    n553,
    n551
  );


  xnor
  g761
  (
    n791,
    n567,
    n493,
    n523,
    n751
  );


  xnor
  g762
  (
    n783,
    n754,
    n512,
    n571,
    n748
  );


  nor
  g763
  (
    n778,
    n525,
    n580,
    n753,
    n517
  );


  nand
  g764
  (
    n761,
    n531,
    n550,
    n504,
    n725
  );


  nor
  g765
  (
    n772,
    n558,
    n751,
    n497,
    n723
  );


  nor
  g766
  (
    n777,
    n754,
    n541,
    n488,
    n496
  );


  xor
  g767
  (
    n788,
    n544,
    n476,
    n575,
    n552
  );


  xnor
  g768
  (
    n759,
    n518,
    n487,
    n748,
    n756
  );


  and
  g769
  (
    n765,
    n478,
    n491,
    n583,
    n510
  );


  and
  g770
  (
    n789,
    n750,
    n754,
    n489,
    n548
  );


  xor
  g771
  (
    n763,
    n747,
    n538,
    n549,
    n503
  );


  nor
  g772
  (
    n768,
    n527,
    n756,
    n526,
    n752
  );


  or
  g773
  (
    n782,
    n485,
    n540,
    n528,
    n543
  );


  xor
  g774
  (
    n801,
    n726,
    n760
  );


  buf
  g775
  (
    n799,
    n727
  );


  or
  g776
  (
    n798,
    n726,
    n726,
    n761,
    n758
  );


  nor
  g777
  (
    n797,
    n727,
    n725
  );


  nand
  g778
  (
    n800,
    n725,
    n759,
    n757,
    n726
  );


  nand
  g779
  (
    n806,
    n799,
    n395
  );


  nand
  g780
  (
    n805,
    n729,
    n798
  );


  nand
  g781
  (
    n802,
    n403,
    n800,
    n407,
    n732
  );


  xor
  g782
  (
    n810,
    n801,
    n766,
    n798,
    n730
  );


  xnor
  g783
  (
    n803,
    n762,
    n400,
    n801,
    n733
  );


  nor
  g784
  (
    n816,
    n800,
    n404,
    n731,
    n110
  );


  and
  g785
  (
    n807,
    n729,
    n799,
    n393,
    n733
  );


  nand
  g786
  (
    n814,
    n729,
    n399,
    n732
  );


  xor
  g787
  (
    n817,
    n798,
    n732,
    n402,
    n730
  );


  or
  g788
  (
    n808,
    n801,
    n800,
    n728,
    n406
  );


  or
  g789
  (
    n811,
    n798,
    n799,
    n764,
    n801
  );


  or
  g790
  (
    n809,
    n405,
    n731,
    n396,
    n401
  );


  or
  g791
  (
    n804,
    n392,
    n765,
    n730,
    n800
  );


  xor
  g792
  (
    n815,
    n398,
    n728,
    n730
  );


  and
  g793
  (
    n813,
    n799,
    n763,
    n731,
    n397
  );


  nor
  g794
  (
    n812,
    n731,
    n729,
    n728,
    n394
  );


  buf
  g795
  (
    n820,
    n785
  );


  buf
  g796
  (
    n826,
    n803
  );


  buf
  g797
  (
    n823,
    n771
  );


  not
  g798
  (
    n830,
    n783
  );


  buf
  g799
  (
    n828,
    n806
  );


  not
  g800
  (
    n824,
    n781
  );


  buf
  g801
  (
    n831,
    n813
  );


  not
  g802
  (
    n825,
    n773
  );


  or
  g803
  (
    n822,
    n811,
    n774,
    n812
  );


  or
  g804
  (
    n821,
    n769,
    n776,
    n813
  );


  xnor
  g805
  (
    KeyWire_0_34,
    n778,
    n808,
    n813
  );


  nand
  g806
  (
    n834,
    n811,
    n784,
    n813
  );


  or
  g807
  (
    n819,
    n782,
    n809,
    n767
  );


  xor
  g808
  (
    n818,
    n802,
    n779,
    n772
  );


  nand
  g809
  (
    n832,
    n775,
    n810,
    n807
  );


  nand
  g810
  (
    n829,
    n805,
    n812,
    n777
  );


  xnor
  g811
  (
    n833,
    n804,
    n780,
    n768,
    n770
  );


  buf
  g812
  (
    n841,
    n819
  );


  buf
  g813
  (
    n852,
    n819
  );


  not
  g814
  (
    KeyWire_0_17,
    n822
  );


  buf
  g815
  (
    n856,
    n822
  );


  not
  g816
  (
    n854,
    n823
  );


  not
  g817
  (
    n835,
    n818
  );


  buf
  g818
  (
    n838,
    n822
  );


  buf
  g819
  (
    n851,
    n822
  );


  not
  g820
  (
    n853,
    n820
  );


  buf
  g821
  (
    n855,
    n821
  );


  not
  g822
  (
    n839,
    n823
  );


  not
  g823
  (
    n850,
    n820
  );


  buf
  g824
  (
    n849,
    n821
  );


  buf
  g825
  (
    n848,
    n820
  );


  not
  g826
  (
    n837,
    n818
  );


  not
  g827
  (
    n846,
    n818
  );


  buf
  g828
  (
    n844,
    n819
  );


  not
  g829
  (
    n836,
    n818
  );


  not
  g830
  (
    n840,
    n819
  );


  buf
  g831
  (
    n842,
    n821
  );


  buf
  g832
  (
    n845,
    n820
  );


  not
  g833
  (
    n847,
    n821
  );


  buf
  g834
  (
    n864,
    n816
  );


  buf
  g835
  (
    n872,
    n823
  );


  not
  g836
  (
    n882,
    n851
  );


  not
  g837
  (
    n893,
    n836
  );


  not
  g838
  (
    n873,
    n824
  );


  not
  g839
  (
    n930,
    n607
  );


  not
  g840
  (
    n943,
    n601
  );


  buf
  g841
  (
    n892,
    n637
  );


  not
  g842
  (
    n890,
    n590
  );


  not
  g843
  (
    n917,
    n845
  );


  not
  g844
  (
    n895,
    n837
  );


  buf
  g845
  (
    KeyWire_0_26,
    n838
  );


  not
  g846
  (
    n939,
    n814
  );


  buf
  g847
  (
    n867,
    n609
  );


  buf
  g848
  (
    n871,
    n619
  );


  buf
  g849
  (
    n906,
    n602
  );


  not
  g850
  (
    n858,
    n855
  );


  not
  g851
  (
    n910,
    n850
  );


  buf
  g852
  (
    n868,
    n734
  );


  not
  g853
  (
    n921,
    n817
  );


  not
  g854
  (
    n905,
    n814
  );


  not
  g855
  (
    n860,
    n587
  );


  buf
  g856
  (
    n874,
    n854
  );


  not
  g857
  (
    n907,
    n824
  );


  buf
  g858
  (
    n880,
    n856
  );


  buf
  g859
  (
    n916,
    n618
  );


  not
  g860
  (
    n898,
    n627
  );


  buf
  g861
  (
    n883,
    n625
  );


  not
  g862
  (
    n926,
    n635
  );


  buf
  g863
  (
    n942,
    n854
  );


  not
  g864
  (
    n870,
    n622
  );


  buf
  g865
  (
    n908,
    n639
  );


  not
  g866
  (
    n887,
    n849
  );


  buf
  g867
  (
    n903,
    n851
  );


  not
  g868
  (
    n859,
    n849
  );


  buf
  g869
  (
    n941,
    n646
  );


  buf
  g870
  (
    n857,
    n856
  );


  not
  g871
  (
    n878,
    n825
  );


  nand
  g872
  (
    n904,
    n855,
    n410,
    n837
  );


  or
  g873
  (
    n894,
    n612,
    n846,
    n836
  );


  xnor
  g874
  (
    n919,
    n852,
    n598,
    n847
  );


  and
  g875
  (
    n925,
    n817,
    n814,
    n848
  );


  nor
  g876
  (
    n901,
    n610,
    n816,
    n851
  );


  xnor
  g877
  (
    n862,
    n630,
    n588,
    n854
  );


  and
  g878
  (
    n900,
    n852,
    n847,
    n733
  );


  nand
  g879
  (
    n922,
    n606,
    n599,
    n611
  );


  xor
  g880
  (
    n937,
    n815,
    n641,
    n624
  );


  nand
  g881
  (
    n931,
    n824,
    n620,
    n584
  );


  xnor
  g882
  (
    n879,
    n632,
    n592,
    n629
  );


  xor
  g883
  (
    n935,
    n837,
    n851,
    n839
  );


  or
  g884
  (
    n913,
    n642,
    n605,
    n841
  );


  xnor
  g885
  (
    n923,
    n600,
    n591,
    n586
  );


  and
  g886
  (
    n889,
    n835,
    n817,
    n849
  );


  nand
  g887
  (
    n912,
    n845,
    n855,
    n413
  );


  nand
  g888
  (
    n944,
    n604,
    n733,
    n848
  );


  and
  g889
  (
    n918,
    n636,
    n854,
    n846
  );


  xor
  g890
  (
    n865,
    n848,
    n838,
    n852
  );


  nor
  g891
  (
    n933,
    n594,
    n852,
    n855
  );


  xnor
  g892
  (
    n896,
    n643,
    n409,
    n825
  );


  and
  g893
  (
    n915,
    n839,
    n846,
    n853
  );


  or
  g894
  (
    n897,
    n853,
    n628,
    n633
  );


  or
  g895
  (
    n909,
    n824,
    n815,
    n408
  );


  xnor
  g896
  (
    n888,
    n615,
    n839,
    n617
  );


  or
  g897
  (
    n891,
    n836,
    n817,
    n596
  );


  nor
  g898
  (
    n920,
    n626,
    n843,
    n853
  );


  nand
  g899
  (
    n940,
    n623,
    n843,
    n608
  );


  nor
  g900
  (
    n899,
    n836,
    n843
  );


  and
  g901
  (
    n877,
    n638,
    n585,
    n840
  );


  nor
  g902
  (
    n902,
    n816,
    n846,
    n837
  );


  xor
  g903
  (
    n876,
    n853,
    n838,
    n840
  );


  xnor
  g904
  (
    n886,
    n835,
    n411,
    n644
  );


  nand
  g905
  (
    n934,
    n734,
    n845,
    n835
  );


  nor
  g906
  (
    n863,
    n844,
    n842,
    n847
  );


  nand
  g907
  (
    n929,
    n841,
    n850,
    n835
  );


  and
  g908
  (
    n927,
    n595,
    n640,
    n840
  );


  xor
  g909
  (
    n869,
    n841,
    n845,
    n850
  );


  nor
  g910
  (
    n928,
    n844,
    n841,
    n631
  );


  nor
  g911
  (
    n936,
    n823,
    n734,
    n815
  );


  xnor
  g912
  (
    n884,
    n634,
    n814,
    n589
  );


  and
  g913
  (
    n875,
    n614,
    n645,
    n597
  );


  nand
  g914
  (
    n881,
    n734,
    n850,
    n847
  );


  xor
  g915
  (
    n924,
    n840,
    n839,
    n856
  );


  or
  g916
  (
    n866,
    n849,
    n848,
    n621
  );


  or
  g917
  (
    n914,
    n842,
    n838,
    n816
  );


  and
  g918
  (
    n861,
    n842,
    n825,
    n616
  );


  or
  g919
  (
    n911,
    n613,
    n603,
    n856
  );


  or
  g920
  (
    n932,
    n842,
    n844
  );


  nor
  g921
  (
    n938,
    n815,
    n412,
    n593
  );


  buf
  g922
  (
    n949,
    n860
  );


  not
  g923
  (
    n950,
    n859
  );


  not
  g924
  (
    n946,
    n827
  );


  not
  g925
  (
    n945,
    n825
  );


  or
  g926
  (
    n952,
    n862,
    n826
  );


  buf
  g927
  (
    n947,
    n826
  );


  xor
  g928
  (
    n951,
    n827,
    n865
  );


  and
  g929
  (
    n953,
    n858,
    n863
  );


  xnor
  g930
  (
    n948,
    n861,
    n864,
    n866,
    n826
  );


  nand
  g931
  (
    n954,
    n950,
    n831,
    n949,
    n832
  );


  nor
  g932
  (
    n955,
    n830,
    n828,
    n832
  );


  or
  g933
  (
    n958,
    n832,
    n946,
    n828,
    n831
  );


  xor
  g934
  (
    n957,
    n830,
    n830,
    n945,
    n951
  );


  or
  g935
  (
    n959,
    n831,
    n831,
    n830,
    n827
  );


  and
  g936
  (
    n956,
    n948,
    n829
  );


  xnor
  g937
  (
    n960,
    n827,
    n947,
    n828,
    n829
  );


  buf
  g938
  (
    n963,
    n958
  );


  not
  g939
  (
    n962,
    n868
  );


  nor
  g940
  (
    n964,
    n867,
    n956
  );


  xnor
  g941
  (
    n961,
    n955,
    n870,
    n869,
    n957
  );


  or
  g942
  (
    n974,
    n872,
    n884,
    n885,
    n880
  );


  xor
  g943
  (
    n978,
    n889,
    n963,
    n886,
    n871
  );


  xnor
  g944
  (
    n972,
    n883,
    n962,
    n961
  );


  nor
  g945
  (
    n975,
    n875,
    n874,
    n883,
    n890
  );


  xor
  g946
  (
    n970,
    n964,
    n964,
    n886,
    n873
  );


  and
  g947
  (
    n965,
    n877,
    n881,
    n889,
    n961
  );


  xnor
  g948
  (
    n967,
    n873,
    n871,
    n882,
    n891
  );


  or
  g949
  (
    n973,
    n872,
    n878,
    n963,
    n962
  );


  xnor
  g950
  (
    n969,
    n881,
    n880,
    n887,
    n964
  );


  xor
  g951
  (
    n976,
    n875,
    n876,
    n874,
    n877
  );


  and
  g952
  (
    n968,
    n890,
    n964,
    n878,
    n888
  );


  xnor
  g953
  (
    n977,
    n884,
    n887,
    n885,
    n963
  );


  xor
  g954
  (
    n966,
    n870,
    n962,
    n879,
    n882
  );


  and
  g955
  (
    n971,
    n879,
    n876,
    n963,
    n888
  );


  xnor
  g956
  (
    n1010,
    n650,
    n970,
    n897,
    n911
  );


  xnor
  g957
  (
    n1031,
    n917,
    n453,
    n918,
    n978
  );


  and
  g958
  (
    n992,
    n735,
    n921,
    n938
  );


  or
  g959
  (
    n1032,
    n938,
    n975,
    n939,
    n910
  );


  and
  g960
  (
    n981,
    n970,
    n654,
    n972,
    n923
  );


  nand
  g961
  (
    n987,
    n973,
    n976,
    n433,
    n897
  );


  nor
  g962
  (
    n1013,
    n929,
    n904,
    n454,
    n736
  );


  xnor
  g963
  (
    n1019,
    n429,
    n926,
    n925,
    n900
  );


  xnor
  g964
  (
    n1002,
    n913,
    n932,
    n903,
    n417
  );


  xnor
  g965
  (
    n997,
    n978,
    n967,
    n917,
    n973
  );


  and
  g966
  (
    n998,
    n927,
    n738,
    n932,
    n892
  );


  and
  g967
  (
    n1015,
    n442,
    n444,
    n934,
    n909
  );


  and
  g968
  (
    n985,
    n904,
    n905,
    n914,
    n968
  );


  xnor
  g969
  (
    n1021,
    n927,
    n911,
    n968,
    n965
  );


  and
  g970
  (
    n1027,
    n912,
    n910,
    n905,
    n965
  );


  or
  g971
  (
    n983,
    n420,
    n647,
    n900,
    n649
  );


  xor
  g972
  (
    n990,
    n738,
    n967
  );


  xor
  g973
  (
    n1023,
    n924,
    n907,
    n893,
    n916
  );


  xnor
  g974
  (
    n1001,
    n972,
    n737,
    n977,
    n447
  );


  and
  g975
  (
    n1012,
    n448,
    n894,
    n432,
    n974
  );


  nand
  g976
  (
    n1000,
    n423,
    n902,
    n965,
    n971
  );


  and
  g977
  (
    n1033,
    n419,
    n440,
    n915,
    n976
  );


  nand
  g978
  (
    n979,
    n935,
    n437,
    n975,
    n895
  );


  xnor
  g979
  (
    n984,
    n972,
    n971,
    n976,
    n908
  );


  nand
  g980
  (
    KeyWire_0_47,
    n735,
    n931,
    n431
  );


  or
  g981
  (
    KeyWire_0_51,
    n446,
    n439,
    n973,
    n435
  );


  nor
  g982
  (
    n995,
    n975,
    n925,
    n969,
    n919
  );


  or
  g983
  (
    n986,
    n939,
    n434,
    n960,
    n936
  );


  and
  g984
  (
    n1007,
    n736,
    n973,
    n930,
    n896
  );


  xor
  g985
  (
    n1003,
    n968,
    n966,
    n924,
    n923
  );


  and
  g986
  (
    n999,
    n937,
    n445,
    n953,
    n906
  );


  nand
  g987
  (
    n1028,
    n928,
    n922,
    n451,
    n735
  );


  xnor
  g988
  (
    n1004,
    n651,
    n430,
    n930,
    n909
  );


  nand
  g989
  (
    n996,
    n898,
    n922,
    n449,
    n899
  );


  or
  g990
  (
    n980,
    n892,
    n977,
    n920,
    n899
  );


  nor
  g991
  (
    n1006,
    n935,
    n418,
    n966,
    n450
  );


  xor
  g992
  (
    n982,
    n425,
    n938,
    n933,
    n969
  );


  xnor
  g993
  (
    n993,
    n736,
    n967,
    n414,
    n966
  );


  nor
  g994
  (
    n1005,
    n933,
    n959,
    n914,
    n901
  );


  and
  g995
  (
    n994,
    n978,
    n436,
    n912,
    n974
  );


  xnor
  g996
  (
    n1018,
    n975,
    n926,
    n907,
    n452
  );


  xnor
  g997
  (
    n1026,
    n969,
    n928,
    n426,
    n648
  );


  and
  g998
  (
    KeyWire_0_31,
    n913,
    n965,
    n416,
    n428
  );


  nor
  g999
  (
    n989,
    n415,
    n934,
    n971,
    n920
  );


  xnor
  g1000
  (
    n1034,
    n921,
    n974,
    n915,
    n438
  );


  nand
  g1001
  (
    KeyWire_0_56,
    n978,
    n966,
    n652,
    n422
  );


  xor
  g1002
  (
    n1020,
    n653,
    n443,
    n421,
    n895
  );


  or
  g1003
  (
    n1011,
    n977,
    n972,
    n737,
    n427
  );


  xnor
  g1004
  (
    n988,
    n937,
    n441,
    n919,
    n971
  );


  or
  g1005
  (
    n1014,
    n970,
    n976,
    n969,
    n896
  );


  nand
  g1006
  (
    n1024,
    n977,
    n918,
    n968,
    n902
  );


  or
  g1007
  (
    n1008,
    n891,
    n737,
    n736,
    n898
  );


  nor
  g1008
  (
    n1029,
    n929,
    n908,
    n424,
    n952
  );


  xnor
  g1009
  (
    n1025,
    n936,
    n903,
    n893,
    n916
  );


  xor
  g1010
  (
    n1030,
    n906,
    n974,
    n970,
    n735
  );


  xnor
  g1011
  (
    n1017,
    n894,
    n737,
    n901,
    n939
  );


  nor
  g1012
  (
    n1078,
    n787,
    n740
  );


  xor
  g1013
  (
    n1070,
    n994,
    n987,
    n789
  );


  xnor
  g1014
  (
    n1041,
    n993,
    n992,
    n678
  );


  xnor
  g1015
  (
    n1045,
    n994,
    n942,
    n990
  );


  xor
  g1016
  (
    n1047,
    n659,
    n984,
    n940
  );


  nor
  g1017
  (
    n1058,
    n834,
    n792
  );


  and
  g1018
  (
    n1039,
    n703,
    n940,
    n671
  );


  nor
  g1019
  (
    n1100,
    n987,
    n705,
    n719
  );


  nor
  g1020
  (
    n1053,
    n740,
    n688,
    n991
  );


  or
  g1021
  (
    n1077,
    n672,
    n656,
    n939
  );


  or
  g1022
  (
    n1096,
    n657,
    n942,
    n987
  );


  xor
  g1023
  (
    n1065,
    n980,
    n787,
    n833
  );


  or
  g1024
  (
    n1098,
    n982,
    n693,
    n986
  );


  nand
  g1025
  (
    n1064,
    n981,
    n996,
    n787
  );


  xor
  g1026
  (
    n1103,
    n994,
    n834,
    n790
  );


  xor
  g1027
  (
    n1060,
    n718,
    n658,
    n791
  );


  nor
  g1028
  (
    n1072,
    n994,
    n791,
    n665
  );


  and
  g1029
  (
    KeyWire_0_3,
    n941,
    n986,
    n791
  );


  nand
  g1030
  (
    n1056,
    n834,
    n674,
    n982
  );


  and
  g1031
  (
    n1049,
    n988,
    n704,
    n679
  );


  xnor
  g1032
  (
    n1094,
    n706,
    n739,
    n983
  );


  or
  g1033
  (
    n1051,
    n787,
    n986,
    n983
  );


  nor
  g1034
  (
    KeyWire_0_18,
    n995,
    n790,
    n708
  );


  nor
  g1035
  (
    n1059,
    n990,
    n833,
    n707
  );


  nor
  g1036
  (
    n1066,
    n943,
    n685,
    n716
  );


  or
  g1037
  (
    n1074,
    n993,
    n680,
    n995
  );


  nand
  g1038
  (
    n1061,
    n670,
    n788,
    n789
  );


  xor
  g1039
  (
    n1085,
    n687,
    n668,
    n663
  );


  and
  g1040
  (
    n1044,
    n983,
    n941,
    n833
  );


  and
  g1041
  (
    n1082,
    n992,
    n792,
    n720
  );


  or
  g1042
  (
    n1088,
    n980,
    n996,
    n667
  );


  or
  g1043
  (
    n1079,
    n701,
    n995,
    n991
  );


  nor
  g1044
  (
    n1038,
    n942,
    n660,
    n988
  );


  or
  g1045
  (
    n1040,
    n833,
    n709,
    n686
  );


  xor
  g1046
  (
    n1086,
    n790,
    n675,
    n989
  );


  xor
  g1047
  (
    n1046,
    n791,
    n990,
    n944
  );


  and
  g1048
  (
    n1080,
    n710,
    n677,
    n740
  );


  xor
  g1049
  (
    n1050,
    n664,
    n673,
    n943
  );


  nor
  g1050
  (
    n1068,
    n984,
    n940,
    n666
  );


  xor
  g1051
  (
    n1102,
    n984,
    n662,
    n981
  );


  xor
  g1052
  (
    n1054,
    n741,
    n991,
    n985
  );


  xnor
  g1053
  (
    n1069,
    n993,
    n943,
    n700
  );


  xnor
  g1054
  (
    n1071,
    n683,
    n987,
    n788
  );


  nor
  g1055
  (
    n1090,
    n741,
    n995,
    n989
  );


  xor
  g1056
  (
    n1043,
    n940,
    n944,
    n786
  );


  or
  g1057
  (
    KeyWire_0_62,
    n786,
    n689,
    n714
  );


  or
  g1058
  (
    n1099,
    n832,
    n989,
    n943
  );


  xnor
  g1059
  (
    n1084,
    n984,
    n996,
    n785
  );


  nand
  g1060
  (
    n1081,
    n982,
    n698,
    n717
  );


  xor
  g1061
  (
    n1093,
    n990,
    n942,
    n711
  );


  or
  g1062
  (
    n1063,
    n741,
    n980,
    n691
  );


  nand
  g1063
  (
    n1083,
    n993,
    n661,
    n985
  );


  nand
  g1064
  (
    n1101,
    n739,
    n741,
    n695
  );


  or
  g1065
  (
    n1036,
    n986,
    n712,
    n789
  );


  xor
  g1066
  (
    n1067,
    n992,
    n985,
    n941
  );


  nand
  g1067
  (
    n1097,
    n694,
    n697,
    n715
  );


  xnor
  g1068
  (
    n1076,
    n786,
    n985,
    n682
  );


  xnor
  g1069
  (
    n1035,
    n669,
    n980,
    n989
  );


  and
  g1070
  (
    n1037,
    n713,
    n790,
    n981
  );


  nor
  g1071
  (
    n1095,
    n738,
    n690,
    n788
  );


  and
  g1072
  (
    n1075,
    n740,
    n944,
    n982
  );


  nor
  g1073
  (
    n1052,
    n992,
    n702,
    n981
  );


  xor
  g1074
  (
    n1048,
    n789,
    n983,
    n988
  );


  nor
  g1075
  (
    n1042,
    n676,
    n739,
    n944
  );


  and
  g1076
  (
    KeyWire_0_58,
    n788,
    n996,
    n655
  );


  or
  g1077
  (
    n1073,
    n834,
    n991,
    n786
  );


  xnor
  g1078
  (
    n1092,
    n988,
    n684,
    n979
  );


  and
  g1079
  (
    n1089,
    n739,
    n941,
    n699
  );


  nor
  g1080
  (
    n1057,
    n681,
    n692,
    n696
  );


  and
  g1081
  (
    n1108,
    n1011,
    n1015,
    n1061,
    n1006
  );


  nand
  g1082
  (
    n1150,
    n1016,
    n1010,
    n1027,
    n1005
  );


  xnor
  g1083
  (
    n1110,
    n1006,
    n997,
    n1078,
    n1020
  );


  nand
  g1084
  (
    n1137,
    n1009,
    n1008,
    n1004
  );


  xnor
  g1085
  (
    n1151,
    n1074,
    n1019,
    n1021,
    n1037
  );


  or
  g1086
  (
    n1130,
    n796,
    n1002,
    n1021,
    n1026
  );


  nand
  g1087
  (
    n1107,
    n1011,
    n794,
    n1075,
    n1018
  );


  and
  g1088
  (
    n1126,
    n794,
    n1035,
    n1008,
    n1081
  );


  xnor
  g1089
  (
    n1153,
    n1039,
    n1000,
    n1029,
    n796
  );


  and
  g1090
  (
    n1142,
    n1023,
    n1027,
    n1014,
    n1049
  );


  xnor
  g1091
  (
    n1136,
    n1066,
    n1024,
    n1076,
    n1022
  );


  and
  g1092
  (
    n1114,
    n1003,
    n1020,
    n795,
    n1044
  );


  xor
  g1093
  (
    n1118,
    n1009,
    n1026,
    n1000,
    n1028
  );


  xnor
  g1094
  (
    n1111,
    n1003,
    n998,
    n1015,
    n1005
  );


  or
  g1095
  (
    n1134,
    n1006,
    n1065,
    n795,
    n1017
  );


  xnor
  g1096
  (
    n1145,
    n1014,
    n795,
    n793,
    n1062
  );


  or
  g1097
  (
    n1109,
    n1001,
    n1029,
    n1007,
    n1012
  );


  and
  g1098
  (
    n1139,
    n1023,
    n997,
    n1022,
    n1045
  );


  and
  g1099
  (
    n1123,
    n1016,
    n1024,
    n1068,
    n1072
  );


  nand
  g1100
  (
    n1127,
    n796,
    n1020,
    n1071,
    n1021
  );


  and
  g1101
  (
    n1120,
    n1059,
    n1046,
    n1027,
    n1016
  );


  xor
  g1102
  (
    n1121,
    n1056,
    n1050,
    n1007,
    n1003
  );


  and
  g1103
  (
    n1146,
    n1000,
    n792,
    n1012,
    n1040
  );


  xnor
  g1104
  (
    n1148,
    n1084,
    n1018,
    n1048,
    n1005
  );


  xor
  g1105
  (
    n1113,
    n1025,
    n1014,
    n1041,
    n1010
  );


  nand
  g1106
  (
    n1147,
    n1010,
    n1014,
    n1025,
    n999
  );


  xnor
  g1107
  (
    n1143,
    n1019,
    n1077,
    n1070,
    n1007
  );


  or
  g1108
  (
    n1122,
    n1069,
    n1073,
    n1036,
    n1023
  );


  or
  g1109
  (
    KeyWire_0_9,
    n1082,
    n1020,
    n1079,
    n1028
  );


  xnor
  g1110
  (
    n1135,
    n1016,
    n793,
    n997,
    n1023
  );


  xor
  g1111
  (
    n1133,
    n1017,
    n998,
    n1024,
    n1053
  );


  nand
  g1112
  (
    n1116,
    n1013,
    n1001,
    n1060,
    n1083
  );


  or
  g1113
  (
    n1105,
    n1029,
    n1015,
    n1028,
    n1008
  );


  nor
  g1114
  (
    n1112,
    n1054,
    n1009,
    n1025,
    n1022
  );


  nand
  g1115
  (
    n1138,
    n1013,
    n1057,
    n793,
    n1022
  );


  nor
  g1116
  (
    n1106,
    n1026,
    n1002,
    n1052,
    n1030
  );


  nand
  g1117
  (
    KeyWire_0_22,
    n1027,
    n1043,
    n1012,
    n1029
  );


  nor
  g1118
  (
    n1104,
    n1011,
    n1004,
    n1024,
    n1063
  );


  xor
  g1119
  (
    n1124,
    n1055,
    n1064,
    n1001,
    n796
  );


  and
  g1120
  (
    n1115,
    n1012,
    n998,
    n1080,
    n999
  );


  and
  g1121
  (
    n1152,
    n1013,
    n1017,
    n998,
    n1010
  );


  xnor
  g1122
  (
    n1128,
    n1017,
    n1051,
    n793,
    n1028
  );


  and
  g1123
  (
    n1117,
    n1067,
    n1004,
    n1019
  );


  nand
  g1124
  (
    n1144,
    n1002,
    n1018,
    n794,
    n1007
  );


  xor
  g1125
  (
    n1140,
    n1005,
    n1001,
    n997,
    n1011
  );


  xor
  g1126
  (
    n1132,
    n999,
    n1038,
    n794,
    n1000
  );


  xnor
  g1127
  (
    n1129,
    n1009,
    n1015,
    n1002,
    n1042
  );


  nand
  g1128
  (
    n1119,
    n1013,
    n999,
    n795,
    n1004
  );


  or
  g1129
  (
    n1131,
    n1047,
    n1006,
    n1003,
    n1058
  );


  and
  g1130
  (
    n1141,
    n1025,
    n1018,
    n1021,
    n1026
  );


  nor
  g1131
  (
    n1171,
    n1109,
    n1138,
    n1087,
    n1148
  );


  and
  g1132
  (
    n1161,
    n1095,
    n1091,
    n1092,
    n1105
  );


  xnor
  g1133
  (
    n1155,
    n1097,
    n1122,
    n1135,
    n1139
  );


  xor
  g1134
  (
    n1157,
    n1108,
    n1134,
    n1140,
    n1121
  );


  xor
  g1135
  (
    n1174,
    n1101,
    n1141,
    n1123,
    n1120
  );


  nand
  g1136
  (
    n1165,
    n1089,
    n1032,
    n1150,
    n1117
  );


  nand
  g1137
  (
    n1158,
    n1127,
    n1146,
    n1118,
    n1137
  );


  and
  g1138
  (
    n1170,
    n1114,
    n1103,
    n1034,
    n1130
  );


  xor
  g1139
  (
    KeyWire_0_15,
    n1144,
    n1153,
    n1034,
    n1133
  );


  xnor
  g1140
  (
    n1162,
    n1125,
    n1152,
    n1104,
    n1098
  );


  and
  g1141
  (
    n1164,
    n1086,
    n1096,
    n1129,
    n1030
  );


  and
  g1142
  (
    n1168,
    n1112,
    n1033,
    n1110,
    n1128
  );


  nand
  g1143
  (
    n1160,
    n1090,
    n1126,
    n1113,
    n1031
  );


  xor
  g1144
  (
    n1175,
    n1033,
    n1031,
    n1100,
    n1030
  );


  nand
  g1145
  (
    n1154,
    n1034,
    n1116,
    n1147,
    n1088
  );


  or
  g1146
  (
    n1156,
    n1093,
    n1106,
    n1031
  );


  and
  g1147
  (
    n1159,
    n1094,
    n1143,
    n1102,
    n1099
  );


  or
  g1148
  (
    n1163,
    n1142,
    n1111,
    n1131,
    n1107
  );


  or
  g1149
  (
    n1169,
    n1124,
    n1030,
    n1032,
    n1085
  );


  nor
  g1150
  (
    n1172,
    n1115,
    n1032,
    n1136,
    n1033
  );


  or
  g1151
  (
    n1173,
    n1151,
    n1034,
    n1033,
    n1145
  );


  xnor
  g1152
  (
    n1167,
    n1032,
    n1149,
    n1132,
    n1119
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n307,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n276,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n618,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1091,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n257,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n546,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n613,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n338,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n679,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1149,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n38,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n771,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n696,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n492,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n284,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1166,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n329,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n843,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n1055,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n282,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n706,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n121,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1125,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n40,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n708,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n494,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n885,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n342,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n787,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n517,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n26,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1016,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n583,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n397,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n827,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n511,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n165,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n507,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n140,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n541,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n316,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n201,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n717,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n147,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n204,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n368,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n702,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n1009,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n52,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n195,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n373,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n1022,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n630,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n500,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n707,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n36,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n991,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n253,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n1062,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n514,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n610,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n244,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n1087,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n295,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

