// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1591_53_6 written by SynthGen on 2021/05/24 19:45:40
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1591_53_6 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18,
 n1045, n1051, n1055, n1053, n1056, n1058, n1048, n1046,
 n1050, n1059, n1057, n1052, n1047, n1123, n1128, n1115,
 n1124, n1227, n1231, n1219, n1228, n1218, n1223, n1230,
 n1609);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18;

output n1045, n1051, n1055, n1053, n1056, n1058, n1048, n1046,
 n1050, n1059, n1057, n1052, n1047, n1123, n1128, n1115,
 n1124, n1227, n1231, n1219, n1228, n1218, n1223, n1230,
 n1609;

wire n19, n20, n21, n22, n23, n24, n25, n26,
 n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n487, n488, n489, n490,
 n491, n492, n493, n494, n495, n496, n497, n498,
 n499, n500, n501, n502, n503, n504, n505, n506,
 n507, n508, n509, n510, n511, n512, n513, n514,
 n515, n516, n517, n518, n519, n520, n521, n522,
 n523, n524, n525, n526, n527, n528, n529, n530,
 n531, n532, n533, n534, n535, n536, n537, n538,
 n539, n540, n541, n542, n543, n544, n545, n546,
 n547, n548, n549, n550, n551, n552, n553, n554,
 n555, n556, n557, n558, n559, n560, n561, n562,
 n563, n564, n565, n566, n567, n568, n569, n570,
 n571, n572, n573, n574, n575, n576, n577, n578,
 n579, n580, n581, n582, n583, n584, n585, n586,
 n587, n588, n589, n590, n591, n592, n593, n594,
 n595, n596, n597, n598, n599, n600, n601, n602,
 n603, n604, n605, n606, n607, n608, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n660, n661, n662, n663, n664, n665, n666,
 n667, n668, n669, n670, n671, n672, n673, n674,
 n675, n676, n677, n678, n679, n680, n681, n682,
 n683, n684, n685, n686, n687, n688, n689, n690,
 n691, n692, n693, n694, n695, n696, n697, n698,
 n699, n700, n701, n702, n703, n704, n705, n706,
 n707, n708, n709, n710, n711, n712, n713, n714,
 n715, n716, n717, n718, n719, n720, n721, n722,
 n723, n724, n725, n726, n727, n728, n729, n730,
 n731, n732, n733, n734, n735, n736, n737, n738,
 n739, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1049, n1054, n1060, n1061, n1062, n1063,
 n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
 n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
 n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
 n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
 n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
 n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
 n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1125, n1126, n1127, n1129, n1130, n1131,
 n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
 n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
 n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
 n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
 n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
 n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
 n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
 n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
 n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
 n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
 n1212, n1213, n1214, n1215, n1216, n1217, n1220, n1221,
 n1222, n1224, n1225, n1226, n1229, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608;

buf  g0 (n48, n13);
buf  g1 (n54, n5);
buf  g2 (n55, n10);
not  g3 (n53, n15);
not  g4 (n21, n12);
not  g5 (n52, n1);
not  g6 (n30, n9);
not  g7 (n79, n16);
not  g8 (n82, n11);
not  g9 (n78, n14);
not  g10 (n85, n8);
buf  g11 (n65, n2);
not  g12 (n47, n3);
buf  g13 (n87, n9);
not  g14 (n75, n2);
buf  g15 (n37, n11);
buf  g16 (n28, n15);
not  g17 (n62, n1);
not  g18 (n58, n8);
buf  g19 (n26, n6);
not  g20 (n76, n15);
buf  g21 (n44, n7);
buf  g22 (n33, n6);
not  g23 (n43, n3);
not  g24 (n77, n4);
buf  g25 (n81, n7);
not  g26 (n32, n10);
buf  g27 (n63, n9);
buf  g28 (n27, n6);
not  g29 (n22, n12);
buf  g30 (n36, n9);
not  g31 (n24, n7);
not  g32 (n20, n2);
buf  g33 (n59, n11);
not  g34 (n74, n16);
not  g35 (n64, n14);
not  g36 (n57, n14);
not  g37 (n86, n4);
not  g38 (n35, n8);
buf  g39 (n72, n7);
buf  g40 (n84, n6);
buf  g41 (n73, n8);
not  g42 (n19, n16);
not  g43 (n39, n10);
not  g44 (n69, n1);
buf  g45 (n68, n17);
not  g46 (n56, n12);
buf  g47 (n51, n10);
buf  g48 (n67, n5);
buf  g49 (n29, n11);
not  g50 (n61, n17);
not  g51 (n40, n16);
buf  g52 (n25, n13);
not  g53 (n42, n18);
not  g54 (n38, n5);
buf  g55 (n31, n14);
buf  g56 (n80, n17);
buf  g57 (n45, n2);
not  g58 (n50, n13);
not  g59 (n71, n4);
buf  g60 (n23, n13);
not  g61 (n66, n15);
not  g62 (n60, n5);
buf  g63 (n49, n3);
buf  g64 (n34, n17);
not  g65 (n41, n12);
buf  g66 (n70, n3);
buf  g67 (n83, n4);
not  g68 (n46, n1);
not  g69 (n88, n21);
buf  g70 (n93, n19);
not  g71 (n91, n19);
buf  g72 (n99, n19);
buf  g73 (n97, n20);
not  g74 (n92, n20);
not  g75 (n90, n20);
buf  g76 (n95, n19);
not  g77 (n89, n20);
buf  g78 (n98, n21);
buf  g79 (n94, n21);
not  g80 (n96, n21);
buf  g81 (n113, n88);
not  g82 (n124, n91);
not  g83 (n121, n92);
not  g84 (n112, n93);
not  g85 (n119, n89);
buf  g86 (n116, n92);
buf  g87 (n114, n94);
not  g88 (n117, n88);
not  g89 (n118, n89);
not  g90 (n127, n90);
not  g91 (n115, n90);
buf  g92 (n122, n90);
not  g93 (n103, n88);
not  g94 (n126, n89);
buf  g95 (n123, n94);
buf  g96 (n101, n94);
not  g97 (n109, n92);
buf  g98 (n120, n89);
buf  g99 (n108, n93);
buf  g100 (n100, n91);
buf  g101 (n107, n91);
buf  g102 (n125, n90);
buf  g103 (n102, n91);
not  g104 (n104, n88);
buf  g105 (n105, n93);
buf  g106 (n106, n94);
buf  g107 (n110, n93);
not  g108 (n111, n92);
buf  g109 (n176, n105);
buf  g110 (n189, n118);
not  g111 (n177, n118);
not  g112 (n200, n58);
not  g113 (n152, n74);
buf  g114 (n211, n115);
not  g115 (n231, n116);
buf  g116 (n179, n25);
not  g117 (n141, n47);
not  g118 (n161, n27);
buf  g119 (n159, n75);
not  g120 (n167, n102);
not  g121 (n154, n71);
not  g122 (n198, n78);
not  g123 (n197, n52);
buf  g124 (n207, n35);
buf  g125 (n187, n98);
not  g126 (n208, n27);
not  g127 (n232, n110);
buf  g128 (n171, n95);
buf  g129 (n156, n65);
buf  g130 (n180, n110);
or   g131 (n199, n106, n44, n55, n104);
xnor g132 (n140, n55, n112, n73, n58);
xnor g133 (n196, n49, n65, n48, n101);
nor  g134 (n185, n75, n26, n51, n35);
nand g135 (n163, n102, n29, n68, n112);
xor  g136 (n220, n124, n31, n105, n26);
nand g137 (n191, n112, n123, n43, n77);
and  g138 (n178, n28, n44, n23, n30);
xor  g139 (n134, n24, n127, n125, n37);
nand g140 (n202, n109, n60, n47, n23);
xnor g141 (n155, n76, n76, n77, n67);
xor  g142 (n192, n70, n25, n127, n113);
or   g143 (n217, n71, n55, n82, n34);
xor  g144 (n144, n127, n104, n114, n58);
xnor g145 (n138, n78, n96, n54, n125);
or   g146 (n132, n117, n67, n124, n40);
nand g147 (n149, n99, n25, n83);
and  g148 (n219, n70, n24, n64, n48);
and  g149 (n131, n53, n64, n69, n74);
xnor g150 (n128, n80, n117, n125, n43);
xnor g151 (n137, n61, n33, n120);
nor  g152 (n135, n81, n26, n82, n54);
nor  g153 (n136, n79, n41, n53, n40);
or   g154 (n143, n124, n59, n73, n118);
and  g155 (n151, n27, n80, n42, n108);
xnor g156 (n215, n68, n100, n114, n127);
nand g157 (n160, n100, n23, n105, n63);
xnor g158 (n186, n103, n119, n60, n47);
xor  g159 (n150, n111, n120, n55, n77);
nand g160 (n175, n63, n116, n112, n102);
and  g161 (n233, n111, n107, n41, n35);
xor  g162 (n234, n126, n99, n71, n116);
and  g163 (n209, n125, n97, n22, n113);
or   g164 (n169, n38, n47, n30, n41);
or   g165 (n146, n66, n38, n123, n97);
xor  g166 (n173, n78, n44, n39);
nand g167 (n157, n32, n97, n64, n109);
and  g168 (n226, n29, n84, n60, n59);
xnor g169 (n158, n107, n43, n74, n23);
nor  g170 (n165, n119, n52, n35, n45);
xnor g171 (n188, n46, n115, n28, n39);
nand g172 (n223, n107, n61, n57, n48);
nand g173 (n201, n70, n36, n68, n49);
or   g174 (n182, n69, n51, n59, n49);
xnor g175 (n212, n117, n107, n100, n115);
and  g176 (n166, n28, n50, n27, n126);
xnor g177 (n214, n73, n126, n75, n62);
nor  g178 (n205, n42, n103, n110, n67);
xnor g179 (n237, n106, n29, n122, n22);
xor  g180 (n239, n109, n28, n81, n53);
nand g181 (n170, n45, n56, n31, n58);
nand g182 (n204, n33, n75, n98, n30);
nand g183 (n235, n56, n108, n73, n103);
nor  g184 (n142, n34, n36, n62, n123);
xor  g185 (n229, n66, n22, n76, n84);
and  g186 (n153, n121, n104, n62, n50);
nand g187 (n190, n114, n111, n51, n124);
xnor g188 (n224, n63, n72, n114, n61);
xnor g189 (n216, n34, n50, n98, n71);
nor  g190 (n228, n81, n123, n116, n41);
xnor g191 (n172, n106, n57, n96);
nor  g192 (n168, n104, n24, n63, n119);
nand g193 (n181, n109, n120, n64, n69);
or   g194 (n145, n60, n46, n36, n32);
xor  g195 (n194, n54, n122, n53, n38);
nor  g196 (n222, n82, n25, n80, n97);
nand g197 (n174, n101, n31, n81, n74);
and  g198 (n236, n49, n78, n32, n121);
xnor g199 (n164, n67, n72, n29, n34);
xnor g200 (n129, n117, n61, n65, n100);
nand g201 (n193, n31, n65, n69, n108);
xnor g202 (n130, n121, n39, n118, n76);
and  g203 (n184, n37, n30, n103, n96);
nand g204 (n195, n51, n33, n46, n82);
and  g205 (n203, n26, n70, n83, n98);
and  g206 (n147, n119, n66, n106, n110);
or   g207 (n148, n42, n95, n52, n79);
xnor g208 (n221, n79, n68, n45, n56);
xor  g209 (n238, n77, n84, n43, n48);
nand g210 (n225, n121, n102, n59, n79);
or   g211 (n213, n95, n122, n52, n42);
or   g212 (n162, n95, n101, n39, n83);
nor  g213 (n230, n57, n122, n96, n99);
nor  g214 (n210, n105, n32, n40, n111);
and  g215 (n183, n72, n33, n54, n38);
and  g216 (n218, n37, n113, n72, n56);
or   g217 (n227, n101, n108, n24, n126);
xnor g218 (n133, n50, n115, n45, n66);
and  g219 (n206, n113, n22, n62, n36);
nor  g220 (n139, n80, n37, n46, n40);
buf  g221 (n246, n157);
not  g222 (n337, n129);
not  g223 (n358, n141);
buf  g224 (n307, n155);
not  g225 (n375, n160);
buf  g226 (n352, n131);
buf  g227 (n269, n144);
not  g228 (n363, n149);
buf  g229 (n353, n158);
not  g230 (n284, n138);
buf  g231 (n289, n129);
buf  g232 (n345, n161);
buf  g233 (n347, n145);
buf  g234 (n311, n149);
buf  g235 (n243, n161);
not  g236 (n362, n136);
not  g237 (n250, n133);
not  g238 (n249, n154);
buf  g239 (n364, n147);
not  g240 (n294, n143);
buf  g241 (n281, n136);
not  g242 (n374, n149);
buf  g243 (n290, n152);
buf  g244 (n321, n129);
not  g245 (n349, n143);
buf  g246 (n320, n141);
not  g247 (n252, n137);
not  g248 (n371, n129);
buf  g249 (n368, n155);
not  g250 (n326, n131);
not  g251 (n355, n146);
not  g252 (n357, n136);
not  g253 (n324, n133);
not  g254 (n322, n144);
not  g255 (n298, n138);
not  g256 (n262, n132);
not  g257 (n265, n150);
not  g258 (n266, n139);
not  g259 (n293, n161);
buf  g260 (n275, n136);
not  g261 (n256, n133);
buf  g262 (n301, n134);
buf  g263 (n297, n145);
not  g264 (n258, n131);
not  g265 (n341, n140);
not  g266 (n268, n148);
not  g267 (n264, n132);
buf  g268 (n306, n160);
buf  g269 (n338, n128);
not  g270 (n248, n130);
buf  g271 (n343, n149);
buf  g272 (n318, n158);
not  g273 (n285, n156);
not  g274 (n312, n150);
buf  g275 (n277, n158);
not  g276 (n270, n153);
not  g277 (n330, n135);
not  g278 (n276, n140);
not  g279 (n305, n142);
buf  g280 (n251, n135);
buf  g281 (n327, n130);
buf  g282 (n302, n131);
not  g283 (n244, n160);
not  g284 (n370, n138);
not  g285 (n314, n147);
buf  g286 (n280, n143);
buf  g287 (n309, n155);
buf  g288 (n273, n132);
not  g289 (n241, n157);
not  g290 (n274, n128);
buf  g291 (n295, n145);
buf  g292 (n304, n134);
not  g293 (n257, n138);
buf  g294 (n272, n143);
not  g295 (n339, n137);
buf  g296 (n360, n151);
buf  g297 (n291, n139);
buf  g298 (n325, n148);
not  g299 (n348, n161);
not  g300 (n310, n133);
not  g301 (n365, n157);
not  g302 (n340, n151);
not  g303 (n282, n142);
buf  g304 (n369, n148);
buf  g305 (n240, n159);
not  g306 (n287, n156);
not  g307 (n346, n159);
buf  g308 (n245, n155);
buf  g309 (n335, n147);
buf  g310 (n263, n154);
buf  g311 (n260, n148);
buf  g312 (n328, n153);
buf  g313 (n247, n137);
not  g314 (n334, n145);
not  g315 (n373, n156);
buf  g316 (n313, n159);
buf  g317 (n342, n137);
buf  g318 (n372, n152);
buf  g319 (n242, n128);
buf  g320 (n292, n153);
not  g321 (n332, n151);
not  g322 (n333, n139);
not  g323 (n288, n142);
buf  g324 (n303, n132);
not  g325 (n329, n152);
buf  g326 (n255, n150);
not  g327 (n359, n158);
buf  g328 (n279, n147);
buf  g329 (n336, n146);
buf  g330 (n308, n135);
not  g331 (n319, n144);
buf  g332 (n300, n150);
buf  g333 (n283, n146);
not  g334 (n315, n152);
not  g335 (n350, n141);
buf  g336 (n317, n141);
not  g337 (n261, n128);
not  g338 (n271, n130);
not  g339 (n278, n134);
buf  g340 (n254, n153);
not  g341 (n286, n144);
buf  g342 (n316, n134);
buf  g343 (n361, n146);
buf  g344 (n366, n162);
not  g345 (n323, n151);
buf  g346 (n296, n159);
buf  g347 (n376, n135);
not  g348 (n344, n142);
not  g349 (n259, n154);
buf  g350 (n367, n157);
buf  g351 (n299, n160);
not  g352 (n351, n130);
buf  g353 (n267, n156);
buf  g354 (n354, n139);
not  g355 (n356, n140);
not  g356 (n253, n154);
not  g357 (n331, n140);
buf  g358 (n446, n261);
buf  g359 (n384, n268);
buf  g360 (n442, n263);
buf  g361 (n461, n250);
buf  g362 (n452, n242);
buf  g363 (n393, n259);
not  g364 (n437, n255);
buf  g365 (n385, n265);
not  g366 (n455, n258);
not  g367 (n394, n265);
buf  g368 (n457, n254);
not  g369 (n443, n266);
buf  g370 (n408, n246);
buf  g371 (n448, n240);
not  g372 (n418, n270);
buf  g373 (n392, n246);
buf  g374 (n423, n240);
not  g375 (n397, n243);
not  g376 (n399, n261);
not  g377 (n378, n245);
not  g378 (n404, n258);
not  g379 (n435, n244);
buf  g380 (n438, n243);
not  g381 (n432, n248);
buf  g382 (n422, n250);
buf  g383 (n451, n268);
not  g384 (n424, n262);
not  g385 (n453, n249);
not  g386 (n421, n241);
not  g387 (n425, n267);
buf  g388 (n462, n256);
not  g389 (n416, n258);
buf  g390 (n403, n269);
not  g391 (n396, n247);
not  g392 (n454, n241);
buf  g393 (n409, n265);
not  g394 (n464, n270);
buf  g395 (n439, n248);
not  g396 (n381, n249);
buf  g397 (n405, n252);
buf  g398 (n413, n267);
buf  g399 (n429, n254);
buf  g400 (n406, n262);
buf  g401 (n456, n252);
buf  g402 (n386, n240);
buf  g403 (n388, n267);
buf  g404 (n440, n257);
buf  g405 (n415, n264);
buf  g406 (n380, n266);
not  g407 (n402, n253);
not  g408 (n427, n260);
buf  g409 (n463, n252);
not  g410 (n410, n245);
buf  g411 (n426, n266);
buf  g412 (n407, n262);
not  g413 (n377, n247);
buf  g414 (n445, n263);
buf  g415 (n434, n247);
buf  g416 (n460, n256);
buf  g417 (n458, n254);
buf  g418 (n428, n259);
buf  g419 (n398, n241);
buf  g420 (n401, n244);
not  g421 (n387, n269);
not  g422 (n389, n248);
buf  g423 (n395, n259);
buf  g424 (n436, n264);
buf  g425 (n390, n255);
not  g426 (n459, n256);
not  g427 (n433, n248);
not  g428 (n420, n251);
nor  g429 (n450, n246, n255, n264);
and  g430 (n382, n267, n249, n268);
nand g431 (n444, n252, n243, n264);
nand g432 (n430, n259, n253, n250);
or   g433 (n411, n241, n257, n260);
nand g434 (n391, n244, n245, n242);
xor  g435 (n431, n245, n247, n251);
and  g436 (n412, n253, n265, n240);
nor  g437 (n417, n255, n263);
xor  g438 (n383, n269, n242, n257);
xor  g439 (n379, n261, n254, n268);
xnor g440 (n447, n257, n260, n256);
or   g441 (n441, n253, n258, n269);
nor  g442 (n419, n262, n246, n251);
xnor g443 (n449, n250, n243, n244);
and  g444 (n400, n266, n251, n242);
xor  g445 (n414, n260, n261, n249);
or   g446 (n542, n336, n308, n189, n354);
nand g447 (n642, n224, n236, n379, n327);
xnor g448 (n469, n236, n226, n394, n277);
xor  g449 (n567, n317, n357, n194, n208);
xor  g450 (n489, n421, n392, n337, n377);
xnor g451 (n557, n357, n170, n272, n215);
nand g452 (n509, n314, n174, n425, n329);
nand g453 (n643, n346, n184, n230, n316);
nand g454 (n688, n415, n408, n289, n216);
or   g455 (n481, n388, n335, n297, n165);
xnor g456 (n528, n168, n316, n300, n320);
nor  g457 (n609, n351, n359, n350, n355);
nor  g458 (n552, n339, n214, n279, n381);
xnor g459 (n654, n166, n339, n411, n221);
or   g460 (n627, n325, n333, n430, n212);
nor  g461 (n564, n227, n185, n204, n272);
nand g462 (n539, n286, n426, n208, n226);
nand g463 (n524, n400, n384, n186, n222);
xnor g464 (n687, n417, n224, n351, n282);
nand g465 (n623, n199, n227, n318, n234);
xnor g466 (n593, n223, n344, n292, n393);
nor  g467 (n631, n297, n197, n358, n273);
or   g468 (n537, n389, n168, n314, n291);
xor  g469 (n558, n275, n188, n186, n343);
nand g470 (n590, n396, n237, n239, n290);
nand g471 (n625, n316, n281, n314, n392);
nand g472 (n570, n229, n204, n396, n214);
xor  g473 (n522, n410, n322, n432, n386);
xnor g474 (n484, n325, n429, n163, n201);
and  g475 (n531, n382, n170, n389, n176);
xnor g476 (n660, n342, n308, n205, n200);
xor  g477 (n587, n288, n434, n225, n421);
xor  g478 (n487, n304, n353, n208, n164);
nand g479 (n685, n357, n298, n353, n338);
nand g480 (n619, n342, n277, n238, n357);
nor  g481 (n596, n227, n304, n403, n382);
xor  g482 (n626, n409, n191, n199, n331);
nor  g483 (n634, n272, n431, n332, n172);
xor  g484 (n667, n188, n200, n404, n385);
xor  g485 (n540, n391, n175, n405, n340);
nor  g486 (n572, n192, n222, n315, n167);
and  g487 (n646, n289, n428, n202, n413);
or   g488 (n617, n430, n429, n341, n291);
or   g489 (n628, n312, n318, n285, n383);
and  g490 (n613, n166, n211, n293, n184);
nor  g491 (n630, n185, n209, n236, n302);
and  g492 (n553, n306, n358, n384, n293);
nand g493 (n541, n406, n224, n302, n327);
or   g494 (n482, n349, n281, n394, n233);
and  g495 (n573, n210, n392, n204, n213);
nor  g496 (n675, n185, n414, n163, n395);
or   g497 (n536, n208, n307, n420, n182);
xor  g498 (n504, n383, n311, n402, n182);
xnor g499 (n598, n273, n403, n360, n387);
or   g500 (n559, n190, n333, n359, n173);
and  g501 (n600, n180, n425, n202, n383);
and  g502 (n467, n317, n203, n396, n281);
or   g503 (n649, n310, n239, n344, n417);
xnor g504 (n525, n414, n348, n275, n169);
xnor g505 (n495, n399, n318, n347, n163);
nand g506 (n673, n228, n355, n299, n182);
nand g507 (n647, n162, n187, n212, n234);
or   g508 (n681, n233, n184, n311, n282);
nand g509 (n611, n298, n310, n425, n324);
xnor g510 (n616, n204, n425, n343, n356);
nand g511 (n580, n218, n320, n391, n378);
and  g512 (n563, n287, n228, n419, n309);
nand g513 (n575, n222, n359, n418, n181);
xor  g514 (n493, n199, n198, n335, n429);
and  g515 (n608, n317, n238, n380, n207);
nand g516 (n682, n275, n183, n338, n353);
xor  g517 (n658, n290, n401, n405, n188);
nor  g518 (n465, n312, n322, n354, n344);
or   g519 (n674, n308, n428, n322, n271);
nand g520 (n543, n380, n203, n287, n329);
or   g521 (n678, n300, n168, n177, n171);
nand g522 (n471, n411, n221, n206, n340);
nor  g523 (n591, n324, n397, n342, n304);
or   g524 (n534, n310, n225, n323, n341);
xnor g525 (n621, n349, n420, n336, n286);
xor  g526 (n526, n223, n330, n198, n232);
nor  g527 (n604, n190, n210, n298, n213);
xnor g528 (n529, n420, n341, n352, n306);
xnor g529 (n523, n309, n278, n412, n307);
nor  g530 (n592, n276, n187, n334, n423);
nor  g531 (n684, n421, n164, n170);
and  g532 (n514, n393, n213, n307, n350);
nor  g533 (n614, n207, n334, n223, n205);
xor  g534 (n690, n427, n274, n413, n193);
nor  g535 (n606, n99, n232, n192, n405);
and  g536 (n648, n313, n393, n282, n324);
xor  g537 (n547, n326, n287, n191, n336);
nor  g538 (n497, n231, n193, n416, n378);
and  g539 (n629, n332, n297, n306, n319);
xor  g540 (n501, n276, n239, n401, n398);
nor  g541 (n510, n180, n323, n354, n310);
xnor g542 (n480, n352, n432, n210, n195);
xnor g543 (n565, n289, n206, n330, n216);
nor  g544 (n490, n216, n196, n340, n418);
xor  g545 (n500, n402, n332, n235, n207);
xnor g546 (n597, n417, n209, n278, n317);
xor  g547 (n546, n180, n235, n217, n214);
and  g548 (n637, n406, n326, n166, n296);
nand g549 (n521, n389, n283, n286, n165);
nand g550 (n498, n189, n200, n419, n163);
xor  g551 (n530, n423, n329, n395, n165);
xor  g552 (n569, n311, n390, n190, n347);
nor  g553 (n636, n189, n220, n170, n400);
nor  g554 (n533, n400, n288, n352, n272);
nor  g555 (n585, n176, n313, n193, n344);
or   g556 (n689, n179, n406, n412, n388);
xnor g557 (n620, n284, n390, n166, n231);
nand g558 (n670, n291, n385, n172, n323);
nor  g559 (n635, n321, n326, n388, n381);
nor  g560 (n491, n236, n290, n403, n422);
nand g561 (n571, n238, n399, n403, n379);
nand g562 (n655, n189, n271, n402, n315);
or   g563 (n601, n313, n378, n179, n296);
xor  g564 (n668, n279, n237, n345, n233);
nand g565 (n665, n321, n201, n355, n346);
xor  g566 (n473, n426, n424, n407, n387);
xor  g567 (n494, n394, n318, n315, n220);
nor  g568 (n653, n321, n225, n337, n424);
xnor g569 (n582, n308, n192, n348, n198);
nand g570 (n513, n176, n191, n424, n219);
and  g571 (n633, n235, n329, n383, n178);
xor  g572 (n479, n346, n336, n312, n184);
nand g573 (n505, n432, n276, n193, n309);
nand g574 (n468, n433, n178, n177, n323);
or   g575 (n663, n178, n195, n238, n327);
xnor g576 (n548, n292, n207, n217, n328);
or   g577 (n566, n274, n221, n179, n168);
xor  g578 (n612, n194, n288, n295, n211);
xnor g579 (n512, n386, n197, n319, n295);
and  g580 (n589, n293, n350, n186, n379);
and  g581 (n661, n380, n359, n379, n278);
nand g582 (n476, n381, n342, n180, n284);
xor  g583 (n652, n224, n401, n225, n274);
nor  g584 (n574, n286, n283, n300, n285);
nor  g585 (n595, n392, n305, n393, n416);
or   g586 (n518, n290, n418, n414, n353);
xnor g587 (n581, n433, n182, n202, n420);
nor  g588 (n560, n406, n228, n347, n230);
or   g589 (n657, n430, n203, n354, n271);
xor  g590 (n578, n215, n391, n292, n299);
or   g591 (n610, n330, n325, n226, n232);
xnor g592 (n666, n305, n309, n231, n348);
and  g593 (n492, n418, n312, n305, n206);
nand g594 (n586, n320, n284, n194, n186);
or   g595 (n641, n294, n332, n358, n423);
or   g596 (n650, n178, n228, n300, n273);
and  g597 (n651, n405, n408, n179, n426);
xnor g598 (n466, n320, n174, n293, n408);
nand g599 (n615, n409, n162, n345, n183);
nand g600 (n680, n196, n190, n294, n219);
nand g601 (n577, n430, n339, n417, n324);
nor  g602 (n503, n296, n280, n215, n195);
xnor g603 (n584, n382, n167, n299, n235);
xnor g604 (n677, n206, n281, n292, n274);
nand g605 (n475, n303, n209, n350, n386);
nand g606 (n638, n434, n212, n171, n314);
and  g607 (n671, n413, n412, n304, n278);
nand g608 (n519, n402, n289, n331, n398);
xnor g609 (n474, n355, n404, n380, n352);
xnor g610 (n632, n426, n328, n382);
xnor g611 (n602, n415, n279, n346, n422);
nor  g612 (n664, n325, n410, n303, n424);
and  g613 (n561, n183, n360, n234, n221);
xnor g614 (n576, n321, n196, n218, n408);
or   g615 (n645, n285, n422, n377, n229);
xnor g616 (n483, n284, n315, n335, n427);
or   g617 (n550, n165, n328, n331, n387);
nand g618 (n605, n388, n301, n385, n294);
nor  g619 (n588, n407, n194, n211, n427);
nand g620 (n508, n347, n399, n171, n427);
xor  g621 (n535, n297, n432, n326, n303);
nand g622 (n662, n219, n229, n316, n285);
nand g623 (n520, n230, n410, n412, n419);
xor  g624 (n618, n164, n415, n395, n397);
xnor g625 (n470, n171, n233, n205, n271);
and  g626 (n672, n230, n288, n345, n386);
xor  g627 (n640, n387, n302, n413, n217);
nand g628 (n599, n377, n348, n337, n237);
xnor g629 (n568, n174, n280, n192, n167);
nand g630 (n659, n301, n343, n183, n433);
xnor g631 (n624, n185, n431, n296, n381);
xnor g632 (n507, n349, n188, n398, n227);
and  g633 (n579, n279, n360, n401, n385);
or   g634 (n607, n339, n407, n411, n181);
or   g635 (n478, n396, n217, n270, n333);
nor  g636 (n488, n231, n187, n428, n273);
nor  g637 (n472, n283, n390, n276, n404);
nor  g638 (n556, n187, n197, n356, n404);
nand g639 (n679, n301, n220, n169, n195);
nor  g640 (n622, n175, n212, n334, n338);
nor  g641 (n551, n275, n173, n169, n177);
or   g642 (n562, n433, n303, n202, n341);
nor  g643 (n477, n216, n291, n429, n351);
xnor g644 (n644, n334, n411, n211, n311);
nand g645 (n486, n295, n306, n349, n287);
xor  g646 (n669, n356, n226, n399, n277);
or   g647 (n603, n360, n331, n218, n395);
xor  g648 (n502, n421, n215, n280, n330);
xor  g649 (n544, n191, n394, n422, n181);
nor  g650 (n683, n337, n400, n172, n298);
xor  g651 (n515, n301, n201, n319, n200);
nand g652 (n516, n397, n181, n327, n205);
xor  g653 (n511, n203, n283, n169, n210);
and  g654 (n545, n229, n409, n431, n173);
xnor g655 (n499, n397, n197, n282, n294);
nand g656 (n517, n333, n222, n213, n305);
and  g657 (n554, n270, n407, n377, n162);
and  g658 (n594, n234, n398, n338, n174);
and  g659 (n506, n358, n280, n345, n219);
and  g660 (n639, n415, n409, n201, n299);
xor  g661 (n656, n237, n198, n414, n175);
and  g662 (n583, n340, n319, n419, n199);
nor  g663 (n549, n172, n173, n378, n177);
nand g664 (n555, n223, n416, n356, n196);
xnor g665 (n485, n307, n416, n391, n390);
nand g666 (n538, n313, n209, n277, n175);
xor  g667 (n686, n214, n232, n384, n343);
xnor g668 (n496, n167, n239, n218, n410);
xor  g669 (n532, n322, n423, n351, n431);
or   g670 (n527, n302, n176, n384, n428);
or   g671 (n676, n389, n335, n295, n220);
xor  g672 (n702, n480, n476, n465, n473);
or   g673 (n703, n466, n478, n470, n476);
nor  g674 (n699, n465, n471, n478, n466);
nand g675 (n706, n483, n481, n472);
xnor g676 (n698, n475, n468, n467, n472);
nor  g677 (n710, n471, n483, n477, n475);
nor  g678 (n691, n468, n481, n480, n483);
xnor g679 (n694, n467, n477, n468, n475);
xor  g680 (n692, n477, n465, n481, n484);
xor  g681 (n700, n470, n465, n473, n471);
nand g682 (n695, n469, n478, n482, n481);
and  g683 (n696, n469, n484, n474, n466);
nor  g684 (n693, n474, n469, n476);
nand g685 (n701, n483, n475, n467, n480);
nor  g686 (n705, n477, n470, n472, n479);
xor  g687 (n709, n471, n479, n478, n480);
or   g688 (n697, n473, n482, n476);
xnor g689 (n707, n474, n474, n467, n470);
nand g690 (n708, n484, n484, n482, n466);
nor  g691 (n704, n473, n479, n468);
and  g692 (n723, n366, n361, n369, n364);
and  g693 (n725, n369, n692, n485, n375);
nand g694 (n722, n374, n364, n361);
xnor g695 (n712, n696, n363, n374, n371);
nand g696 (n715, n367, n693, n486, n361);
xnor g697 (n726, n372, n693, n485);
xor  g698 (n732, n370, n696, n693, n375);
nand g699 (n719, n695, n368, n376, n367);
xnor g700 (n713, n371, n692, n696, n365);
xnor g701 (n717, n694, n365, n373, n366);
xnor g702 (n720, n362, n372, n367, n376);
and  g703 (n733, n368, n363, n370, n376);
nor  g704 (n718, n366, n694, n697, n373);
nor  g705 (n727, n375, n486, n372, n363);
nor  g706 (n714, n691, n374, n370, n695);
or   g707 (n716, n692, n691, n372, n371);
xnor g708 (n721, n368, n486, n371, n374);
nor  g709 (n711, n376, n487, n365);
xor  g710 (n729, n362, n693, n364);
nor  g711 (n734, n695, n373, n486, n362);
and  g712 (n728, n365, n487, n695, n369);
or   g713 (n735, n694, n696, n366, n375);
xnor g714 (n731, n692, n691, n373, n485);
xnor g715 (n724, n370, n691, n368, n694);
xnor g716 (n730, n369, n362, n367, n363);
and  g717 (n773, n719, n716, n514, n500);
xnor g718 (n780, n495, n500, n522, n516);
nand g719 (n756, n491, n497, n509, n714);
or   g720 (n779, n717, n513, n489, n509);
xor  g721 (n757, n501, n519, n506, n513);
xnor g722 (n777, n721, n495, n489, n503);
xnor g723 (n741, n510, n520, n488, n502);
xor  g724 (n750, n499, n508, n714, n489);
and  g725 (n739, n515, n501, n505, n711);
nor  g726 (n782, n504, n720, n515, n505);
xnor g727 (n744, n492, n513, n500, n503);
nor  g728 (n760, n499, n721, n720, n522);
and  g729 (n765, n507, n722, n504);
nor  g730 (n749, n713, n723, n506, n517);
or   g731 (n736, n725, n511, n488, n502);
or   g732 (n775, n488, n726, n522, n498);
nand g733 (n762, n522, n492, n712, n505);
nor  g734 (n737, n503, n724, n498, n490);
nor  g735 (n763, n512, n498, n494, n721);
nor  g736 (n770, n727, n492, n520, n496);
xnor g737 (n745, n497, n495, n502, n722);
nand g738 (n742, n491, n493, n725);
or   g739 (n766, n500, n521, n519, n508);
xor  g740 (n776, n519, n520, n509, n726);
xor  g741 (n771, n512, n493, n494, n722);
and  g742 (n740, n510, n512, n490, n511);
xnor g743 (n767, n499, n504, n514, n496);
nand g744 (n769, n493, n495, n498, n724);
and  g745 (n738, n521, n511, n488, n724);
or   g746 (n743, n507, n516, n514, n521);
and  g747 (n755, n723, n720, n511, n715);
xor  g748 (n747, n499, n497, n513, n518);
or   g749 (n781, n718, n517, n491);
nand g750 (n759, n507, n508, n518, n494);
xor  g751 (n772, n518, n506, n515, n722);
or   g752 (n752, n719, n726, n509);
or   g753 (n751, n487, n501, n508, n724);
nor  g754 (n746, n510, n490, n512, n723);
nand g755 (n778, n721, n503, n502, n490);
xnor g756 (n761, n716, n496, n711);
nor  g757 (n758, n517, n507, n489, n519);
or   g758 (n753, n516, n514, n718, n520);
or   g759 (n748, n725, n715, n497, n720);
xnor g760 (n768, n723, n506, n505, n712);
nand g761 (n764, n510, n493, n501, n521);
or   g762 (n774, n492, n518, n517, n516);
and  g763 (n754, n713, n494, n515, n717);
nand g764 (n879, n624, n610, n768, n588);
xor  g765 (n870, n645, n649, n596, n619);
or   g766 (n810, n537, n615, n648, n624);
xor  g767 (n951, n546, n563, n640, n611);
nand g768 (n872, n655, n609, n628, n617);
nor  g769 (n922, n765, n588, n780, n630);
or   g770 (n787, n779, n556, n615, n755);
and  g771 (n900, n747, n575, n533, n618);
xnor g772 (n793, n638, n563, n762);
xnor g773 (n871, n661, n572, n583, n575);
xnor g774 (n893, n757, n641, n549, n555);
nor  g775 (n876, n609, n631, n540, n613);
xor  g776 (n851, n545, n558, n564, n536);
nand g777 (n947, n765, n571, n640, n542);
xnor g778 (n929, n641, n749, n756, n598);
xnor g779 (n895, n574, n581, n662, n750);
and  g780 (n819, n601, n565, n639, n659);
xnor g781 (n902, n738, n588, n638, n523);
and  g782 (n839, n566, n553, n530, n548);
nor  g783 (n822, n771, n752, n552, n741);
nor  g784 (n959, n616, n632, n603, n531);
nor  g785 (n835, n524, n629, n649, n654);
and  g786 (n956, n549, n623, n777, n575);
xnor g787 (n901, n582, n621, n620, n647);
or   g788 (n830, n741, n584, n638, n590);
xnor g789 (n783, n540, n768, n614, n596);
xnor g790 (n904, n616, n594, n596, n611);
xnor g791 (n909, n523, n537, n646, n544);
or   g792 (n933, n577, n541, n639, n761);
nand g793 (n911, n629, n615, n549, n761);
xnor g794 (n815, n740, n530, n591, n754);
xnor g795 (n866, n598, n740, n534, n567);
xor  g796 (n837, n586, n630, n538, n595);
xnor g797 (n965, n586, n559, n632, n556);
and  g798 (n784, n561, n642, n776, n746);
or   g799 (n955, n543, n555, n532, n582);
xor  g800 (n948, n573, n579, n534, n635);
nand g801 (n898, n552, n663, n736, n644);
xnor g802 (n953, n593, n539, n764, n773);
nor  g803 (n915, n632, n525, n755, n557);
xnor g804 (n889, n538, n524, n566, n600);
nand g805 (n926, n766, n621, n769, n657);
xnor g806 (n944, n658, n539, n776, n549);
or   g807 (n791, n773, n567, n607, n608);
xnor g808 (n849, n535, n624, n637, n561);
nor  g809 (n875, n562, n639, n640, n750);
xnor g810 (n908, n585, n561, n752, n606);
nand g811 (n836, n643, n626, n736, n655);
and  g812 (n840, n628, n782, n560, n654);
nand g813 (n916, n571, n743, n614, n764);
nand g814 (n934, n753, n656, n592, n627);
and  g815 (n824, n615, n636, n599, n564);
nor  g816 (n788, n662, n780, n621, n558);
nand g817 (n921, n606, n526, n602, n560);
xor  g818 (n790, n736, n527, n634, n569);
xor  g819 (n852, n748, n646, n554, n607);
or   g820 (n949, n746, n551, n640, n594);
xnor g821 (n785, n583, n618, n645, n749);
nand g822 (n925, n539, n743, n629, n537);
nor  g823 (n885, n597, n579, n562, n626);
nor  g824 (n930, n751, n659, n553, n650);
and  g825 (n857, n565, n609, n639, n655);
or   g826 (n968, n662, n595, n546, n627);
and  g827 (n843, n651, n601, n576, n774);
xnor g828 (n935, n557, n607, n587, n622);
xnor g829 (n932, n766, n552, n594, n749);
and  g830 (n903, n748, n568, n741, n648);
or   g831 (n863, n573, n598, n551, n541);
nor  g832 (n821, n572, n573, n570, n557);
nand g833 (n906, n760, n602, n569, n641);
xor  g834 (n842, n605, n660, n770, n769);
xor  g835 (n806, n602, n772, n545, n635);
nand g836 (n865, n650, n642, n762, n629);
nor  g837 (n844, n611, n652, n531, n622);
and  g838 (n816, n599, n753, n552, n532);
xor  g839 (n800, n547, n581, n622, n578);
or   g840 (n847, n600, n660, n776, n636);
nor  g841 (n808, n570, n581, n573, n770);
nor  g842 (n864, n737, n662, n525, n781);
nor  g843 (n884, n567, n527, n547, n744);
xnor g844 (n805, n580, n648, n529, n528);
and  g845 (n940, n646, n758, n579, n769);
and  g846 (n854, n544, n747, n595, n560);
nand g847 (n950, n653, n659, n569, n533);
nand g848 (n832, n606, n535, n603, n645);
xor  g849 (n818, n602, n566, n622, n753);
and  g850 (n804, n614, n605, n527, n528);
xor  g851 (n964, n551, n543, n540, n771);
nor  g852 (n919, n745, n576, n535, n658);
xnor g853 (n860, n763, n770, n570, n647);
or   g854 (n896, n774, n618, n619, n765);
nand g855 (n946, n756, n764, n657, n563);
xnor g856 (n960, n563, n626, n758, n586);
xor  g857 (n883, n608, n579, n531, n652);
xnor g858 (n823, n632, n564, n538, n631);
or   g859 (n858, n589, n610, n547, n751);
xnor g860 (n942, n641, n778, n775, n644);
and  g861 (n888, n653, n580, n564, n610);
nor  g862 (n937, n757, n637, n562, n760);
xor  g863 (n918, n550, n749, n578, n589);
nand g864 (n877, n587, n743, n583, n623);
nor  g865 (n868, n742, n560, n574, n535);
nor  g866 (n966, n759, n634, n614, n571);
xor  g867 (n862, n630, n595, n751, n766);
and  g868 (n923, n553, n781, n603, n736);
and  g869 (n910, n601, n571, n646, n753);
nor  g870 (n855, n634, n550, n737, n644);
nand g871 (n891, n623, n738, n652, n541);
nand g872 (n945, n765, n771, n558, n763);
nand g873 (n917, n542, n656, n764, n592);
xnor g874 (n789, n545, n661, n591, n559);
xor  g875 (n943, n581, n756, n759, n590);
and  g876 (n803, n577, n648, n778, n575);
or   g877 (n905, n628, n554, n758, n772);
xor  g878 (n848, n637, n636, n537, n529);
or   g879 (n828, n578, n758, n745, n617);
xnor g880 (n856, n544, n528, n577, n601);
and  g881 (n799, n780, n577, n591, n613);
nand g882 (n867, n663, n657, n762, n619);
xnor g883 (n927, n523, n556, n545);
xnor g884 (n845, n584, n604, n567, n754);
xor  g885 (n882, n779, n598, n625, n760);
and  g886 (n920, n767, n550, n555, n526);
nor  g887 (n786, n782, n559, n739);
or   g888 (n859, n546, n747, n612, n763);
nor  g889 (n961, n580, n660, n599, n659);
nand g890 (n801, n626, n744, n530, n778);
nor  g891 (n807, n746, n608, n760, n603);
nand g892 (n846, n527, n652, n772, n647);
xor  g893 (n826, n561, n613, n534, n661);
nor  g894 (n924, n658, n585, n554, n526);
xor  g895 (n931, n613, n634, n637, n582);
or   g896 (n825, n554, n633, n747, n625);
nand g897 (n820, n533, n755, n781, n773);
nor  g898 (n907, n532, n742, n776, n779);
or   g899 (n886, n643, n750, n625, n761);
or   g900 (n794, n775, n584, n620, n600);
and  g901 (n938, n770, n597, n744, n627);
and  g902 (n796, n649, n543, n585, n643);
nor  g903 (n827, n774, n739, n775, n534);
nand g904 (n853, n526, n656, n654, n593);
nor  g905 (n811, n663, n584, n576, n572);
and  g906 (n831, n757, n548, n570, n600);
and  g907 (n969, n568, n609, n645, n745);
xnor g908 (n970, n656, n586, n525, n631);
xor  g909 (n954, n769, n740, n612, n658);
nor  g910 (n814, n620, n550, n752, n737);
or   g911 (n874, n742, n739, n582, n568);
and  g912 (n850, n568, n643, n647, n628);
xor  g913 (n841, n772, n616, n661, n532);
and  g914 (n967, n748, n555, n597, n528);
nand g915 (n899, n642, n590, n546, n636);
xnor g916 (n958, n757, n604, n616, n651);
nand g917 (n802, n635, n529, n539, n638);
and  g918 (n957, n605, n565, n777, n536);
or   g919 (n838, n612, n763, n745, n542);
or   g920 (n878, n737, n593, n771, n583);
or   g921 (n892, n617, n738, n624, n587);
nand g922 (n797, n653, n608, n774, n580);
xor  g923 (n894, n533, n585, n589, n536);
xnor g924 (n936, n548, n591, n593, n642);
and  g925 (n829, n759, n596, n777, n569);
nand g926 (n880, n777, n768, n754, n599);
and  g927 (n809, n543, n649, n750, n606);
xor  g928 (n812, n743, n633, n755, n562);
nor  g929 (n890, n592, n524, n779, n612);
or   g930 (n817, n541, n620, n651, n588);
nor  g931 (n928, n572, n557, n551, n536);
or   g932 (n798, n751, n523, n592, n529);
xnor g933 (n873, n566, n631, n740, n663);
nor  g934 (n914, n633, n650, n782);
xor  g935 (n913, n767, n635, n544, n590);
xor  g936 (n941, n578, n619, n542, n767);
xnor g937 (n834, n617, n644, n547, n589);
xnor g938 (n963, n553, n604, n605, n754);
and  g939 (n833, n574, n761, n594, n773);
nor  g940 (n897, n775, n587, n660, n782);
or   g941 (n887, n611, n548, n742, n759);
nor  g942 (n795, n627, n607, n780, n531);
xnor g943 (n869, n538, n768, n778, n748);
nor  g944 (n861, n576, n524, n781, n746);
xor  g945 (n792, n540, n525, n530, n766);
xnor g946 (n813, n655, n739, n657, n654);
and  g947 (n962, n574, n597, n752, n756);
xnor g948 (n912, n625, n604, n738, n744);
or   g949 (n881, n558, n767, n633, n741);
xnor g950 (n952, n651, n565, n623, n653);
nand g951 (n939, n610, n630, n621, n618);
xor  g952 (n977, n881, n856, n847, n829);
nand g953 (n992, n864, n830, n799, n865);
nor  g954 (n983, n909, n861, n853, n825);
xor  g955 (n978, n823, n805, n802, n859);
nand g956 (n993, n868, n880, n863, n785);
nand g957 (n975, n883, n795, n903, n866);
nor  g958 (n994, n820, n907, n867, n812);
nand g959 (n973, n909, n869, n879, n874);
xnor g960 (n989, n909, n857, n875, n819);
xor  g961 (n985, n893, n888, n846, n824);
xor  g962 (n986, n811, n876, n844, n848);
and  g963 (n984, n813, n904, n895);
nand g964 (n1006, n884, n790, n908, n882);
nor  g965 (n997, n862, n860, n850, n902);
xor  g966 (n998, n892, n808, n870, n783);
or   g967 (n995, n800, n877, n818, n843);
nand g968 (n980, n797, n834, n664, n903);
xor  g969 (n1007, n842, n901, n910, n835);
xor  g970 (n1001, n793, n809, n845, n788);
or   g971 (n1004, n796, n902, n854, n898);
nand g972 (n990, n828, n887, n837, n886);
and  g973 (n1005, n794, n807, n907, n872);
and  g974 (n976, n901, n899, n889, n831);
nor  g975 (n999, n901, n900, n852, n896);
and  g976 (n1003, n840, n849, n786, n814);
nand g977 (n1000, n903, n804, n836, n904);
xnor g978 (n987, n902, n839, n841, n908);
xor  g979 (n974, n838, n792, n907, n822);
and  g980 (n972, n851, n906, n817, n905);
xnor g981 (n981, n905, n906, n815);
nand g982 (n991, n803, n833, n789, n891);
xnor g983 (n982, n871, n806, n826, n873);
nand g984 (n1002, n858, n801, n897, n894);
xor  g985 (n988, n827, n821, n908, n885);
or   g986 (n971, n787, n791, n798, n784);
xor  g987 (n979, n664, n878, n810, n816);
xnor g988 (n996, n832, n855, n890, n905);
not  g989 (n1009, n728);
or   g990 (n1010, n975, n728);
nand g991 (n1012, n727, n971, n729, n728);
or   g992 (n1008, n974, n729, n972);
xnor g993 (n1011, n729, n973, n727);
buf  g994 (n1020, n1010);
not  g995 (n1014, n911);
not  g996 (n1021, n912);
buf  g997 (n1018, n1009);
not  g998 (n1013, n911);
not  g999 (n1016, n1008);
buf  g1000 (n1017, n1008);
not  g1001 (n1023, n910);
not  g1002 (n1015, n911);
nand g1003 (n1019, n1009, n1010);
and  g1004 (n1024, n1009, n912, n1010, n910);
xnor g1005 (n1022, n1009, n1008, n912);
buf  g1006 (n1038, n915);
buf  g1007 (n1027, n914);
not  g1008 (n1035, n913);
buf  g1009 (n1031, n916);
buf  g1010 (n1039, n915);
not  g1011 (n1034, n1016);
buf  g1012 (n1033, n1014);
buf  g1013 (n1032, n914);
not  g1014 (n1026, n913);
not  g1015 (n1036, n1016);
buf  g1016 (n1030, n914);
not  g1017 (n1037, n916);
nand g1018 (n1040, n1015, n1013);
xnor g1019 (n1028, n916, n1014);
nor  g1020 (n1029, n915, n1016, n913, n1015);
nand g1021 (n1025, n1015, n1016, n1013);
buf  g1022 (n1044, n1025);
buf  g1023 (n1041, n1025);
not  g1024 (n1043, n1025);
buf  g1025 (n1042, n1025);
or   g1026 (n1052, n1011, n993, n1041, n1042);
nor  g1027 (n1055, n981, n1018, n991, n1041);
nor  g1028 (n1051, n1018, n1012, n1004, n1017);
nand g1029 (n1053, n1044, n1002, n987, n1011);
and  g1030 (n1050, n1006, n978, n999, n1003);
xor  g1031 (n1059, n994, n1043, n979);
or   g1032 (n1054, n998, n1042, n1017, n1044);
nor  g1033 (n1056, n997, n976, n1017);
and  g1034 (n1058, n984, n988, n1001, n1042);
xor  g1035 (n1046, n992, n1043, n1012, n985);
nor  g1036 (n1047, n1042, n1044, n1041, n1005);
or   g1037 (n1045, n982, n977, n980, n1043);
or   g1038 (n1049, n986, n1011, n989, n917);
and  g1039 (n1057, n996, n1007, n995, n983);
nor  g1040 (n1048, n990, n1000, n1011, n1044);
buf  g1041 (n1060, n1018);
or   g1042 (n1061, n1059, n1058);
xnor g1043 (n1065, n1019, n1020, n1060);
and  g1044 (n1063, n1021, n1061, n1060);
and  g1045 (n1064, n1022, n1021, n1024, n1019);
or   g1046 (n1066, n1019, n1022, n1021);
and  g1047 (n1069, n1061, n1021, n1023, n1060);
or   g1048 (n1068, n1024, n1023, n1018);
xnor g1049 (n1067, n1022, n1020, n1023, n1024);
nand g1050 (n1062, n1061, n1019, n1020);
buf  g1051 (n1089, n1068);
buf  g1052 (n1092, n1034);
buf  g1053 (n1099, n1028);
buf  g1054 (n1075, n1062);
buf  g1055 (n1082, n1067);
buf  g1056 (n1097, n1063);
buf  g1057 (n1083, n1028);
not  g1058 (n1084, n1063);
buf  g1059 (n1070, n1030);
not  g1060 (n1098, n1068);
not  g1061 (n1088, n1031);
buf  g1062 (n1078, n1030);
not  g1063 (n1081, n1030);
or   g1064 (n1096, n1069, n1036, n1038);
and  g1065 (n1076, n1067, n1068, n664, n1063);
xnor g1066 (n1072, n1065, n1035, n1027, n1066);
xnor g1067 (n1077, n1036, n1029, n1034, n1035);
nor  g1068 (n1071, n1032, n1065, n1026, n1067);
xnor g1069 (n1094, n1064, n1036, n1037, n1032);
nor  g1070 (n1074, n1029, n1062, n1031);
nand g1071 (n1091, n1064, n1027, n1034, n1035);
or   g1072 (n1093, n664, n1066, n1029, n1034);
and  g1073 (n1095, n1066, n1069, n1032, n1038);
xnor g1074 (n1090, n1033, n1035, n1031, n1068);
nor  g1075 (n1080, n1027, n1026, n1028, n1064);
and  g1076 (n1100, n1066, n1069, n1063, n1032);
or   g1077 (n1101, n1026, n1062, n1038, n1037);
and  g1078 (n1073, n1064, n1039, n1067, n1037);
xor  g1079 (n1079, n1062, n665, n1037, n1065);
and  g1080 (n1087, n1027, n1038, n1036, n1029);
or   g1081 (n1085, n1033, n1065, n1069, n1030);
nor  g1082 (n1086, n1028, n1033, n1026);
not  g1083 (n1107, n1070);
nor  g1084 (n1114, n1075, n1072, n1074);
xor  g1085 (n1113, n1078, n1071, n666);
xnor g1086 (n1105, n1070, n1071, n1073);
xor  g1087 (n1109, n1077, n666, n1073);
xnor g1088 (n1106, n1073, n1074, n1075);
nor  g1089 (n1111, n1073, n1071, n665);
xnor g1090 (n1104, n1076, n666, n1078);
nand g1091 (n1108, n1077, n1076);
nand g1092 (n1112, n1070, n1074, n1076);
xnor g1093 (n1102, n1075, n665, n1071, n1072);
xnor g1094 (n1110, n1072, n665, n1074, n1077);
or   g1095 (n1103, n1075, n1077, n1070, n1072);
or   g1096 (n1123, n1081, n1109, n1106);
xnor g1097 (n1124, n1108, n1108, n1112, n1111);
nand g1098 (n1126, n1107, n1082, n1079, n1102);
xnor g1099 (n1121, n1103, n1105, n1110);
nand g1100 (n1129, n1105, n1104, n1112, n1111);
nor  g1101 (n1125, n1108, n1103, n1106, n1102);
xnor g1102 (n1117, n1079, n1110, n1108);
or   g1103 (n1118, n1106, n1078, n1109, n1102);
nor  g1104 (n1127, n1110, n1111, n666, n1109);
xor  g1105 (n1120, n1102, n1080, n1106);
xor  g1106 (n1115, n1080, n1103, n1079);
xor  g1107 (n1116, n1081, n1109, n1104, n1105);
nand g1108 (n1122, n1081, n1079, n1082, n1104);
nand g1109 (n1128, n1078, n1104, n1111, n1107);
xnor g1110 (n1119, n1080, n1081, n1107);
xnor g1111 (n1136, n1123, n1088);
not  g1112 (n1132, n1084);
nand g1113 (n1135, n1087, n1119);
or   g1114 (n1133, n1083, n1127, n1126);
and  g1115 (n1139, n1084, n1087, n1086);
or   g1116 (n1130, n1087, n1086, n1082, n1085);
nand g1117 (n1137, n1124, n1122, n1128, n1125);
xnor g1118 (n1140, n1083, n1086, n1120);
xor  g1119 (n1138, n1088, n1085, n1121);
nor  g1120 (n1131, n1083, n1129, n1082, n1087);
nor  g1121 (n1134, n1084, n1085, n1083, n1088);
nor  g1122 (n1145, n1097, n1096, n1091, n1133);
and  g1123 (n1149, n1131, n1096, n1098);
and  g1124 (n1154, n1099, n1133, n1089, n1131);
nand g1125 (n1150, n1095, n1095, n1133, n1091);
or   g1126 (n1152, n1094, n1097, n1132, n1089);
xor  g1127 (n1144, n1098, n1092, n1130);
nor  g1128 (n1146, n1095, n1099, n1132, n1092);
xnor g1129 (n1142, n1090, n1133, n1093, n1091);
nand g1130 (n1147, n1132, n1130, n1092, n1089);
nor  g1131 (n1153, n1100, n1130, n1094, n1093);
xor  g1132 (n1143, n1097, n1088, n1095, n1090);
nand g1133 (n1151, n1099, n1096, n1097, n1100);
xnor g1134 (n1141, n1131, n1096, n1098, n1089);
nor  g1135 (n1156, n1134, n1132, n1090);
nor  g1136 (n1148, n1094, n1099, n1091, n1100);
and  g1137 (n1155, n1131, n1094, n1093);
buf  g1138 (n1158, n1144);
buf  g1139 (n1165, n1101);
buf  g1140 (n1166, n1145);
not  g1141 (n1157, n1101);
not  g1142 (n1164, n1141);
buf  g1143 (n1163, n1101);
not  g1144 (n1159, n1143);
not  g1145 (n1167, n1101);
buf  g1146 (n1168, n1112);
nand g1147 (n1161, n1144, n1113, n1112);
nor  g1148 (n1162, n1141, n1144, n1143, n1142);
or   g1149 (n1160, n1100, n1143, n1142);
buf  g1150 (n1171, n1158);
not  g1151 (n1172, n1113);
nand g1152 (n1173, n1113, n1135, n1157);
nor  g1153 (n1169, n1157, n1114, n1134);
and  g1154 (n1170, n1134, n1157, n1113);
xnor g1155 (n1174, n1158, n1134, n1114);
nand g1156 (n1196, n1173, n1151, n1137, n1170);
nor  g1157 (n1184, n1155, n1150, n1154, n1138);
xnor g1158 (n1191, n667, n1149, n1140, n1152);
and  g1159 (n1185, n1138, n1139, n1136, n1149);
nor  g1160 (n1194, n1138, n1169, n1136, n668);
and  g1161 (n1195, n1155, n1137, n1169, n1145);
nor  g1162 (n1190, n1155, n668, n1170, n1150);
and  g1163 (n1178, n1136, n1171, n1156, n1169);
or   g1164 (n1177, n1148, n1153, n667, n1152);
xor  g1165 (n1179, n1154, n1135, n1171, n1139);
nor  g1166 (n1187, n1145, n1169, n1149, n1153);
nor  g1167 (n1192, n1172, n1137, n1152, n1148);
nor  g1168 (n1183, n1147, n1151, n1172);
and  g1169 (n1181, n1173, n668, n1156);
or   g1170 (n1180, n1171, n1138, n1147, n1151);
or   g1171 (n1186, n1136, n1172, n1139, n1173);
xor  g1172 (n1176, n1146, n1146, n1148, n667);
nand g1173 (n1188, n1174, n1135, n917, n1137);
or   g1174 (n1175, n1153, n1170, n1139);
nand g1175 (n1189, n1146, n1173, n1171, n1140);
or   g1176 (n1193, n1147, n1140, n1150, n1156);
nand g1177 (n1182, n1140, n1154, n1174, n667);
not  g1178 (n1199, n1176);
buf  g1179 (n1198, n1175);
not  g1180 (n1200, n1176);
xnor g1181 (n1197, n1176, n1175);
or   g1182 (n1205, n1197, n1163, n1161, n1158);
or   g1183 (n1207, n1165, n1159, n1200, n1198);
xor  g1184 (n1202, n1161, n1174, n1162);
xnor g1185 (n1211, n1159, n1167, n1200, n1197);
nand g1186 (n1216, n1197, n1164, n1161, n1165);
nor  g1187 (n1209, n1161, n1160, n1197, n1166);
or   g1188 (n1208, n1166, n1200, n1177);
and  g1189 (n1204, n1162, n1177, n1166, n1198);
and  g1190 (n1206, n1168, n1177, n1163, n1164);
nor  g1191 (n1212, n1199, n1167, n1160, n1174);
xor  g1192 (n1203, n1160, n1163, n1168, n1176);
nand g1193 (n1215, n1168, n1159, n1167);
nor  g1194 (n1201, n1162, n1160, n1165, n1167);
xor  g1195 (n1210, n1165, n1199, n1164);
and  g1196 (n1214, n1199, n1166, n1198, n1168);
nor  g1197 (n1213, n1199, n1163, n1158, n1198);
or   g1198 (n1219, n1202, n1187, n1201, n1177);
nand g1199 (n1229, n1188, n1182, n1185, n1205);
xor  g1200 (n1220, n1180, n1186, n1185);
and  g1201 (n1225, n1187, n1203, n1181, n1180);
and  g1202 (n1228, n1184, n1183, n1187, n1178);
or   g1203 (n1218, n1202, n1183, n1205, n1179);
nand g1204 (n1231, n1181, n1181, n1201, n1203);
or   g1205 (n1226, n1182, n1184, n1178, n1203);
and  g1206 (n1222, n1179, n1182, n1201, n1178);
xor  g1207 (n1230, n1178, n1186, n1204, n1188);
xor  g1208 (n1217, n1186, n1184, n1182, n1202);
nor  g1209 (n1221, n1185, n1188, n1179, n1184);
and  g1210 (n1227, n1188, n1179, n1204, n1180);
xor  g1211 (n1223, n1205, n1187, n1186, n1181);
and  g1212 (n1224, n1180, n1204, n1183);
nand g1213 (n1236, n1228, n1190, n1191);
nor  g1214 (n1237, n1189, n1190, n1225, n1192);
and  g1215 (n1232, n1193, n1191, n1192, n1229);
and  g1216 (n1233, n1224, n1189, n1192, n1190);
nor  g1217 (n1235, n1189, n1191, n1227, n1226);
and  g1218 (n1234, n1192, n1191, n1190, n1189);
xor  g1219 (n1241, n1233, n1208, n1206, n1207);
and  g1220 (n1238, n1195, n1207, n1194, n1232);
nand g1221 (n1239, n1193, n1194, n1206, n1195);
or   g1222 (n1242, n1206, n1195, n1196);
or   g1223 (n1244, n1196, n1232, n1195, n1194);
xnor g1224 (n1240, n1232, n1194, n1193);
xnor g1225 (n1243, n1207, n1233, n1232);
buf  g1226 (n1252, n1242);
buf  g1227 (n1246, n1238);
not  g1228 (n1251, n1242);
not  g1229 (n1250, n1240);
buf  g1230 (n1254, n1243);
buf  g1231 (n1245, n1208);
buf  g1232 (n1249, n1239);
not  g1233 (n1247, n1243);
buf  g1234 (n1253, n1241);
nand g1235 (n1248, n1244, n1241);
nor  g1236 (n1258, n672, n673, n669, n1213);
nand g1237 (n1265, n1246, n1247, n1210);
xor  g1238 (n1260, n672, n1248, n1208, n1214);
nand g1239 (n1268, n1213, n674, n1211, n1247);
and  g1240 (n1264, n671, n670, n1248, n1209);
xor  g1241 (n1259, n1248, n672, n670);
or   g1242 (n1261, n671, n1214, n1212, n1210);
xor  g1243 (n1256, n1214, n1245, n669, n1248);
nand g1244 (n1266, n671, n1246, n669);
nor  g1245 (n1255, n1210, n1211, n671, n672);
nor  g1246 (n1262, n1246, n673, n1213, n1209);
or   g1247 (n1257, n1216, n1246, n1209, n673);
nand g1248 (n1263, n1216, n1247, n1211, n1245);
or   g1249 (n1267, n1215, n1212, n670, n1245);
or   g1250 (n1269, n1212, n1215, n673);
nand g1251 (n1304, n458, n454, n436, n459);
xnor g1252 (n1288, n462, n455, n1267, n453);
nor  g1253 (n1291, n434, n439, n450, n437);
nand g1254 (n1302, n1234, n456, n1235, n1262);
and  g1255 (n1293, n459, n1266, n458, n457);
xor  g1256 (n1283, n1233, n443, n1266, n439);
and  g1257 (n1308, n442, n461, n1235);
or   g1258 (n1278, n447, n452, n1235, n441);
or   g1259 (n1299, n1268, n438, n1260);
and  g1260 (n1305, n454, n453, n1268, n442);
nand g1261 (n1295, n1262, n1268, n441, n454);
xnor g1262 (n1310, n435, n1236, n455, n460);
xnor g1263 (n1271, n464, n1236, n443, n1262);
xor  g1264 (n1300, n449, n457, n439, n1265);
xor  g1265 (n1297, n435, n444, n437, n451);
nand g1266 (n1275, n437, n453, n1269, n440);
nand g1267 (n1306, n1264, n1260, n1261, n1263);
xor  g1268 (n1276, n1258, n1267, n443, n435);
nor  g1269 (n1307, n1263, n436, n439, n461);
or   g1270 (n1279, n463, n463, n1267, n443);
or   g1271 (n1315, n463, n460, n457, n1266);
nor  g1272 (n1282, n1255, n436, n1265, n1269);
nand g1273 (n1274, n438, n452, n1261, n459);
nor  g1274 (n1285, n456, n458, n441, n445);
or   g1275 (n1284, n438, n450, n462, n445);
xor  g1276 (n1286, n463, n1265, n444, n458);
xor  g1277 (n1311, n450, n453, n1237, n456);
nor  g1278 (n1270, n440, n454, n1268, n445);
and  g1279 (n1280, n440, n451, n460, n1264);
nor  g1280 (n1309, n459, n455, n1237, n436);
and  g1281 (n1296, n447, n1256, n1257, n1237);
and  g1282 (n1314, n448, n462, n434, n1236);
nor  g1283 (n1303, n447, n440, n1259, n441);
nand g1284 (n1292, n449, n446, n1266, n460);
or   g1285 (n1313, n1264, n462, n1257, n1269);
or   g1286 (n1294, n447, n1263, n446, n448);
nor  g1287 (n1281, n1234, n1237, n449, n445);
xnor g1288 (n1312, n1231, n1256, n446, n1265);
xnor g1289 (n1290, n1263, n1267, n435, n455);
nand g1290 (n1277, n452, n451, n449, n444);
xnor g1291 (n1272, n1234, n451, n1264, n1235);
nand g1292 (n1298, n448, n1262, n461, n1259);
xor  g1293 (n1301, n442, n446, n448, n450);
xnor g1294 (n1273, n444, n442, n1269, n437);
xnor g1295 (n1289, n1236, n456, n457, n1255);
nor  g1296 (n1287, n1258, n452, n1230, n1234);
nor  g1297 (n1329, n679, n1250, n682, n1272);
and  g1298 (n1335, n1278, n675, n1270, n1274);
and  g1299 (n1344, n688, n681, n1272, n1251);
xnor g1300 (n1334, n1276, n686, n1275);
nand g1301 (n1353, n1273, n685, n675, n734);
xnor g1302 (n1352, n690, n733, n681, n735);
xnor g1303 (n1319, n684, n677, n1273, n733);
or   g1304 (n1322, n677, n735, n680, n685);
nand g1305 (n1327, n676, n735, n689, n734);
and  g1306 (n1347, n1274, n687, n685, n674);
xnor g1307 (n1351, n732, n1251, n1249, n687);
nor  g1308 (n1330, n680, n683, n1278, n686);
xor  g1309 (n1326, n685, n677, n687, n1250);
nand g1310 (n1320, n1250, n1254, n1253, n1270);
and  g1311 (n1333, n730, n1250, n689, n674);
xnor g1312 (n1342, n1271, n1272, n1252);
nand g1313 (n1325, n1249, n684, n1274, n680);
nand g1314 (n1349, n1270, n690, n678, n731);
xnor g1315 (n1340, n678, n1277, n683, n733);
xnor g1316 (n1332, n1275, n689, n690, n678);
and  g1317 (n1343, n1277, n674, n687, n1276);
nor  g1318 (n1338, n735, n1252, n1251, n679);
and  g1319 (n1336, n732, n1273, n1253, n680);
and  g1320 (n1345, n734, n683, n688);
nor  g1321 (n1328, n1277, n1278, n676, n1249);
nor  g1322 (n1331, n730, n684, n1253, n681);
or   g1323 (n1348, n676, n682, n1254, n1279);
nand g1324 (n1318, n734, n1276, n1249, n1251);
xnor g1325 (n1350, n1273, n1270, n730, n1272);
xnor g1326 (n1321, n675, n1254, n678, n1271);
nor  g1327 (n1341, n1252, n731, n1274, n730);
nor  g1328 (n1337, n1276, n686, n731);
nand g1329 (n1346, n679, n1279, n732, n1277);
xnor g1330 (n1317, n677, n733, n1254, n688);
nand g1331 (n1323, n676, n682, n679);
xor  g1332 (n1316, n1278, n1271, n1275, n686);
xor  g1333 (n1339, n684, n689, n688, n1271);
xnor g1334 (n1324, n1253, n675, n681, n732);
nand g1335 (n1374, n1285, n698, n1284, n699);
nor  g1336 (n1376, n1323, n1286, n1283, n1285);
and  g1337 (n1355, n698, n708, n709, n704);
and  g1338 (n1360, n699, n1333, n700);
nand g1339 (n1369, n1334, n1279, n1284, n698);
xnor g1340 (n1382, n707, n709, n1283, n1285);
and  g1341 (n1361, n698, n1343, n703, n1282);
xnor g1342 (n1364, n1320, n1321, n1281);
and  g1343 (n1354, n699, n1336, n1244, n1286);
or   g1344 (n1359, n1283, n702, n1324, n703);
nor  g1345 (n1375, n1281, n1280, n707, n701);
xnor g1346 (n1365, n710, n1280, n702, n706);
xor  g1347 (n1380, n1345, n708, n1328, n702);
xor  g1348 (n1378, n1330, n1327, n705, n1337);
and  g1349 (n1356, n1282, n701, n1340);
and  g1350 (n1368, n710, n1287, n1279, n705);
nor  g1351 (n1370, n1283, n1339, n1332, n1284);
xor  g1352 (n1373, n1319, n701, n699, n697);
or   g1353 (n1357, n707, n1281, n1342, n709);
or   g1354 (n1367, n1335, n704, n1338, n1287);
xnor g1355 (n1372, n1316, n1286, n697, n708);
xnor g1356 (n1383, n704, n1317, n1318, n706);
nor  g1357 (n1363, n917, n1344, n706, n710);
and  g1358 (n1366, n697, n706, n1280, n700);
or   g1359 (n1362, n1280, n707, n1285, n1286);
xnor g1360 (n1377, n1326, n702, n1341, n708);
and  g1361 (n1381, n1325, n700, n1329, n705);
nand g1362 (n1371, n1282, n705, n703, n1322);
xnor g1363 (n1358, n1284, n710, n1282, n704);
or   g1364 (n1379, n703, n1287, n1331, n709);
nand g1365 (n1394, n927, n1358, n919, n1362);
xor  g1366 (n1389, n918, n1355, n1364, n927);
xor  g1367 (n1391, n923, n1363, n1360, n1357);
and  g1368 (n1390, n919, n927, n924, n923);
nand g1369 (n1392, n1354, n923, n925, n928);
and  g1370 (n1386, n921, n919, n918, n926);
nand g1371 (n1393, n921, n928, n926);
or   g1372 (n1388, n922, n920);
nor  g1373 (n1384, n918, n924, n921, n925);
nand g1374 (n1387, n922, n1359, n926, n924);
xnor g1375 (n1385, n1356, n1361, n925, n920);
xor  g1376 (n1413, n1302, n1305, n1391, n1297);
nor  g1377 (n1407, n1394, n1311, n1364, n1384);
and  g1378 (n1426, n1300, n1389, n1309, n1297);
or   g1379 (n1405, n1312, n1394, n1307);
and  g1380 (n1432, n1291, n1306, n1302, n1388);
nor  g1381 (n1412, n1299, n1392, n1290, n1306);
nor  g1382 (n1414, n1310, n1387, n1305);
or   g1383 (n1430, n1298, n1295, n1288, n1296);
and  g1384 (n1396, n1387, n1301, n1309, n1303);
or   g1385 (n1420, n1288, n1296, n1385, n1384);
xor  g1386 (n1419, n1313, n1314, n1300, n1309);
xor  g1387 (n1416, n1312, n1300, n1291, n1386);
nor  g1388 (n1431, n1299, n1313, n1294, n1390);
or   g1389 (n1399, n1390, n1308, n1393, n1288);
nor  g1390 (n1433, n1297, n1309, n1287, n1289);
xor  g1391 (n1423, n1295, n1297, n1393, n1385);
xnor g1392 (n1418, n1294, n1305, n1304, n1312);
or   g1393 (n1404, n1394, n1310, n1292, n1299);
xnor g1394 (n1428, n1303, n1311, n1387, n1392);
nand g1395 (n1409, n1315, n1296, n1301, n1293);
or   g1396 (n1400, n1304, n1386, n1298, n1302);
and  g1397 (n1427, n1315, n1314, n1393, n1293);
nand g1398 (n1421, n1391, n1308, n1293, n1290);
and  g1399 (n1397, n1304, n1298, n1303, n1299);
nand g1400 (n1403, n1307, n1315, n1301, n1314);
xnor g1401 (n1406, n1296, n1390, n1304, n1313);
or   g1402 (n1395, n1288, n1313, n1291, n1289);
xor  g1403 (n1402, n1310, n1295, n1298, n1365);
and  g1404 (n1425, n1305, n1308, n1300, n1389);
xor  g1405 (n1415, n1295, n1391, n1389, n1366);
nand g1406 (n1422, n1289, n1302, n1393, n1386);
nand g1407 (n1411, n1391, n1294, n1365, n1312);
xnor g1408 (n1429, n1394, n1315, n1388, n1292);
xor  g1409 (n1424, n1292, n1311, n1306, n1303);
nor  g1410 (n1410, n1290, n1311, n1307, n1388);
xor  g1411 (n1398, n1390, n1291, n1292, n1310);
and  g1412 (n1417, n1289, n1294, n1389, n1392);
or   g1413 (n1408, n1290, n1314, n1308, n1392);
nor  g1414 (n1401, n1301, n1293, n1306, n1388);
nor  g1415 (n1475, n932, n963, n1420, n938);
or   g1416 (n1477, n949, n1425, n936, n1367);
and  g1417 (n1446, n965, n955, n1413, n941);
xnor g1418 (n1455, n948, n930, n957, n959);
nand g1419 (n1450, n1432, n962, n954, n1370);
or   g1420 (n1445, n1409, n956, n1400, n1406);
xnor g1421 (n1453, n951, n961, n1433, n943);
or   g1422 (n1471, n933, n1408, n967, n946);
or   g1423 (n1447, n1415, n948, n1371, n935);
and  g1424 (n1469, n966, n969, n947, n953);
nand g1425 (n1462, n1405, n942, n945, n929);
and  g1426 (n1435, n968, n949, n960, n939);
nor  g1427 (n1452, n947, n964, n1428, n961);
and  g1428 (n1456, n1431, n969, n943, n941);
xnor g1429 (n1440, n943, n962, n970, n955);
nand g1430 (n1466, n1417, n1395, n1430, n940);
nand g1431 (n1436, n958, n1427, n953, n934);
or   g1432 (n1451, n1421, n941, n963, n958);
nor  g1433 (n1468, n946, n1367, n931, n968);
nor  g1434 (n1474, n962, n1430, n1432, n966);
or   g1435 (n1449, n1403, n956, n955, n1396);
nor  g1436 (n1441, n1416, n1399, n931, n933);
nor  g1437 (n1437, n929, n957, n950, n1370);
xor  g1438 (n1448, n1366, n1404, n964, n1426);
xnor g1439 (n1470, n944, n951, n965, n942);
or   g1440 (n1459, n931, n1398, n932, n1431);
and  g1441 (n1463, n959, n939, n936, n1418);
xnor g1442 (n1473, n952, n956, n965, n1397);
and  g1443 (n1454, n1368, n938, n939, n949);
xor  g1444 (n1443, n967, n937, n952);
nor  g1445 (n1465, n1401, n961, n1422, n930);
nand g1446 (n1439, n1412, n1414, n934, n966);
xnor g1447 (n1434, n954, n1407, n1411, n930);
nor  g1448 (n1442, n1423, n940, n954, n937);
nand g1449 (n1476, n958, n1410, n944, n952);
or   g1450 (n1478, n946, n1419, n1369, n933);
xnor g1451 (n1472, n969, n945, n959, n948);
xor  g1452 (n1460, n967, n944, n942, n936);
xnor g1453 (n1438, n964, n1429, n951, n957);
xor  g1454 (n1444, n1369, n953, n1368, n929);
xnor g1455 (n1457, n934, n963, n938, n1402);
or   g1456 (n1458, n945, n1424, n950, n947);
and  g1457 (n1461, n935, n1428, n970, n932);
xnor g1458 (n1467, n1433, n950, n960, n940);
nor  g1459 (n1464, n1429, n968, n935, n960);
xor  g1460 (n1479, n1371, n1372, n1434);
and  g1461 (n1481, n1375, n1373, n1374);
nor  g1462 (n1480, n1373, n1375, n1479);
buf  g1463 (n1483, n1480);
buf  g1464 (n1484, n1435);
buf  g1465 (n1482, n1480);
nor  g1466 (n1485, n1435, n1434);
and  g1467 (n1495, n1381, n1378, n1484, n1479);
or   g1468 (n1487, n1482, n1483, n1040);
nor  g1469 (n1491, n1377, n1382, n1349, n1040);
xor  g1470 (n1492, n1484, n1346, n1039, n1383);
nor  g1471 (n1490, n1376, n1352, n1485, n1381);
or   g1472 (n1497, n1040, n1479, n1481);
nor  g1473 (n1493, n1347, n1196, n690, n1376);
xnor g1474 (n1488, n1482, n1483, n1481);
nor  g1475 (n1500, n1216, n1382, n1378, n1350);
nor  g1476 (n1486, n1380, n1353, n1383, n1485);
xor  g1477 (n1494, n1379, n1039, n1380);
xor  g1478 (n1498, n1482, n1012, n1348, n1377);
or   g1479 (n1496, n1484, n1481, n1351, n1485);
nor  g1480 (n1489, n1040, n1024, n1482, n970);
nor  g1481 (n1499, n1379, n1012, n1485, n1484);
and  g1482 (n1537, n1436, n1486, n1465, n1440);
and  g1483 (n1502, n1490, n1441, n1498, n1466);
and  g1484 (n1539, n1488, n1478, n1473, n1498);
or   g1485 (n1503, n1496, n1458, n1459, n1461);
nor  g1486 (n1535, n1476, n1473, n1450, n1475);
and  g1487 (n1546, n1436, n1465, n1472, n1487);
nand g1488 (n1522, n1497, n1497, n1473, n1455);
xnor g1489 (n1527, n1442, n1435, n1477, n1438);
xor  g1490 (n1545, n1447, n1459, n1488);
and  g1491 (n1513, n1477, n1492, n1468, n1489);
or   g1492 (n1504, n1436, n1494, n1493, n1456);
nand g1493 (n1538, n1476, n1439, n1473, n1442);
nand g1494 (n1514, n1477, n1498, n1467, n1460);
nand g1495 (n1533, n1449, n1459, n1471, n1470);
nor  g1496 (n1518, n1453, n1448, n1463, n1457);
xnor g1497 (n1548, n1447, n1491, n1461, n1452);
nand g1498 (n1517, n1442, n1451, n1457, n1474);
and  g1499 (n1523, n1445, n1500, n1462, n1469);
and  g1500 (n1515, n1477, n1498, n1465, n1478);
xor  g1501 (n1510, n1439, n1489, n1487, n1456);
xnor g1502 (n1509, n1468, n1453, n1475, n1472);
or   g1503 (n1521, n1476, n1446, n1448, n1454);
nand g1504 (n1547, n1443, n1441, n1478, n1493);
xor  g1505 (n1541, n1451, n1447, n1465, n1486);
nor  g1506 (n1543, n1467, n1467, n1462, n1446);
nand g1507 (n1529, n1437, n1494, n1476);
nor  g1508 (n1531, n1437, n1450, n1460, n1487);
nor  g1509 (n1532, n1472, n1495, n1471);
and  g1510 (n1528, n1472, n1469, n1475, n1493);
or   g1511 (n1525, n1439, n1489, n1462, n1470);
nand g1512 (n1516, n1500, n1491, n1469, n1490);
or   g1513 (n1507, n1438, n1466, n1458, n1470);
and  g1514 (n1540, n1499, n1490, n1450, n1443);
nand g1515 (n1536, n1443, n1457, n1449, n1454);
nand g1516 (n1505, n1474, n1471, n1440, n1445);
and  g1517 (n1506, n1478, n1464, n1449, n1453);
and  g1518 (n1530, n1444, n1492, n1475, n1486);
and  g1519 (n1542, n1440, n1446, n1474, n1456);
xnor g1520 (n1512, n1460, n1458, n1461, n1471);
and  g1521 (n1508, n1451, n1452, n1500, n1438);
xnor g1522 (n1501, n1466, n1495, n1464, n1445);
nor  g1523 (n1520, n1467, n1463, n1437, n1444);
xor  g1524 (n1511, n1464, n1474, n1491, n1455);
and  g1525 (n1544, n1497, n1468, n1496, n1463);
nand g1526 (n1534, n1452, n1444, n1466, n1499);
xor  g1527 (n1526, n1500, n1496, n1448, n1470);
xor  g1528 (n1524, n1469, n1455, n1499);
or   g1529 (n1519, n1441, n1468, n1454, n1492);
and  g1530 (n1560, n1535, n1525, n1544, n1521);
and  g1531 (n1557, n1523, n18, n85, n86);
or   g1532 (n1584, n1540, n1516, n1501, n1533);
and  g1533 (n1555, n1543, n1510, n1544, n1533);
and  g1534 (n1579, n1526, n86, n1531, n1548);
xor  g1535 (n1553, n1523, n1503, n1527, n1534);
or   g1536 (n1568, n87, n86, n1526, n1508);
xor  g1537 (n1562, n1522, n1507, n1520, n1544);
and  g1538 (n1550, n1512, n1509, n1502);
or   g1539 (n1556, n1530, n1536, n1542);
and  g1540 (n1573, n1532, n1547, n1521, n1543);
nand g1541 (n1574, n1507, n1537, n1527, n1511);
nand g1542 (n1570, n1547, n1519, n1531, n1533);
nand g1543 (n1582, n1532, n1548, n1501, n1502);
xnor g1544 (n1551, n87, n1528, n1529, n1541);
nand g1545 (n1577, n1547, n1537, n1531, n1513);
xnor g1546 (n1583, n1535, n1536, n18, n1515);
nor  g1547 (n1561, n1503, n1542, n1530, n1529);
nor  g1548 (n1567, n1524, n1546, n1514, n1520);
nand g1549 (n1586, n1543, n1539, n1538);
xor  g1550 (n1563, n1504, n1546, n1506, n1545);
or   g1551 (n1580, n87, n1513, n1548, n1516);
and  g1552 (n1588, n1538, n1545, n1529, n1541);
or   g1553 (n1578, n1540, n1548, n1519, n1527);
nand g1554 (n1581, n1540, n84, n1505, n1541);
xnor g1555 (n1549, n85, n1543, n1547, n1524);
or   g1556 (n1572, n1510, n1533, n1528, n1545);
and  g1557 (n1571, n1546, n1505, n1525, n86);
nand g1558 (n1566, n1538, n1530, n1524, n1515);
or   g1559 (n1575, n1545, n1532, n1512, n1517);
nor  g1560 (n1587, n87, n1508, n1537, n1534);
and  g1561 (n1552, n1504, n1514, n18, n1544);
and  g1562 (n1559, n1534, n1537, n1522, n1535);
nor  g1563 (n1558, n1530, n1535, n1506, n1539);
or   g1564 (n1585, n1534, n1523, n1532, n1546);
or   g1565 (n1565, n1527, n1528, n1517, n1542);
and  g1566 (n1554, n1528, n1511, n1536);
nor  g1567 (n1569, n85, n1518, n1540, n1538);
nor  g1568 (n1564, n1518, n1529, n1541, n1526);
xnor g1569 (n1576, n85, n1539, n1531, n1525);
or   g1570 (n1591, n1552, n1551);
or   g1571 (n1589, n1554, n1549);
xnor g1572 (n1590, n1550, n1553);
xor  g1573 (n1592, n1555, n1556, n1589);
xnor g1574 (n1593, n1559, n1592, n1560, n1558);
xnor g1575 (n1594, n1561, n1557, n1592, n1562);
buf  g1576 (n1595, n1563);
and  g1577 (n1596, n1593, n1564, n1594);
xor  g1578 (n1600, n1596, n1587, n1573, n1576);
xor  g1579 (n1597, n1588, n1575, n1568, n1570);
nand g1580 (n1598, n1577, n1574, n1567, n1566);
xor  g1581 (n1601, n1580, n1571, n1578, n1581);
nand g1582 (n1602, n1596, n1582, n1583, n1569);
xnor g1583 (n1599, n1596, n1586, n1585, n1565);
xnor g1584 (n1604, n1579, n1595, n1572);
or   g1585 (n1603, n1584, n1596, n1595);
nand g1586 (n1608, n1602, n464, n1599, n1597);
xnor g1587 (n1606, n1603, n1591, n1598);
and  g1588 (n1607, n1591, n1601, n1590, n1600);
xnor g1589 (n1605, n1590, n464, n1604);
and  g1590 (n1609, n1607, n1606, n1608, n1605);
endmodule
