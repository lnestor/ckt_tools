

module Stat_2920_932
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n45,
  n46,
  n47,
  n48,
  n49,
  n1080,
  n1082,
  n1957,
  n1958,
  n1956,
  n1960,
  n2618,
  n2619,
  n2616,
  n2963,
  n2960,
  n2958,
  n2957,
  n2956,
  n2968,
  n2961,
  n2964,
  n2969,
  n2966,
  n2959,
  n2954,
  n2967,
  n2955,
  n2965,
  n2962,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input n33;
  input n34;
  input n35;
  input n36;
  input n37;
  input n38;
  input n39;
  input n40;
  input n41;
  input n42;
  input n43;
  input n44;
  input n45;
  input n46;
  input n47;
  input n48;
  input n49;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n1080;
  output n1082;
  output n1957;
  output n1958;
  output n1956;
  output n1960;
  output n2618;
  output n2619;
  output n2616;
  output n2963;
  output n2960;
  output n2958;
  output n2957;
  output n2956;
  output n2968;
  output n2961;
  output n2964;
  output n2969;
  output n2966;
  output n2959;
  output n2954;
  output n2967;
  output n2955;
  output n2965;
  output n2962;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1081;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1959;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2617;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n74,
    n1
  );


  nand
  g1
  (
    n75,
    n17,
    n28,
    n23,
    n32
  );


  nand
  g2
  (
    n50,
    n38,
    n23,
    n21,
    n12
  );


  or
  g3
  (
    n87,
    n24,
    n8,
    n11,
    n25
  );


  or
  g4
  (
    n73,
    n30,
    n7,
    n3,
    n11
  );


  xnor
  g5
  (
    n83,
    n19,
    n31,
    n6,
    n12
  );


  and
  g6
  (
    n65,
    n31,
    n21,
    n10,
    n34
  );


  or
  g7
  (
    n66,
    n28,
    n37,
    n18,
    n14
  );


  nor
  g8
  (
    n62,
    n24,
    n28,
    n32,
    n12
  );


  xnor
  g9
  (
    n60,
    n14,
    n30,
    n19,
    n16
  );


  nand
  g10
  (
    n71,
    n29,
    n7,
    n26,
    n4
  );


  xor
  g11
  (
    n52,
    n22,
    n1,
    n13,
    n36
  );


  xor
  g12
  (
    n55,
    n20,
    n31,
    n25,
    n14
  );


  xnor
  g13
  (
    n77,
    n18,
    n37,
    n33,
    n5
  );


  nand
  g14
  (
    n85,
    n34,
    n13,
    n26,
    n21
  );


  and
  g15
  (
    n79,
    n17,
    n4,
    n22,
    n13
  );


  or
  g16
  (
    n78,
    n9,
    n25,
    n14,
    n5
  );


  xnor
  g17
  (
    n69,
    n37,
    n16,
    n26,
    n20
  );


  nor
  g18
  (
    n86,
    n24,
    n3,
    n17,
    n5
  );


  nor
  g19
  (
    n53,
    n5,
    n10,
    n6,
    n35
  );


  nand
  g20
  (
    n72,
    n15,
    n35,
    n27,
    n36
  );


  or
  g21
  (
    n81,
    n2,
    n16,
    n29,
    n32
  );


  or
  g22
  (
    n59,
    n1,
    n19,
    n12,
    n30
  );


  xnor
  g23
  (
    n56,
    n23,
    n22,
    n19,
    n4
  );


  nand
  g24
  (
    n84,
    n27,
    n30,
    n36,
    n26
  );


  and
  g25
  (
    n57,
    n3,
    n9,
    n7,
    n15
  );


  nand
  g26
  (
    n70,
    n18,
    n33,
    n11,
    n22
  );


  xor
  g27
  (
    n58,
    n15,
    n33,
    n29,
    n20
  );


  or
  g28
  (
    n64,
    n32,
    n10,
    n20,
    n23
  );


  xnor
  g29
  (
    n51,
    n10,
    n9,
    n15,
    n37
  );


  xor
  g30
  (
    n76,
    n4,
    n6,
    n24,
    n17
  );


  xor
  g31
  (
    n63,
    n7,
    n2,
    n35,
    n13
  );


  xnor
  g32
  (
    n61,
    n35,
    n31,
    n34,
    n27
  );


  and
  g33
  (
    n54,
    n27,
    n28,
    n29,
    n6
  );


  xor
  g34
  (
    n82,
    n25,
    n11,
    n2,
    n8
  );


  or
  g35
  (
    n67,
    n2,
    n21,
    n8,
    n33
  );


  xnor
  g36
  (
    n68,
    n3,
    n36,
    n8,
    n1
  );


  nor
  g37
  (
    KeyWire_0_39,
    n34,
    n16,
    n9,
    n18
  );


  buf
  g38
  (
    n88,
    n50
  );


  not
  g39
  (
    n89,
    n88
  );


  buf
  g40
  (
    n92,
    n88
  );


  buf
  g41
  (
    n90,
    n88
  );


  buf
  g42
  (
    n91,
    n88
  );


  buf
  g43
  (
    n94,
    n89
  );


  buf
  g44
  (
    n98,
    n41
  );


  not
  g45
  (
    n93,
    n39
  );


  not
  g46
  (
    n99,
    n42
  );


  not
  g47
  (
    n103,
    n91
  );


  not
  g48
  (
    n96,
    n92
  );


  not
  g49
  (
    n106,
    n40
  );


  not
  g50
  (
    n97,
    n41
  );


  not
  g51
  (
    n102,
    n91
  );


  xor
  g52
  (
    n101,
    n91,
    n90,
    n39
  );


  xnor
  g53
  (
    n95,
    n91,
    n92,
    n40,
    n41
  );


  nand
  g54
  (
    n107,
    n38,
    n89,
    n40,
    n90
  );


  xor
  g55
  (
    n105,
    n90,
    n92,
    n38
  );


  and
  g56
  (
    n104,
    n92,
    n90,
    n89,
    n39
  );


  or
  g57
  (
    n100,
    n41,
    n39,
    n89,
    n40
  );


  buf
  g58
  (
    n130,
    n96
  );


  buf
  g59
  (
    n123,
    n97
  );


  not
  g60
  (
    n161,
    n105
  );


  buf
  g61
  (
    n110,
    n94
  );


  buf
  g62
  (
    n108,
    n104
  );


  not
  g63
  (
    n138,
    n97
  );


  buf
  g64
  (
    n109,
    n106
  );


  buf
  g65
  (
    n141,
    n99
  );


  buf
  g66
  (
    n131,
    n103
  );


  buf
  g67
  (
    n142,
    n93
  );


  buf
  g68
  (
    n153,
    n95
  );


  buf
  g69
  (
    n118,
    n93
  );


  buf
  g70
  (
    n143,
    n93
  );


  not
  g71
  (
    n152,
    n104
  );


  not
  g72
  (
    n136,
    n104
  );


  not
  g73
  (
    n129,
    n98
  );


  buf
  g74
  (
    n116,
    n97
  );


  buf
  g75
  (
    n148,
    n106
  );


  buf
  g76
  (
    n156,
    n98
  );


  not
  g77
  (
    KeyWire_0_2,
    n94
  );


  not
  g78
  (
    n134,
    n100
  );


  not
  g79
  (
    n121,
    n99
  );


  not
  g80
  (
    n155,
    n105
  );


  buf
  g81
  (
    n158,
    n100
  );


  not
  g82
  (
    n128,
    n96
  );


  not
  g83
  (
    n163,
    n103
  );


  not
  g84
  (
    n137,
    n101
  );


  not
  g85
  (
    n132,
    n102
  );


  buf
  g86
  (
    n147,
    n101
  );


  buf
  g87
  (
    n154,
    n103
  );


  buf
  g88
  (
    n144,
    n94
  );


  not
  g89
  (
    n115,
    n99
  );


  buf
  g90
  (
    n120,
    n104
  );


  buf
  g91
  (
    n133,
    n103
  );


  buf
  g92
  (
    n151,
    n95
  );


  buf
  g93
  (
    n127,
    n96
  );


  buf
  g94
  (
    n162,
    n95
  );


  not
  g95
  (
    n157,
    n106
  );


  buf
  g96
  (
    n150,
    n100
  );


  not
  g97
  (
    n124,
    n95
  );


  buf
  g98
  (
    n139,
    n102
  );


  buf
  g99
  (
    KeyWire_0_62,
    n98
  );


  not
  g100
  (
    n114,
    n101
  );


  not
  g101
  (
    n160,
    n97
  );


  buf
  g102
  (
    n125,
    n102
  );


  buf
  g103
  (
    n159,
    n93
  );


  not
  g104
  (
    n113,
    n106
  );


  buf
  g105
  (
    n140,
    n99
  );


  buf
  g106
  (
    n117,
    n102
  );


  not
  g107
  (
    n135,
    n105
  );


  buf
  g108
  (
    n122,
    n94
  );


  not
  g109
  (
    n119,
    n101
  );


  buf
  g110
  (
    n146,
    n96
  );


  not
  g111
  (
    n149,
    n98
  );


  not
  g112
  (
    n111,
    n100
  );


  buf
  g113
  (
    n126,
    n105
  );


  not
  g114
  (
    n218,
    n125
  );


  not
  g115
  (
    n164,
    n113
  );


  not
  g116
  (
    n239,
    n124
  );


  buf
  g117
  (
    n194,
    n50
  );


  buf
  g118
  (
    n169,
    n50
  );


  buf
  g119
  (
    n167,
    n108
  );


  not
  g120
  (
    n235,
    n112
  );


  buf
  g121
  (
    n198,
    n117
  );


  buf
  g122
  (
    n238,
    n122
  );


  buf
  g123
  (
    n210,
    n119
  );


  buf
  g124
  (
    n192,
    n111
  );


  not
  g125
  (
    n176,
    n108
  );


  buf
  g126
  (
    n200,
    n118
  );


  not
  g127
  (
    n230,
    n121
  );


  not
  g128
  (
    n196,
    n124
  );


  not
  g129
  (
    n207,
    n126
  );


  buf
  g130
  (
    n240,
    n114
  );


  buf
  g131
  (
    n225,
    n109
  );


  buf
  g132
  (
    n188,
    n126
  );


  buf
  g133
  (
    n177,
    n115
  );


  not
  g134
  (
    n234,
    n113
  );


  not
  g135
  (
    n186,
    n127
  );


  not
  g136
  (
    n213,
    n119
  );


  not
  g137
  (
    n228,
    n114
  );


  buf
  g138
  (
    n195,
    n115
  );


  buf
  g139
  (
    n184,
    n111
  );


  not
  g140
  (
    n172,
    n110
  );


  buf
  g141
  (
    n226,
    n113
  );


  buf
  g142
  (
    n209,
    n110
  );


  not
  g143
  (
    n175,
    n116
  );


  buf
  g144
  (
    n191,
    n112
  );


  buf
  g145
  (
    n232,
    n114
  );


  buf
  g146
  (
    n178,
    n117
  );


  not
  g147
  (
    n219,
    n124
  );


  not
  g148
  (
    n212,
    n123
  );


  buf
  g149
  (
    n229,
    n123
  );


  buf
  g150
  (
    n216,
    n125
  );


  buf
  g151
  (
    n180,
    n123
  );


  not
  g152
  (
    n221,
    n116
  );


  buf
  g153
  (
    n204,
    n118
  );


  not
  g154
  (
    n173,
    n50
  );


  not
  g155
  (
    n166,
    n109
  );


  buf
  g156
  (
    n199,
    n114
  );


  not
  g157
  (
    n170,
    n118
  );


  buf
  g158
  (
    n222,
    n120
  );


  buf
  g159
  (
    KeyWire_0_0,
    n126
  );


  not
  g160
  (
    n174,
    n118
  );


  buf
  g161
  (
    n205,
    n110
  );


  buf
  g162
  (
    n211,
    n116
  );


  buf
  g163
  (
    n189,
    n116
  );


  buf
  g164
  (
    n181,
    n124
  );


  not
  g165
  (
    n231,
    n125
  );


  not
  g166
  (
    n223,
    n108
  );


  not
  g167
  (
    n237,
    n121
  );


  not
  g168
  (
    n214,
    n122
  );


  buf
  g169
  (
    n179,
    n123
  );


  not
  g170
  (
    n168,
    n120
  );


  buf
  g171
  (
    n165,
    n121
  );


  not
  g172
  (
    n236,
    n108
  );


  buf
  g173
  (
    n202,
    n126
  );


  not
  g174
  (
    n224,
    n117
  );


  not
  g175
  (
    n187,
    n110
  );


  buf
  g176
  (
    n233,
    n111
  );


  not
  g177
  (
    n227,
    n122
  );


  buf
  g178
  (
    n193,
    n117
  );


  buf
  g179
  (
    n197,
    n115
  );


  not
  g180
  (
    n217,
    n125
  );


  buf
  g181
  (
    n190,
    n113
  );


  not
  g182
  (
    n208,
    n112
  );


  buf
  g183
  (
    n171,
    n115
  );


  not
  g184
  (
    n206,
    n111
  );


  not
  g185
  (
    n183,
    n120
  );


  buf
  g186
  (
    n185,
    n109
  );


  buf
  g187
  (
    n220,
    n119
  );


  not
  g188
  (
    n203,
    n119
  );


  not
  g189
  (
    n201,
    n122
  );


  xnor
  g190
  (
    n215,
    n109,
    n120,
    n121,
    n112
  );


  buf
  g191
  (
    n257,
    n170
  );


  buf
  g192
  (
    n246,
    n164
  );


  not
  g193
  (
    n256,
    n166
  );


  buf
  g194
  (
    n264,
    n165
  );


  not
  g195
  (
    n248,
    n169
  );


  not
  g196
  (
    n250,
    n169
  );


  buf
  g197
  (
    n262,
    n168
  );


  not
  g198
  (
    n241,
    n167
  );


  buf
  g199
  (
    n242,
    n168
  );


  not
  g200
  (
    n247,
    n165
  );


  not
  g201
  (
    n259,
    n164
  );


  not
  g202
  (
    n249,
    n164
  );


  buf
  g203
  (
    n263,
    n165
  );


  not
  g204
  (
    n245,
    n164
  );


  buf
  g205
  (
    n243,
    n169
  );


  not
  g206
  (
    n255,
    n166
  );


  not
  g207
  (
    n258,
    n169
  );


  buf
  g208
  (
    n261,
    n166
  );


  not
  g209
  (
    n252,
    n167
  );


  not
  g210
  (
    n265,
    n167
  );


  buf
  g211
  (
    n253,
    n165
  );


  not
  g212
  (
    n254,
    n167
  );


  buf
  g213
  (
    n244,
    n166
  );


  not
  g214
  (
    n260,
    n168
  );


  buf
  g215
  (
    n251,
    n168
  );


  xnor
  g216
  (
    n282,
    n242,
    n184,
    n201,
    n203
  );


  and
  g217
  (
    n347,
    n172,
    n198,
    n175,
    n261
  );


  nor
  g218
  (
    n284,
    n214,
    n194,
    n42,
    n184
  );


  xor
  g219
  (
    n276,
    n185,
    n220,
    n45,
    n204
  );


  nand
  g220
  (
    n308,
    n258,
    n211,
    n191,
    n247
  );


  nor
  g221
  (
    n344,
    n218,
    n173,
    n209,
    n225
  );


  nand
  g222
  (
    n300,
    n223,
    n236,
    n187,
    n252
  );


  xnor
  g223
  (
    n352,
    n197,
    n259,
    n234,
    n255
  );


  or
  g224
  (
    n269,
    n206,
    n44,
    n255,
    n170
  );


  xnor
  g225
  (
    n338,
    n239,
    n252,
    n242,
    n179
  );


  xor
  g226
  (
    n280,
    n201,
    n255,
    n254,
    n203
  );


  xor
  g227
  (
    n295,
    n207,
    n192,
    n189,
    n215
  );


  nand
  g228
  (
    n362,
    n181,
    n261,
    n199,
    n182
  );


  and
  g229
  (
    n340,
    n192,
    n243,
    n194,
    n46
  );


  xnor
  g230
  (
    n279,
    n262,
    n262,
    n207,
    n257
  );


  nor
  g231
  (
    n354,
    n223,
    n225,
    n260,
    n202
  );


  nor
  g232
  (
    n345,
    n43,
    n221,
    n224,
    n248
  );


  xor
  g233
  (
    n274,
    n47,
    n199,
    n197,
    n201
  );


  xnor
  g234
  (
    n322,
    n174,
    n43,
    n212,
    n239
  );


  nor
  g235
  (
    n358,
    n174,
    n238,
    n264,
    n202
  );


  nor
  g236
  (
    n311,
    n186,
    n170,
    n261,
    n265
  );


  xor
  g237
  (
    n291,
    n249,
    n198,
    n194,
    n239
  );


  xnor
  g238
  (
    n277,
    n209,
    n205,
    n217,
    n208
  );


  or
  g239
  (
    n312,
    n251,
    n195,
    n44,
    n227
  );


  nand
  g240
  (
    n273,
    n183,
    n235,
    n263,
    n248
  );


  or
  g241
  (
    n301,
    n245,
    n225,
    n246,
    n175
  );


  xnor
  g242
  (
    n297,
    n223,
    n215,
    n214,
    n188
  );


  xor
  g243
  (
    n333,
    n199,
    n222,
    n237,
    n232
  );


  xnor
  g244
  (
    n314,
    n186,
    n216,
    n42,
    n262
  );


  xnor
  g245
  (
    n350,
    n204,
    n180,
    n221,
    n186
  );


  nor
  g246
  (
    n287,
    n238,
    n238,
    n244,
    n174
  );


  xor
  g247
  (
    n309,
    n250,
    n190,
    n202,
    n228
  );


  and
  g248
  (
    n343,
    n44,
    n227,
    n215,
    n245
  );


  and
  g249
  (
    n267,
    n213,
    n172,
    n194,
    n43
  );


  xor
  g250
  (
    n348,
    n260,
    n185,
    n258,
    n249
  );


  or
  g251
  (
    n326,
    n214,
    n222,
    n212,
    n238
  );


  or
  g252
  (
    n294,
    n236,
    n256,
    n172,
    n210
  );


  xor
  g253
  (
    n275,
    n198,
    n216,
    n241,
    n254
  );


  xnor
  g254
  (
    n361,
    n256,
    n214,
    n204,
    n246
  );


  xnor
  g255
  (
    n310,
    n195,
    n180,
    n254,
    n208
  );


  nor
  g256
  (
    n330,
    n235,
    n178,
    n244,
    n184
  );


  nand
  g257
  (
    n351,
    n181,
    n215,
    n256,
    n191
  );


  nand
  g258
  (
    n335,
    n47,
    n252,
    n250,
    n197
  );


  xor
  g259
  (
    n290,
    n249,
    n226,
    n236,
    n248
  );


  nand
  g260
  (
    n365,
    n233,
    n183,
    n229,
    n193
  );


  xor
  g261
  (
    n325,
    n225,
    n218,
    n179,
    n205
  );


  nand
  g262
  (
    n319,
    n190,
    n175,
    n45,
    n217
  );


  nor
  g263
  (
    n268,
    n210,
    n180,
    n184,
    n188
  );


  xnor
  g264
  (
    n271,
    n209,
    n253,
    n193,
    n254
  );


  nor
  g265
  (
    n337,
    n190,
    n251,
    n241,
    n43
  );


  and
  g266
  (
    n321,
    n218,
    n196,
    n189,
    n241
  );


  nor
  g267
  (
    n342,
    n234,
    n183,
    n181,
    n260
  );


  nor
  g268
  (
    n289,
    n187,
    n228,
    n197,
    n262
  );


  nor
  g269
  (
    n329,
    n243,
    n263,
    n200,
    n45
  );


  xor
  g270
  (
    n307,
    n191,
    n219,
    n261,
    n224
  );


  or
  g271
  (
    n328,
    n224,
    n187,
    n230,
    n227
  );


  or
  g272
  (
    n357,
    n213,
    n206,
    n217,
    n218
  );


  xnor
  g273
  (
    n332,
    n264,
    n232,
    n207,
    n176
  );


  nor
  g274
  (
    n316,
    n263,
    n245,
    n224,
    n265
  );


  or
  g275
  (
    n356,
    n230,
    n233,
    n235,
    n199
  );


  xor
  g276
  (
    n341,
    n173,
    n226,
    n176,
    n196
  );


  xnor
  g277
  (
    n302,
    n210,
    n265,
    n200,
    n230
  );


  and
  g278
  (
    n304,
    n177,
    n232,
    n212,
    n217
  );


  xor
  g279
  (
    n296,
    n196,
    n256,
    n234,
    n176
  );


  and
  g280
  (
    n293,
    n200,
    n220,
    n189,
    n212
  );


  nand
  g281
  (
    n339,
    n211,
    n192,
    n232,
    n259
  );


  xor
  g282
  (
    n327,
    n251,
    n259,
    n203,
    n208
  );


  nand
  g283
  (
    n355,
    n221,
    n231,
    n182,
    n205
  );


  xnor
  g284
  (
    n346,
    n188,
    n208,
    n229,
    n246
  );


  xor
  g285
  (
    n285,
    n177,
    n173,
    n235,
    n223
  );


  xor
  g286
  (
    n286,
    n250,
    n234,
    n45,
    n248
  );


  and
  g287
  (
    n278,
    n177,
    n251,
    n229,
    n204
  );


  or
  g288
  (
    n363,
    n246,
    n237,
    n195,
    n193
  );


  xnor
  g289
  (
    n364,
    n178,
    n177,
    n195,
    n47
  );


  and
  g290
  (
    n349,
    n252,
    n171,
    n230
  );


  and
  g291
  (
    n317,
    n242,
    n181,
    n222,
    n231
  );


  nand
  g292
  (
    n306,
    n206,
    n201,
    n205,
    n180
  );


  and
  g293
  (
    n360,
    n190,
    n237,
    n263,
    n176
  );


  xnor
  g294
  (
    n323,
    n219,
    n257,
    n253,
    n247
  );


  and
  g295
  (
    n305,
    n260,
    n226,
    n220,
    n171
  );


  nand
  g296
  (
    n324,
    n42,
    n257,
    n210,
    n237
  );


  or
  g297
  (
    n334,
    n231,
    n173,
    n192,
    n249
  );


  nor
  g298
  (
    n270,
    n46,
    n207,
    n213,
    n245
  );


  and
  g299
  (
    n336,
    n175,
    n253,
    n198,
    n46
  );


  and
  g300
  (
    n303,
    n226,
    n222,
    n189,
    n265
  );


  and
  g301
  (
    n359,
    n187,
    n228,
    n209,
    n191
  );


  or
  g302
  (
    n313,
    n243,
    n264,
    n172,
    n182
  );


  nand
  g303
  (
    n288,
    n183,
    n253,
    n220,
    n227
  );


  and
  g304
  (
    n320,
    n182,
    n250,
    n200,
    n231
  );


  xnor
  g305
  (
    n318,
    n185,
    n247,
    n257,
    n178
  );


  and
  g306
  (
    n283,
    n46,
    n247,
    n211,
    n258
  );


  or
  g307
  (
    n281,
    n264,
    n203,
    n219,
    n229
  );


  or
  g308
  (
    n292,
    n188,
    n179,
    n185,
    n219
  );


  xnor
  g309
  (
    n315,
    n244,
    n243,
    n211,
    n258
  );


  or
  g310
  (
    n353,
    n178,
    n193,
    n216,
    n228
  );


  and
  g311
  (
    n272,
    n206,
    n170,
    n179,
    n241
  );


  nor
  g312
  (
    n266,
    n233,
    n259,
    n242,
    n255
  );


  and
  g313
  (
    n298,
    n233,
    n202,
    n213,
    n221
  );


  or
  g314
  (
    n331,
    n44,
    n236,
    n186,
    n196
  );


  or
  g315
  (
    n299,
    n244,
    n171,
    n174,
    n216
  );


  not
  g316
  (
    n378,
    n269
  );


  not
  g317
  (
    n366,
    n127
  );


  not
  g318
  (
    n374,
    n267
  );


  buf
  g319
  (
    n372,
    n269
  );


  buf
  g320
  (
    n368,
    n266
  );


  not
  g321
  (
    n376,
    n267
  );


  not
  g322
  (
    n375,
    n270
  );


  buf
  g323
  (
    n370,
    n127
  );


  buf
  g324
  (
    n380,
    n128
  );


  buf
  g325
  (
    n373,
    n266
  );


  not
  g326
  (
    n371,
    n267
  );


  not
  g327
  (
    n377,
    n268
  );


  xnor
  g328
  (
    KeyWire_0_13,
    n269,
    n128,
    n266,
    n267
  );


  and
  g329
  (
    n367,
    n266,
    n268
  );


  xor
  g330
  (
    n369,
    n269,
    n128,
    n127
  );


  and
  g331
  (
    n383,
    n132,
    n134,
    n135
  );


  xor
  g332
  (
    n387,
    n367,
    n130,
    n131,
    n129
  );


  xor
  g333
  (
    n385,
    n132,
    n131,
    n366,
    n134
  );


  and
  g334
  (
    n384,
    n367,
    n135,
    n131,
    n129
  );


  nand
  g335
  (
    n382,
    n131,
    n132,
    n366
  );


  xnor
  g336
  (
    n386,
    n130,
    n129,
    n133
  );


  nand
  g337
  (
    n388,
    n130,
    n367,
    n134,
    n133
  );


  and
  g338
  (
    n381,
    n130,
    n366,
    n133
  );


  and
  g339
  (
    n389,
    n368,
    n367,
    n133,
    n134
  );


  xor
  g340
  (
    n398,
    n57,
    n58,
    n240,
    n387
  );


  xor
  g341
  (
    n421,
    n388,
    n64,
    n63,
    n386
  );


  xnor
  g342
  (
    n401,
    n64,
    n66,
    n384,
    n62
  );


  nor
  g343
  (
    n408,
    n385,
    n73,
    n51
  );


  and
  g344
  (
    n412,
    n240,
    n61,
    n54,
    n53
  );


  nand
  g345
  (
    n420,
    n73,
    n389,
    n381,
    n71
  );


  or
  g346
  (
    n416,
    n61,
    n384,
    n385,
    n71
  );


  nor
  g347
  (
    n392,
    n385,
    n52,
    n382,
    n64
  );


  xor
  g348
  (
    n402,
    n385,
    n51,
    n65,
    n71
  );


  xor
  g349
  (
    n390,
    n53,
    n67,
    n69,
    n58
  );


  nand
  g350
  (
    n414,
    n68,
    n72,
    n60
  );


  nand
  g351
  (
    n409,
    n383,
    n382,
    n58,
    n57
  );


  or
  g352
  (
    n417,
    n66,
    n66,
    n60,
    n384
  );


  xnor
  g353
  (
    n406,
    n383,
    n55,
    n59,
    n72
  );


  xor
  g354
  (
    n415,
    n386,
    n56,
    n57
  );


  xor
  g355
  (
    n393,
    n384,
    n55,
    n67
  );


  nand
  g356
  (
    n400,
    n386,
    n69,
    n65,
    n68
  );


  and
  g357
  (
    n394,
    n70,
    n60,
    n388,
    n65
  );


  and
  g358
  (
    n395,
    n62,
    n239,
    n383,
    n53
  );


  nand
  g359
  (
    n397,
    n72,
    n52,
    n68,
    n60
  );


  and
  g360
  (
    KeyWire_0_14,
    n56,
    n58,
    n54,
    n52
  );


  and
  g361
  (
    n404,
    n64,
    n388,
    n382,
    n54
  );


  xnor
  g362
  (
    n403,
    n70,
    n70,
    n59,
    n67
  );


  or
  g363
  (
    KeyWire_0_22,
    n383,
    n69,
    n57,
    n71
  );


  xnor
  g364
  (
    n391,
    n56,
    n240,
    n62
  );


  xnor
  g365
  (
    n419,
    n51,
    n389,
    n59,
    n68
  );


  nand
  g366
  (
    n407,
    n53,
    n55,
    n382,
    n59
  );


  xor
  g367
  (
    n405,
    n61,
    n66,
    n69,
    n387
  );


  and
  g368
  (
    n411,
    n54,
    n389,
    n388,
    n387
  );


  nand
  g369
  (
    n396,
    n386,
    n62,
    n61,
    n387
  );


  nor
  g370
  (
    n399,
    n70,
    n52,
    n63,
    n65
  );


  or
  g371
  (
    n413,
    n73,
    n63,
    n67
  );


  not
  g372
  (
    n438,
    n400
  );


  buf
  g373
  (
    n484,
    n419
  );


  buf
  g374
  (
    n447,
    n407
  );


  buf
  g375
  (
    n480,
    n420
  );


  not
  g376
  (
    KeyWire_0_58,
    n400
  );


  not
  g377
  (
    n434,
    n404
  );


  buf
  g378
  (
    n486,
    n401
  );


  not
  g379
  (
    n435,
    n408
  );


  not
  g380
  (
    n445,
    n421
  );


  not
  g381
  (
    n492,
    n389
  );


  not
  g382
  (
    n454,
    n393
  );


  buf
  g383
  (
    n457,
    n416
  );


  not
  g384
  (
    n430,
    n398
  );


  buf
  g385
  (
    n446,
    n420
  );


  buf
  g386
  (
    n466,
    n397
  );


  not
  g387
  (
    n443,
    n410
  );


  buf
  g388
  (
    n433,
    n419
  );


  not
  g389
  (
    n487,
    n397
  );


  not
  g390
  (
    n470,
    n417
  );


  not
  g391
  (
    n441,
    n409
  );


  not
  g392
  (
    n449,
    n407
  );


  not
  g393
  (
    n475,
    n417
  );


  buf
  g394
  (
    n453,
    n402
  );


  buf
  g395
  (
    n490,
    n417
  );


  not
  g396
  (
    n479,
    n416
  );


  not
  g397
  (
    n462,
    n412
  );


  not
  g398
  (
    n473,
    n391
  );


  buf
  g399
  (
    n431,
    n419
  );


  not
  g400
  (
    n478,
    n418
  );


  buf
  g401
  (
    n463,
    n419
  );


  buf
  g402
  (
    n437,
    n415
  );


  not
  g403
  (
    n436,
    n412
  );


  buf
  g404
  (
    n429,
    n403
  );


  not
  g405
  (
    n476,
    n392
  );


  buf
  g406
  (
    n493,
    n410
  );


  not
  g407
  (
    n468,
    n392
  );


  buf
  g408
  (
    n461,
    n421
  );


  not
  g409
  (
    n489,
    n417
  );


  buf
  g410
  (
    n427,
    n418
  );


  not
  g411
  (
    n477,
    n398
  );


  not
  g412
  (
    n460,
    n408
  );


  not
  g413
  (
    n483,
    n411
  );


  buf
  g414
  (
    n428,
    n406
  );


  not
  g415
  (
    n440,
    n416
  );


  buf
  g416
  (
    n451,
    n402
  );


  buf
  g417
  (
    KeyWire_0_59,
    n411
  );


  buf
  g418
  (
    n448,
    n409
  );


  buf
  g419
  (
    n494,
    n395
  );


  buf
  g420
  (
    n474,
    n421
  );


  not
  g421
  (
    n425,
    n399
  );


  not
  g422
  (
    n481,
    n396
  );


  not
  g423
  (
    n424,
    n413
  );


  not
  g424
  (
    n488,
    n393
  );


  not
  g425
  (
    n485,
    n394
  );


  not
  g426
  (
    n452,
    n395
  );


  buf
  g427
  (
    n469,
    n399
  );


  not
  g428
  (
    n450,
    n420
  );


  not
  g429
  (
    n459,
    n390
  );


  not
  g430
  (
    n482,
    n405
  );


  not
  g431
  (
    n442,
    n420
  );


  not
  g432
  (
    n456,
    n404
  );


  buf
  g433
  (
    n426,
    n416
  );


  not
  g434
  (
    n432,
    n418
  );


  buf
  g435
  (
    n423,
    n403
  );


  not
  g436
  (
    n439,
    n405
  );


  buf
  g437
  (
    n458,
    n406
  );


  not
  g438
  (
    KeyWire_0_3,
    n413
  );


  buf
  g439
  (
    n455,
    n394
  );


  buf
  g440
  (
    n472,
    n414
  );


  not
  g441
  (
    n471,
    n401
  );


  buf
  g442
  (
    n464,
    n396
  );


  not
  g443
  (
    n465,
    n418
  );


  and
  g444
  (
    n467,
    n415,
    n414
  );


  xor
  g445
  (
    n503,
    n304,
    n288,
    n302,
    n336
  );


  nor
  g446
  (
    n546,
    n321,
    n305,
    n314,
    n271
  );


  nand
  g447
  (
    n565,
    n324,
    n439,
    n336
  );


  xnor
  g448
  (
    n574,
    n293,
    n422,
    n274,
    n343
  );


  nand
  g449
  (
    KeyWire_0_44,
    n278,
    n279,
    n437,
    n301
  );


  nor
  g450
  (
    n564,
    n307,
    n306,
    n277,
    n338
  );


  nand
  g451
  (
    n521,
    n298,
    n280,
    n288,
    n310
  );


  and
  g452
  (
    n524,
    n328,
    n333,
    n428,
    n300
  );


  xor
  g453
  (
    n526,
    n422,
    n330,
    n290,
    n289
  );


  nor
  g454
  (
    n566,
    n295,
    n302,
    n300,
    n334
  );


  and
  g455
  (
    n523,
    n331,
    n313,
    n299,
    n286
  );


  xor
  g456
  (
    n540,
    n330,
    n343,
    n332,
    n270
  );


  nand
  g457
  (
    n535,
    n294,
    n427,
    n431,
    n430
  );


  xor
  g458
  (
    n508,
    n277,
    n332,
    n436,
    n278
  );


  xor
  g459
  (
    n561,
    n306,
    n286,
    n302,
    n293
  );


  or
  g460
  (
    n582,
    n440,
    n270,
    n273,
    n312
  );


  nor
  g461
  (
    n568,
    n271,
    n323,
    n439,
    n274
  );


  and
  g462
  (
    n578,
    n283,
    n338,
    n426,
    n443
  );


  and
  g463
  (
    n542,
    n300,
    n424,
    n427,
    n430
  );


  xor
  g464
  (
    n507,
    n340,
    n344,
    n441,
    n307
  );


  and
  g465
  (
    n588,
    n435,
    n294,
    n307,
    n428
  );


  and
  g466
  (
    n576,
    n425,
    n324,
    n426,
    n439
  );


  or
  g467
  (
    n528,
    n306,
    n322,
    n329,
    n315
  );


  or
  g468
  (
    n562,
    n281,
    n280,
    n292,
    n428
  );


  nor
  g469
  (
    n570,
    n310,
    n332,
    n315,
    n284
  );


  xnor
  g470
  (
    n555,
    n335,
    n322,
    n306,
    n286
  );


  nand
  g471
  (
    n584,
    n287,
    n440,
    n434,
    n432
  );


  nand
  g472
  (
    n533,
    n309,
    n443,
    n321,
    n296
  );


  and
  g473
  (
    n573,
    n310,
    n422,
    n297,
    n329
  );


  xor
  g474
  (
    n539,
    n437,
    n431,
    n323,
    n282
  );


  and
  g475
  (
    n513,
    n273,
    n337,
    n294,
    n339
  );


  xor
  g476
  (
    n512,
    n328,
    n303,
    n329,
    n442
  );


  xnor
  g477
  (
    n520,
    n443,
    n312,
    n327,
    n328
  );


  or
  g478
  (
    n544,
    n446,
    n436,
    n335,
    n283
  );


  xnor
  g479
  (
    n518,
    n281,
    n275,
    n343,
    n319
  );


  nor
  g480
  (
    n495,
    n423,
    n291,
    n320,
    n318
  );


  nor
  g481
  (
    n559,
    n323,
    n337,
    n274,
    n318
  );


  or
  g482
  (
    n591,
    n276,
    n282,
    n311,
    n283
  );


  or
  g483
  (
    n511,
    n446,
    n422,
    n304,
    n436
  );


  nand
  g484
  (
    n497,
    n334,
    n322,
    n297,
    n428
  );


  nor
  g485
  (
    n531,
    n314,
    n434,
    n293,
    n443
  );


  and
  g486
  (
    n548,
    n323,
    n290,
    n441,
    n318
  );


  xor
  g487
  (
    n530,
    n433,
    n442,
    n332,
    n292
  );


  nor
  g488
  (
    n505,
    n340,
    n302,
    n299,
    n276
  );


  nor
  g489
  (
    n587,
    n321,
    n342,
    n317,
    n292
  );


  xor
  g490
  (
    n592,
    n271,
    n432,
    n341,
    n314
  );


  nor
  g491
  (
    n529,
    n337,
    n432,
    n280,
    n424
  );


  xor
  g492
  (
    n527,
    n304,
    n296,
    n297,
    n325
  );


  xor
  g493
  (
    n577,
    n438,
    n325,
    n280,
    n286
  );


  or
  g494
  (
    n514,
    n335,
    n341,
    n272,
    n288
  );


  nand
  g495
  (
    n572,
    n433,
    n299,
    n423,
    n315
  );


  nor
  g496
  (
    n589,
    n272,
    n282,
    n431,
    n291
  );


  nor
  g497
  (
    n586,
    n444,
    n435,
    n291,
    n312
  );


  xor
  g498
  (
    n550,
    n290,
    n441,
    n325,
    n339
  );


  nand
  g499
  (
    n590,
    n301,
    n343,
    n308,
    n327
  );


  xor
  g500
  (
    n532,
    n311,
    n272,
    n426,
    n299
  );


  nor
  g501
  (
    n536,
    n309,
    n270,
    n331,
    n279
  );


  xor
  g502
  (
    n580,
    n435,
    n329,
    n310,
    n336
  );


  and
  g503
  (
    n545,
    n314,
    n294,
    n342,
    n298
  );


  nor
  g504
  (
    n553,
    n277,
    n326,
    n316,
    n308
  );


  nand
  g505
  (
    n557,
    n316,
    n324,
    n273,
    n341
  );


  xor
  g506
  (
    n558,
    n297,
    n330,
    n311,
    n445
  );


  xnor
  g507
  (
    n551,
    n328,
    n285,
    n316,
    n335
  );


  nor
  g508
  (
    n569,
    n296,
    n424,
    n326,
    n275
  );


  nor
  g509
  (
    n499,
    n315,
    n444,
    n284
  );


  xnor
  g510
  (
    n506,
    n321,
    n429,
    n320,
    n313
  );


  xor
  g511
  (
    n549,
    n295,
    n427,
    n425,
    n316
  );


  nand
  g512
  (
    n579,
    n441,
    n430,
    n438,
    n337
  );


  nor
  g513
  (
    n502,
    n276,
    n287,
    n289
  );


  or
  g514
  (
    n501,
    n438,
    n291,
    n285,
    n279
  );


  nor
  g515
  (
    n541,
    n444,
    n334,
    n308,
    n327
  );


  nor
  g516
  (
    n552,
    n340,
    n303,
    n436,
    n425
  );


  nor
  g517
  (
    n583,
    n325,
    n424,
    n275,
    n331
  );


  xnor
  g518
  (
    n500,
    n292,
    n426,
    n344,
    n311
  );


  and
  g519
  (
    n510,
    n301,
    n319,
    n305,
    n272
  );


  or
  g520
  (
    n516,
    n342,
    n429,
    n339,
    n331
  );


  xor
  g521
  (
    n563,
    n445,
    n276,
    n334,
    n423
  );


  xor
  g522
  (
    n498,
    n435,
    n303,
    n440,
    n279
  );


  nand
  g523
  (
    n554,
    n437,
    n305,
    n338,
    n283
  );


  nor
  g524
  (
    n517,
    n433,
    n340,
    n423,
    n444
  );


  or
  g525
  (
    n567,
    n273,
    n282,
    n309,
    n330
  );


  and
  g526
  (
    n496,
    n288,
    n303,
    n313,
    n434
  );


  nor
  g527
  (
    n581,
    n312,
    n277,
    n442,
    n287
  );


  nand
  g528
  (
    n504,
    n296,
    n285,
    n326,
    n313
  );


  or
  g529
  (
    n575,
    n298,
    n319,
    n295,
    n429
  );


  nand
  g530
  (
    n593,
    n317,
    n308,
    n289,
    n320
  );


  nand
  g531
  (
    n515,
    n293,
    n341,
    n298,
    n300
  );


  nand
  g532
  (
    n534,
    n320,
    n338,
    n304,
    n430
  );


  xnor
  g533
  (
    n571,
    n437,
    n278,
    n427,
    n290
  );


  xor
  g534
  (
    n537,
    n425,
    n278,
    n285,
    n446
  );


  or
  g535
  (
    n585,
    n318,
    n438,
    n431,
    n289
  );


  xor
  g536
  (
    n525,
    n301,
    n284,
    n326,
    n322
  );


  and
  g537
  (
    n560,
    n281,
    n433,
    n275,
    n324
  );


  and
  g538
  (
    n556,
    n295,
    n432,
    n442,
    n274
  );


  and
  g539
  (
    n543,
    n309,
    n319,
    n342,
    n445
  );


  xnor
  g540
  (
    n519,
    n281,
    n317,
    n271,
    n333
  );


  xnor
  g541
  (
    n538,
    n429,
    n305,
    n445,
    n434
  );


  nand
  g542
  (
    n509,
    n327,
    n307,
    n333,
    n440
  );


  xor
  g543
  (
    n522,
    n317,
    n333,
    n336,
    n339
  );


  not
  g544
  (
    n594,
    n499
  );


  not
  g545
  (
    n608,
    n502
  );


  not
  g546
  (
    n613,
    n501
  );


  not
  g547
  (
    KeyWire_0_19,
    n497
  );


  buf
  g548
  (
    KeyWire_0_27,
    n503
  );


  buf
  g549
  (
    n614,
    n495
  );


  buf
  g550
  (
    n622,
    n496
  );


  not
  g551
  (
    n597,
    n498
  );


  buf
  g552
  (
    n599,
    n498
  );


  buf
  g553
  (
    n625,
    n496
  );


  not
  g554
  (
    n629,
    n504
  );


  not
  g555
  (
    n623,
    n498
  );


  not
  g556
  (
    n621,
    n502
  );


  not
  g557
  (
    n628,
    n499
  );


  buf
  g558
  (
    n609,
    n501
  );


  buf
  g559
  (
    n600,
    n502
  );


  buf
  g560
  (
    KeyWire_0_53,
    n503
  );


  buf
  g561
  (
    n616,
    n500
  );


  not
  g562
  (
    n607,
    n500
  );


  buf
  g563
  (
    n601,
    n503
  );


  not
  g564
  (
    n602,
    n495
  );


  buf
  g565
  (
    n598,
    n503
  );


  not
  g566
  (
    n619,
    n496
  );


  buf
  g567
  (
    n605,
    n502
  );


  buf
  g568
  (
    n595,
    n501
  );


  not
  g569
  (
    n606,
    n500
  );


  not
  g570
  (
    n618,
    n497
  );


  not
  g571
  (
    n627,
    n497
  );


  not
  g572
  (
    n604,
    n501
  );


  not
  g573
  (
    n630,
    n500
  );


  not
  g574
  (
    n596,
    n495
  );


  buf
  g575
  (
    n624,
    n495
  );


  not
  g576
  (
    n612,
    n496
  );


  buf
  g577
  (
    n620,
    n497
  );


  buf
  g578
  (
    n617,
    n499
  );


  buf
  g579
  (
    n603,
    n498
  );


  not
  g580
  (
    n615,
    n499
  );


  buf
  g581
  (
    n647,
    n74
  );


  buf
  g582
  (
    n698,
    n77
  );


  not
  g583
  (
    n675,
    n148
  );


  buf
  g584
  (
    n709,
    n599
  );


  not
  g585
  (
    n641,
    n604
  );


  buf
  g586
  (
    n670,
    n143
  );


  buf
  g587
  (
    KeyWire_0_9,
    n597
  );


  not
  g588
  (
    n655,
    n601
  );


  not
  g589
  (
    n676,
    n613
  );


  not
  g590
  (
    n699,
    n607
  );


  not
  g591
  (
    n661,
    n144
  );


  not
  g592
  (
    n660,
    n608
  );


  not
  g593
  (
    n686,
    n596
  );


  not
  g594
  (
    n706,
    n150
  );


  not
  g595
  (
    n653,
    n603
  );


  not
  g596
  (
    n632,
    n137
  );


  buf
  g597
  (
    n673,
    n80
  );


  not
  g598
  (
    n667,
    n141
  );


  not
  g599
  (
    n682,
    n79
  );


  buf
  g600
  (
    n650,
    n142
  );


  buf
  g601
  (
    n648,
    n142
  );


  buf
  g602
  (
    n689,
    n598
  );


  buf
  g603
  (
    n683,
    n148
  );


  buf
  g604
  (
    n631,
    n140
  );


  buf
  g605
  (
    n703,
    n77
  );


  not
  g606
  (
    n642,
    n75
  );


  not
  g607
  (
    n690,
    n75
  );


  not
  g608
  (
    n678,
    n606
  );


  buf
  g609
  (
    n693,
    n77
  );


  buf
  g610
  (
    n664,
    n76
  );


  buf
  g611
  (
    n704,
    n149
  );


  not
  g612
  (
    n702,
    n138
  );


  buf
  g613
  (
    n712,
    n78
  );


  not
  g614
  (
    n711,
    n78
  );


  buf
  g615
  (
    n636,
    n151
  );


  buf
  g616
  (
    n634,
    n605
  );


  buf
  g617
  (
    n656,
    n138
  );


  buf
  g618
  (
    n662,
    n604
  );


  not
  g619
  (
    n645,
    n149
  );


  buf
  g620
  (
    n679,
    n597
  );


  buf
  g621
  (
    n700,
    n145
  );


  buf
  g622
  (
    KeyWire_0_52,
    n150
  );


  buf
  g623
  (
    n640,
    n144
  );


  buf
  g624
  (
    n657,
    n607
  );


  buf
  g625
  (
    n697,
    n146
  );


  buf
  g626
  (
    n663,
    n78
  );


  not
  g627
  (
    n637,
    n140
  );


  not
  g628
  (
    n643,
    n144
  );


  not
  g629
  (
    n685,
    n607
  );


  buf
  g630
  (
    n635,
    n151
  );


  buf
  g631
  (
    n666,
    n146
  );


  buf
  g632
  (
    n710,
    n144
  );


  not
  g633
  (
    n708,
    n140
  );


  buf
  g634
  (
    n646,
    n135
  );


  xnor
  g635
  (
    n695,
    n594,
    n608,
    n150,
    n606
  );


  or
  g636
  (
    n713,
    n145,
    n609,
    n74,
    n600
  );


  nor
  g637
  (
    n669,
    n609,
    n613,
    n137,
    n75
  );


  xnor
  g638
  (
    n644,
    n597,
    n605,
    n75,
    n142
  );


  and
  g639
  (
    n687,
    n136,
    n594,
    n596,
    n76
  );


  xnor
  g640
  (
    n696,
    n606,
    n600,
    n140,
    n143
  );


  xor
  g641
  (
    n668,
    n608,
    n147,
    n138,
    n598
  );


  and
  g642
  (
    n654,
    n610,
    n76,
    n596,
    n599
  );


  and
  g643
  (
    n691,
    n611,
    n141,
    n610,
    n612
  );


  nand
  g644
  (
    n705,
    n600,
    n78,
    n604,
    n607
  );


  xnor
  g645
  (
    n681,
    n143,
    n602,
    n139,
    n601
  );


  or
  g646
  (
    n651,
    n146,
    n603,
    n147,
    n79
  );


  nor
  g647
  (
    n665,
    n136,
    n73,
    n147,
    n600
  );


  xnor
  g648
  (
    n680,
    n137,
    n79,
    n603,
    n602
  );


  xnor
  g649
  (
    n638,
    n596,
    n595,
    n614,
    n139
  );


  nand
  g650
  (
    n649,
    n74,
    n602,
    n149,
    n613
  );


  and
  g651
  (
    n694,
    n609,
    n149,
    n614,
    n605
  );


  xor
  g652
  (
    n639,
    n598,
    n142,
    n148,
    n147
  );


  xnor
  g653
  (
    n674,
    n601,
    n614,
    n611,
    n597
  );


  or
  g654
  (
    n707,
    n613,
    n612,
    n139,
    n143
  );


  and
  g655
  (
    n714,
    n610,
    n594,
    n595,
    n151
  );


  or
  g656
  (
    n659,
    n79,
    n150,
    n137,
    n595
  );


  or
  g657
  (
    n633,
    n136,
    n611,
    n614,
    n610
  );


  xor
  g658
  (
    n658,
    n602,
    n139,
    n595,
    n141
  );


  xnor
  g659
  (
    n672,
    n145,
    n611,
    n599,
    n608
  );


  xor
  g660
  (
    n684,
    n138,
    n148,
    n609,
    n141
  );


  nand
  g661
  (
    n671,
    n145,
    n146,
    n605,
    n601
  );


  nor
  g662
  (
    n688,
    n603,
    n612,
    n594,
    n76
  );


  xnor
  g663
  (
    n692,
    n604,
    n606,
    n136,
    n599
  );


  nand
  g664
  (
    n652,
    n74,
    n598,
    n77,
    n612
  );


  not
  g665
  (
    n720,
    n631
  );


  not
  g666
  (
    n716,
    n632
  );


  buf
  g667
  (
    n719,
    n631
  );


  xnor
  g668
  (
    n718,
    n631,
    n632,
    n421,
    n634
  );


  xor
  g669
  (
    n715,
    n632,
    n633
  );


  and
  g670
  (
    n717,
    n634,
    n632,
    n631,
    n633
  );


  or
  g671
  (
    n723,
    n375,
    n369,
    n82,
    n368
  );


  nor
  g672
  (
    n732,
    n720,
    n371,
    n449,
    n715
  );


  xnor
  g673
  (
    n730,
    n718,
    n717,
    n370,
    n447
  );


  nand
  g674
  (
    n721,
    n720,
    n716,
    n80
  );


  and
  g675
  (
    n722,
    n371,
    n84,
    n720,
    n372
  );


  and
  g676
  (
    n731,
    n372,
    n716,
    n83,
    n376
  );


  nand
  g677
  (
    n741,
    n717,
    n372,
    n447,
    n718
  );


  nor
  g678
  (
    n733,
    n373,
    n375,
    n447,
    n374
  );


  xor
  g679
  (
    n738,
    n374,
    n81,
    n716,
    n718
  );


  xor
  g680
  (
    n725,
    n373,
    n720,
    n369,
    n719
  );


  nand
  g681
  (
    n728,
    n81,
    n371,
    n374,
    n375
  );


  nor
  g682
  (
    n737,
    n83,
    n83,
    n84,
    n369
  );


  or
  g683
  (
    n727,
    n368,
    n84,
    n82
  );


  nor
  g684
  (
    n739,
    n719,
    n719,
    n370,
    n448
  );


  nand
  g685
  (
    n734,
    n373,
    n369,
    n717,
    n81
  );


  or
  g686
  (
    n736,
    n373,
    n448,
    n447,
    n376
  );


  and
  g687
  (
    n729,
    n82,
    n80,
    n81,
    n719
  );


  nor
  g688
  (
    n735,
    n374,
    n376,
    n372,
    n370
  );


  nand
  g689
  (
    n740,
    n370,
    n448,
    n83,
    n718
  );


  xnor
  g690
  (
    n724,
    n80,
    n371,
    n717,
    n376
  );


  xnor
  g691
  (
    n726,
    n446,
    n448,
    n375,
    n368
  );


  not
  g692
  (
    n747,
    n724
  );


  not
  g693
  (
    n746,
    n721
  );


  not
  g694
  (
    n744,
    n721
  );


  buf
  g695
  (
    n745,
    n725
  );


  buf
  g696
  (
    n742,
    n724
  );


  not
  g697
  (
    n756,
    n724
  );


  buf
  g698
  (
    n751,
    n724
  );


  buf
  g699
  (
    n754,
    n723
  );


  buf
  g700
  (
    n743,
    n725
  );


  not
  g701
  (
    KeyWire_0_31,
    n721
  );


  buf
  g702
  (
    n752,
    n721
  );


  not
  g703
  (
    n758,
    n723
  );


  not
  g704
  (
    n748,
    n722
  );


  not
  g705
  (
    n757,
    n722
  );


  not
  g706
  (
    n759,
    n722
  );


  buf
  g707
  (
    n755,
    n725
  );


  not
  g708
  (
    n749,
    n723
  );


  buf
  g709
  (
    n760,
    n722
  );


  buf
  g710
  (
    n753,
    n723
  );


  xor
  g711
  (
    n774,
    n377,
    n377,
    n745,
    n157
  );


  xor
  g712
  (
    n775,
    n743,
    n377,
    n153,
    n154
  );


  xor
  g713
  (
    n766,
    n158,
    n157,
    n378
  );


  nand
  g714
  (
    n772,
    n154,
    n156,
    n152,
    n151
  );


  or
  g715
  (
    n761,
    n744,
    n152,
    n746
  );


  nand
  g716
  (
    n764,
    n377,
    n155,
    n634,
    n158
  );


  xnor
  g717
  (
    n773,
    n744,
    n156,
    n159,
    n378
  );


  and
  g718
  (
    KeyWire_0_12,
    n155,
    n743,
    n379,
    n745
  );


  xnor
  g719
  (
    n771,
    n153,
    n379,
    n744,
    n745
  );


  xnor
  g720
  (
    n762,
    n155,
    n380,
    n154,
    n379
  );


  or
  g721
  (
    n763,
    n745,
    n153,
    n742,
    n156
  );


  nor
  g722
  (
    n770,
    n156,
    n743,
    n152
  );


  nor
  g723
  (
    KeyWire_0_57,
    n157,
    n744,
    n158,
    n380
  );


  nand
  g724
  (
    n768,
    n152,
    n153,
    n154,
    n158
  );


  xor
  g725
  (
    n767,
    n379,
    n155,
    n378
  );


  nand
  g726
  (
    n791,
    n655,
    n659,
    n643,
    n647
  );


  xnor
  g727
  (
    KeyWire_0_23,
    n647,
    n644,
    n635
  );


  xor
  g728
  (
    n788,
    n766,
    n657,
    n655,
    n645
  );


  xor
  g729
  (
    n815,
    n637,
    n638,
    n650,
    n771
  );


  and
  g730
  (
    n817,
    n641,
    n661,
    n649,
    n773
  );


  and
  g731
  (
    n821,
    n775,
    n636,
    n770,
    n643
  );


  xnor
  g732
  (
    n799,
    n764,
    n768,
    n765,
    n664
  );


  xor
  g733
  (
    n783,
    n654,
    n671,
    n659,
    n636
  );


  nand
  g734
  (
    n790,
    n771,
    n667,
    n657,
    n663
  );


  nor
  g735
  (
    n810,
    n662,
    n771,
    n635,
    n657
  );


  and
  g736
  (
    n824,
    n655,
    n658,
    n669,
    n667
  );


  nand
  g737
  (
    n795,
    n668,
    n641,
    n635,
    n774
  );


  nor
  g738
  (
    n819,
    n768,
    n656,
    n774,
    n641
  );


  xnor
  g739
  (
    n825,
    n644,
    n649,
    n654,
    n774
  );


  xnor
  g740
  (
    n794,
    n769,
    n669,
    n636,
    n768
  );


  xor
  g741
  (
    n777,
    n644,
    n770,
    n648,
    n661
  );


  xor
  g742
  (
    n798,
    n670,
    n666,
    n652,
    n659
  );


  and
  g743
  (
    n823,
    n771,
    n637,
    n773
  );


  nor
  g744
  (
    n818,
    n775,
    n775,
    n653,
    n670
  );


  xor
  g745
  (
    n808,
    n641,
    n652,
    n764,
    n663
  );


  nor
  g746
  (
    n826,
    n657,
    n665,
    n648,
    n672
  );


  xnor
  g747
  (
    n781,
    n661,
    n648,
    n663,
    n668
  );


  nor
  g748
  (
    n785,
    n639,
    n658,
    n638,
    n774
  );


  or
  g749
  (
    n778,
    n664,
    n772,
    n646,
    n767
  );


  nand
  g750
  (
    n804,
    n763,
    n766,
    n652,
    n671
  );


  nand
  g751
  (
    n803,
    n640,
    n653,
    n664,
    n639
  );


  nor
  g752
  (
    n782,
    n669,
    n638,
    n651,
    n666
  );


  nand
  g753
  (
    n814,
    n767,
    n647,
    n646
  );


  xor
  g754
  (
    n809,
    n766,
    n658,
    n662,
    n654
  );


  xor
  g755
  (
    n812,
    n661,
    n655,
    n653,
    n658
  );


  xnor
  g756
  (
    n805,
    n773,
    n646,
    n672,
    n639
  );


  xnor
  g757
  (
    n789,
    n642,
    n645,
    n651,
    n650
  );


  and
  g758
  (
    n800,
    n667,
    n643,
    n644,
    n671
  );


  nor
  g759
  (
    n822,
    n772,
    n640,
    n660,
    n637
  );


  xnor
  g760
  (
    n793,
    n659,
    n669,
    n769,
    n768
  );


  nand
  g761
  (
    n787,
    n650,
    n770,
    n765
  );


  or
  g762
  (
    n802,
    n649,
    n642,
    n638,
    n647
  );


  and
  g763
  (
    n784,
    n769,
    n656,
    n648,
    n761
  );


  nor
  g764
  (
    n807,
    n652,
    n772,
    n762,
    n662
  );


  xor
  g765
  (
    n816,
    n651,
    n651,
    n640,
    n660
  );


  and
  g766
  (
    n792,
    n672,
    n665,
    n767,
    n645
  );


  xor
  g767
  (
    n820,
    n766,
    n665,
    n660
  );


  and
  g768
  (
    n786,
    n664,
    n767,
    n670,
    n637
  );


  and
  g769
  (
    n797,
    n775,
    n666,
    n671,
    n672
  );


  xor
  g770
  (
    n811,
    n656,
    n640,
    n765,
    n649
  );


  nor
  g771
  (
    n780,
    n643,
    n668,
    n665,
    n634
  );


  or
  g772
  (
    n813,
    n639,
    n642,
    n654,
    n666
  );


  nand
  g773
  (
    n801,
    n668,
    n670,
    n663,
    n763
  );


  nor
  g774
  (
    n806,
    n765,
    n667,
    n645,
    n642
  );


  xor
  g775
  (
    KeyWire_0_35,
    n772,
    n636,
    n653,
    n650
  );


  or
  g776
  (
    n776,
    n762,
    n769,
    n662,
    n656
  );


  buf
  g777
  (
    n843,
    n811
  );


  not
  g778
  (
    n837,
    n790
  );


  not
  g779
  (
    n864,
    n799
  );


  not
  g780
  (
    n841,
    n791
  );


  buf
  g781
  (
    n853,
    n800
  );


  not
  g782
  (
    n861,
    n810
  );


  not
  g783
  (
    n839,
    n787
  );


  not
  g784
  (
    n849,
    n796
  );


  not
  g785
  (
    n827,
    n785
  );


  buf
  g786
  (
    n844,
    n794
  );


  buf
  g787
  (
    n835,
    n777
  );


  not
  g788
  (
    n840,
    n807
  );


  not
  g789
  (
    n863,
    n813
  );


  not
  g790
  (
    n854,
    n781
  );


  not
  g791
  (
    n833,
    n778
  );


  buf
  g792
  (
    n828,
    n792
  );


  not
  g793
  (
    n855,
    n808
  );


  not
  g794
  (
    n830,
    n776
  );


  buf
  g795
  (
    n866,
    n789
  );


  buf
  g796
  (
    n852,
    n805
  );


  buf
  g797
  (
    n856,
    n793
  );


  not
  g798
  (
    n846,
    n783
  );


  not
  g799
  (
    n848,
    n815
  );


  not
  g800
  (
    n836,
    n795
  );


  buf
  g801
  (
    n857,
    n806
  );


  buf
  g802
  (
    n862,
    n780
  );


  buf
  g803
  (
    n834,
    n788
  );


  not
  g804
  (
    n845,
    n802
  );


  not
  g805
  (
    n860,
    n812
  );


  buf
  g806
  (
    n831,
    n786
  );


  buf
  g807
  (
    n859,
    n809
  );


  buf
  g808
  (
    n847,
    n779
  );


  not
  g809
  (
    n858,
    n804
  );


  not
  g810
  (
    n838,
    n784
  );


  buf
  g811
  (
    n842,
    n814
  );


  not
  g812
  (
    n851,
    n782
  );


  not
  g813
  (
    n865,
    n797
  );


  not
  g814
  (
    n850,
    n801
  );


  buf
  g815
  (
    n829,
    n803
  );


  buf
  g816
  (
    n832,
    n798
  );


  or
  g817
  (
    n874,
    n357,
    n728,
    n351,
    n835
  );


  or
  g818
  (
    n879,
    n735,
    n834,
    n728,
    n357
  );


  and
  g819
  (
    n881,
    n833,
    n729,
    n835,
    n346
  );


  xor
  g820
  (
    n884,
    n830,
    n359,
    n352,
    n828
  );


  nand
  g821
  (
    n891,
    n345,
    n356,
    n351,
    n359
  );


  xor
  g822
  (
    n887,
    n354,
    n358,
    n735,
    n350
  );


  xnor
  g823
  (
    n897,
    n830,
    n350,
    n829,
    n727
  );


  or
  g824
  (
    n885,
    n827,
    n737,
    n835,
    n344
  );


  nand
  g825
  (
    n873,
    n731,
    n354,
    n347,
    n828
  );


  and
  g826
  (
    n867,
    n346,
    n359,
    n356,
    n832
  );


  or
  g827
  (
    n868,
    n358,
    n354,
    n730,
    n345
  );


  or
  g828
  (
    n892,
    n732,
    n350,
    n829,
    n349
  );


  and
  g829
  (
    n895,
    n354,
    n345,
    n831,
    n827
  );


  nand
  g830
  (
    n889,
    n832,
    n736,
    n353,
    n348
  );


  xnor
  g831
  (
    n903,
    n357,
    n726,
    n832,
    n731
  );


  xnor
  g832
  (
    n871,
    n731,
    n360,
    n733,
    n348
  );


  xor
  g833
  (
    n902,
    n730,
    n355,
    n835,
    n736
  );


  and
  g834
  (
    n898,
    n355,
    n729,
    n347,
    n344
  );


  nor
  g835
  (
    n894,
    n730,
    n346,
    n359,
    n352
  );


  or
  g836
  (
    n882,
    n348,
    n347,
    n725,
    n352
  );


  nor
  g837
  (
    n875,
    n358,
    n831,
    n736,
    n353
  );


  nor
  g838
  (
    n901,
    n731,
    n733,
    n732,
    n349
  );


  or
  g839
  (
    n872,
    n829,
    n831,
    n836,
    n832
  );


  and
  g840
  (
    n878,
    n349,
    n833,
    n734,
    n737
  );


  xor
  g841
  (
    n888,
    n831,
    n349,
    n830,
    n356
  );


  xor
  g842
  (
    n869,
    n351,
    n346,
    n828,
    n734
  );


  and
  g843
  (
    n890,
    n732,
    n727,
    n726,
    n350
  );


  and
  g844
  (
    n883,
    n358,
    n353,
    n828,
    n356
  );


  and
  g845
  (
    KeyWire_0_29,
    n728,
    n732,
    n736,
    n737
  );


  nand
  g846
  (
    n876,
    n728,
    n352,
    n733,
    n730
  );


  nor
  g847
  (
    n896,
    n357,
    n351,
    n834
  );


  and
  g848
  (
    n886,
    n345,
    n347,
    n348,
    n735
  );


  xor
  g849
  (
    n893,
    n833,
    n353,
    n727,
    n735
  );


  nor
  g850
  (
    n900,
    n729,
    n733,
    n726,
    n827
  );


  and
  g851
  (
    n870,
    n827,
    n830,
    n734,
    n355
  );


  xor
  g852
  (
    n880,
    n834,
    n833,
    n734,
    n727
  );


  xnor
  g853
  (
    n877,
    n355,
    n729,
    n726,
    n829
  );


  nand
  g854
  (
    n924,
    n676,
    n509,
    n514,
    n675
  );


  nor
  g855
  (
    n926,
    n509,
    n514,
    n506,
    n513
  );


  and
  g856
  (
    n910,
    n867,
    n870,
    n884,
    n883
  );


  or
  g857
  (
    KeyWire_0_48,
    n673,
    n675,
    n515
  );


  nand
  g858
  (
    n904,
    n673,
    n507,
    n747,
    n504
  );


  xnor
  g859
  (
    n925,
    n882,
    n508,
    n515,
    n881
  );


  nor
  g860
  (
    n918,
    n872,
    n507,
    n675,
    n513
  );


  or
  g861
  (
    n911,
    n504,
    n514,
    n505,
    n511
  );


  nand
  g862
  (
    n909,
    n507,
    n746,
    n888,
    n513
  );


  and
  g863
  (
    n913,
    n516,
    n512,
    n509,
    n505
  );


  xnor
  g864
  (
    n906,
    n506,
    n674,
    n876,
    n516
  );


  or
  g865
  (
    n916,
    n516,
    n508,
    n512
  );


  nand
  g866
  (
    n905,
    n511,
    n874,
    n506,
    n877
  );


  xnor
  g867
  (
    n907,
    n510,
    n674,
    n673,
    n509
  );


  xnor
  g868
  (
    n921,
    n505,
    n885,
    n676,
    n504
  );


  nor
  g869
  (
    n914,
    n869,
    n513,
    n746,
    n510
  );


  xor
  g870
  (
    n920,
    n507,
    n505,
    n511,
    n871
  );


  nor
  g871
  (
    n908,
    n506,
    n873,
    n889,
    n508
  );


  xor
  g872
  (
    n917,
    n886,
    n676,
    n673,
    n515
  );


  and
  g873
  (
    n915,
    n674,
    n510,
    n880,
    n878
  );


  xnor
  g874
  (
    n923,
    n510,
    n868,
    n875,
    n514
  );


  xor
  g875
  (
    n912,
    n674,
    n887,
    n879,
    n516
  );


  or
  g876
  (
    n919,
    n508,
    n511,
    n512,
    n515
  );


  not
  g877
  (
    KeyWire_0_50,
    n906
  );


  buf
  g878
  (
    n928,
    n904
  );


  buf
  g879
  (
    n927,
    n907
  );


  buf
  g880
  (
    n929,
    n905
  );


  xor
  g881
  (
    n933,
    n929,
    n678,
    n927
  );


  nand
  g882
  (
    n937,
    n928,
    n681,
    n684,
    n738
  );


  xor
  g883
  (
    n941,
    n679,
    n677,
    n682,
    n678
  );


  xnor
  g884
  (
    n934,
    n928,
    n684,
    n680,
    n678
  );


  xor
  g885
  (
    n939,
    n682,
    n928,
    n683,
    n930
  );


  nor
  g886
  (
    n940,
    n679,
    n677,
    n684,
    n685
  );


  xor
  g887
  (
    n931,
    n677,
    n738,
    n927,
    n685
  );


  xnor
  g888
  (
    n942,
    n738,
    n683,
    n928,
    n680
  );


  nor
  g889
  (
    n936,
    n929,
    n684,
    n677,
    n681
  );


  nand
  g890
  (
    n943,
    n927,
    n683,
    n676
  );


  xor
  g891
  (
    n935,
    n685,
    n681,
    n680
  );


  and
  g892
  (
    n944,
    n738,
    n679,
    n682
  );


  and
  g893
  (
    n932,
    n681,
    n678,
    n685,
    n929
  );


  nand
  g894
  (
    n938,
    n929,
    n737,
    n679,
    n930
  );


  nor
  g895
  (
    n985,
    n936,
    n849,
    n943,
    n939
  );


  nor
  g896
  (
    n973,
    n450,
    n750,
    n850,
    n853
  );


  xor
  g897
  (
    n984,
    n449,
    n942,
    n750,
    n933
  );


  xnor
  g898
  (
    n949,
    n855,
    n851,
    n861,
    n838
  );


  xnor
  g899
  (
    n974,
    n862,
    n943,
    n838,
    n748
  );


  nand
  g900
  (
    n980,
    n846,
    n863,
    n855,
    n836
  );


  xor
  g901
  (
    n991,
    n850,
    n849,
    n843,
    n752
  );


  nor
  g902
  (
    n961,
    n940,
    n751,
    n840,
    n857
  );


  or
  g903
  (
    n950,
    n858,
    n863,
    n852,
    n854
  );


  or
  g904
  (
    KeyWire_0_17,
    n944,
    n856,
    n840,
    n450
  );


  xnor
  g905
  (
    n955,
    n860,
    n855,
    n857
  );


  or
  g906
  (
    n953,
    n942,
    n848,
    n847,
    n861
  );


  xnor
  g907
  (
    n946,
    n940,
    n753,
    n942,
    n748
  );


  and
  g908
  (
    n959,
    n838,
    n858,
    n932,
    n939
  );


  or
  g909
  (
    n947,
    n845,
    n837,
    n451
  );


  and
  g910
  (
    n945,
    n839,
    n939,
    n450,
    n862
  );


  or
  g911
  (
    n970,
    n843,
    n938,
    n839,
    n935
  );


  nor
  g912
  (
    n957,
    n941,
    n853,
    n852,
    n943
  );


  xnor
  g913
  (
    n951,
    n934,
    n937,
    n854,
    n842
  );


  xor
  g914
  (
    n983,
    n854,
    n842,
    n843,
    n856
  );


  nand
  g915
  (
    n981,
    n847,
    n937,
    n846,
    n856
  );


  and
  g916
  (
    n978,
    n931,
    n842,
    n751,
    n836
  );


  xnor
  g917
  (
    n987,
    n939,
    n940,
    n847,
    n942
  );


  or
  g918
  (
    n977,
    n941,
    n842,
    n850,
    n852
  );


  nand
  g919
  (
    n965,
    n859,
    n861,
    n837,
    n844
  );


  nor
  g920
  (
    n969,
    n747,
    n748,
    n941
  );


  or
  g921
  (
    n976,
    n862,
    n844,
    n449,
    n849
  );


  nor
  g922
  (
    n967,
    n936,
    n750,
    n853,
    n851
  );


  xor
  g923
  (
    n954,
    n451,
    n938,
    n936,
    n838
  );


  xor
  g924
  (
    n966,
    n860,
    n848,
    n934,
    n935
  );


  or
  g925
  (
    n990,
    n840,
    n944,
    n860,
    n751
  );


  or
  g926
  (
    n958,
    n848,
    n858,
    n938,
    n937
  );


  xnor
  g927
  (
    n975,
    n860,
    n837,
    n849,
    n749
  );


  xnor
  g928
  (
    n972,
    n859,
    n846,
    n839,
    n844
  );


  nor
  g929
  (
    n962,
    n839,
    n859,
    n938,
    n941
  );


  or
  g930
  (
    n979,
    n852,
    n940,
    n848,
    n836
  );


  nor
  g931
  (
    n992,
    n857,
    n935,
    n747,
    n851
  );


  nor
  g932
  (
    n948,
    n935,
    n861,
    n854,
    n840
  );


  or
  g933
  (
    n952,
    n844,
    n752,
    n845,
    n751
  );


  or
  g934
  (
    n968,
    n862,
    n846,
    n934,
    n841
  );


  and
  g935
  (
    n964,
    n841,
    n752,
    n845,
    n855
  );


  nor
  g936
  (
    n988,
    n863,
    n937,
    n944,
    n943
  );


  nand
  g937
  (
    n963,
    n859,
    n863,
    n845,
    n856
  );


  nor
  g938
  (
    n986,
    n847,
    n841,
    n449,
    n858
  );


  or
  g939
  (
    n971,
    n850,
    n853,
    n933,
    n851
  );


  nor
  g940
  (
    n956,
    n450,
    n936,
    n747,
    n750
  );


  and
  g941
  (
    n989,
    n934,
    n749,
    n944
  );


  nand
  g942
  (
    n982,
    n841,
    n843,
    n749,
    n752
  );


  buf
  g943
  (
    n995,
    n945
  );


  buf
  g944
  (
    n996,
    n945
  );


  not
  g945
  (
    n994,
    n945
  );


  buf
  g946
  (
    n993,
    n945
  );


  buf
  g947
  (
    n1003,
    n993
  );


  not
  g948
  (
    n1002,
    n755
  );


  buf
  g949
  (
    KeyWire_0_26,
    n994
  );


  buf
  g950
  (
    n1009,
    n756
  );


  buf
  g951
  (
    n1000,
    n994
  );


  buf
  g952
  (
    n998,
    n996
  );


  not
  g953
  (
    n1008,
    n946
  );


  or
  g954
  (
    n1010,
    n757,
    n994,
    n995
  );


  xnor
  g955
  (
    n1007,
    n758,
    n946,
    n755
  );


  nor
  g956
  (
    n1001,
    n757,
    n993,
    n995,
    n996
  );


  nor
  g957
  (
    n1011,
    n754,
    n756,
    n758,
    n947
  );


  nand
  g958
  (
    n997,
    n946,
    n995,
    n754,
    n996
  );


  nand
  g959
  (
    n1004,
    n753,
    n756
  );


  xor
  g960
  (
    n999,
    n755,
    n993,
    n996
  );


  and
  g961
  (
    n1005,
    n757,
    n754,
    n753
  );


  xor
  g962
  (
    n1006,
    n758,
    n995,
    n757,
    n755
  );


  nand
  g963
  (
    n1026,
    n687,
    n690,
    n1002,
    n692
  );


  xnor
  g964
  (
    n1024,
    n689,
    n686,
    n1003,
    n688
  );


  nor
  g965
  (
    n1022,
    n689,
    n692,
    n997,
    n691
  );


  nor
  g966
  (
    n1020,
    n998,
    n692,
    n688,
    n999
  );


  or
  g967
  (
    n1023,
    n1001,
    n689,
    n694,
    n1002
  );


  or
  g968
  (
    n1021,
    n693,
    n693,
    n686,
    n998
  );


  or
  g969
  (
    n1027,
    n1000,
    n687,
    n1001,
    n999
  );


  nand
  g970
  (
    n1015,
    n690,
    n686,
    n692,
    n688
  );


  and
  g971
  (
    n1019,
    n999,
    n997,
    n694
  );


  and
  g972
  (
    n1013,
    n689,
    n690,
    n693,
    n687
  );


  xnor
  g973
  (
    n1014,
    n1000,
    n1002,
    n691
  );


  nor
  g974
  (
    n1018,
    n690,
    n999,
    n1004,
    n691
  );


  or
  g975
  (
    n1017,
    n1002,
    n686,
    n694,
    n1003
  );


  xor
  g976
  (
    n1016,
    n693,
    n1003,
    n997,
    n1001
  );


  xor
  g977
  (
    n1028,
    n998,
    n688,
    n1000,
    n1003
  );


  xor
  g978
  (
    n1025,
    n1000,
    n687,
    n1001,
    n998
  );


  not
  g979
  (
    n1029,
    n1025
  );


  buf
  g980
  (
    n1035,
    n1027
  );


  buf
  g981
  (
    n1040,
    n1025
  );


  not
  g982
  (
    n1055,
    n1028
  );


  not
  g983
  (
    n1054,
    n1013
  );


  not
  g984
  (
    n1056,
    n1019
  );


  buf
  g985
  (
    n1038,
    n1019
  );


  not
  g986
  (
    n1043,
    n1018
  );


  buf
  g987
  (
    n1031,
    n1023
  );


  not
  g988
  (
    n1046,
    n1016
  );


  buf
  g989
  (
    n1033,
    n1017
  );


  not
  g990
  (
    n1036,
    n1017
  );


  buf
  g991
  (
    n1039,
    n1022
  );


  buf
  g992
  (
    n1041,
    n1020
  );


  buf
  g993
  (
    n1044,
    n1026
  );


  buf
  g994
  (
    n1047,
    n1027
  );


  not
  g995
  (
    n1045,
    n1018
  );


  buf
  g996
  (
    n1048,
    n1015
  );


  buf
  g997
  (
    n1050,
    n1028
  );


  not
  g998
  (
    n1032,
    n1020
  );


  buf
  g999
  (
    n1030,
    n1026
  );


  buf
  g1000
  (
    n1049,
    n1024
  );


  not
  g1001
  (
    n1052,
    n1014
  );


  buf
  g1002
  (
    n1037,
    n1021
  );


  buf
  g1003
  (
    n1034,
    n1021
  );


  buf
  g1004
  (
    n1051,
    n1023
  );


  not
  g1005
  (
    n1053,
    n1022
  );


  not
  g1006
  (
    n1042,
    n1024
  );


  not
  g1007
  (
    n1060,
    n739
  );


  buf
  g1008
  (
    n1065,
    n740
  );


  not
  g1009
  (
    n1062,
    n740
  );


  buf
  g1010
  (
    n1059,
    n739
  );


  not
  g1011
  (
    n1061,
    n1030
  );


  not
  g1012
  (
    n1057,
    n1031
  );


  buf
  g1013
  (
    n1064,
    n1030
  );


  nand
  g1014
  (
    n1058,
    n1030,
    n739,
    n1029
  );


  xnor
  g1015
  (
    n1063,
    n739,
    n1029,
    n1030
  );


  xor
  g1016
  (
    n1067,
    n1057,
    n760
  );


  xor
  g1017
  (
    n1070,
    n760,
    n759
  );


  or
  g1018
  (
    n1066,
    n1031,
    n1057
  );


  xor
  g1019
  (
    n1068,
    n1057,
    n759
  );


  nand
  g1020
  (
    n1069,
    n758,
    n760,
    n1058
  );


  buf
  g1021
  (
    n1071,
    n1067
  );


  not
  g1022
  (
    n1077,
    n1066
  );


  buf
  g1023
  (
    n1074,
    n1068
  );


  buf
  g1024
  (
    n1073,
    n1070
  );


  not
  g1025
  (
    n1078,
    n1070
  );


  buf
  g1026
  (
    n1076,
    n1070
  );


  not
  g1027
  (
    n1075,
    n1069
  );


  buf
  g1028
  (
    n1072,
    n1070
  );


  and
  g1029
  (
    n1083,
    n948,
    n950,
    n951,
    n949
  );


  xor
  g1030
  (
    n1079,
    n1072,
    n951,
    n1075,
    n1073
  );


  and
  g1031
  (
    n1088,
    n947,
    n1074,
    n952,
    n1072
  );


  nor
  g1032
  (
    n1086,
    n947,
    n948,
    n950,
    n1071
  );


  nor
  g1033
  (
    n1084,
    n948,
    n1071,
    n1075,
    n951
  );


  nor
  g1034
  (
    n1081,
    n1071,
    n949,
    n1072
  );


  nor
  g1035
  (
    n1085,
    n1071,
    n1074,
    n952,
    n1073
  );


  or
  g1036
  (
    n1080,
    n948,
    n952,
    n947,
    n949
  );


  xnor
  g1037
  (
    n1082,
    n1072,
    n1073,
    n950
  );


  nor
  g1038
  (
    n1087,
    n1073,
    n1074,
    n951
  );


  buf
  g1039
  (
    n1092,
    n1059
  );


  buf
  g1040
  (
    n1096,
    n1059
  );


  not
  g1041
  (
    n1093,
    n1059
  );


  not
  g1042
  (
    n1095,
    n1083
  );


  not
  g1043
  (
    n1089,
    n1058
  );


  nor
  g1044
  (
    n1094,
    n1084,
    n1058,
    n1060,
    n1088
  );


  xnor
  g1045
  (
    n1090,
    n1058,
    n1086,
    n1085,
    n1087
  );


  and
  g1046
  (
    n1091,
    n1081,
    n1082,
    n1059,
    n1031
  );


  buf
  g1047
  (
    n1106,
    n959
  );


  or
  g1048
  (
    n1101,
    n1090,
    n959,
    n952
  );


  or
  g1049
  (
    n1111,
    n957,
    n1092,
    n956
  );


  xnor
  g1050
  (
    n1098,
    n955,
    n954
  );


  xor
  g1051
  (
    n1099,
    n953,
    n958,
    n956
  );


  and
  g1052
  (
    n1102,
    n1089,
    n1092
  );


  nor
  g1053
  (
    n1112,
    n1092,
    n954,
    n955
  );


  and
  g1054
  (
    n1105,
    n956,
    n1091,
    n959
  );


  xor
  g1055
  (
    n1103,
    n1090,
    n958,
    n1091
  );


  and
  g1056
  (
    n1110,
    n957,
    n958,
    n960
  );


  nand
  g1057
  (
    n1104,
    n1089,
    n1091,
    n1090
  );


  xor
  g1058
  (
    n1109,
    n1090,
    n953,
    n956
  );


  or
  g1059
  (
    n1097,
    n958,
    n953,
    n1089
  );


  nand
  g1060
  (
    n1107,
    n954,
    n1089,
    n957
  );


  nand
  g1061
  (
    n1100,
    n955,
    n957,
    n1091
  );


  nor
  g1062
  (
    n1108,
    n955,
    n959,
    n953
  );


  xnor
  g1063
  (
    n1113,
    n1097,
    n360
  );


  not
  g1064
  (
    n1116,
    n1113
  );


  not
  g1065
  (
    n1114,
    n1113
  );


  buf
  g1066
  (
    n1115,
    n1113
  );


  buf
  g1067
  (
    n1117,
    n1113
  );


  buf
  g1068
  (
    n1118,
    n1114
  );


  buf
  g1069
  (
    n1126,
    n1116
  );


  buf
  g1070
  (
    n1123,
    n1116
  );


  not
  g1071
  (
    n1128,
    n1114
  );


  not
  g1072
  (
    n1120,
    n1115
  );


  not
  g1073
  (
    n1125,
    n1115
  );


  not
  g1074
  (
    n1130,
    n1116
  );


  buf
  g1075
  (
    n1124,
    n1114
  );


  buf
  g1076
  (
    n1129,
    n1116
  );


  not
  g1077
  (
    n1119,
    n1115
  );


  not
  g1078
  (
    n1127,
    n1117
  );


  buf
  g1079
  (
    n1121,
    n1114
  );


  buf
  g1080
  (
    n1122,
    n1115
  );


  xor
  g1081
  (
    n1169,
    n975,
    n1130,
    n1048,
    n1128
  );


  nor
  g1082
  (
    n1131,
    n970,
    n963,
    n1043,
    n974
  );


  nand
  g1083
  (
    n1159,
    n1033,
    n964,
    n1128,
    n963
  );


  nand
  g1084
  (
    n1141,
    n1045,
    n967,
    n1119,
    n1036
  );


  xor
  g1085
  (
    n1144,
    n1040,
    n1035,
    n1125,
    n1037
  );


  nor
  g1086
  (
    n1149,
    n969,
    n971,
    n1124
  );


  nor
  g1087
  (
    n1152,
    n961,
    n1039,
    n1035,
    n1119
  );


  nand
  g1088
  (
    n1174,
    n1126,
    n961,
    n1037,
    n1123
  );


  and
  g1089
  (
    n1146,
    n960,
    n1042,
    n1122,
    n1129
  );


  nand
  g1090
  (
    n1135,
    n1035,
    n1125,
    n1043,
    n965
  );


  xnor
  g1091
  (
    n1163,
    n964,
    n972,
    n1047,
    n1032
  );


  nand
  g1092
  (
    n1148,
    n970,
    n1032,
    n967,
    n1039
  );


  or
  g1093
  (
    n1171,
    n1032,
    n1041,
    n969,
    n1130
  );


  xnor
  g1094
  (
    KeyWire_0_1,
    n975,
    n1048,
    n968
  );


  nand
  g1095
  (
    n1170,
    n1121,
    n974,
    n1126,
    n1124
  );


  nand
  g1096
  (
    n1132,
    n1034,
    n1042,
    n1125,
    n969
  );


  or
  g1097
  (
    n1158,
    n1129,
    n970,
    n960,
    n1047
  );


  xor
  g1098
  (
    n1167,
    n970,
    n1129,
    n1036,
    n1034
  );


  or
  g1099
  (
    n1175,
    n1043,
    n975,
    n964,
    n962
  );


  nor
  g1100
  (
    n1164,
    n1042,
    n1038,
    n1044,
    n1118
  );


  or
  g1101
  (
    n1150,
    n1038,
    n1124,
    n975,
    n967
  );


  xor
  g1102
  (
    n1168,
    n1125,
    n1033,
    n1046,
    n1123
  );


  xnor
  g1103
  (
    KeyWire_0_47,
    n965,
    n973,
    n974,
    n966
  );


  xor
  g1104
  (
    n1147,
    n968,
    n1129,
    n962,
    n973
  );


  xnor
  g1105
  (
    n1145,
    n966,
    n1040,
    n1044,
    n1038
  );


  nand
  g1106
  (
    n1157,
    n965,
    n1127,
    n1038
  );


  xnor
  g1107
  (
    n1153,
    n1043,
    n966,
    n1121
  );


  and
  g1108
  (
    n1133,
    n964,
    n967,
    n1049,
    n962
  );


  nor
  g1109
  (
    n1143,
    n1039,
    n972,
    n1122
  );


  xnor
  g1110
  (
    n1160,
    n1041,
    n1033,
    n971,
    n1046
  );


  and
  g1111
  (
    n1156,
    n976,
    n1046,
    n963,
    n1041
  );


  xnor
  g1112
  (
    n1162,
    n973,
    n1126,
    n1122,
    n1034
  );


  xor
  g1113
  (
    n1154,
    n1034,
    n1035,
    n1036,
    n965
  );


  and
  g1114
  (
    n1151,
    n974,
    n1120,
    n972,
    n1040
  );


  xnor
  g1115
  (
    n1134,
    n1126,
    n969,
    n1036,
    n1039
  );


  xor
  g1116
  (
    n1173,
    n1033,
    n1031,
    n1037,
    n1121
  );


  xor
  g1117
  (
    n1166,
    n961,
    n1127,
    n1130,
    n1032
  );


  and
  g1118
  (
    n1137,
    n961,
    n1120,
    n1121,
    n1044
  );


  nor
  g1119
  (
    n1140,
    n960,
    n1045,
    n971
  );


  nand
  g1120
  (
    n1142,
    n1037,
    n973,
    n1128,
    n1127
  );


  or
  g1121
  (
    n1139,
    n968,
    n1123,
    n1128,
    n1042
  );


  nand
  g1122
  (
    n1172,
    n968,
    n1123,
    n1047,
    n1045
  );


  nand
  g1123
  (
    n1155,
    n1122,
    n1040,
    n1046,
    n1044
  );


  and
  g1124
  (
    n1136,
    n976,
    n1124,
    n1130,
    n963
  );


  xnor
  g1125
  (
    n1165,
    n1048,
    n1041,
    n1047,
    n962
  );


  not
  g1126
  (
    n1179,
    n1061
  );


  buf
  g1127
  (
    n1177,
    n1061
  );


  xor
  g1128
  (
    n1178,
    n1060,
    n1131,
    n1061
  );


  nor
  g1129
  (
    KeyWire_0_43,
    n1131,
    n1060
  );


  or
  g1130
  (
    n1192,
    n1005,
    n1177,
    n1007,
    n1008
  );


  nand
  g1131
  (
    n1187,
    n978,
    n976,
    n979,
    n1010
  );


  and
  g1132
  (
    n1185,
    n1176,
    n1179,
    n1007,
    n1004
  );


  and
  g1133
  (
    n1194,
    n1009,
    n1004,
    n1005,
    n1010
  );


  xnor
  g1134
  (
    n1186,
    n1008,
    n1006,
    n1010,
    n1009
  );


  nor
  g1135
  (
    n1193,
    n1007,
    n977,
    n1006
  );


  or
  g1136
  (
    n1184,
    n976,
    n1177,
    n1005
  );


  nand
  g1137
  (
    n1190,
    n1178,
    n1177,
    n1179,
    n978
  );


  and
  g1138
  (
    n1191,
    n979,
    n978,
    n1179,
    n1006
  );


  nor
  g1139
  (
    n1181,
    n1010,
    n977,
    n1176,
    n1009
  );


  or
  g1140
  (
    n1180,
    n1177,
    n1011,
    n977,
    n979
  );


  xnor
  g1141
  (
    n1183,
    n1008,
    n1011,
    n1178
  );


  xor
  g1142
  (
    n1189,
    n1004,
    n979,
    n1178,
    n1176
  );


  nand
  g1143
  (
    n1188,
    n1006,
    n1179,
    n1011
  );


  and
  g1144
  (
    n1182,
    n1008,
    n978,
    n1009,
    n1007
  );


  buf
  g1145
  (
    n1195,
    n1180
  );


  not
  g1146
  (
    n1196,
    n1195
  );


  buf
  g1147
  (
    n1197,
    n1195
  );


  not
  g1148
  (
    n1198,
    n1196
  );


  not
  g1149
  (
    n1200,
    n1198
  );


  buf
  g1150
  (
    n1199,
    n1198
  );


  and
  g1151
  (
    n1207,
    n1182,
    n1200,
    n1180
  );


  nor
  g1152
  (
    n1205,
    n1181,
    n1183,
    n1200
  );


  xnor
  g1153
  (
    n1202,
    n1182,
    n1075,
    n1181,
    n1183
  );


  and
  g1154
  (
    n1203,
    n1076,
    n1076,
    n1183,
    n1182
  );


  nand
  g1155
  (
    n1201,
    n1182,
    n1077,
    n1181,
    n1199
  );


  xnor
  g1156
  (
    n1208,
    n1076,
    n1076,
    n1199,
    n1200
  );


  nand
  g1157
  (
    n1206,
    n1181,
    n1075,
    n1077
  );


  xnor
  g1158
  (
    n1204,
    n1180,
    n1200,
    n1199
  );


  and
  g1159
  (
    n1218,
    n1204,
    n1195,
    n1202,
    n1205
  );


  and
  g1160
  (
    n1219,
    n1203,
    n1061,
    n821,
    n826
  );


  nand
  g1161
  (
    n1217,
    n825,
    n818,
    n1202,
    n821
  );


  and
  g1162
  (
    n1225,
    n818,
    n1203,
    n817,
    n820
  );


  or
  g1163
  (
    n1220,
    n823,
    n1202,
    n817,
    n1203
  );


  nor
  g1164
  (
    n1224,
    n1205,
    n815,
    n822,
    n824
  );


  nor
  g1165
  (
    n1215,
    n822,
    n1201,
    n823
  );


  and
  g1166
  (
    n1214,
    n1201,
    n1204,
    n820
  );


  xor
  g1167
  (
    n1212,
    n826,
    n816,
    n1206
  );


  nand
  g1168
  (
    n1222,
    n1201,
    n816,
    n47,
    n824
  );


  xnor
  g1169
  (
    n1213,
    n824,
    n823,
    n822
  );


  nor
  g1170
  (
    n1211,
    n816,
    n817,
    n819,
    n1205
  );


  xor
  g1171
  (
    n1221,
    n1203,
    n825,
    n819,
    n1205
  );


  xor
  g1172
  (
    n1209,
    n815,
    n818,
    n821
  );


  nor
  g1173
  (
    n1223,
    n817,
    n820,
    n819
  );


  nand
  g1174
  (
    n1216,
    n816,
    n825,
    n1195,
    n819
  );


  xor
  g1175
  (
    n1226,
    n822,
    n818,
    n815,
    n825
  );


  and
  g1176
  (
    n1227,
    n826,
    n826,
    n1117,
    n1202
  );


  nand
  g1177
  (
    n1210,
    n1204,
    n1117,
    n824
  );


  not
  g1178
  (
    n1255,
    n1226
  );


  not
  g1179
  (
    n1240,
    n1223
  );


  not
  g1180
  (
    n1237,
    n1216
  );


  buf
  g1181
  (
    n1261,
    n86
  );


  not
  g1182
  (
    n1253,
    n1078
  );


  not
  g1183
  (
    n1256,
    n87
  );


  not
  g1184
  (
    n1238,
    n1093
  );


  buf
  g1185
  (
    n1266,
    n1209
  );


  buf
  g1186
  (
    n1233,
    n1226
  );


  buf
  g1187
  (
    n1247,
    n1214
  );


  not
  g1188
  (
    n1252,
    n1218
  );


  not
  g1189
  (
    n1262,
    n1210
  );


  buf
  g1190
  (
    n1265,
    n1226
  );


  not
  g1191
  (
    n1246,
    n85
  );


  buf
  g1192
  (
    n1268,
    n1209
  );


  buf
  g1193
  (
    n1229,
    n1221
  );


  not
  g1194
  (
    n1254,
    n1216
  );


  not
  g1195
  (
    n1245,
    n1078
  );


  buf
  g1196
  (
    n1264,
    n86
  );


  not
  g1197
  (
    n1239,
    n1219
  );


  not
  g1198
  (
    n1234,
    n1220
  );


  buf
  g1199
  (
    n1236,
    n1227
  );


  buf
  g1200
  (
    n1258,
    n1213
  );


  not
  g1201
  (
    n1250,
    n361
  );


  buf
  g1202
  (
    n1249,
    n1225
  );


  not
  g1203
  (
    n1241,
    n1226
  );


  not
  g1204
  (
    n1269,
    n1213
  );


  not
  g1205
  (
    n1260,
    n86
  );


  buf
  g1206
  (
    n1263,
    n1215
  );


  not
  g1207
  (
    n1228,
    n1211
  );


  not
  g1208
  (
    n1257,
    n1196
  );


  not
  g1209
  (
    n1232,
    n84
  );


  xnor
  g1210
  (
    n1231,
    n1211,
    n1220,
    n87
  );


  nand
  g1211
  (
    n1248,
    n1212,
    n1077,
    n87
  );


  xor
  g1212
  (
    n1242,
    n87,
    n1227,
    n1218
  );


  or
  g1213
  (
    n1259,
    n1214,
    n85,
    n1217
  );


  xor
  g1214
  (
    n1243,
    n1225,
    n1227,
    n1222
  );


  xor
  g1215
  (
    n1244,
    n1217,
    n1222,
    n1078
  );


  or
  g1216
  (
    n1235,
    n1224,
    n1212,
    n1210
  );


  and
  g1217
  (
    n1267,
    n1227,
    n1223,
    n1224
  );


  and
  g1218
  (
    n1230,
    n1215,
    n85
  );


  xnor
  g1219
  (
    n1251,
    n1221,
    n86,
    n1219
  );


  nand
  g1220
  (
    n1426,
    n471,
    n1099,
    n453,
    n1252
  );


  xor
  g1221
  (
    n1383,
    n1249,
    n1151,
    n1231,
    n462
  );


  xnor
  g1222
  (
    n1382,
    n1167,
    n902,
    n1160,
    n615
  );


  xnor
  g1223
  (
    n1290,
    n1265,
    n1245,
    n1263,
    n1189
  );


  or
  g1224
  (
    n1367,
    n472,
    n1100,
    n1170,
    n1103
  );


  nor
  g1225
  (
    n1423,
    n1232,
    n1245,
    n1266,
    n1152
  );


  nand
  g1226
  (
    n1340,
    n457,
    n467,
    n1188,
    n1193
  );


  nor
  g1227
  (
    n1334,
    n1162,
    n1140,
    n472,
    n1151
  );


  nor
  g1228
  (
    n1387,
    n1144,
    n482,
    n457,
    n470
  );


  or
  g1229
  (
    n1316,
    n1148,
    n457,
    n1266,
    n1259
  );


  and
  g1230
  (
    n1338,
    n1163,
    n470,
    n473,
    n1256
  );


  nor
  g1231
  (
    n1434,
    n1111,
    n1167,
    n477,
    n484
  );


  nor
  g1232
  (
    n1366,
    n473,
    n469,
    n624,
    n1194
  );


  or
  g1233
  (
    KeyWire_0_10,
    n1145,
    n474,
    n1110,
    n1267
  );


  xor
  g1234
  (
    n1302,
    n470,
    n1260,
    n1261,
    n475
  );


  nand
  g1235
  (
    n1325,
    n1243,
    n892,
    n1108,
    n864
  );


  xnor
  g1236
  (
    n1371,
    n459,
    n1147,
    n629,
    n452
  );


  nor
  g1237
  (
    n1359,
    n1187,
    n483,
    n1256,
    n1191
  );


  xnor
  g1238
  (
    n1411,
    n477,
    n107,
    n1230,
    n1146
  );


  and
  g1239
  (
    n1282,
    n1170,
    n1243,
    n1152,
    n1186
  );


  nand
  g1240
  (
    n1277,
    n461,
    n1184,
    n1154,
    n1147
  );


  nor
  g1241
  (
    n1395,
    n619,
    n1250,
    n622,
    n1135
  );


  and
  g1242
  (
    n1413,
    n617,
    n616,
    n1153,
    n493
  );


  and
  g1243
  (
    n1272,
    n1186,
    n898,
    n1193,
    n479
  );


  xnor
  g1244
  (
    n1410,
    n482,
    n460,
    n1258,
    n484
  );


  xnor
  g1245
  (
    n1375,
    n1163,
    n1265,
    n1246,
    n1151
  );


  and
  g1246
  (
    n1317,
    n618,
    n463,
    n477,
    n1235
  );


  and
  g1247
  (
    n1284,
    n1261,
    n478,
    n1253,
    n481
  );


  or
  g1248
  (
    n1429,
    n1165,
    n1238,
    n1139,
    n1264
  );


  xnor
  g1249
  (
    n1273,
    n1254,
    n1149,
    n899,
    n469
  );


  and
  g1250
  (
    n1418,
    n617,
    n1228,
    n619,
    n1112
  );


  or
  g1251
  (
    n1378,
    n1232,
    n459,
    n1268,
    n463
  );


  xor
  g1252
  (
    n1309,
    n1235,
    n1229,
    n490,
    n1228
  );


  or
  g1253
  (
    n1304,
    n1141,
    n1192,
    n1245,
    n1171
  );


  nand
  g1254
  (
    n1271,
    n463,
    n903,
    n1150,
    n1133
  );


  or
  g1255
  (
    n1274,
    n1244,
    n466,
    n616,
    n490
  );


  xnor
  g1256
  (
    n1341,
    n456,
    n627,
    n1159,
    n626
  );


  and
  g1257
  (
    n1335,
    n1158,
    n476,
    n1254,
    n478
  );


  nor
  g1258
  (
    n1360,
    n618,
    n1132,
    n1150,
    n462
  );


  xnor
  g1259
  (
    n1376,
    n457,
    n630,
    n1268,
    n1264
  );


  and
  g1260
  (
    n1403,
    n1193,
    n1160,
    n623,
    n1240
  );


  nor
  g1261
  (
    n1305,
    n1249,
    n618,
    n1132,
    n479
  );


  or
  g1262
  (
    KeyWire_0_7,
    n1240,
    n864,
    n1172,
    n1157
  );


  nand
  g1263
  (
    n1430,
    n1251,
    n1258,
    n460,
    n453
  );


  xnor
  g1264
  (
    n1389,
    n1165,
    n1166,
    n620,
    n454
  );


  nand
  g1265
  (
    n1356,
    n1246,
    n466,
    n1188,
    n451
  );


  xnor
  g1266
  (
    n1422,
    n1241,
    n896,
    n1159,
    n1237
  );


  nor
  g1267
  (
    n1431,
    n453,
    n1169,
    n1163,
    n456
  );


  nand
  g1268
  (
    n1433,
    n454,
    n1269,
    n468,
    n1164
  );


  xor
  g1269
  (
    n1346,
    n466,
    n1187,
    n1168,
    n490
  );


  and
  g1270
  (
    n1286,
    n1233,
    n629,
    n619,
    n487
  );


  xor
  g1271
  (
    n1318,
    n1267,
    n629,
    n487,
    n1165
  );


  and
  g1272
  (
    n1415,
    n1172,
    n890,
    n462,
    n1135
  );


  nor
  g1273
  (
    n1307,
    n1153,
    n1234,
    n459,
    n1239
  );


  nand
  g1274
  (
    n1355,
    n1241,
    n1247,
    n1254,
    n625
  );


  nor
  g1275
  (
    n1347,
    n1257,
    n1156,
    n482,
    n621
  );


  xnor
  g1276
  (
    n1275,
    n455,
    n1229,
    n1244,
    n1241
  );


  or
  g1277
  (
    n1308,
    n475,
    n1134,
    n628,
    n1137
  );


  or
  g1278
  (
    n1285,
    n492,
    n1242,
    n1241,
    n1138
  );


  nand
  g1279
  (
    n1311,
    n1143,
    n470,
    n1232,
    n461
  );


  nand
  g1280
  (
    n1337,
    n1140,
    n1263,
    n107,
    n1192
  );


  nor
  g1281
  (
    n1437,
    n625,
    n1269,
    n1184,
    n1134
  );


  and
  g1282
  (
    n1390,
    n900,
    n1151,
    n1256
  );


  nand
  g1283
  (
    n1419,
    n458,
    n1101,
    n1267,
    n1145
  );


  nand
  g1284
  (
    n1280,
    n1261,
    n466,
    n622,
    n1143
  );


  xor
  g1285
  (
    n1399,
    n1252,
    n478,
    n1078,
    n1262
  );


  or
  g1286
  (
    n1393,
    n494,
    n1172,
    n615,
    n1161
  );


  nand
  g1287
  (
    n1386,
    n901,
    n1156,
    n1251,
    n469
  );


  xor
  g1288
  (
    n1379,
    n1145,
    n1148,
    n628,
    n1268
  );


  and
  g1289
  (
    n1343,
    n456,
    n1135,
    n1138,
    n1142
  );


  xor
  g1290
  (
    n1295,
    n493,
    n1167,
    n1146,
    n616
  );


  nor
  g1291
  (
    n1327,
    n1153,
    n486,
    n1239,
    n893
  );


  nor
  g1292
  (
    n1414,
    n1269,
    n464,
    n1160,
    n1265
  );


  nor
  g1293
  (
    n1402,
    n620,
    n902,
    n1243,
    n1169
  );


  nand
  g1294
  (
    n1345,
    n486,
    n1190,
    n1164,
    n1187
  );


  or
  g1295
  (
    n1372,
    n1158,
    n1154,
    n489,
    n1166
  );


  xor
  g1296
  (
    n1324,
    n1161,
    n630,
    n629,
    n453
  );


  and
  g1297
  (
    n1293,
    n622,
    n464,
    n494,
    n1247
  );


  xor
  g1298
  (
    n1432,
    n484,
    n485,
    n1190,
    n451
  );


  nor
  g1299
  (
    n1373,
    n1236,
    n1146,
    n480,
    n1171
  );


  and
  g1300
  (
    n1336,
    n623,
    n1140,
    n476,
    n1248
  );


  xnor
  g1301
  (
    n1436,
    n626,
    n493,
    n455,
    n468
  );


  or
  g1302
  (
    n1314,
    n494,
    n1233,
    n1238,
    n1246
  );


  nor
  g1303
  (
    n1350,
    n1191,
    n1188,
    n1144,
    n1234
  );


  nand
  g1304
  (
    n1394,
    n1250,
    n902,
    n901,
    n621
  );


  and
  g1305
  (
    n1332,
    n1238,
    n1141,
    n488,
    n483
  );


  xnor
  g1306
  (
    n1369,
    n1133,
    n1192,
    n107,
    n1184
  );


  xor
  g1307
  (
    n1401,
    n476,
    n1150,
    n1156,
    n491
  );


  xor
  g1308
  (
    n1331,
    n489,
    n1262,
    n626,
    n1252
  );


  or
  g1309
  (
    n1270,
    n380,
    n894,
    n1269,
    n1255
  );


  nand
  g1310
  (
    n1385,
    n1267,
    n1185,
    n1194,
    n1161
  );


  xor
  g1311
  (
    n1339,
    n1247,
    n1162,
    n479,
    n895
  );


  xor
  g1312
  (
    n1291,
    n1147,
    n1190,
    n492,
    n1247
  );


  xnor
  g1313
  (
    n1288,
    n1152,
    n483,
    n1250,
    n488
  );


  xnor
  g1314
  (
    n1278,
    n474,
    n492,
    n1186,
    n1169
  );


  or
  g1315
  (
    n1333,
    n493,
    n1230,
    n1264,
    n471
  );


  xor
  g1316
  (
    n1400,
    n1184,
    n468,
    n474,
    n1266
  );


  xnor
  g1317
  (
    n1298,
    n491,
    n1261,
    n458,
    n1112
  );


  nor
  g1318
  (
    n1427,
    n1253,
    n1250,
    n1229,
    n462
  );


  xor
  g1319
  (
    n1276,
    n480,
    n1167,
    n1174,
    n903
  );


  nand
  g1320
  (
    n1299,
    n1242,
    n1186,
    n1136,
    n1158
  );


  nand
  g1321
  (
    n1364,
    n484,
    n472,
    n1141,
    n1257
  );


  nor
  g1322
  (
    n1405,
    n1258,
    n478,
    n455,
    n1172
  );


  nor
  g1323
  (
    n1424,
    n1243,
    n1259,
    n1190,
    n452
  );


  nand
  g1324
  (
    n1416,
    n454,
    n1137,
    n1264,
    n1253
  );


  xnor
  g1325
  (
    n1391,
    n1147,
    n1154,
    n1106,
    n1164
  );


  xnor
  g1326
  (
    n1292,
    n1169,
    n458,
    n1132,
    n461
  );


  or
  g1327
  (
    n1370,
    n1248,
    n1228,
    n1139,
    n1160
  );


  nor
  g1328
  (
    n1396,
    n1254,
    n1153,
    n1253,
    n903
  );


  xor
  g1329
  (
    n1377,
    n458,
    n467,
    n1136,
    n1268
  );


  and
  g1330
  (
    n1363,
    n1242,
    n1109,
    n452,
    n1150
  );


  xnor
  g1331
  (
    n1296,
    n1157,
    n1262,
    n1145,
    n487
  );


  xor
  g1332
  (
    n1421,
    n628,
    n1146,
    n480,
    n621
  );


  nand
  g1333
  (
    n1428,
    n459,
    n380,
    n1136,
    n1234
  );


  nand
  g1334
  (
    n1319,
    n1168,
    n1239,
    n464,
    n1134
  );


  nor
  g1335
  (
    n1279,
    n1171,
    n474,
    n1257,
    n494
  );


  nor
  g1336
  (
    n1328,
    n1133,
    n1132,
    n1236,
    n1260
  );


  and
  g1337
  (
    n1409,
    n1193,
    n618,
    n476,
    n107
  );


  nand
  g1338
  (
    n1281,
    n1142,
    n1166,
    n1148,
    n1171
  );


  or
  g1339
  (
    n1306,
    n489,
    n1255,
    n491,
    n1240
  );


  xor
  g1340
  (
    n1351,
    n1158,
    n1266,
    n1231,
    n1185
  );


  or
  g1341
  (
    n1344,
    n1236,
    n1231,
    n1229,
    n1111
  );


  and
  g1342
  (
    n1408,
    n900,
    n473,
    n1237,
    n1162
  );


  xnor
  g1343
  (
    n1313,
    n1255,
    n485,
    n1230,
    n1244
  );


  or
  g1344
  (
    n1353,
    n1232,
    n1139,
    n480,
    n627
  );


  and
  g1345
  (
    n1388,
    n456,
    n1198,
    n1248,
    n1236
  );


  or
  g1346
  (
    n1374,
    n621,
    n1148,
    n467,
    n463
  );


  nor
  g1347
  (
    n1362,
    n1235,
    n1249,
    n1258
  );


  or
  g1348
  (
    n1380,
    n1105,
    n1107,
    n897,
    n491
  );


  nand
  g1349
  (
    n1354,
    n1166,
    n1263,
    n1159,
    n903
  );


  nor
  g1350
  (
    n1361,
    n864,
    n488,
    n1159,
    n1137
  );


  nor
  g1351
  (
    n1368,
    n1237,
    n465,
    n1173,
    n469
  );


  or
  g1352
  (
    n1406,
    n1263,
    n1138,
    n1157,
    n1233
  );


  and
  g1353
  (
    n1301,
    n1137,
    n1246,
    n1133,
    n1251
  );


  nor
  g1354
  (
    n1297,
    n1149,
    n1162,
    n623,
    n620
  );


  or
  g1355
  (
    n1365,
    n1192,
    n1188,
    n1149,
    n471
  );


  or
  g1356
  (
    n1289,
    n1185,
    n460,
    n1237,
    n1260
  );


  xnor
  g1357
  (
    n1381,
    n1185,
    n1248,
    n492,
    n473
  );


  xnor
  g1358
  (
    n1321,
    n1189,
    n475,
    n864,
    n1102
  );


  nand
  g1359
  (
    n1392,
    n1238,
    n1251,
    n471,
    n630
  );


  and
  g1360
  (
    n1342,
    n455,
    n1155,
    n627,
    n468
  );


  xor
  g1361
  (
    n1287,
    n1187,
    n461,
    n1260,
    n1144
  );


  and
  g1362
  (
    n1294,
    n479,
    n1191,
    n624,
    n1173
  );


  xnor
  g1363
  (
    n1420,
    n1245,
    n1135,
    n1168,
    n486
  );


  xor
  g1364
  (
    n1310,
    n1240,
    n1231,
    n628,
    n1239
  );


  or
  g1365
  (
    n1323,
    n452,
    n481,
    n622,
    n488
  );


  xnor
  g1366
  (
    n1435,
    n625,
    n902,
    n626,
    n485
  );


  or
  g1367
  (
    n1283,
    n1173,
    n1194,
    n481,
    n1161
  );


  or
  g1368
  (
    n1326,
    n1141,
    n1265,
    n465,
    n1164
  );


  xor
  g1369
  (
    n1358,
    n1233,
    n1098,
    n489,
    n1168
  );


  xnor
  g1370
  (
    n1352,
    n1149,
    n630,
    n1191,
    n1257
  );


  xor
  g1371
  (
    n1329,
    n1140,
    n1170,
    n475,
    n482
  );


  and
  g1372
  (
    n1330,
    n1173,
    n464,
    n1242,
    n465
  );


  or
  g1373
  (
    n1398,
    n490,
    n1255,
    n1152,
    n617
  );


  nand
  g1374
  (
    n1300,
    n467,
    n624,
    n1154,
    n1155
  );


  nor
  g1375
  (
    n1322,
    n1136,
    n1189,
    n1139,
    n627
  );


  or
  g1376
  (
    n1357,
    n1142,
    n615,
    n1262,
    n1155
  );


  nand
  g1377
  (
    n1425,
    n1198,
    n1155,
    n1244,
    n472
  );


  xor
  g1378
  (
    n1404,
    n891,
    n619,
    n623,
    n1194
  );


  and
  g1379
  (
    n1412,
    n1163,
    n454,
    n1104,
    n460
  );


  and
  g1380
  (
    n1407,
    n1144,
    n1170,
    n481,
    n477
  );


  xnor
  g1381
  (
    n1384,
    n625,
    n1230,
    n620,
    n624
  );


  nor
  g1382
  (
    n1312,
    n485,
    n1234,
    n1259,
    n487
  );


  nand
  g1383
  (
    n1348,
    n486,
    n1189,
    n1228,
    n1143
  );


  and
  g1384
  (
    n1320,
    n483,
    n1165,
    n1134,
    n1157
  );


  xor
  g1385
  (
    n1349,
    n465,
    n1235,
    n1252,
    n1110
  );


  and
  g1386
  (
    n1303,
    n1138,
    n615,
    n1142,
    n1156
  );


  xor
  g1387
  (
    n1397,
    n1259,
    n616,
    n1143,
    n617
  );


  nor
  g1388
  (
    n1626,
    n697,
    n696,
    n1270,
    n524
  );


  nor
  g1389
  (
    n1566,
    n1317,
    n1339,
    n1387,
    n1398
  );


  and
  g1390
  (
    n1466,
    n1365,
    n560,
    n581,
    n554
  );


  or
  g1391
  (
    n1438,
    n1271,
    n1344,
    n554,
    n582
  );


  xnor
  g1392
  (
    n1511,
    n542,
    n580,
    n523,
    n714
  );


  nand
  g1393
  (
    n1523,
    n1347,
    n1380,
    n529,
    n592
  );


  xnor
  g1394
  (
    n1526,
    n1358,
    n1429,
    n1314,
    n1093
  );


  xnor
  g1395
  (
    n1674,
    n574,
    n569,
    n1345,
    n1279
  );


  nor
  g1396
  (
    KeyWire_0_45,
    n567,
    n1274,
    n1428,
    n1337
  );


  or
  g1397
  (
    n1561,
    n1370,
    n1355,
    n531,
    n578
  );


  or
  g1398
  (
    n1683,
    n1283,
    n524,
    n1328,
    n571
  );


  nor
  g1399
  (
    n1604,
    n581,
    n528,
    n1295,
    n1425
  );


  xor
  g1400
  (
    n1633,
    n571,
    n1358,
    n709,
    n1317
  );


  and
  g1401
  (
    n1634,
    n539,
    n559,
    n711,
    n1329
  );


  xor
  g1402
  (
    n1585,
    n1315,
    n1360,
    n1339,
    n589
  );


  and
  g1403
  (
    n1642,
    n1394,
    n544,
    n1360,
    n550
  );


  nand
  g1404
  (
    n1679,
    n1416,
    n1332,
    n702,
    n582
  );


  xnor
  g1405
  (
    n1457,
    n518,
    n557,
    n551,
    n703
  );


  xor
  g1406
  (
    n1572,
    n1328,
    n1096,
    n1381,
    n1421
  );


  xor
  g1407
  (
    n1580,
    n912,
    n917,
    n530,
    n916
  );


  and
  g1408
  (
    n1592,
    n1404,
    n1270,
    n1407,
    n539
  );


  xor
  g1409
  (
    n1474,
    n1344,
    n546,
    n1422,
    n1308
  );


  and
  g1410
  (
    n1599,
    n1403,
    n1389,
    n1302,
    n1406
  );


  nor
  g1411
  (
    n1593,
    n1284,
    n1274,
    n517,
    n1368
  );


  xnor
  g1412
  (
    n1546,
    n566,
    n576,
    n1420,
    n547
  );


  and
  g1413
  (
    n1606,
    n1356,
    n559,
    n1341,
    n1359
  );


  nand
  g1414
  (
    n1571,
    n1373,
    n1311,
    n525,
    n1304
  );


  or
  g1415
  (
    n1530,
    n1276,
    n1327,
    n541,
    n582
  );


  or
  g1416
  (
    n1468,
    n1321,
    n159,
    n553,
    n1301
  );


  xor
  g1417
  (
    KeyWire_0_33,
    n909,
    n555,
    n1411,
    n1347
  );


  nand
  g1418
  (
    n1516,
    n1272,
    n517,
    n593,
    n562
  );


  nand
  g1419
  (
    n1608,
    n1325,
    n570,
    n709,
    n1381
  );


  xor
  g1420
  (
    n1518,
    n1287,
    n1338,
    n1278,
    n526
  );


  and
  g1421
  (
    n1672,
    n1416,
    n565,
    n585,
    n713
  );


  nand
  g1422
  (
    n1534,
    n1362,
    n1310,
    n1291
  );


  nor
  g1423
  (
    n1455,
    n1280,
    n1297,
    n593,
    n706
  );


  xnor
  g1424
  (
    n1491,
    n1291,
    n1424,
    n1357,
    n921
  );


  and
  g1425
  (
    n1689,
    n1283,
    n1378,
    n1394,
    n1385
  );


  and
  g1426
  (
    n1453,
    n711,
    n1408,
    n1336,
    n705
  );


  xnor
  g1427
  (
    n1677,
    n710,
    n1323,
    n1273,
    n1278
  );


  nand
  g1428
  (
    n1506,
    n1338,
    n1396,
    n532,
    n556
  );


  and
  g1429
  (
    n1521,
    n1395,
    n537,
    n1354,
    n1298
  );


  and
  g1430
  (
    n1496,
    n1351,
    n561,
    n1382,
    n1305
  );


  or
  g1431
  (
    n1616,
    n593,
    n1094,
    n1419,
    n1290
  );


  nand
  g1432
  (
    n1476,
    n1271,
    n1372,
    n1327,
    n1366
  );


  nand
  g1433
  (
    n1471,
    n583,
    n1277,
    n534,
    n1289
  );


  or
  g1434
  (
    n1560,
    n1292,
    n1414,
    n1353,
    n1355
  );


  xor
  g1435
  (
    n1478,
    n1340,
    n1384,
    n1281,
    n576
  );


  or
  g1436
  (
    n1623,
    n1351,
    n550,
    n1418,
    n1275
  );


  nand
  g1437
  (
    n1535,
    n1318,
    n1375,
    n1420,
    n540
  );


  and
  g1438
  (
    n1682,
    n1332,
    n523,
    n546,
    n1346
  );


  xor
  g1439
  (
    n1690,
    n553,
    n1273,
    n1304,
    n1362
  );


  or
  g1440
  (
    n1567,
    n1310,
    n560,
    n557,
    n1410
  );


  nor
  g1441
  (
    KeyWire_0_24,
    n549,
    n1353,
    n702,
    n566
  );


  xor
  g1442
  (
    n1536,
    n1319,
    n1095,
    n1367,
    n575
  );


  or
  g1443
  (
    n1644,
    n590,
    n574,
    n551,
    n1410
  );


  xor
  g1444
  (
    n1452,
    n1413,
    n520,
    n548,
    n584
  );


  nand
  g1445
  (
    n1697,
    n1346,
    n712,
    n1408,
    n1366
  );


  nor
  g1446
  (
    n1448,
    n588,
    n1094,
    n1326,
    n1294
  );


  and
  g1447
  (
    n1620,
    n1286,
    n1427,
    n1382,
    n1327
  );


  nand
  g1448
  (
    n1552,
    n1303,
    n1302,
    n555,
    n1326
  );


  nand
  g1449
  (
    n1639,
    n561,
    n1366,
    n534,
    n1419
  );


  or
  g1450
  (
    n1481,
    n696,
    n1381,
    n1404,
    n1346
  );


  nor
  g1451
  (
    n1461,
    n1336,
    n1291,
    n713,
    n1274
  );


  and
  g1452
  (
    n1532,
    n533,
    n1341,
    n1411,
    n537
  );


  xor
  g1453
  (
    n1512,
    n1332,
    n520,
    n700,
    n1388
  );


  nand
  g1454
  (
    n1696,
    n1270,
    n1290,
    n1336,
    n517
  );


  nor
  g1455
  (
    n1544,
    n1279,
    n1329,
    n1303,
    n1324
  );


  xor
  g1456
  (
    n1628,
    n1363,
    n1331,
    n700,
    n1375
  );


  nand
  g1457
  (
    n1612,
    n564,
    n1356,
    n578,
    n550
  );


  xnor
  g1458
  (
    n1637,
    n1405,
    n536,
    n545,
    n1377
  );


  xnor
  g1459
  (
    n1641,
    n519,
    n1323,
    n524,
    n569
  );


  nor
  g1460
  (
    n1450,
    n1343,
    n1334,
    n1387,
    n1328
  );


  xor
  g1461
  (
    n1702,
    n711,
    n583,
    n590,
    n537
  );


  nand
  g1462
  (
    n1675,
    n592,
    n586,
    n1272,
    n580
  );


  nor
  g1463
  (
    n1600,
    n1369,
    n1301,
    n562,
    n1314
  );


  xnor
  g1464
  (
    n1494,
    n1385,
    n1420,
    n706,
    n526
  );


  nor
  g1465
  (
    n1464,
    n563,
    n1389,
    n1393
  );


  and
  g1466
  (
    n1598,
    n531,
    n1426,
    n1424,
    n1330
  );


  xnor
  g1467
  (
    n1447,
    n1378,
    n566,
    n556,
    n1417
  );


  nand
  g1468
  (
    n1531,
    n1334,
    n523,
    n1402,
    n1418
  );


  xor
  g1469
  (
    n1666,
    n518,
    n592,
    n1409,
    n520
  );


  or
  g1470
  (
    n1640,
    n1422,
    n1386,
    n1285,
    n1308
  );


  or
  g1471
  (
    n1581,
    n527,
    n591,
    n1324,
    n525
  );


  xor
  g1472
  (
    n1444,
    n542,
    n1282,
    n1308,
    n531
  );


  or
  g1473
  (
    n1627,
    n1370,
    n574,
    n578,
    n547
  );


  xor
  g1474
  (
    n1470,
    n1361,
    n1420,
    n579,
    n1425
  );


  xor
  g1475
  (
    n1681,
    n1392,
    n1293,
    n1342
  );


  xor
  g1476
  (
    n1582,
    n1403,
    n713,
    n1380,
    n1311
  );


  xor
  g1477
  (
    n1563,
    n1281,
    n1316,
    n544,
    n1278
  );


  or
  g1478
  (
    n1595,
    n547,
    n695,
    n541,
    n1412
  );


  and
  g1479
  (
    n1483,
    n551,
    n1344,
    n1280,
    n1343
  );


  nand
  g1480
  (
    n1662,
    n698,
    n577,
    n532,
    n1391
  );


  nor
  g1481
  (
    n1649,
    n1407,
    n545,
    n1281,
    n550
  );


  nor
  g1482
  (
    n1497,
    n1379,
    n534,
    n1347,
    n1387
  );


  nand
  g1483
  (
    n1484,
    n1406,
    n1321,
    n705,
    n526
  );


  or
  g1484
  (
    n1510,
    n1287,
    n1314,
    n587,
    n1352
  );


  or
  g1485
  (
    n1584,
    n1303,
    n535,
    n1361,
    n1349
  );


  nand
  g1486
  (
    n1501,
    n542,
    n1417,
    n523,
    n552
  );


  or
  g1487
  (
    n1685,
    n1400,
    n517,
    n704,
    n529
  );


  and
  g1488
  (
    n1556,
    n1403,
    n1394,
    n526,
    n708
  );


  or
  g1489
  (
    n1446,
    n1354,
    n911,
    n1326,
    n1392
  );


  xor
  g1490
  (
    n1482,
    n1422,
    n1404,
    n581,
    n920
  );


  xnor
  g1491
  (
    n1579,
    n1423,
    n1404,
    n1283,
    n1354
  );


  and
  g1492
  (
    n1469,
    n518,
    n1388,
    n1382,
    n555
  );


  nor
  g1493
  (
    n1473,
    n527,
    n1416,
    n700,
    n1315
  );


  or
  g1494
  (
    n1659,
    n1095,
    n537,
    n532,
    n1319
  );


  xor
  g1495
  (
    n1617,
    n538,
    n1325,
    n1320,
    n1375
  );


  nor
  g1496
  (
    n1575,
    n1348,
    n1094,
    n1336,
    n542
  );


  nor
  g1497
  (
    n1670,
    n1409,
    n1320,
    n1311,
    n1344
  );


  and
  g1498
  (
    n1622,
    n593,
    n1414,
    n1401,
    n1345
  );


  xnor
  g1499
  (
    n1533,
    n1398,
    n1350,
    n1379,
    n1393
  );


  nand
  g1500
  (
    KeyWire_0_63,
    n1321,
    n1388,
    n913,
    n714
  );


  xnor
  g1501
  (
    n1643,
    n1270,
    n1322,
    n703,
    n1359
  );


  nor
  g1502
  (
    n1503,
    n1284,
    n1350,
    n1323,
    n703
  );


  xor
  g1503
  (
    n1520,
    n1367,
    n1366,
    n585,
    n1331
  );


  or
  g1504
  (
    n1467,
    n1399,
    n1429,
    n577,
    n910
  );


  xor
  g1505
  (
    n1680,
    n573,
    n570,
    n1297,
    n704
  );


  and
  g1506
  (
    n1485,
    n1412,
    n1397,
    n1426,
    n1285
  );


  or
  g1507
  (
    n1698,
    n1384,
    n554,
    n1424,
    n1405
  );


  nor
  g1508
  (
    n1658,
    n566,
    n1301,
    n1337,
    n1419
  );


  nor
  g1509
  (
    n1538,
    n1299,
    n1274,
    n914,
    n1330
  );


  or
  g1510
  (
    n1619,
    n533,
    n591,
    n1384,
    n535
  );


  or
  g1511
  (
    n1502,
    n540,
    n588,
    n1349,
    n1368
  );


  and
  g1512
  (
    n1499,
    n1272,
    n1382,
    n1285,
    n1331
  );


  nor
  g1513
  (
    n1583,
    n1418,
    n1323,
    n527,
    n1333
  );


  nor
  g1514
  (
    n1542,
    n1389,
    n1401,
    n1427,
    n1360
  );


  xnor
  g1515
  (
    n1454,
    n530,
    n1386,
    n1385,
    n561
  );


  xnor
  g1516
  (
    n1610,
    n1308,
    n1402,
    n1297,
    n1339
  );


  or
  g1517
  (
    n1480,
    n1397,
    n543,
    n695,
    n1322
  );


  and
  g1518
  (
    n1687,
    n1307,
    n919,
    n1367,
    n1398
  );


  or
  g1519
  (
    n1573,
    n1325,
    n1380,
    n519,
    n1343
  );


  nor
  g1520
  (
    n1458,
    n1386,
    n1423,
    n1392,
    n1096
  );


  xnor
  g1521
  (
    n1553,
    n1300,
    n591,
    n699,
    n1295
  );


  nor
  g1522
  (
    n1653,
    n1391,
    n1309,
    n521,
    n698
  );


  nand
  g1523
  (
    n1442,
    n708,
    n562,
    n924,
    n588
  );


  xnor
  g1524
  (
    n1660,
    n1352,
    n573,
    n1369,
    n519
  );


  nor
  g1525
  (
    n1588,
    n1271,
    n1094,
    n1277,
    n1378
  );


  xnor
  g1526
  (
    n1631,
    n1293,
    n1413,
    n1358,
    n1307
  );


  xor
  g1527
  (
    n1570,
    n586,
    n536,
    n532,
    n1275
  );


  nor
  g1528
  (
    n1691,
    n698,
    n559,
    n568,
    n1370
  );


  nand
  g1529
  (
    n1463,
    n1342,
    n1318,
    n1427,
    n1387
  );


  nor
  g1530
  (
    n1465,
    n525,
    n541,
    n1373,
    n586
  );


  nor
  g1531
  (
    n1551,
    n1341,
    n1348,
    n1292,
    n548
  );


  xnor
  g1532
  (
    n1625,
    n530,
    n1326,
    n1355,
    n586
  );


  nand
  g1533
  (
    n1489,
    n1372,
    n536,
    n1348
  );


  and
  g1534
  (
    n1661,
    n1396,
    n1298,
    n1286,
    n1399
  );


  xnor
  g1535
  (
    n1540,
    n544,
    n1413,
    n524
  );


  or
  g1536
  (
    n1671,
    n1286,
    n592,
    n1415,
    n1288
  );


  xor
  g1537
  (
    n1493,
    n567,
    n1307,
    n1310,
    n1276
  );


  nor
  g1538
  (
    n1508,
    n707,
    n1374,
    n1349,
    n1410
  );


  or
  g1539
  (
    n1647,
    n1309,
    n1408,
    n1355,
    n1335
  );


  or
  g1540
  (
    n1549,
    n1425,
    n1374,
    n1301,
    n565
  );


  or
  g1541
  (
    n1594,
    n1384,
    n1304,
    n529,
    n1383
  );


  nor
  g1542
  (
    n1654,
    n1330,
    n1345,
    n577,
    n541
  );


  xnor
  g1543
  (
    n1605,
    n1376,
    n530,
    n583,
    n707
  );


  xnor
  g1544
  (
    n1439,
    n558,
    n709,
    n582,
    n1417
  );


  and
  g1545
  (
    n1507,
    n1284,
    n1288,
    n1371,
    n589
  );


  xnor
  g1546
  (
    n1564,
    n1342,
    n538,
    n1386,
    n543
  );


  nand
  g1547
  (
    n1543,
    n699,
    n1394,
    n573,
    n1364
  );


  or
  g1548
  (
    n1688,
    n527,
    n1324,
    n548,
    n1405
  );


  nand
  g1549
  (
    n1514,
    n564,
    n1412,
    n1350,
    n1360
  );


  xor
  g1550
  (
    n1621,
    n1282,
    n540,
    n1298
  );


  or
  g1551
  (
    n1636,
    n1405,
    n1329,
    n533,
    n1350
  );


  xor
  g1552
  (
    n1517,
    n1414,
    n572,
    n1417,
    n1294
  );


  and
  g1553
  (
    n1562,
    n1316,
    n1280,
    n697,
    n1429
  );


  or
  g1554
  (
    n1651,
    n1409,
    n1388,
    n1290,
    n1421
  );


  nand
  g1555
  (
    n1490,
    n1296,
    n1338,
    n1304,
    n1359
  );


  nand
  g1556
  (
    n1475,
    n579,
    n710,
    n1293,
    n1364
  );


  or
  g1557
  (
    n1576,
    n1414,
    n1400,
    n591,
    n1313
  );


  nor
  g1558
  (
    n1477,
    n573,
    n696,
    n701,
    n1340
  );


  xnor
  g1559
  (
    n1441,
    n1333,
    n1279,
    n1277,
    n577
  );


  or
  g1560
  (
    n1522,
    n1349,
    n1335,
    n1312,
    n706
  );


  xnor
  g1561
  (
    n1545,
    n568,
    n710,
    n1278,
    n1307
  );


  nor
  g1562
  (
    n1449,
    n559,
    n1320,
    n1322,
    n1383
  );


  or
  g1563
  (
    n1618,
    n1391,
    n705,
    n522,
    n1370
  );


  or
  g1564
  (
    n1537,
    n549,
    n1422,
    n1415,
    n569
  );


  or
  g1565
  (
    n1462,
    n1272,
    n1377,
    n1396,
    n1340
  );


  nand
  g1566
  (
    n1665,
    n1306,
    n569,
    n1348,
    n918
  );


  and
  g1567
  (
    n1645,
    n1380,
    n922,
    n556,
    n1313
  );


  nand
  g1568
  (
    n1495,
    n1408,
    n1338,
    n1354,
    n1363
  );


  or
  g1569
  (
    n1451,
    n1358,
    n528,
    n1095,
    n525
  );


  and
  g1570
  (
    n1498,
    n1406,
    n1289,
    n583,
    n1335
  );


  and
  g1571
  (
    n1487,
    n584,
    n1357,
    n551,
    n531
  );


  xnor
  g1572
  (
    n1638,
    n1356,
    n1343,
    n1271,
    n1426
  );


  or
  g1573
  (
    n1558,
    n1391,
    n584,
    n1400,
    n545
  );


  xor
  g1574
  (
    n1568,
    n1281,
    n533,
    n587,
    n1409
  );


  xor
  g1575
  (
    n1574,
    n1313,
    n575,
    n557,
    n1292
  );


  xor
  g1576
  (
    n1472,
    n555,
    n701,
    n544,
    n1320
  );


  and
  g1577
  (
    n1657,
    n558,
    n1309,
    n556,
    n522
  );


  or
  g1578
  (
    n1700,
    n538,
    n699,
    n1367,
    n1381
  );


  or
  g1579
  (
    n1440,
    n1377,
    n1415,
    n1399,
    n1397
  );


  xnor
  g1580
  (
    n1692,
    n1282,
    n701,
    n1371,
    n571
  );


  or
  g1581
  (
    n1515,
    n1364,
    n1383,
    n1293,
    n711
  );


  xor
  g1582
  (
    n1590,
    n1390,
    n1351,
    n1296,
    n572
  );


  xnor
  g1583
  (
    n1650,
    n1093,
    n1363,
    n560,
    n1375
  );


  xnor
  g1584
  (
    n1500,
    n1276,
    n546,
    n1332,
    n1341
  );


  or
  g1585
  (
    n1701,
    n1352,
    n1300,
    n1331,
    n1275
  );


  xnor
  g1586
  (
    n1652,
    n1361,
    n1291,
    n570,
    n1359
  );


  nor
  g1587
  (
    n1486,
    n704,
    n1329,
    n1425,
    n694
  );


  and
  g1588
  (
    n1656,
    n1290,
    n574,
    n1288,
    n1346
  );


  xnor
  g1589
  (
    n1547,
    n1347,
    n714,
    n588,
    n1397
  );


  nor
  g1590
  (
    n1646,
    n1399,
    n708,
    n1395,
    n552
  );


  or
  g1591
  (
    n1676,
    n549,
    n1345,
    n1390,
    n1361
  );


  nor
  g1592
  (
    n1577,
    n1299,
    n576,
    n707,
    n1412
  );


  or
  g1593
  (
    n1539,
    n708,
    n1317,
    n585,
    n702
  );


  nand
  g1594
  (
    n1527,
    n1393,
    n565,
    n1315,
    n1421
  );


  and
  g1595
  (
    n1678,
    n1096,
    n1327,
    n1334,
    n707
  );


  and
  g1596
  (
    n1505,
    n1371,
    n1402,
    n1285,
    n1374
  );


  xor
  g1597
  (
    n1460,
    n521,
    n1419,
    n580
  );


  nand
  g1598
  (
    n1557,
    n1296,
    n528,
    n1424,
    n1093
  );


  or
  g1599
  (
    n1528,
    n1353,
    n572,
    n1377,
    n1403
  );


  nand
  g1600
  (
    n1525,
    n519,
    n923,
    n1334,
    n534
  );


  nand
  g1601
  (
    n1695,
    n1313,
    n547,
    n1363,
    n1357
  );


  or
  g1602
  (
    KeyWire_0_55,
    n700,
    n1312,
    n1317,
    n1368
  );


  and
  g1603
  (
    n1554,
    n561,
    n1401,
    n1300,
    n553
  );


  nor
  g1604
  (
    n1443,
    n1418,
    n705,
    n706,
    n1305
  );


  or
  g1605
  (
    n1614,
    n564,
    n712,
    n1328,
    n568
  );


  and
  g1606
  (
    n1456,
    n1312,
    n1423,
    n587,
    n1383
  );


  and
  g1607
  (
    n1655,
    n1395,
    n1297,
    n1385,
    n1306
  );


  xor
  g1608
  (
    n1630,
    n1373,
    n1402,
    n1407,
    n709
  );


  xnor
  g1609
  (
    n1529,
    n699,
    n562,
    n697,
    n1340
  );


  and
  g1610
  (
    n1589,
    n1362,
    n565,
    n1287,
    n1415
  );


  xnor
  g1611
  (
    n1648,
    n1379,
    n1321,
    n704,
    n1365
  );


  xnor
  g1612
  (
    n1624,
    n1371,
    n1284,
    n579,
    n1295
  );


  xnor
  g1613
  (
    n1635,
    n1400,
    n712,
    n1303,
    n590
  );


  or
  g1614
  (
    n1596,
    n558,
    n522,
    n1372,
    n1302
  );


  or
  g1615
  (
    n1578,
    n1288,
    n695,
    n1393,
    n1277
  );


  and
  g1616
  (
    n1541,
    n1406,
    n521,
    n1426,
    n1299
  );


  xor
  g1617
  (
    n1694,
    n1372,
    n1379,
    n1289,
    n1294
  );


  xnor
  g1618
  (
    n1555,
    n1305,
    n1324,
    n1275,
    n1428
  );


  and
  g1619
  (
    n1548,
    n552,
    n1401,
    n560,
    n1428
  );


  or
  g1620
  (
    n1686,
    n1292,
    n1365,
    n1337,
    n1305
  );


  or
  g1621
  (
    n1684,
    n1368,
    n1356,
    n159,
    n1353
  );


  xnor
  g1622
  (
    n1587,
    n578,
    n557,
    n576,
    n564
  );


  and
  g1623
  (
    n1607,
    n1300,
    n563,
    n908,
    n1362
  );


  xor
  g1624
  (
    n1611,
    n558,
    n546,
    n1339,
    n1376
  );


  xor
  g1625
  (
    n1663,
    n1318,
    n553,
    n1374,
    n924
  );


  or
  g1626
  (
    n1601,
    n696,
    n1314,
    n1322,
    n713
  );


  xor
  g1627
  (
    n1509,
    n575,
    n710,
    n529,
    n567
  );


  xor
  g1628
  (
    n1615,
    n538,
    n1352,
    n571,
    n1395
  );


  nor
  g1629
  (
    n1632,
    n1306,
    n1316,
    n1289
  );


  and
  g1630
  (
    n1668,
    n1279,
    n1302,
    n520,
    n1333
  );


  xnor
  g1631
  (
    n1586,
    n1423,
    n545,
    n575,
    n549
  );


  or
  g1632
  (
    n1703,
    n1369,
    n554,
    n518,
    n1390
  );


  or
  g1633
  (
    n1693,
    n563,
    n1319,
    n1407,
    n521
  );


  and
  g1634
  (
    n1550,
    n584,
    n1421,
    n703,
    n1318
  );


  nand
  g1635
  (
    n1591,
    n1319,
    n1335,
    n915,
    n1410
  );


  or
  g1636
  (
    n1479,
    n552,
    n1273,
    n1306,
    n1286
  );


  nand
  g1637
  (
    n1513,
    n539,
    n695,
    n1273,
    n1295
  );


  and
  g1638
  (
    n1504,
    n1096,
    n589,
    n1364,
    n1315
  );


  xor
  g1639
  (
    n1597,
    n548,
    n1416,
    n581,
    n585
  );


  nor
  g1640
  (
    n1603,
    n1390,
    n1299,
    n714,
    n587
  );


  and
  g1641
  (
    n1609,
    n1376,
    n1396,
    n568,
    n1357
  );


  nand
  g1642
  (
    n1667,
    n1369,
    n590,
    n1427,
    n1378
  );


  nand
  g1643
  (
    n1445,
    n1282,
    n1312,
    n701,
    n697
  );


  and
  g1644
  (
    n1559,
    n698,
    n1283,
    n1309,
    n579
  );


  nand
  g1645
  (
    n1488,
    n1351,
    n1392,
    n1411,
    n1330
  );


  nor
  g1646
  (
    n1699,
    n1311,
    n1411,
    n1095,
    n1296
  );


  xor
  g1647
  (
    n1673,
    n1365,
    n1337,
    n540,
    n543
  );


  or
  g1648
  (
    n1459,
    n567,
    n1333,
    n1429,
    n1428
  );


  xnor
  g1649
  (
    n1669,
    n522,
    n539,
    n572,
    n712
  );


  xnor
  g1650
  (
    n1629,
    n1376,
    n535,
    n1280,
    n528
  );


  nor
  g1651
  (
    n1519,
    n1294,
    n543,
    n570,
    n1287
  );


  or
  g1652
  (
    n1602,
    n535,
    n1373,
    n1276,
    n1325
  );


  and
  g1653
  (
    n1664,
    n589,
    n563,
    n702,
    n1398
  );


  nand
  g1654
  (
    KeyWire_0_36,
    n1559,
    n1591,
    n1641,
    n1537
  );


  nor
  g1655
  (
    n1796,
    n1545,
    n1536,
    n1540,
    n1480
  );


  xor
  g1656
  (
    n1878,
    n1558,
    n1547,
    n1598,
    n1469
  );


  xnor
  g1657
  (
    n1787,
    n1647,
    n1633,
    n1446,
    n1471
  );


  nand
  g1658
  (
    n1750,
    n1633,
    n1586,
    n1497,
    n1557
  );


  xnor
  g1659
  (
    n1935,
    n1433,
    n1625,
    n1550,
    n1604
  );


  or
  g1660
  (
    n1714,
    n1592,
    n1649,
    n1481,
    n1644
  );


  or
  g1661
  (
    n1863,
    n1508,
    n1441,
    n1487,
    n1579
  );


  and
  g1662
  (
    n1899,
    n1541,
    n1629,
    n1509,
    n1514
  );


  and
  g1663
  (
    KeyWire_0_61,
    n1590,
    n1207,
    n1616,
    n1649
  );


  nor
  g1664
  (
    n1883,
    n1615,
    n1575,
    n1515,
    n1548
  );


  and
  g1665
  (
    KeyWire_0_11,
    n1557,
    n1661,
    n1505,
    n1500
  );


  nor
  g1666
  (
    n1917,
    n1590,
    n1606,
    n1562,
    n1667
  );


  nand
  g1667
  (
    n1821,
    n1488,
    n1450,
    n1547,
    n1624
  );


  or
  g1668
  (
    n1791,
    n1596,
    n1541,
    n1208,
    n1589
  );


  nand
  g1669
  (
    KeyWire_0_16,
    n1464,
    n1591,
    n1499,
    n1510
  );


  nand
  g1670
  (
    n1886,
    n1656,
    n1641,
    n1440,
    n1543
  );


  and
  g1671
  (
    n1833,
    n1577,
    n1585,
    n1574,
    n1668
  );


  nand
  g1672
  (
    n1776,
    n1206,
    n1496,
    n1538,
    n1521
  );


  or
  g1673
  (
    n1716,
    n1508,
    n1663,
    n1530,
    n1671
  );


  xnor
  g1674
  (
    n1810,
    n1529,
    n1459,
    n1542,
    n1567
  );


  and
  g1675
  (
    n1782,
    n1673,
    n1457,
    n1437,
    n1208
  );


  xor
  g1676
  (
    n1851,
    n1608,
    n1576,
    n1599,
    n1616
  );


  or
  g1677
  (
    n1875,
    n1592,
    n1666,
    n1501
  );


  xor
  g1678
  (
    n1845,
    n1649,
    n1605,
    n1622,
    n1670
  );


  nand
  g1679
  (
    n1809,
    n1439,
    n1511,
    n1479,
    n1671
  );


  xor
  g1680
  (
    n1839,
    n1655,
    n1627,
    n1587,
    n1644
  );


  xor
  g1681
  (
    n1908,
    n1613,
    n1466,
    n1439,
    n1507
  );


  nand
  g1682
  (
    n1759,
    n1522,
    n1660,
    n1506,
    n1550
  );


  xor
  g1683
  (
    n1721,
    n1546,
    n1614,
    n1548,
    n1653
  );


  and
  g1684
  (
    n1783,
    n1669,
    n1436,
    n1472,
    n1438
  );


  and
  g1685
  (
    n1947,
    n1587,
    n1582,
    n1650,
    n1473
  );


  and
  g1686
  (
    n1726,
    n1433,
    n1548,
    n1535,
    n1662
  );


  and
  g1687
  (
    n1814,
    n1207,
    n1530,
    n1651,
    n1666
  );


  nor
  g1688
  (
    n1815,
    n1568,
    n1638,
    n1604,
    n1533
  );


  or
  g1689
  (
    n1837,
    n1659,
    n1612,
    n1485,
    n1539
  );


  nor
  g1690
  (
    n1874,
    n1448,
    n1630,
    n1654,
    n1516
  );


  xnor
  g1691
  (
    n1806,
    n1506,
    n1526,
    n1563
  );


  and
  g1692
  (
    n1857,
    n1461,
    n1573,
    n1628,
    n1634
  );


  and
  g1693
  (
    n1732,
    n1549,
    n1553,
    n1670,
    n1585
  );


  nor
  g1694
  (
    n1803,
    n1492,
    n1440,
    n1601,
    n1589
  );


  xor
  g1695
  (
    n1744,
    n1617,
    n1606,
    n1611,
    n1517
  );


  or
  g1696
  (
    n1948,
    n1485,
    n1634,
    n1474,
    n1526
  );


  or
  g1697
  (
    n1887,
    n1489,
    n1458,
    n1450,
    n1522
  );


  or
  g1698
  (
    n1927,
    n1635,
    n1574,
    n1607,
    n1619
  );


  xor
  g1699
  (
    n1895,
    n1490,
    n1636,
    n1618,
    n1438
  );


  nor
  g1700
  (
    n1755,
    n1558,
    n1659,
    n1660,
    n1670
  );


  xor
  g1701
  (
    n1751,
    n1544,
    n1642,
    n1437,
    n1672
  );


  nand
  g1702
  (
    n1774,
    n1636,
    n1624,
    n1526,
    n1578
  );


  nand
  g1703
  (
    n1784,
    n1433,
    n1667,
    n1538,
    n1657
  );


  nand
  g1704
  (
    n1792,
    n1641,
    n1645,
    n1524,
    n1477
  );


  nor
  g1705
  (
    n1747,
    n1466,
    n1568,
    n1494,
    n1448
  );


  nor
  g1706
  (
    n1890,
    n1489,
    n1513,
    n1449,
    n1615
  );


  or
  g1707
  (
    n1812,
    n1449,
    n1508,
    n1493,
    n1439
  );


  xnor
  g1708
  (
    n1775,
    n1522,
    n1479,
    n1588,
    n1515
  );


  xnor
  g1709
  (
    n1804,
    n1570,
    n1591,
    n1582,
    n1460
  );


  nor
  g1710
  (
    n1892,
    n1497,
    n1623,
    n1505,
    n1593
  );


  or
  g1711
  (
    n1754,
    n1207,
    n1604,
    n1649,
    n1516
  );


  xor
  g1712
  (
    n1842,
    n1580,
    n1614,
    n1592,
    n1595
  );


  or
  g1713
  (
    n1773,
    n1441,
    n1646,
    n1523,
    n1547
  );


  xor
  g1714
  (
    n1933,
    n1509,
    n1578,
    n1563,
    n1620
  );


  nor
  g1715
  (
    n1934,
    n1566,
    n1432,
    n1630,
    n1511
  );


  xor
  g1716
  (
    n1818,
    n1669,
    n1512,
    n1455,
    n1483
  );


  nor
  g1717
  (
    n1752,
    n1460,
    n1435,
    n1631,
    n1462
  );


  xnor
  g1718
  (
    n1885,
    n1468,
    n1570,
    n1544,
    n1644
  );


  xor
  g1719
  (
    n1820,
    n1456,
    n1516,
    n1617,
    n1664
  );


  nor
  g1720
  (
    n1847,
    n1533,
    n1661,
    n1551,
    n1569
  );


  nand
  g1721
  (
    n1718,
    n1606,
    n1571,
    n1539,
    n1556
  );


  xor
  g1722
  (
    n1719,
    n1470,
    n1467,
    n1628,
    n1490
  );


  xor
  g1723
  (
    n1938,
    n1584,
    n1652,
    n1494,
    n1461
  );


  and
  g1724
  (
    n1789,
    n1617,
    n1559,
    n1196,
    n1573
  );


  xor
  g1725
  (
    n1835,
    n1563,
    n1486,
    n1534,
    n1430
  );


  nor
  g1726
  (
    n1849,
    n1664,
    n1457,
    n1612,
    n1553
  );


  xor
  g1727
  (
    n1765,
    n1603,
    n1647,
    n1597,
    n1537
  );


  nor
  g1728
  (
    n1936,
    n1591,
    n1445,
    n1609,
    n1659
  );


  xor
  g1729
  (
    n1746,
    n1517,
    n1605,
    n1435,
    n1604
  );


  xnor
  g1730
  (
    n1788,
    n1491,
    n1600,
    n1520,
    n1665
  );


  xnor
  g1731
  (
    n1930,
    n1619,
    n1674,
    n1645,
    n1545
  );


  and
  g1732
  (
    n1888,
    n1491,
    n1622,
    n1488,
    n1561
  );


  xnor
  g1733
  (
    n1760,
    n1658,
    n1528,
    n1471,
    n1456
  );


  and
  g1734
  (
    n1757,
    n1562,
    n1480,
    n1519,
    n1611
  );


  nor
  g1735
  (
    n1801,
    n1615,
    n1635,
    n1627,
    n1586
  );


  and
  g1736
  (
    n1816,
    n1635,
    n1646,
    n1467,
    n1480
  );


  nand
  g1737
  (
    n1846,
    n1583,
    n1492,
    n1629,
    n1557
  );


  nand
  g1738
  (
    n1922,
    n1490,
    n1498,
    n1430,
    n1671
  );


  xnor
  g1739
  (
    n1704,
    n1592,
    n1621,
    n1581,
    n1473
  );


  nor
  g1740
  (
    n1722,
    n1663,
    n1598,
    n1462,
    n1622
  );


  and
  g1741
  (
    n1799,
    n1581,
    n1484,
    n1630,
    n1507
  );


  nand
  g1742
  (
    n1943,
    n1560,
    n1478,
    n1628,
    n1430
  );


  nand
  g1743
  (
    n1769,
    n1631,
    n1538,
    n1564,
    n1559
  );


  nor
  g1744
  (
    n1738,
    n1525,
    n1549,
    n1587,
    n1551
  );


  or
  g1745
  (
    n1944,
    n1579,
    n1459,
    n1638,
    n1447
  );


  xnor
  g1746
  (
    n1850,
    n1492,
    n1504,
    n1539,
    n1582
  );


  or
  g1747
  (
    n1884,
    n1475,
    n1527,
    n1631,
    n1444
  );


  and
  g1748
  (
    n1872,
    n1430,
    n1599,
    n1654,
    n1485
  );


  xnor
  g1749
  (
    n1828,
    n1495,
    n1542,
    n1500,
    n1206
  );


  xnor
  g1750
  (
    n1731,
    n1558,
    n1597,
    n1672,
    n1496
  );


  nor
  g1751
  (
    n1709,
    n1535,
    n1673,
    n1568,
    n1564
  );


  or
  g1752
  (
    n1767,
    n1648,
    n1634,
    n1531,
    n1545
  );


  xnor
  g1753
  (
    n1909,
    n1655,
    n1546,
    n1463,
    n1473
  );


  xnor
  g1754
  (
    n1761,
    n1588,
    n1672,
    n1506,
    n1543
  );


  nor
  g1755
  (
    n1913,
    n1515,
    n1542,
    n1637,
    n1639
  );


  and
  g1756
  (
    n1891,
    n1497,
    n1576,
    n1606,
    n1642
  );


  xnor
  g1757
  (
    n1902,
    n1634,
    n1536,
    n1518,
    n1466
  );


  nand
  g1758
  (
    n1705,
    n1435,
    n1431,
    n1482,
    n1467
  );


  and
  g1759
  (
    n1853,
    n1653,
    n1512,
    n1566,
    n1658
  );


  nor
  g1760
  (
    n1932,
    n1473,
    n1504,
    n1534,
    n1603
  );


  xor
  g1761
  (
    n1728,
    n1441,
    n1465,
    n1479,
    n1644
  );


  nor
  g1762
  (
    n1869,
    n1566,
    n1505,
    n1664,
    n1443
  );


  xnor
  g1763
  (
    n1770,
    n1598,
    n1513,
    n1588,
    n1650
  );


  and
  g1764
  (
    n1861,
    n1503,
    n1600,
    n1571,
    n1491
  );


  nand
  g1765
  (
    n1827,
    n1207,
    n1669,
    n1619,
    n1612
  );


  xor
  g1766
  (
    n1779,
    n1657,
    n1607,
    n1467,
    n1672
  );


  nor
  g1767
  (
    n1912,
    n1446,
    n1518,
    n1563,
    n1514
  );


  xor
  g1768
  (
    n1873,
    n1510,
    n1555,
    n1515,
    n1608
  );


  and
  g1769
  (
    n1858,
    n1588,
    n1455,
    n1465,
    n1481
  );


  xnor
  g1770
  (
    n1717,
    n1524,
    n1556,
    n1590,
    n1514
  );


  nor
  g1771
  (
    n1802,
    n1523,
    n1670,
    n1625,
    n1441
  );


  and
  g1772
  (
    n1838,
    n1458,
    n1569,
    n1452,
    n1600
  );


  xor
  g1773
  (
    n1949,
    n1530,
    n1196,
    n1436,
    n1489
  );


  or
  g1774
  (
    n1727,
    n1527,
    n1471,
    n1503,
    n1436
  );


  nor
  g1775
  (
    n1832,
    n1652,
    n1594,
    n1482,
    n1442
  );


  or
  g1776
  (
    n1894,
    n1453,
    n1661,
    n1556,
    n1521
  );


  and
  g1777
  (
    n1919,
    n1517,
    n1614,
    n1462,
    n1560
  );


  or
  g1778
  (
    n1711,
    n1595,
    n1609,
    n1558,
    n1434
  );


  and
  g1779
  (
    n1910,
    n1567,
    n1575,
    n1545,
    n1641
  );


  nand
  g1780
  (
    n1707,
    n1576,
    n1197,
    n1485,
    n1464
  );


  xor
  g1781
  (
    n1798,
    n1576,
    n1539,
    n1470,
    n1435
  );


  xnor
  g1782
  (
    n1817,
    n1499,
    n1564,
    n1535,
    n1671
  );


  xnor
  g1783
  (
    n1739,
    n1642,
    n1587,
    n1560,
    n1574
  );


  xnor
  g1784
  (
    n1906,
    n1498,
    n1442,
    n1560,
    n1537
  );


  nor
  g1785
  (
    n1748,
    n1493,
    n1605,
    n1594,
    n1451
  );


  nor
  g1786
  (
    n1925,
    n1637,
    n1632,
    n1654,
    n1628
  );


  nand
  g1787
  (
    n1915,
    n1621,
    n1643,
    n1590,
    n1600
  );


  and
  g1788
  (
    n1900,
    n1633,
    n1579,
    n1518,
    n1443
  );


  nor
  g1789
  (
    n1733,
    n1548,
    n1554,
    n1562,
    n1667
  );


  and
  g1790
  (
    n1905,
    n1555,
    n1540,
    n1593,
    n1611
  );


  nand
  g1791
  (
    n1942,
    n1645,
    n1501,
    n1651,
    n1583
  );


  nor
  g1792
  (
    n1785,
    n1498,
    n1472,
    n1585,
    n1629
  );


  xnor
  g1793
  (
    n1764,
    n1472,
    n1474,
    n1622,
    n930
  );


  xnor
  g1794
  (
    n1800,
    n1620,
    n1493,
    n1640,
    n1584
  );


  nand
  g1795
  (
    n1781,
    n1486,
    n1484,
    n1637,
    n1488
  );


  or
  g1796
  (
    n1826,
    n1455,
    n1639,
    n1669,
    n1582
  );


  nor
  g1797
  (
    n1929,
    n1550,
    n1513,
    n1673,
    n1505
  );


  xnor
  g1798
  (
    n1829,
    n1519,
    n1626,
    n930,
    n1509
  );


  and
  g1799
  (
    n1825,
    n1551,
    n1479,
    n1646,
    n1637
  );


  or
  g1800
  (
    n1706,
    n1525,
    n1570,
    n1471,
    n1478
  );


  xnor
  g1801
  (
    n1896,
    n1208,
    n1561,
    n1495,
    n1597
  );


  xor
  g1802
  (
    n1946,
    n1474,
    n1495,
    n1454,
    n1608
  );


  xnor
  g1803
  (
    n1766,
    n1583,
    n1517,
    n1535,
    n1609
  );


  xnor
  g1804
  (
    n1824,
    n1623,
    n1657,
    n1448,
    n1543
  );


  xor
  g1805
  (
    n1745,
    n1445,
    n1663,
    n1464,
    n1661
  );


  and
  g1806
  (
    n1893,
    n1498,
    n1638,
    n1434,
    n1554
  );


  xor
  g1807
  (
    n1939,
    n1580,
    n1478,
    n1520,
    n1546
  );


  nor
  g1808
  (
    n1881,
    n1559,
    n1453,
    n1660,
    n1502
  );


  xor
  g1809
  (
    KeyWire_0_18,
    n1482,
    n1554,
    n1618,
    n1533
  );


  and
  g1810
  (
    n1871,
    n1472,
    n1487,
    n1447,
    n1453
  );


  nand
  g1811
  (
    n1848,
    n1432,
    n1603,
    n1528,
    n1662
  );


  nand
  g1812
  (
    n1823,
    n1611,
    n1546,
    n1617,
    n1439
  );


  xnor
  g1813
  (
    n1777,
    n1468,
    n1444,
    n1461,
    n1449
  );


  or
  g1814
  (
    n1911,
    n1603,
    n1536,
    n1457,
    n1450
  );


  and
  g1815
  (
    n1737,
    n1613,
    n1567,
    n1609,
    n1469
  );


  xnor
  g1816
  (
    n1822,
    n1626,
    n1491,
    n1500,
    n1469
  );


  or
  g1817
  (
    n1805,
    n1502,
    n1550,
    n1431,
    n1610
  );


  nand
  g1818
  (
    n1901,
    n1574,
    n1477,
    n1521,
    n1451
  );


  xnor
  g1819
  (
    n1795,
    n1486,
    n1665,
    n1562,
    n1540
  );


  xnor
  g1820
  (
    n1921,
    n1593,
    n1577,
    n1594,
    n1508
  );


  or
  g1821
  (
    n1730,
    n1639,
    n1519,
    n1443,
    n1518
  );


  nor
  g1822
  (
    n1876,
    n1470,
    n1647,
    n1489,
    n1474
  );


  xor
  g1823
  (
    n1808,
    n1459,
    n1573,
    n1542,
    n1463
  );


  xnor
  g1824
  (
    n1903,
    n1488,
    n1490,
    n1636,
    n1657
  );


  xnor
  g1825
  (
    n1740,
    n1496,
    n1627,
    n1636,
    n1666
  );


  nand
  g1826
  (
    n1797,
    n1476,
    n1525,
    n1571,
    n1556
  );


  nand
  g1827
  (
    n1811,
    n1527,
    n1532,
    n1504,
    n1442
  );


  nor
  g1828
  (
    n1831,
    n1621,
    n1510,
    n1602,
    n1197
  );


  xor
  g1829
  (
    n1840,
    n1506,
    n1552,
    n1484,
    n1616
  );


  or
  g1830
  (
    n1843,
    n1596,
    n1532,
    n1623,
    n1553
  );


  and
  g1831
  (
    n1786,
    n1656,
    n1614,
    n1494,
    n1594
  );


  xor
  g1832
  (
    n1841,
    n1610,
    n1507,
    n1643,
    n1583
  );


  or
  g1833
  (
    n1852,
    n1638,
    n1432,
    n1483,
    n1520
  );


  or
  g1834
  (
    n1844,
    n1601,
    n1437,
    n1477,
    n1596
  );


  or
  g1835
  (
    n1855,
    n1541,
    n1524,
    n1652,
    n1531
  );


  xor
  g1836
  (
    n1931,
    n1470,
    n1581,
    n1500,
    n1630
  );


  xor
  g1837
  (
    n1813,
    n1660,
    n1651,
    n1533,
    n1648
  );


  nor
  g1838
  (
    n1904,
    n1468,
    n1432,
    n1572,
    n1668
  );


  nor
  g1839
  (
    n1794,
    n1444,
    n1442,
    n1525,
    n1619
  );


  xnor
  g1840
  (
    n1836,
    n1448,
    n1534,
    n1519,
    n1466
  );


  xor
  g1841
  (
    n1715,
    n1493,
    n1640,
    n1569,
    n1632
  );


  nor
  g1842
  (
    n1763,
    n1444,
    n1565,
    n1446,
    n1532
  );


  nor
  g1843
  (
    n1819,
    n1438,
    n1524,
    n1477,
    n1531
  );


  xnor
  g1844
  (
    n1952,
    n1618,
    n1564,
    n1431,
    n1447
  );


  nand
  g1845
  (
    n1898,
    n1577,
    n1626,
    n1452,
    n1632
  );


  nor
  g1846
  (
    n1877,
    n1580,
    n1487,
    n1571,
    n1437
  );


  nand
  g1847
  (
    n1768,
    n1512,
    n1667,
    n1561,
    n1624
  );


  nand
  g1848
  (
    n1790,
    n1475,
    n1598,
    n1643,
    n1534
  );


  xor
  g1849
  (
    n1734,
    n1484,
    n1573,
    n1452,
    n1554
  );


  or
  g1850
  (
    n1923,
    n1593,
    n1599,
    n1665,
    n1589
  );


  nand
  g1851
  (
    n1941,
    n1551,
    n1452,
    n1569,
    n1468
  );


  or
  g1852
  (
    n1758,
    n1572,
    n1541,
    n1673,
    n1602
  );


  nor
  g1853
  (
    n1870,
    n1476,
    n1595,
    n1465,
    n1668
  );


  or
  g1854
  (
    n1868,
    n1570,
    n1501,
    n1462,
    n1543
  );


  nand
  g1855
  (
    n1862,
    n1601,
    n1618,
    n1664,
    n1655
  );


  nand
  g1856
  (
    n1713,
    n1450,
    n1575,
    n1633,
    n1481
  );


  nor
  g1857
  (
    n1741,
    n1568,
    n1476,
    n1449,
    n1663
  );


  nand
  g1858
  (
    n1924,
    n1453,
    n1648,
    n1516,
    n1504
  );


  nor
  g1859
  (
    KeyWire_0_5,
    n1613,
    n1455,
    n1512,
    n1537
  );


  nor
  g1860
  (
    n1735,
    n1566,
    n1538,
    n1555,
    n1631
  );


  or
  g1861
  (
    n1951,
    n1445,
    n1659,
    n1596,
    n1510
  );


  xor
  g1862
  (
    n1854,
    n1658,
    n1495,
    n1499,
    n1433
  );


  or
  g1863
  (
    n1743,
    n1527,
    n1469,
    n1478,
    n1577
  );


  nor
  g1864
  (
    n1920,
    n1475,
    n1458,
    n1578,
    n1446
  );


  or
  g1865
  (
    n1897,
    n1544,
    n1584,
    n1436,
    n1456
  );


  or
  g1866
  (
    n1928,
    n1465,
    n1514,
    n1503,
    n1458
  );


  xor
  g1867
  (
    n1926,
    n1658,
    n1656,
    n1197,
    n1607
  );


  or
  g1868
  (
    n1880,
    n1561,
    n1650,
    n1623,
    n1457
  );


  nand
  g1869
  (
    n1720,
    n1612,
    n1552,
    n1584,
    n1639
  );


  or
  g1870
  (
    n1710,
    n1579,
    n1581,
    n1544,
    n1645
  );


  or
  g1871
  (
    n1860,
    n1653,
    n1475,
    n1549,
    n1586
  );


  xnor
  g1872
  (
    n1712,
    n1601,
    n1655,
    n1461,
    n1674
  );


  and
  g1873
  (
    n1749,
    n1552,
    n1463,
    n1499,
    n1454
  );


  xor
  g1874
  (
    KeyWire_0_15,
    n1443,
    n1602,
    n1578,
    n1197
  );


  xnor
  g1875
  (
    n1778,
    n1653,
    n1528,
    n1459,
    n1595
  );


  or
  g1876
  (
    n1725,
    n1434,
    n1487,
    n1625,
    n1553
  );


  nor
  g1877
  (
    n1879,
    n1642,
    n1650,
    n1511,
    n1665
  );


  nand
  g1878
  (
    n1736,
    n1431,
    n1620,
    n1586,
    n1529
  );


  nand
  g1879
  (
    n1708,
    n1608,
    n1625,
    n1530,
    n1565
  );


  nor
  g1880
  (
    n1723,
    n1521,
    n1451,
    n1610,
    n1532
  );


  nand
  g1881
  (
    n1772,
    n1632,
    n1540,
    n1621,
    n1476
  );


  and
  g1882
  (
    n1907,
    n1610,
    n1494,
    n1572,
    n1486
  );


  and
  g1883
  (
    n1859,
    n1529,
    n1640,
    n1531,
    n1481
  );


  xnor
  g1884
  (
    n1753,
    n1662,
    n1536,
    n1668,
    n1646
  );


  xnor
  g1885
  (
    n1830,
    n1567,
    n1523,
    n1624,
    n1607
  );


  or
  g1886
  (
    n1834,
    n1616,
    n1580,
    n1597,
    n1523
  );


  xor
  g1887
  (
    n1940,
    n1620,
    n1613,
    n1451,
    n1547
  );


  xnor
  g1888
  (
    n1724,
    n1549,
    n1647,
    n1463,
    n1208
  );


  or
  g1889
  (
    n1950,
    n1492,
    n1585,
    n1438,
    n1497
  );


  xnor
  g1890
  (
    n1793,
    n1434,
    n1501,
    n1602,
    n1507
  );


  nand
  g1891
  (
    n1866,
    n1656,
    n1513,
    n1643,
    n1464
  );


  nor
  g1892
  (
    n1916,
    n1529,
    n1605,
    n1447,
    n1503
  );


  and
  g1893
  (
    n1856,
    n1482,
    n1652,
    n1572,
    n1496
  );


  or
  g1894
  (
    n1807,
    n1456,
    n1520,
    n1615,
    n1552
  );


  xor
  g1895
  (
    n1742,
    n1483,
    n1460,
    n1565,
    n1480
  );


  xnor
  g1896
  (
    n1882,
    n1599,
    n1440,
    n1445
  );


  or
  g1897
  (
    n1865,
    n1483,
    n1454,
    n1565,
    n1557
  );


  xor
  g1898
  (
    n1889,
    n1555,
    n1511,
    n1522,
    n1654
  );


  nand
  g1899
  (
    n1937,
    n1648,
    n1502,
    n1640,
    n1627
  );


  xnor
  g1900
  (
    n1914,
    n1635,
    n1509,
    n1662,
    n1629
  );


  or
  g1901
  (
    n1945,
    n1502,
    n1460,
    n1651,
    n1575
  );


  and
  g1902
  (
    n1918,
    n1626,
    n1454,
    n1589,
    n1528
  );


  nand
  g1903
  (
    n1953,
    n1705,
    n1706
  );


  xor
  g1904
  (
    n1954,
    n1706,
    n1705,
    n1704
  );


  and
  g1905
  (
    n1955,
    n1706,
    n1707
  );


  nor
  g1906
  (
    n1963,
    n1955,
    n1953,
    n1954,
    n1709
  );


  xnor
  g1907
  (
    n1961,
    n1710,
    n1709,
    n1713,
    n1708
  );


  xor
  g1908
  (
    n1962,
    n1712,
    n1708,
    n1710
  );


  xnor
  g1909
  (
    n1964,
    n1713,
    n1953,
    n1708,
    n1711
  );


  xnor
  g1910
  (
    n1960,
    n1709,
    n1712,
    n1707,
    n1714
  );


  xor
  g1911
  (
    n1957,
    n1953,
    n1712,
    n1714,
    n1954
  );


  and
  g1912
  (
    n1959,
    n1712,
    n1709,
    n1708,
    n1710
  );


  xor
  g1913
  (
    n1958,
    n1954,
    n1711,
    n1713
  );


  xnor
  g1914
  (
    n1956,
    n1953,
    n1711,
    n1954,
    n1713
  );


  buf
  g1915
  (
    KeyWire_0_4,
    n1715
  );


  not
  g1916
  (
    n1966,
    n1714
  );


  not
  g1917
  (
    n1969,
    n1960
  );


  and
  g1918
  (
    n1965,
    n1714,
    n1963,
    n1961
  );


  xnor
  g1919
  (
    n1967,
    n1962,
    n1964,
    n1715
  );


  or
  g1920
  (
    n1982,
    n1727,
    n1727,
    n1719,
    n1718
  );


  nand
  g1921
  (
    n1985,
    n1966,
    n1729,
    n1726
  );


  xor
  g1922
  (
    n1983,
    n1723,
    n1719,
    n1722
  );


  and
  g1923
  (
    n1987,
    n1716,
    n1967,
    n1965
  );


  xor
  g1924
  (
    n1979,
    n1968,
    n1721,
    n1716,
    n1715
  );


  xor
  g1925
  (
    n1978,
    n1720,
    n1716,
    n1726,
    n1727
  );


  or
  g1926
  (
    n1976,
    n1965,
    n1715,
    n1728
  );


  nand
  g1927
  (
    n1977,
    n1717,
    n1729,
    n1969,
    n1968
  );


  nand
  g1928
  (
    n1972,
    n1726,
    n1969,
    n1723,
    n1722
  );


  nor
  g1929
  (
    n1980,
    n1727,
    n1724,
    n1730
  );


  xnor
  g1930
  (
    n1984,
    n1724,
    n1967,
    n1720,
    n1716
  );


  and
  g1931
  (
    n1975,
    n1730,
    n1723,
    n1966,
    n1725
  );


  xor
  g1932
  (
    n1974,
    n1723,
    n1728,
    n1720,
    n1965
  );


  nor
  g1933
  (
    n1989,
    n1966,
    n1717,
    n1725
  );


  or
  g1934
  (
    n1988,
    n1718,
    n1725,
    n1726,
    n1967
  );


  and
  g1935
  (
    n1973,
    n1969,
    n1719,
    n1728,
    n1968
  );


  nand
  g1936
  (
    n1970,
    n1966,
    n1719,
    n1721,
    n1729
  );


  xor
  g1937
  (
    n1986,
    n1967,
    n1718,
    n1721,
    n1720
  );


  nand
  g1938
  (
    n1971,
    n1721,
    n1969,
    n1722,
    n1718
  );


  and
  g1939
  (
    n1981,
    n1717,
    n1724,
    n1968,
    n1725
  );


  nor
  g1940
  (
    n2043,
    n1756,
    n1747,
    n1772,
    n1755
  );


  nand
  g1941
  (
    n2046,
    n1975,
    n1761,
    n1970,
    n1775
  );


  and
  g1942
  (
    n1994,
    n1786,
    n1739,
    n1737,
    n1730
  );


  or
  g1943
  (
    n2037,
    n1738,
    n1758,
    n1764,
    n1975
  );


  xor
  g1944
  (
    n2014,
    n1984,
    n1733,
    n1759,
    n1972
  );


  xnor
  g1945
  (
    n2056,
    n1765,
    n1777,
    n1787,
    n1784
  );


  xor
  g1946
  (
    n1998,
    n1776,
    n1757,
    n1758,
    n1987
  );


  or
  g1947
  (
    n2023,
    n1773,
    n1986,
    n1972,
    n1780
  );


  nand
  g1948
  (
    n2007,
    n1742,
    n1984,
    n1758,
    n1741
  );


  nand
  g1949
  (
    n2063,
    n1753,
    n1986,
    n1786,
    n1777
  );


  xor
  g1950
  (
    n2006,
    n1978,
    n1785,
    n1762,
    n1775
  );


  or
  g1951
  (
    n2066,
    n1760,
    n1978,
    n1768,
    n1752
  );


  and
  g1952
  (
    n2047,
    n1744,
    n1748,
    n1742,
    n1733
  );


  xor
  g1953
  (
    n2048,
    n1754,
    n1743,
    n1988,
    n1737
  );


  xor
  g1954
  (
    n2040,
    n1771,
    n1780,
    n1736,
    n1757
  );


  or
  g1955
  (
    n2042,
    n1987,
    n1730,
    n1761,
    n1785
  );


  nor
  g1956
  (
    n2044,
    n1751,
    n1977,
    n1786,
    n1752
  );


  and
  g1957
  (
    n2001,
    n1785,
    n1767,
    n1746,
    n1979
  );


  nor
  g1958
  (
    n1999,
    n1732,
    n1984,
    n1747,
    n1771
  );


  or
  g1959
  (
    n2050,
    n1979,
    n1989,
    n1779,
    n1740
  );


  and
  g1960
  (
    n2064,
    n1988,
    n1732,
    n1756,
    n1750
  );


  xnor
  g1961
  (
    n2039,
    n1738,
    n1983,
    n1981,
    n1747
  );


  nor
  g1962
  (
    n2016,
    n1784,
    n1768,
    n1779,
    n1787
  );


  xor
  g1963
  (
    n2067,
    n1790,
    n1759,
    n1750,
    n1788
  );


  or
  g1964
  (
    n2000,
    n1971,
    n1762,
    n1753,
    n1741
  );


  xor
  g1965
  (
    n2025,
    n1788,
    n1778,
    n1741,
    n1988
  );


  nand
  g1966
  (
    n2019,
    n1784,
    n1975,
    n1777,
    n1764
  );


  nand
  g1967
  (
    n2018,
    n1783,
    n1743,
    n1776,
    n1779
  );


  nand
  g1968
  (
    n2003,
    n1765,
    n1783,
    n1982,
    n1761
  );


  xor
  g1969
  (
    n2055,
    n1980,
    n1735,
    n1744,
    n1757
  );


  nor
  g1970
  (
    n1991,
    n1979,
    n1770,
    n1740,
    n1972
  );


  xor
  g1971
  (
    n2017,
    n1731,
    n1753,
    n1756,
    n1987
  );


  nor
  g1972
  (
    n2029,
    n1774,
    n1971,
    n1733,
    n1977
  );


  and
  g1973
  (
    n2033,
    n1775,
    n1983,
    n1973,
    n1782
  );


  xnor
  g1974
  (
    n2036,
    n1982,
    n1775,
    n1768,
    n1773
  );


  or
  g1975
  (
    n2057,
    n1736,
    n1759,
    n1774,
    n1745
  );


  xor
  g1976
  (
    n2002,
    n1735,
    n1740,
    n1747,
    n1786
  );


  xor
  g1977
  (
    n2026,
    n1752,
    n1978,
    n1985,
    n1739
  );


  and
  g1978
  (
    n2013,
    n1976,
    n1789,
    n1765,
    n1734
  );


  xor
  g1979
  (
    n1990,
    n1758,
    n1770,
    n1746,
    n1973
  );


  and
  g1980
  (
    n2052,
    n1732,
    n1985,
    n1778
  );


  xnor
  g1981
  (
    n2015,
    n1731,
    n1782,
    n1743,
    n1734
  );


  xnor
  g1982
  (
    n2069,
    n1970,
    n1737,
    n1767,
    n1989
  );


  and
  g1983
  (
    n2024,
    n1745,
    n1981,
    n1757,
    n1783
  );


  or
  g1984
  (
    n2010,
    n1749,
    n1980,
    n1789,
    n1748
  );


  xnor
  g1985
  (
    n2045,
    n1781,
    n1974,
    n1744,
    n1971
  );


  and
  g1986
  (
    n2058,
    n1976,
    n1986,
    n1731,
    n1760
  );


  xnor
  g1987
  (
    n1996,
    n1741,
    n1782,
    n1755,
    n1773
  );


  nor
  g1988
  (
    n2060,
    n1977,
    n1754,
    n1769,
    n1742
  );


  xor
  g1989
  (
    n1995,
    n1987,
    n1763,
    n1979,
    n1981
  );


  and
  g1990
  (
    n2031,
    n1769,
    n1970,
    n1754,
    n1731
  );


  and
  g1991
  (
    n2022,
    n1762,
    n1980,
    n1744,
    n1973
  );


  xor
  g1992
  (
    n2051,
    n1759,
    n1755,
    n1749,
    n1753
  );


  nand
  g1993
  (
    n2038,
    n1782,
    n1778,
    n1971,
    n1749
  );


  and
  g1994
  (
    n1993,
    n1983,
    n1977,
    n1745,
    n1738
  );


  nand
  g1995
  (
    n2061,
    n1740,
    n1781,
    n1739
  );


  nor
  g1996
  (
    n2032,
    n1766,
    n1756,
    n1779,
    n1750
  );


  nor
  g1997
  (
    n2009,
    n1772,
    n1746,
    n1787,
    n1742
  );


  or
  g1998
  (
    KeyWire_0_60,
    n1982,
    n1776,
    n1760,
    n1763
  );


  or
  g1999
  (
    n2005,
    n1785,
    n1739,
    n1738,
    n1751
  );


  and
  g2000
  (
    n2011,
    n1972,
    n1737,
    n1745,
    n1974
  );


  or
  g2001
  (
    n2059,
    n1770,
    n1751,
    n1746,
    n1767
  );


  xor
  g2002
  (
    n2035,
    n1766,
    n1773,
    n1988,
    n1982
  );


  xnor
  g2003
  (
    n2053,
    n1978,
    n1781,
    n1772,
    n1975
  );


  xnor
  g2004
  (
    n2030,
    n1983,
    n1765,
    n1766,
    n1734
  );


  and
  g2005
  (
    n2004,
    n1787,
    n1974,
    n1976,
    n1771
  );


  nor
  g2006
  (
    n2027,
    n1986,
    n1769,
    n1774,
    n1749
  );


  xor
  g2007
  (
    n2020,
    n1735,
    n1764,
    n1733,
    n1754
  );


  xnor
  g2008
  (
    n2008,
    n1767,
    n1770,
    n1780,
    n1752
  );


  or
  g2009
  (
    n2054,
    n1743,
    n1760,
    n1734,
    n1774
  );


  and
  g2010
  (
    n2034,
    n1981,
    n1783,
    n1784,
    n1763
  );


  xnor
  g2011
  (
    n2028,
    n1973,
    n1789,
    n1985
  );


  and
  g2012
  (
    n2049,
    n1976,
    n1970,
    n1735,
    n1776
  );


  xnor
  g2013
  (
    n1997,
    n1751,
    n1989,
    n1750,
    n1761
  );


  or
  g2014
  (
    n2012,
    n1790,
    n1771,
    n1768,
    n1736
  );


  and
  g2015
  (
    n2021,
    n1755,
    n1772,
    n1769,
    n1780
  );


  or
  g2016
  (
    n1992,
    n1732,
    n1974,
    n1766,
    n1777
  );


  and
  g2017
  (
    n2068,
    n1984,
    n1748,
    n1778
  );


  nand
  g2018
  (
    n2041,
    n1980,
    n1788,
    n1763,
    n1989
  );


  and
  g2019
  (
    n2065,
    n1764,
    n1762,
    n1736,
    n1788
  );


  xor
  g2020
  (
    n2075,
    n1050,
    n1052,
    n1054,
    n1051
  );


  xnor
  g2021
  (
    n2077,
    n1991,
    n1053
  );


  or
  g2022
  (
    n2073,
    n1049,
    n1050,
    n1051
  );


  and
  g2023
  (
    n2072,
    n1052,
    n1050,
    n1990,
    n1991
  );


  xnor
  g2024
  (
    n2071,
    n1054,
    n1052,
    n1990
  );


  xnor
  g2025
  (
    n2074,
    n1053,
    n1990,
    n1049,
    n1054
  );


  nor
  g2026
  (
    n2076,
    n1053,
    n1049,
    n1992,
    n1990
  );


  and
  g2027
  (
    n2070,
    n1050,
    n1051,
    n1054,
    n1991
  );


  and
  g2028
  (
    n2102,
    n2071,
    n1994,
    n2077,
    n1993
  );


  or
  g2029
  (
    n2094,
    n2077,
    n1999,
    n2003,
    n2000
  );


  xnor
  g2030
  (
    n2109,
    n2002,
    n1992,
    n1794,
    n1675
  );


  xor
  g2031
  (
    n2084,
    n1992,
    n2003,
    n1995,
    n2075
  );


  nand
  g2032
  (
    n2097,
    n1794,
    n2000,
    n1795,
    n2005
  );


  nand
  g2033
  (
    n2108,
    n2073,
    n1675,
    n2071,
    n2002
  );


  xor
  g2034
  (
    n2100,
    n1997,
    n1793,
    n1994,
    n2074
  );


  or
  g2035
  (
    n2106,
    n1796,
    n1798,
    n2005,
    n1793
  );


  and
  g2036
  (
    n2095,
    n2074,
    n1795,
    n1997,
    n2070
  );


  xnor
  g2037
  (
    n2099,
    n2076,
    n1992,
    n2072,
    n2075
  );


  nand
  g2038
  (
    n2107,
    n2004,
    n2002,
    n1674,
    n2001
  );


  and
  g2039
  (
    n2093,
    n1797,
    n2001,
    n1676
  );


  nand
  g2040
  (
    n2105,
    n2074,
    n2000,
    n2072,
    n1995
  );


  nand
  g2041
  (
    n2081,
    n2071,
    n1796,
    n2073,
    n2004
  );


  nand
  g2042
  (
    n2101,
    n1798,
    n1793,
    n1796
  );


  or
  g2043
  (
    n2098,
    n2074,
    n1791,
    n2070,
    n1998
  );


  xnor
  g2044
  (
    KeyWire_0_46,
    n1791,
    n1996,
    n1795,
    n1994
  );


  nor
  g2045
  (
    n2078,
    n1798,
    n2005,
    n1797,
    n1799
  );


  nor
  g2046
  (
    n2096,
    n2076,
    n1796,
    n1995,
    n1997
  );


  or
  g2047
  (
    KeyWire_0_32,
    n1996,
    n1995,
    n1997,
    n1993
  );


  or
  g2048
  (
    n2087,
    n1998,
    n2073,
    n1795,
    n2072
  );


  nor
  g2049
  (
    n2089,
    n2004,
    n1998,
    n2077,
    n2076
  );


  nand
  g2050
  (
    n2083,
    n2002,
    n2070,
    n2077,
    n1998
  );


  xor
  g2051
  (
    n2086,
    n1999,
    n1996,
    n1994,
    n1790
  );


  nor
  g2052
  (
    n2092,
    n1993,
    n1675,
    n1792,
    n1790
  );


  nand
  g2053
  (
    n2088,
    n1798,
    n1792,
    n1791,
    n2003
  );


  or
  g2054
  (
    n2082,
    n2001,
    n2000,
    n1674,
    n2072
  );


  and
  g2055
  (
    n2103,
    n2003,
    n1797,
    n1792,
    n1675
  );


  nor
  g2056
  (
    n2104,
    n2071,
    n1996,
    n2070,
    n2004
  );


  xor
  g2057
  (
    n2090,
    n1792,
    n1797,
    n2076,
    n1999
  );


  nor
  g2058
  (
    n2079,
    n1791,
    n2073,
    n1999,
    n1794
  );


  nor
  g2059
  (
    n2091,
    n1993,
    n1794,
    n2075
  );


  nor
  g2060
  (
    n2123,
    n2105,
    n1799,
    n2109,
    n2099
  );


  or
  g2061
  (
    n2111,
    n1822,
    n1818,
    n1803,
    n2103
  );


  nor
  g2062
  (
    n2128,
    n1805,
    n1801,
    n1820,
    n1800
  );


  nand
  g2063
  (
    n2141,
    n2087,
    n1816,
    n1800,
    n2088
  );


  nand
  g2064
  (
    n2136,
    n1808,
    n1810,
    n1807,
    n1809
  );


  or
  g2065
  (
    n2115,
    n1810,
    n1802,
    n1812,
    n2086
  );


  or
  g2066
  (
    n2140,
    n2079,
    n1808,
    n2091,
    n1820
  );


  nor
  g2067
  (
    n2114,
    n2106,
    n1803,
    n1800,
    n2098
  );


  or
  g2068
  (
    n2137,
    n1805,
    n1816,
    n1799,
    n1803
  );


  and
  g2069
  (
    n2118,
    n1823,
    n2096,
    n2089,
    n1818
  );


  or
  g2070
  (
    n2139,
    n2094,
    n1807,
    n1804,
    n2092
  );


  and
  g2071
  (
    n2125,
    n2108,
    n1813,
    n1819,
    n1801
  );


  xor
  g2072
  (
    n2113,
    n1811,
    n2090,
    n1818,
    n1801
  );


  xnor
  g2073
  (
    n2120,
    n1812,
    n1813,
    n1820,
    n2082
  );


  and
  g2074
  (
    n2133,
    n1806,
    n1817,
    n1811,
    n1815
  );


  xor
  g2075
  (
    n2110,
    n1803,
    n1804,
    n1813,
    n2080
  );


  xnor
  g2076
  (
    n2135,
    n2100,
    n1812,
    n1802,
    n1804
  );


  xnor
  g2077
  (
    n2132,
    n1802,
    n1816,
    n1822,
    n1810
  );


  nand
  g2078
  (
    n2121,
    n2104,
    n2095,
    n1815,
    n1814
  );


  and
  g2079
  (
    n2129,
    n1819,
    n2102,
    n2097,
    n1817
  );


  and
  g2080
  (
    n2122,
    n2084,
    n1814,
    n1821,
    n1801
  );


  nand
  g2081
  (
    n2119,
    n1822,
    n1812,
    n2101,
    n1807
  );


  or
  g2082
  (
    n2131,
    n1814,
    n1814,
    n1815,
    n1806
  );


  xnor
  g2083
  (
    n2138,
    n1806,
    n1817,
    n1816,
    n1821
  );


  nor
  g2084
  (
    n2127,
    n2078,
    n1815,
    n1809
  );


  nor
  g2085
  (
    n2112,
    n1805,
    n2085,
    n1821,
    n1804
  );


  or
  g2086
  (
    n2116,
    n2093,
    n1820,
    n1799,
    n1800
  );


  xor
  g2087
  (
    n2124,
    n1819,
    n1805,
    n1802,
    n1810
  );


  xnor
  g2088
  (
    n2117,
    n1813,
    n1822,
    n1811
  );


  or
  g2089
  (
    n2134,
    n1807,
    n2107,
    n1819,
    n1817
  );


  and
  g2090
  (
    n2126,
    n1821,
    n1808,
    n2081
  );


  xor
  g2091
  (
    n2130,
    n2083,
    n1809,
    n1818,
    n1806
  );


  or
  g2092
  (
    n2152,
    n2065,
    n2051,
    n1686,
    n2121
  );


  nor
  g2093
  (
    n2246,
    n2052,
    n1678,
    n2123,
    n1698
  );


  nor
  g2094
  (
    n2269,
    n2018,
    n1689,
    n2057,
    n2009
  );


  and
  g2095
  (
    KeyWire_0_28,
    n2013,
    n1680,
    n2134,
    n1676
  );


  nand
  g2096
  (
    n2260,
    n2026,
    n2113,
    n2020,
    n2005
  );


  nor
  g2097
  (
    n2234,
    n2139,
    n1702,
    n2054,
    n1677
  );


  xor
  g2098
  (
    n2158,
    n2126,
    n2049,
    n2037,
    n2011
  );


  nand
  g2099
  (
    n2238,
    n2038,
    n2038,
    n2019,
    n2113
  );


  xnor
  g2100
  (
    n2229,
    n2061,
    n49,
    n1955,
    n2122
  );


  and
  g2101
  (
    n2157,
    n2055,
    n2137,
    n2058,
    n2049
  );


  nor
  g2102
  (
    n2206,
    n1676,
    n2034,
    n2053,
    n2062
  );


  nor
  g2103
  (
    n2201,
    n2043,
    n2051,
    n2135,
    n2059
  );


  nand
  g2104
  (
    n2214,
    n2141,
    n1682,
    n2011,
    n2114
  );


  nor
  g2105
  (
    n2209,
    n2015,
    n1681,
    n2007,
    n2012
  );


  or
  g2106
  (
    n2223,
    n1692,
    n2062,
    n1689,
    n2010
  );


  nor
  g2107
  (
    n2154,
    n2056,
    n1688,
    n2035,
    n2060
  );


  nor
  g2108
  (
    n2212,
    n2014,
    n1677,
    n2007,
    n2031
  );


  xor
  g2109
  (
    n2187,
    n2063,
    n2127,
    n2050,
    n1699
  );


  or
  g2110
  (
    n2222,
    n2114,
    n2017,
    n2119,
    n48
  );


  or
  g2111
  (
    n2261,
    n1690,
    n2126,
    n1677,
    n1698
  );


  xnor
  g2112
  (
    n2257,
    n2115,
    n1678,
    n1687,
    n2067
  );


  xor
  g2113
  (
    n2268,
    n2025,
    n2116,
    n2055,
    n361
  );


  xor
  g2114
  (
    n2190,
    n1697,
    n2023,
    n2067,
    n2114
  );


  or
  g2115
  (
    n2241,
    n2060,
    n2066,
    n2039,
    n2014
  );


  or
  g2116
  (
    n2151,
    n1694,
    n1690,
    n2063,
    n2053
  );


  xnor
  g2117
  (
    n2153,
    n2030,
    n2013,
    n1676,
    n2021
  );


  xor
  g2118
  (
    n2156,
    n2137,
    n2139,
    n2061
  );


  or
  g2119
  (
    n2161,
    n2060,
    n2112,
    n2131
  );


  nor
  g2120
  (
    n2247,
    n1703,
    n2128,
    n1682,
    n2056
  );


  nor
  g2121
  (
    n2164,
    n2051,
    n2128,
    n2057,
    n2059
  );


  xnor
  g2122
  (
    n2263,
    n2061,
    n2008,
    n2037,
    n2126
  );


  xnor
  g2123
  (
    n2203,
    n161,
    n2129,
    n2042
  );


  nand
  g2124
  (
    n2237,
    n2130,
    n1693,
    n2117,
    n2025
  );


  xor
  g2125
  (
    n2147,
    n2055,
    n2009,
    n2114,
    n2040
  );


  and
  g2126
  (
    n2219,
    n2054,
    n1696,
    n2047,
    n2035
  );


  nand
  g2127
  (
    n2194,
    n2115,
    n2140,
    n2120,
    n2064
  );


  or
  g2128
  (
    KeyWire_0_21,
    n2048,
    n2054,
    n2024,
    n2141
  );


  xnor
  g2129
  (
    n2244,
    n2017,
    n2111,
    n2030,
    n48
  );


  nand
  g2130
  (
    n2191,
    n159,
    n2035,
    n2060,
    n2015
  );


  and
  g2131
  (
    n2226,
    n2011,
    n2027,
    n2131,
    n2047
  );


  and
  g2132
  (
    n2239,
    n2130,
    n1682,
    n2134,
    n2124
  );


  nand
  g2133
  (
    KeyWire_0_30,
    n2055,
    n1684,
    n2043,
    n2059
  );


  or
  g2134
  (
    n2227,
    n2048,
    n1700,
    n2136,
    n2119
  );


  or
  g2135
  (
    n2146,
    n2140,
    n1700,
    n2009,
    n2029
  );


  xnor
  g2136
  (
    n2189,
    n2014,
    n2041,
    n1691,
    n2131
  );


  nor
  g2137
  (
    n2230,
    n2121,
    n1695,
    n1679,
    n2065
  );


  xor
  g2138
  (
    n2216,
    n1679,
    n1677,
    n2056,
    n1678
  );


  xnor
  g2139
  (
    n2208,
    n2028,
    n2141,
    n1687,
    n2029
  );


  xor
  g2140
  (
    n2163,
    n1688,
    n1690,
    n49
  );


  xnor
  g2141
  (
    n2266,
    n1697,
    n2123,
    n2118,
    n160
  );


  nor
  g2142
  (
    n2207,
    n2122,
    n2140,
    n362,
    n2011
  );


  nand
  g2143
  (
    n2221,
    n2027,
    n2007,
    n2041,
    n1702
  );


  xor
  g2144
  (
    n2228,
    n1686,
    n2110,
    n2122,
    n1695
  );


  xnor
  g2145
  (
    n2177,
    n1701,
    n2134,
    n1686,
    n2015
  );


  xnor
  g2146
  (
    n2232,
    n2010,
    n2025,
    n2113,
    n1688
  );


  and
  g2147
  (
    n2249,
    n2117,
    n2120,
    n1698,
    n1684
  );


  nand
  g2148
  (
    n2167,
    n1696,
    n2016,
    n2138,
    n2039
  );


  xnor
  g2149
  (
    n2174,
    n2050,
    n2127,
    n2058,
    n2111
  );


  nand
  g2150
  (
    n2173,
    n2127,
    n2136,
    n2010,
    n2062
  );


  xor
  g2151
  (
    n2259,
    n1691,
    n2026,
    n2023,
    n2064
  );


  or
  g2152
  (
    n2256,
    n2018,
    n2115,
    n2019,
    n1701
  );


  xor
  g2153
  (
    n2170,
    n2125,
    n2057,
    n2113,
    n2064
  );


  or
  g2154
  (
    n2142,
    n2046,
    n2010,
    n2033,
    n2138
  );


  xnor
  g2155
  (
    n2148,
    n2135,
    n2049,
    n160,
    n1702
  );


  nor
  g2156
  (
    n2210,
    n2125,
    n2131,
    n2052,
    n1695
  );


  nor
  g2157
  (
    n2250,
    n2124,
    n2118,
    n2046,
    n2041
  );


  nor
  g2158
  (
    n2184,
    n160,
    n2123,
    n2036,
    n2052
  );


  or
  g2159
  (
    n2145,
    n2014,
    n2127,
    n2039,
    n1694
  );


  nand
  g2160
  (
    n2180,
    n2044,
    n2120,
    n2046,
    n1679
  );


  nor
  g2161
  (
    n2235,
    n2117,
    n2056,
    n1687,
    n2046
  );


  xor
  g2162
  (
    n2155,
    n2021,
    n1689,
    n1694,
    n1685
  );


  xor
  g2163
  (
    n2240,
    n2024,
    n2031,
    n2029,
    n1703
  );


  nor
  g2164
  (
    n2245,
    n2037,
    n1692,
    n2067,
    n2047
  );


  nand
  g2165
  (
    n2178,
    n2050,
    n361,
    n1691,
    n2136
  );


  nand
  g2166
  (
    n2258,
    n1682,
    n2066,
    n2023,
    n2045
  );


  nand
  g2167
  (
    n2202,
    n361,
    n2028,
    n2132,
    n2021
  );


  nor
  g2168
  (
    n2182,
    n49,
    n2038,
    n2016,
    n2024
  );


  and
  g2169
  (
    n2220,
    n2141,
    n2007,
    n1685,
    n2008
  );


  nor
  g2170
  (
    n2262,
    n1691,
    n2111,
    n1693,
    n1685
  );


  nand
  g2171
  (
    n2159,
    n1700,
    n2021,
    n2123,
    n1701
  );


  or
  g2172
  (
    n2265,
    n2020,
    n2117,
    n2017,
    n1955
  );


  nand
  g2173
  (
    n2160,
    n2026,
    n1679,
    n1699,
    n2024
  );


  nand
  g2174
  (
    n2183,
    n2033,
    n2048,
    n2132,
    n2118
  );


  and
  g2175
  (
    n2267,
    n2115,
    n2015,
    n49,
    n2006
  );


  and
  g2176
  (
    n2205,
    n2121,
    n2133,
    n2110,
    n2020
  );


  xnor
  g2177
  (
    n2204,
    n2064,
    n2028,
    n2030,
    n2135
  );


  or
  g2178
  (
    n2188,
    n2118,
    n2006,
    n2134,
    n1696
  );


  and
  g2179
  (
    n2168,
    n2133,
    n1698,
    n2033,
    n1703
  );


  nand
  g2180
  (
    n2196,
    n2033,
    n1684,
    n2016,
    n2121
  );


  or
  g2181
  (
    n2225,
    n1697,
    n2022,
    n2116,
    n2112
  );


  xnor
  g2182
  (
    n2166,
    n1680,
    n1699,
    n2124,
    n2022
  );


  nand
  g2183
  (
    n2193,
    n2137,
    n2027,
    n1955
  );


  nor
  g2184
  (
    n2192,
    n2043,
    n2013,
    n1703,
    n2062
  );


  or
  g2185
  (
    n2213,
    n2058,
    n2135,
    n2067,
    n2139
  );


  xnor
  g2186
  (
    n2165,
    n2008,
    n2116,
    n2025
  );


  or
  g2187
  (
    n2217,
    n2031,
    n2052,
    n2059,
    n2034
  );


  xnor
  g2188
  (
    n2251,
    n1685,
    n2140,
    n160,
    n2133
  );


  nor
  g2189
  (
    n2169,
    n2132,
    n1686,
    n2032
  );


  nor
  g2190
  (
    n2185,
    n2129,
    n1681,
    n2065,
    n2053
  );


  and
  g2191
  (
    n2175,
    n2022,
    n2028,
    n2047,
    n1692
  );


  or
  g2192
  (
    n2143,
    n2126,
    n1687,
    n2128,
    n2044
  );


  xor
  g2193
  (
    n2215,
    n2133,
    n2026,
    n2119,
    n1683
  );


  xnor
  g2194
  (
    n2150,
    n2120,
    n2110,
    n2129,
    n2125
  );


  xnor
  g2195
  (
    n2181,
    n2019,
    n48,
    n2045,
    n1693
  );


  xnor
  g2196
  (
    n2264,
    n2045,
    n2006,
    n2051,
    n2042
  );


  xnor
  g2197
  (
    n2248,
    n2043,
    n2042,
    n2022,
    n1693
  );


  and
  g2198
  (
    n2233,
    n2040,
    n2130,
    n2030,
    n2012
  );


  xor
  g2199
  (
    n2200,
    n48,
    n2039,
    n2019,
    n2013
  );


  or
  g2200
  (
    n2236,
    n2034,
    n2049,
    n2012,
    n2066
  );


  xnor
  g2201
  (
    n2253,
    n2063,
    n1699,
    n2036,
    n2124
  );


  or
  g2202
  (
    n2186,
    n2065,
    n1683,
    n1701,
    n2020
  );


  or
  g2203
  (
    n2176,
    n2061,
    n2050,
    n2054,
    n2110
  );


  nor
  g2204
  (
    n2252,
    n1688,
    n2136,
    n2130,
    n2138
  );


  nand
  g2205
  (
    n2218,
    n2036,
    n1695,
    n1697,
    n1684
  );


  xnor
  g2206
  (
    n2198,
    n2038,
    n1700,
    n2040,
    n2048
  );


  or
  g2207
  (
    n2254,
    n1683,
    n2016,
    n2125,
    n161
  );


  and
  g2208
  (
    n2172,
    n2044,
    n2032,
    n2041,
    n2018
  );


  nand
  g2209
  (
    n2149,
    n2042,
    n1692,
    n2012,
    n1702
  );


  xnor
  g2210
  (
    n2211,
    n2037,
    n2063,
    n2029,
    n2053
  );


  nand
  g2211
  (
    n2171,
    n2066,
    n1689,
    n2031,
    n2122
  );


  and
  g2212
  (
    n2179,
    n1694,
    n2112,
    n1696,
    n1678
  );


  xor
  g2213
  (
    n2195,
    n2058,
    n1823,
    n2119,
    n1681
  );


  nand
  g2214
  (
    n2197,
    n2036,
    n2032,
    n1681,
    n1680
  );


  and
  g2215
  (
    n2231,
    n2040,
    n2128,
    n2057,
    n2023
  );


  xnor
  g2216
  (
    n2224,
    n2009,
    n362,
    n1680,
    n2035
  );


  and
  g2217
  (
    n2162,
    n2008,
    n2006,
    n2111,
    n2045
  );


  and
  g2218
  (
    n2243,
    n2132,
    n2018,
    n2034,
    n1683
  );


  or
  g2219
  (
    n2199,
    n2044,
    n2137,
    n2017,
    n2138
  );


  nor
  g2220
  (
    n2475,
    n1916,
    n981,
    n1921
  );


  nand
  g2221
  (
    n2521,
    n1924,
    n2187,
    n2159
  );


  and
  g2222
  (
    n2444,
    n2254,
    n2167,
    n1866
  );


  nand
  g2223
  (
    n2299,
    n1893,
    n2180,
    n2175
  );


  or
  g2224
  (
    n2443,
    n1825,
    n1850,
    n1934
  );


  or
  g2225
  (
    KeyWire_0_49,
    n1892,
    n2242,
    n2207
  );


  xor
  g2226
  (
    n2375,
    n1929,
    n1880,
    n1848
  );


  nand
  g2227
  (
    n2325,
    n1922,
    n1834,
    n2243
  );


  nand
  g2228
  (
    n2307,
    n2161,
    n1846,
    n991
  );


  xor
  g2229
  (
    n2469,
    n1907,
    n2202,
    n2166
  );


  and
  g2230
  (
    n2508,
    n1896,
    n2160,
    n2144
  );


  and
  g2231
  (
    n2441,
    n1882,
    n1849,
    n2208
  );


  xnor
  g2232
  (
    n2402,
    n2182,
    n1852,
    n2219
  );


  nor
  g2233
  (
    n2423,
    n1855,
    n1869,
    n2164
  );


  nor
  g2234
  (
    n2294,
    n2160,
    n2178,
    n2184
  );


  xnor
  g2235
  (
    n2532,
    n1888,
    n1879,
    n1830
  );


  nor
  g2236
  (
    n2528,
    n2248,
    n1923,
    n2142
  );


  nor
  g2237
  (
    n2295,
    n1858,
    n1892,
    n2247
  );


  and
  g2238
  (
    n2483,
    n1913,
    n2193,
    n2162
  );


  xnor
  g2239
  (
    n2530,
    n2187,
    n2190,
    n2203
  );


  xnor
  g2240
  (
    n2488,
    n1913,
    n2197,
    n1870
  );


  nand
  g2241
  (
    n2420,
    n1844,
    n2181,
    n2188
  );


  and
  g2242
  (
    n2514,
    n2256,
    n1923,
    n1875
  );


  nand
  g2243
  (
    n2397,
    n2153,
    n1823,
    n1922
  );


  xor
  g2244
  (
    n2355,
    n2250,
    n1912,
    n1849
  );


  nand
  g2245
  (
    n2484,
    n2192,
    n988,
    n2161
  );


  xor
  g2246
  (
    n2446,
    n989,
    n1861,
    n2171
  );


  or
  g2247
  (
    n2512,
    n2262,
    n1910,
    n2162
  );


  or
  g2248
  (
    n2385,
    n985,
    n2262,
    n2156,
    n2069
  );


  nand
  g2249
  (
    n2418,
    n1933,
    n2154,
    n2179,
    n1911
  );


  or
  g2250
  (
    n2474,
    n1860,
    n985,
    n2167,
    n1905
  );


  or
  g2251
  (
    n2425,
    n364,
    n2259,
    n1890,
    n2254
  );


  or
  g2252
  (
    n2324,
    n1866,
    n1889,
    n1881,
    n1844
  );


  nand
  g2253
  (
    n2279,
    n2237,
    n987,
    n1902,
    n1877
  );


  or
  g2254
  (
    n2305,
    n2158,
    n2170,
    n2207,
    n2187
  );


  nand
  g2255
  (
    n2524,
    n1885,
    n1867,
    n2168,
    n2241
  );


  xor
  g2256
  (
    n2431,
    n1864,
    n2168,
    n2252,
    n2239
  );


  or
  g2257
  (
    n2478,
    n1823,
    n2239,
    n1833,
    n2251
  );


  xnor
  g2258
  (
    n2445,
    n1924,
    n2208,
    n2142,
    n2193
  );


  nand
  g2259
  (
    n2400,
    n2184,
    n365,
    n2155,
    n1863
  );


  nand
  g2260
  (
    n2353,
    n2226,
    n2182,
    n2181,
    n1901
  );


  nand
  g2261
  (
    n2343,
    n2230,
    n2186,
    n983,
    n990
  );


  xnor
  g2262
  (
    n2471,
    n2162,
    n2205,
    n2165,
    n2160
  );


  nand
  g2263
  (
    n2510,
    n1835,
    n1832,
    n2189,
    n2232
  );


  nor
  g2264
  (
    n2292,
    n2210,
    n2145,
    n2259,
    n2152
  );


  and
  g2265
  (
    n2470,
    n1884,
    n2196,
    n1868,
    n1932
  );


  nor
  g2266
  (
    n2366,
    n2227,
    n1938,
    n1933,
    n2237
  );


  nand
  g2267
  (
    n2289,
    n2221,
    n2213,
    n2222,
    n2182
  );


  nor
  g2268
  (
    n2274,
    n1914,
    n1914,
    n2205,
    n1874
  );


  nand
  g2269
  (
    n2370,
    n1856,
    n2238,
    n1920,
    n1883
  );


  xnor
  g2270
  (
    n2298,
    n2261,
    n1836,
    n2263,
    n1918
  );


  and
  g2271
  (
    n2513,
    n2249,
    n1924,
    n1868,
    n1891
  );


  nand
  g2272
  (
    n2413,
    n986,
    n2178,
    n2186,
    n1840
  );


  xor
  g2273
  (
    n2403,
    n1927,
    n2153,
    n2169,
    n1891
  );


  or
  g2274
  (
    n2395,
    n2227,
    n2213,
    n1872,
    n2189
  );


  xnor
  g2275
  (
    n2500,
    n1905,
    n2232,
    n1898,
    n1908
  );


  or
  g2276
  (
    n2509,
    n2187,
    n363,
    n2269,
    n2164
  );


  or
  g2277
  (
    n2316,
    n1937,
    n2158,
    n2244,
    n1890
  );


  xor
  g2278
  (
    n2365,
    n2177,
    n2190,
    n1866,
    n2194
  );


  xor
  g2279
  (
    n2497,
    n2211,
    n2183,
    n2227,
    n2255
  );


  xor
  g2280
  (
    n2498,
    n1914,
    n1841,
    n1919,
    n2245
  );


  nor
  g2281
  (
    n2270,
    n1853,
    n1881,
    n1935,
    n2251
  );


  nor
  g2282
  (
    n2363,
    n1900,
    n986,
    n2265,
    n1919
  );


  or
  g2283
  (
    n2293,
    n1873,
    n1855,
    n1833,
    n1896
  );


  xnor
  g2284
  (
    n2520,
    n1888,
    n2236,
    n1879,
    n1850
  );


  xor
  g2285
  (
    n2318,
    n981,
    n1869,
    n1847,
    n1925
  );


  and
  g2286
  (
    n2384,
    n2206,
    n2202,
    n2191,
    n2220
  );


  and
  g2287
  (
    n2281,
    n1928,
    n984,
    n1845,
    n362
  );


  nand
  g2288
  (
    n2329,
    n2261,
    n1865,
    n1930,
    n2256
  );


  or
  g2289
  (
    n2278,
    n2152,
    n2238,
    n2205,
    n1826
  );


  nand
  g2290
  (
    n2301,
    n2188,
    n1831,
    n1896,
    n2235
  );


  nand
  g2291
  (
    n2522,
    n2197,
    n990,
    n2253,
    n1878
  );


  xor
  g2292
  (
    n2495,
    n2191,
    n2231,
    n1884,
    n1834
  );


  xor
  g2293
  (
    n2439,
    n991,
    n1863,
    n1901,
    n1825
  );


  nand
  g2294
  (
    n2482,
    n1851,
    n1921,
    n1835,
    n2248
  );


  or
  g2295
  (
    n2427,
    n2180,
    n2212,
    n980,
    n1830
  );


  xor
  g2296
  (
    n2409,
    n1893,
    n1897,
    n1838,
    n1850
  );


  and
  g2297
  (
    n2472,
    n2194,
    n1858,
    n1838,
    n2243
  );


  or
  g2298
  (
    n2393,
    n1928,
    n1860,
    n1911,
    n2148
  );


  xor
  g2299
  (
    n2473,
    n1939,
    n1888,
    n1831,
    n1903
  );


  xnor
  g2300
  (
    n2436,
    n2171,
    n989,
    n1861,
    n1853
  );


  xnor
  g2301
  (
    n2280,
    n1829,
    n1854,
    n1931,
    n1840
  );


  xor
  g2302
  (
    n2376,
    n2196,
    n988,
    n1876,
    n1889
  );


  nand
  g2303
  (
    n2531,
    n1882,
    n2212,
    n1916,
    n2261
  );


  and
  g2304
  (
    n2290,
    n2157,
    n1857,
    n1861,
    n1931
  );


  nor
  g2305
  (
    n2306,
    n2230,
    n1842,
    n1878
  );


  and
  g2306
  (
    n2330,
    n1897,
    n2145,
    n1869,
    n2197
  );


  xnor
  g2307
  (
    n2372,
    n983,
    n1840,
    n2262,
    n2248
  );


  nor
  g2308
  (
    n2358,
    n2196,
    n2229,
    n2264,
    n1914
  );


  nor
  g2309
  (
    n2391,
    n2239,
    n1879,
    n2249,
    n2159
  );


  xnor
  g2310
  (
    KeyWire_0_25,
    n2201,
    n1831,
    n2183,
    n1855
  );


  nor
  g2311
  (
    n2388,
    n1827,
    n2234,
    n1831,
    n2151
  );


  xor
  g2312
  (
    n2492,
    n1827,
    n2173,
    n1848,
    n2068
  );


  or
  g2313
  (
    n2504,
    n2191,
    n1838,
    n2268,
    n1920
  );


  xor
  g2314
  (
    n2417,
    n2218,
    n2214,
    n2182,
    n2175
  );


  xnor
  g2315
  (
    n2369,
    n2249,
    n1910,
    n2267,
    n1897
  );


  xor
  g2316
  (
    n2311,
    n1837,
    n2268,
    n1876,
    n2233
  );


  and
  g2317
  (
    n2455,
    n1934,
    n2185,
    n983,
    n2169
  );


  nand
  g2318
  (
    n2435,
    n1865,
    n1864,
    n1894,
    n2269
  );


  and
  g2319
  (
    n2379,
    n2199,
    n2212,
    n2147,
    n2242
  );


  nand
  g2320
  (
    n2422,
    n2167,
    n2267,
    n2175,
    n2160
  );


  xnor
  g2321
  (
    n2407,
    n1837,
    n2179,
    n1851,
    n1825
  );


  and
  g2322
  (
    n2414,
    n2151,
    n2266,
    n1839,
    n1892
  );


  and
  g2323
  (
    n2377,
    n2157,
    n2166,
    n1900,
    n2216
  );


  and
  g2324
  (
    n2399,
    n1860,
    n2229,
    n2220,
    n2224
  );


  xnor
  g2325
  (
    n2456,
    n1892,
    n1832,
    n2221,
    n2246
  );


  nor
  g2326
  (
    n2354,
    n2242,
    n2183,
    n2172,
    n2165
  );


  xor
  g2327
  (
    n2309,
    n2176,
    n1916,
    n2152,
    n2248
  );


  nor
  g2328
  (
    n2516,
    n1857,
    n2252,
    n2237,
    n2144
  );


  xnor
  g2329
  (
    n2338,
    n2172,
    n1874,
    n1908,
    n2255
  );


  xor
  g2330
  (
    n2421,
    n1880,
    n985,
    n2144,
    n2210
  );


  and
  g2331
  (
    n2382,
    n1919,
    n1868,
    n2168,
    n2206
  );


  or
  g2332
  (
    n2493,
    n2240,
    n2244,
    n1926,
    n1840
  );


  nand
  g2333
  (
    n2442,
    n1874,
    n2244,
    n1929,
    n1918
  );


  xor
  g2334
  (
    n2273,
    n2185,
    n2195,
    n1830,
    n2158
  );


  nand
  g2335
  (
    n2538,
    n1882,
    n2166,
    n2215,
    n1902
  );


  and
  g2336
  (
    n2347,
    n2162,
    n2257,
    n2146,
    n2200
  );


  xor
  g2337
  (
    n2272,
    n1875,
    n992,
    n1886,
    n2172
  );


  nor
  g2338
  (
    n2428,
    n2268,
    n2200,
    n1918,
    n2150
  );


  xor
  g2339
  (
    n2464,
    n1863,
    n1938,
    n1927,
    n2244
  );


  xor
  g2340
  (
    n2450,
    n1904,
    n2154,
    n2231,
    n2219
  );


  nand
  g2341
  (
    n2405,
    n365,
    n365,
    n2171,
    n1909
  );


  or
  g2342
  (
    n2537,
    n1936,
    n1874,
    n1915,
    n1922
  );


  xor
  g2343
  (
    n2394,
    n1828,
    n1883,
    n2174,
    n1846
  );


  and
  g2344
  (
    n2433,
    n1843,
    n2153,
    n1877,
    n1847
  );


  and
  g2345
  (
    n2386,
    n2189,
    n1923,
    n2257,
    n1937
  );


  nor
  g2346
  (
    n2378,
    n1877,
    n2201,
    n2170,
    n1895
  );


  and
  g2347
  (
    n2312,
    n2265,
    n1899,
    n1878,
    n1859
  );


  xnor
  g2348
  (
    n2460,
    n2234,
    n2156,
    n2154,
    n2255
  );


  nand
  g2349
  (
    n2503,
    n1847,
    n2206,
    n982,
    n2179
  );


  xor
  g2350
  (
    n2357,
    n2173,
    n2247,
    n2186,
    n2228
  );


  xor
  g2351
  (
    n2398,
    n1862,
    n2223,
    n1883,
    n2258
  );


  and
  g2352
  (
    n2406,
    n2264,
    n1885,
    n1887,
    n992
  );


  xor
  g2353
  (
    KeyWire_0_41,
    n2228,
    n987,
    n1843,
    n2143
  );


  nor
  g2354
  (
    n2506,
    n2155,
    n1830,
    n1899,
    n1923
  );


  nor
  g2355
  (
    n2302,
    n2177,
    n981,
    n2207,
    n1935
  );


  nand
  g2356
  (
    n2315,
    n1873,
    n2212,
    n2204,
    n2068
  );


  and
  g2357
  (
    n2360,
    n2253,
    n1869,
    n2150,
    n2238
  );


  nand
  g2358
  (
    n2486,
    n2223,
    n1913,
    n2238,
    n2151
  );


  and
  g2359
  (
    n2396,
    n2148,
    n2198,
    n1891,
    n2257
  );


  xor
  g2360
  (
    n2313,
    n1838,
    n2225,
    n982,
    n2143
  );


  xnor
  g2361
  (
    n2415,
    n2163,
    n2264,
    n1917,
    n2195
  );


  nand
  g2362
  (
    n2437,
    n2252,
    n1926,
    n2235,
    n2161
  );


  nor
  g2363
  (
    n2291,
    n2192,
    n2256,
    n2237,
    n2235
  );


  or
  g2364
  (
    n2317,
    n985,
    n2145,
    n364,
    n2165
  );


  nand
  g2365
  (
    n2449,
    n2146,
    n1870,
    n1871,
    n2195
  );


  nor
  g2366
  (
    n2319,
    n2146,
    n2156,
    n2165,
    n2232
  );


  xnor
  g2367
  (
    n2332,
    n2169,
    n1826,
    n984,
    n1912
  );


  xor
  g2368
  (
    n2519,
    n2179,
    n1916,
    n2199,
    n2215
  );


  nand
  g2369
  (
    n2477,
    n1882,
    n1934,
    n1854,
    n1890
  );


  xnor
  g2370
  (
    n2285,
    n2194,
    n2243,
    n1875,
    n2157
  );


  xnor
  g2371
  (
    n2368,
    n2269,
    n2202,
    n1827,
    n1858
  );


  nor
  g2372
  (
    KeyWire_0_54,
    n2211,
    n1833,
    n980,
    n2258
  );


  nor
  g2373
  (
    n2333,
    n2245,
    n2177,
    n2163,
    n989
  );


  and
  g2374
  (
    n2434,
    n1859,
    n1887,
    n1824,
    n2263
  );


  nand
  g2375
  (
    n2462,
    n1836,
    n2149,
    n2175,
    n2185
  );


  xnor
  g2376
  (
    n2481,
    n1880,
    n2186,
    n1929,
    n1850
  );


  xnor
  g2377
  (
    n2381,
    n2204,
    n1921,
    n2225,
    n1936
  );


  xnor
  g2378
  (
    n2539,
    n2192,
    n982,
    n2223,
    n1922
  );


  xnor
  g2379
  (
    n2430,
    n2188,
    n2150,
    n1832,
    n1894
  );


  xnor
  g2380
  (
    n2392,
    n1893,
    n2266,
    n2246,
    n1877
  );


  xnor
  g2381
  (
    n2374,
    n1828,
    n2149,
    n1824,
    n1912
  );


  or
  g2382
  (
    n2467,
    n2226,
    n2261,
    n1841,
    n1862
  );


  xnor
  g2383
  (
    n2331,
    n1865,
    n2247,
    n2159,
    n1828
  );


  xor
  g2384
  (
    n2457,
    n1886,
    n1844,
    n2147,
    n1870
  );


  xnor
  g2385
  (
    n2371,
    n1835,
    n990,
    n1906,
    n1871
  );


  and
  g2386
  (
    n2502,
    n1826,
    n2181,
    n2185,
    n1858
  );


  xor
  g2387
  (
    n2340,
    n2197,
    n1837,
    n1911,
    n1905
  );


  and
  g2388
  (
    n2485,
    n1900,
    n2166,
    n2265,
    n365
  );


  or
  g2389
  (
    n2297,
    n2158,
    n2224,
    n1933,
    n2230
  );


  xnor
  g2390
  (
    n2344,
    n2220,
    n1933,
    n1907,
    n1901
  );


  nand
  g2391
  (
    n2527,
    n1847,
    n2247,
    n2225,
    n2267
  );


  and
  g2392
  (
    n2401,
    n2170,
    n1834,
    n1903,
    n2147
  );


  and
  g2393
  (
    n2380,
    n1900,
    n1881,
    n2196,
    n2200
  );


  nand
  g2394
  (
    n2507,
    n2203,
    n1886,
    n1825,
    n1934
  );


  nand
  g2395
  (
    n2494,
    n2231,
    n1867,
    n1857,
    n2217
  );


  xnor
  g2396
  (
    n2341,
    n1839,
    n2181,
    n1865,
    n2213
  );


  nand
  g2397
  (
    n2505,
    n1824,
    n1868,
    n1937
  );


  and
  g2398
  (
    n2518,
    n2069,
    n1940,
    n2234,
    n2207
  );


  and
  g2399
  (
    n2308,
    n2258,
    n2233,
    n1908,
    n1837
  );


  or
  g2400
  (
    n2349,
    n2161,
    n1913,
    n2229,
    n1928
  );


  nand
  g2401
  (
    n2416,
    n1841,
    n1844,
    n1939,
    n1829
  );


  xnor
  g2402
  (
    n2359,
    n2152,
    n2217,
    n2251,
    n2260
  );


  xor
  g2403
  (
    n2303,
    n2169,
    n1845,
    n2233,
    n1863
  );


  or
  g2404
  (
    n2461,
    n363,
    n1897,
    n2199,
    n1927
  );


  nor
  g2405
  (
    n2286,
    n2221,
    n1911,
    n1893,
    n2260
  );


  or
  g2406
  (
    n2335,
    n362,
    n1894,
    n1906,
    n2228
  );


  xor
  g2407
  (
    n2334,
    n2260,
    n1932,
    n1845,
    n2233
  );


  xnor
  g2408
  (
    n2468,
    n2204,
    n2148,
    n991,
    n2199
  );


  xnor
  g2409
  (
    n2491,
    n992,
    n980,
    n1930,
    n1919
  );


  xor
  g2410
  (
    n2389,
    n2234,
    n2190,
    n1836,
    n1866
  );


  and
  g2411
  (
    n2271,
    n1871,
    n2254,
    n1851,
    n980
  );


  xor
  g2412
  (
    n2487,
    n1883,
    n1859,
    n2211,
    n2176
  );


  xor
  g2413
  (
    n2459,
    n2201,
    n2225,
    n2155,
    n2240
  );


  nand
  g2414
  (
    n2523,
    n2184,
    n2216,
    n1904,
    n2263
  );


  nand
  g2415
  (
    n2517,
    n1878,
    n2221,
    n2214,
    n2258
  );


  or
  g2416
  (
    n2304,
    n2253,
    n1936,
    n1896,
    n1846
  );


  and
  g2417
  (
    n2387,
    n1870,
    n1920,
    n2180,
    n2256
  );


  nand
  g2418
  (
    n2511,
    n1939,
    n2214,
    n1843,
    n2236
  );


  nor
  g2419
  (
    n2501,
    n2164,
    n1829,
    n1849,
    n2246
  );


  xor
  g2420
  (
    n2300,
    n2174,
    n2229,
    n2173,
    n1856
  );


  xnor
  g2421
  (
    n2529,
    n2249,
    n990,
    n2250,
    n2174
  );


  and
  g2422
  (
    n2327,
    n2178,
    n2206,
    n982,
    n1899
  );


  nand
  g2423
  (
    n2276,
    n2163,
    n1898,
    n1871,
    n2240
  );


  or
  g2424
  (
    n2282,
    n1915,
    n1939,
    n2215,
    n2159
  );


  or
  g2425
  (
    n2411,
    n1891,
    n2188,
    n1867,
    n1880
  );


  xnor
  g2426
  (
    n2465,
    n2222,
    n2257,
    n1885,
    n2242
  );


  nand
  g2427
  (
    n2350,
    n1902,
    n2149,
    n1846,
    n986
  );


  xnor
  g2428
  (
    n2339,
    n2243,
    n1932,
    n1841,
    n2216
  );


  xor
  g2429
  (
    n2367,
    n992,
    n2262,
    n1859,
    n1864
  );


  nand
  g2430
  (
    n2453,
    n1879,
    n2266,
    n1898,
    n1915
  );


  nor
  g2431
  (
    n2348,
    n1888,
    n1867,
    n2172,
    n1902
  );


  nand
  g2432
  (
    n2479,
    n2265,
    n1926,
    n1842,
    n2142
  );


  and
  g2433
  (
    n2328,
    n1872,
    n2218,
    n2266,
    n2193
  );


  or
  g2434
  (
    n2408,
    n2230,
    n986,
    n1908,
    n2232
  );


  nand
  g2435
  (
    n2536,
    n2254,
    n2068,
    n1848,
    n1845
  );


  xor
  g2436
  (
    n2438,
    n1854,
    n2145,
    n2176,
    n2198
  );


  and
  g2437
  (
    n2424,
    n2224,
    n1853,
    n2240,
    n2210
  );


  or
  g2438
  (
    n2489,
    n2194,
    n1856,
    n2146,
    n1855
  );


  nand
  g2439
  (
    n2351,
    n1886,
    n1852,
    n984,
    n2268
  );


  or
  g2440
  (
    n2288,
    n2180,
    n2219,
    n2208,
    n1872
  );


  nor
  g2441
  (
    n2346,
    n2189,
    n1890,
    n1938,
    n1921
  );


  xnor
  g2442
  (
    n2452,
    n363,
    n2228,
    n1852,
    n2208
  );


  xor
  g2443
  (
    n2526,
    n1930,
    n1889,
    n1904,
    n1895
  );


  nor
  g2444
  (
    n2337,
    n1904,
    n1924,
    n2250,
    n1936
  );


  xor
  g2445
  (
    n2451,
    n1848,
    n1938,
    n1931,
    n2202
  );


  and
  g2446
  (
    n2454,
    n2149,
    n1903,
    n1920,
    n1887
  );


  xor
  g2447
  (
    n2535,
    n2191,
    n2259,
    n2220,
    n1917
  );


  xnor
  g2448
  (
    n2533,
    n2198,
    n2260,
    n2153,
    n2144
  );


  xnor
  g2449
  (
    n2373,
    n1876,
    n1925,
    n2245,
    n1899
  );


  and
  g2450
  (
    n2364,
    n1852,
    n1909,
    n1833,
    n1826
  );


  xnor
  g2451
  (
    n2448,
    n2236,
    n1928,
    n2143,
    n991
  );


  nand
  g2452
  (
    n2419,
    n1895,
    n1903,
    n2222,
    n1864
  );


  nor
  g2453
  (
    n2336,
    n2251,
    n2193,
    n2204,
    n1905
  );


  xnor
  g2454
  (
    n2310,
    n2209,
    n1857,
    n1832,
    n2241
  );


  xor
  g2455
  (
    n2432,
    n2219,
    n1827,
    n2236,
    n1917
  );


  nor
  g2456
  (
    n2326,
    n1887,
    n2209,
    n2069
  );


  xor
  g2457
  (
    n2410,
    n1861,
    n1927,
    n1898,
    n1925
  );


  xnor
  g2458
  (
    n2383,
    n1884,
    n2213,
    n1834,
    n2210
  );


  nand
  g2459
  (
    n2440,
    n2171,
    n1930,
    n1894,
    n1876
  );


  nor
  g2460
  (
    n2362,
    n2178,
    n981,
    n2215,
    n1935
  );


  nor
  g2461
  (
    n2345,
    n2176,
    n987,
    n2226,
    n2241
  );


  nand
  g2462
  (
    n2283,
    n989,
    n2252,
    n364,
    n1931
  );


  xnor
  g2463
  (
    n2277,
    n1851,
    n1872,
    n1907,
    n984
  );


  or
  g2464
  (
    n2515,
    n2231,
    n1824,
    n2156,
    n2150
  );


  nor
  g2465
  (
    n2321,
    n1854,
    n2198,
    n1895,
    n2155
  );


  and
  g2466
  (
    n2466,
    n2154,
    n987,
    n1839,
    n1849
  );


  xor
  g2467
  (
    n2296,
    n2170,
    n2227,
    n2209,
    n988
  );


  or
  g2468
  (
    n2342,
    n2192,
    n2201,
    n2190,
    n2174
  );


  xor
  g2469
  (
    n2287,
    n1835,
    n1918,
    n2168,
    n1910
  );


  xor
  g2470
  (
    n2463,
    n2164,
    n2218,
    n1917,
    n363
  );


  xnor
  g2471
  (
    n2525,
    n1925,
    n983,
    n2195,
    n2223
  );


  nor
  g2472
  (
    n2390,
    n1862,
    n1829,
    n2148,
    n1873
  );


  xnor
  g2473
  (
    n2323,
    n1885,
    n2147,
    n2241,
    n2151
  );


  xnor
  g2474
  (
    n2534,
    n2239,
    n1926,
    n2163,
    n2250
  );


  nand
  g2475
  (
    n2480,
    n2218,
    n2224,
    n1909,
    n1906
  );


  nor
  g2476
  (
    n2314,
    n1932,
    n1915,
    n2203,
    n2217
  );


  nand
  g2477
  (
    n2476,
    n2167,
    n1842,
    n1836,
    n1884
  );


  or
  g2478
  (
    n2356,
    n1853,
    n1875,
    n2203,
    n2222
  );


  nand
  g2479
  (
    n2426,
    n2246,
    n1907,
    n2205,
    n2157
  );


  nand
  g2480
  (
    n2284,
    n1860,
    n2259,
    n2211,
    n2217
  );


  or
  g2481
  (
    n2458,
    n2184,
    n1839,
    n1909,
    n1901
  );


  or
  g2482
  (
    n2404,
    n2142,
    n2245,
    n2253,
    n1889
  );


  or
  g2483
  (
    n2412,
    n2255,
    n1843,
    n2200,
    n2263
  );


  and
  g2484
  (
    n2429,
    n1912,
    n1856,
    n2267,
    n1873
  );


  and
  g2485
  (
    n2320,
    n364,
    n2264,
    n2235,
    n1910
  );


  nand
  g2486
  (
    n2490,
    n1862,
    n2173,
    n2068,
    n1828
  );


  nor
  g2487
  (
    n2361,
    n2216,
    n2226,
    n2269,
    n2177
  );


  nor
  g2488
  (
    n2322,
    n2183,
    n1929,
    n2143,
    n1881
  );


  and
  g2489
  (
    n2499,
    n1935,
    n1906,
    n2214,
    n988
  );


  buf
  g2490
  (
    n2557,
    n2315
  );


  not
  g2491
  (
    n2560,
    n2285
  );


  not
  g2492
  (
    n2563,
    n2298
  );


  buf
  g2493
  (
    n2541,
    n2276
  );


  buf
  g2494
  (
    n2558,
    n2283
  );


  buf
  g2495
  (
    n2555,
    n2297
  );


  buf
  g2496
  (
    n2553,
    n2305
  );


  buf
  g2497
  (
    n2552,
    n2310
  );


  buf
  g2498
  (
    n2561,
    n2288
  );


  buf
  g2499
  (
    n2540,
    n2316
  );


  not
  g2500
  (
    n2543,
    n2313
  );


  buf
  g2501
  (
    n2547,
    n2307
  );


  not
  g2502
  (
    n2546,
    n2317
  );


  buf
  g2503
  (
    n2545,
    n2272
  );


  not
  g2504
  (
    n2550,
    n2271
  );


  not
  g2505
  (
    n2559,
    n2312
  );


  xnor
  g2506
  (
    n2548,
    n2304,
    n2292,
    n2306,
    n2278
  );


  and
  g2507
  (
    n2544,
    n2290,
    n2311,
    n2299,
    n2284
  );


  or
  g2508
  (
    n2551,
    n2294,
    n2280,
    n2279,
    n2314
  );


  xnor
  g2509
  (
    n2542,
    n2303,
    n2302,
    n2286,
    n2301
  );


  nor
  g2510
  (
    n2549,
    n2287,
    n2270,
    n2309,
    n2293
  );


  and
  g2511
  (
    n2554,
    n2291,
    n2282,
    n2275,
    n2273
  );


  or
  g2512
  (
    n2562,
    n2281,
    n2308,
    n2277,
    n2274
  );


  xor
  g2513
  (
    n2556,
    n2296,
    n2300,
    n2289,
    n2295
  );


  nor
  g2514
  (
    n2565,
    n2541,
    n2326,
    n2540,
    n2321
  );


  xnor
  g2515
  (
    n2566,
    n2319,
    n2325,
    n2327,
    n2320
  );


  nor
  g2516
  (
    n2567,
    n2318,
    n2328,
    n2329,
    n2542
  );


  and
  g2517
  (
    n2564,
    n2324,
    n2543,
    n2322,
    n2323
  );


  and
  g2518
  (
    n2574,
    n2554,
    n2550,
    n2548,
    n2546
  );


  and
  g2519
  (
    n2572,
    n2565,
    n2566,
    n2555
  );


  xnor
  g2520
  (
    n2570,
    n2552,
    n2555,
    n2554,
    n2565
  );


  and
  g2521
  (
    n2571,
    n2545,
    n2547,
    n2555,
    n2553
  );


  or
  g2522
  (
    n2569,
    n2544,
    n2567,
    n2553,
    n2564
  );


  and
  g2523
  (
    n2568,
    n2553,
    n2553,
    n2549,
    n2551
  );


  or
  g2524
  (
    n2573,
    n2567,
    n2554,
    n2566
  );


  xnor
  g2525
  (
    n2588,
    n2333,
    n2365,
    n2362,
    n2388
  );


  xnor
  g2526
  (
    n2583,
    n2388,
    n2373,
    n2375,
    n2391
  );


  or
  g2527
  (
    n2601,
    n2570,
    n2374,
    n2574,
    n2572
  );


  xor
  g2528
  (
    n2592,
    n2569,
    n2381,
    n2350
  );


  nor
  g2529
  (
    n2598,
    n2389,
    n2380,
    n2382,
    n2374
  );


  xor
  g2530
  (
    KeyWire_0_6,
    n2348,
    n2367,
    n2353,
    n2361
  );


  xnor
  g2531
  (
    n2587,
    n2334,
    n2377,
    n2574,
    n2383
  );


  nand
  g2532
  (
    n2584,
    n2337,
    n2345,
    n2382,
    n2379
  );


  xor
  g2533
  (
    n2591,
    n2338,
    n2573,
    n2569,
    n2375
  );


  xnor
  g2534
  (
    n2599,
    n2354,
    n2360,
    n2570,
    n2389
  );


  or
  g2535
  (
    n2576,
    n2358,
    n2340,
    n2570,
    n2569
  );


  nor
  g2536
  (
    n2596,
    n2387,
    n2383,
    n2371,
    n2372
  );


  xor
  g2537
  (
    n2597,
    n2572,
    n2356,
    n2343,
    n2330
  );


  xnor
  g2538
  (
    n2594,
    n2572,
    n2377,
    n2573,
    n2369
  );


  or
  g2539
  (
    n2577,
    n2363,
    n2571,
    n2376,
    n2573
  );


  nor
  g2540
  (
    n2578,
    n2346,
    n2368,
    n2571,
    n2372
  );


  nor
  g2541
  (
    n2585,
    n2347,
    n2573,
    n2385,
    n2331
  );


  xor
  g2542
  (
    n2581,
    n2344,
    n2380,
    n2568
  );


  and
  g2543
  (
    n2582,
    n2390,
    n2378,
    n2568,
    n2572
  );


  nor
  g2544
  (
    KeyWire_0_42,
    n2359,
    n2370,
    n2339,
    n2351
  );


  or
  g2545
  (
    n2579,
    n2376,
    n2341,
    n2574,
    n2357
  );


  and
  g2546
  (
    n2600,
    n2384,
    n2570,
    n2574,
    n2390
  );


  nand
  g2547
  (
    n2575,
    n2370,
    n2569,
    n2384,
    n2352
  );


  xor
  g2548
  (
    KeyWire_0_20,
    n2364,
    n2366,
    n2349,
    n2391
  );


  xnor
  g2549
  (
    n2586,
    n2355,
    n2342,
    n2332,
    n2386
  );


  and
  g2550
  (
    n2589,
    n2385,
    n2373,
    n2371,
    n2571
  );


  nor
  g2551
  (
    n2602,
    n2378,
    n2379,
    n2336,
    n2387
  );


  xor
  g2552
  (
    n2590,
    n2335,
    n2568,
    n2571,
    n2386
  );


  buf
  g2553
  (
    n2604,
    n2577
  );


  xor
  g2554
  (
    n2603,
    n2392,
    n2576
  );


  and
  g2555
  (
    n2605,
    n2392,
    n2575
  );


  xnor
  g2556
  (
    n2607,
    n2603,
    n2557,
    n2556
  );


  nand
  g2557
  (
    n2606,
    n2557,
    n2556,
    n2604
  );


  or
  g2558
  (
    n2612,
    n2607,
    n163
  );


  xor
  g2559
  (
    n2611,
    n161,
    n162,
    n2394
  );


  xor
  g2560
  (
    n2610,
    n2606,
    n2393,
    n162
  );


  nor
  g2561
  (
    n2608,
    n163,
    n2607,
    n162
  );


  xor
  g2562
  (
    n2609,
    n161,
    n2393,
    n163,
    n2607
  );


  or
  g2563
  (
    n2614,
    n2395,
    n2609,
    n2396
  );


  nand
  g2564
  (
    n2615,
    n2608,
    n2400,
    n2399,
    n2402
  );


  xnor
  g2565
  (
    n2613,
    n2402,
    n2397
  );


  or
  g2566
  (
    n2617,
    n2398,
    n2401,
    n2400
  );


  xor
  g2567
  (
    n2616,
    n2403,
    n2402,
    n2608,
    n2609
  );


  or
  g2568
  (
    n2619,
    n2398,
    n2609,
    n2608,
    n2403
  );


  and
  g2569
  (
    n2618,
    n2395,
    n2394,
    n2399,
    n2608
  );


  or
  g2570
  (
    n2620,
    n2558,
    n2616,
    n2557,
    n2619
  );


  xor
  g2571
  (
    n2623,
    n2618,
    n2559
  );


  xnor
  g2572
  (
    n2622,
    n2617,
    n2560,
    n2558
  );


  nor
  g2573
  (
    n2621,
    n2559,
    n2558,
    n2557
  );


  nor
  g2574
  (
    n2625,
    n2621,
    n2404,
    n2405
  );


  nand
  g2575
  (
    n2624,
    n2620,
    n2403,
    n2404
  );


  xnor
  g2576
  (
    n2626,
    n2622,
    n2404,
    n2405
  );


  nor
  g2577
  (
    n2627,
    n2561,
    n2624,
    n2560
  );


  xnor
  g2578
  (
    n2628,
    n2627,
    n2627,
    n2580,
    n2589
  );


  nand
  g2579
  (
    n2630,
    n2587,
    n2588,
    n2627,
    n2581
  );


  nor
  g2580
  (
    n2629,
    n2627,
    n2579,
    n2578,
    n2585
  );


  or
  g2581
  (
    n2631,
    n2583,
    n2582,
    n2584,
    n2586
  );


  xnor
  g2582
  (
    n2633,
    n2630,
    n2631,
    n2628,
    n2629
  );


  xnor
  g2583
  (
    n2632,
    n2631,
    n2629,
    n2630
  );


  nand
  g2584
  (
    n2634,
    n2629,
    n2629,
    n2590,
    n2630
  );


  nand
  g2585
  (
    n2636,
    n2405,
    n2407,
    n2406
  );


  or
  g2586
  (
    n2635,
    n2406,
    n2406,
    n2633,
    n2632
  );


  or
  g2587
  (
    n2638,
    n2562,
    n2635,
    n2563,
    n2561
  );


  or
  g2588
  (
    n2637,
    n2561,
    n2562,
    n2563
  );


  or
  g2589
  (
    n2639,
    n2562,
    n2636,
    n2561
  );


  or
  g2590
  (
    n2640,
    n2637,
    n2638,
    n2407
  );


  nand
  g2591
  (
    n2641,
    n2407,
    n2408
  );


  and
  g2592
  (
    n2642,
    n2640,
    n2563
  );


  or
  g2593
  (
    n2644,
    n1940,
    n1941,
    n2642
  );


  nand
  g2594
  (
    n2643,
    n1941,
    n1940,
    n2642
  );


  or
  g2595
  (
    n2648,
    n925,
    n2643,
    n1942,
    n1941
  );


  xor
  g2596
  (
    n2646,
    n1943,
    n1942,
    n2643
  );


  or
  g2597
  (
    n2645,
    n1942,
    n926,
    n1012
  );


  xnor
  g2598
  (
    n2647,
    n1943,
    n2643,
    n1942,
    n925
  );


  xnor
  g2599
  (
    n2651,
    n2600,
    n2592,
    n2594,
    n2597
  );


  xnor
  g2600
  (
    n2650,
    n2598,
    n2595,
    n2591,
    n2599
  );


  xnor
  g2601
  (
    n2652,
    n2593,
    n2646,
    n2600,
    n2645
  );


  nand
  g2602
  (
    n2649,
    n2648,
    n2639,
    n2647,
    n2596
  );


  or
  g2603
  (
    n2665,
    n741,
    n2612,
    n1056,
    n2610
  );


  xnor
  g2604
  (
    n2662,
    n2601,
    n2610,
    n2650,
    n2602
  );


  nand
  g2605
  (
    n2656,
    n1012,
    n2605,
    n1056,
    n2611
  );


  xor
  g2606
  (
    n2653,
    n2602,
    n2602,
    n2649,
    n865
  );


  nor
  g2607
  (
    n2661,
    n2612,
    n866,
    n740
  );


  nor
  g2608
  (
    n2655,
    n1055,
    n2641,
    n2601,
    n2602
  );


  xor
  g2609
  (
    n2663,
    n2612,
    n866,
    n2652
  );


  and
  g2610
  (
    n2666,
    n2651,
    n2650,
    n741
  );


  xor
  g2611
  (
    n2659,
    n2651,
    n1055,
    n2650,
    n865
  );


  and
  g2612
  (
    KeyWire_0_51,
    n2609,
    n2610,
    n2651,
    n2652
  );


  xor
  g2613
  (
    n2658,
    n2611,
    n1055,
    n2610,
    n2634
  );


  nand
  g2614
  (
    n2668,
    n1012,
    n2652,
    n2649
  );


  nand
  g2615
  (
    n2654,
    n866,
    n2650,
    n1012,
    n865
  );


  and
  g2616
  (
    n2657,
    n865,
    n1055,
    n2601
  );


  xor
  g2617
  (
    n2660,
    n2611,
    n2651,
    n2612,
    n741
  );


  nor
  g2618
  (
    n2667,
    n2649,
    n2649,
    n2611,
    n2563
  );


  nand
  g2619
  (
    n2669,
    n2655,
    n2654,
    n2656,
    n2653
  );


  xnor
  g2620
  (
    n2670,
    n2658,
    n2657,
    n2631
  );


  or
  g2621
  (
    n2671,
    n2623,
    n2670,
    n2644,
    n2659
  );


  and
  g2622
  (
    n2672,
    n2669,
    n2644
  );


  xor
  g2623
  (
    n2677,
    n2671,
    n2671,
    n1063,
    n1056
  );


  and
  g2624
  (
    n2676,
    n2667,
    n2666,
    n1064,
    n1056
  );


  nand
  g2625
  (
    n2679,
    n2664,
    n1063,
    n2672
  );


  nor
  g2626
  (
    n2673,
    n2069,
    n1062,
    n2660,
    n2626
  );


  xnor
  g2627
  (
    n2678,
    n2668,
    n1063,
    n2662,
    n2408
  );


  nor
  g2628
  (
    n2675,
    n2671,
    n2672,
    n1062
  );


  nor
  g2629
  (
    n2674,
    n2671,
    n2661,
    n1062
  );


  xor
  g2630
  (
    n2680,
    n2663,
    n2625,
    n2665,
    n2672
  );


  buf
  g2631
  (
    n2681,
    n2675
  );


  not
  g2632
  (
    n2683,
    n2673
  );


  not
  g2633
  (
    n2682,
    n2674
  );


  buf
  g2634
  (
    n2684,
    n2676
  );


  xnor
  g2635
  (
    n2690,
    n1951,
    n1943,
    n1949
  );


  xor
  g2636
  (
    n2687,
    n2683,
    n1945,
    n2682
  );


  or
  g2637
  (
    n2688,
    n2677,
    n1950,
    n1952,
    n2682
  );


  nor
  g2638
  (
    n2695,
    n2680,
    n1948,
    n1947
  );


  and
  g2639
  (
    n2693,
    n2681,
    n2681,
    n2683,
    n1950
  );


  xor
  g2640
  (
    n2692,
    n1945,
    n2679,
    n2681,
    n1951
  );


  xnor
  g2641
  (
    n2685,
    n1949,
    n1946,
    n1948
  );


  xnor
  g2642
  (
    n2698,
    n2682,
    n1946,
    n2684
  );


  or
  g2643
  (
    n2697,
    n1945,
    n1945,
    n1949,
    n2683
  );


  nand
  g2644
  (
    n2694,
    n2678,
    n1952,
    n1944
  );


  xor
  g2645
  (
    n2686,
    n1948,
    n2679,
    n2677
  );


  nand
  g2646
  (
    n2691,
    n1947,
    n2679,
    n1946,
    n2684
  );


  xnor
  g2647
  (
    n2699,
    n1944,
    n1944,
    n2680,
    n1946
  );


  xor
  g2648
  (
    n2700,
    n1947,
    n1951,
    n2683,
    n2684
  );


  nor
  g2649
  (
    n2689,
    n2678,
    n1952,
    n1944,
    n1943
  );


  or
  g2650
  (
    n2696,
    n1951,
    n1950,
    n2681
  );


  not
  g2651
  (
    n2706,
    n1175
  );


  not
  g2652
  (
    n2707,
    n1174
  );


  nor
  g2653
  (
    n2705,
    n1175,
    n1174
  );


  xor
  g2654
  (
    n2704,
    n1174,
    n2688
  );


  nand
  g2655
  (
    KeyWire_0_56,
    n2689,
    n2693
  );


  xnor
  g2656
  (
    n2702,
    n2692,
    n2691
  );


  or
  g2657
  (
    n2708,
    n1175,
    n2686
  );


  xor
  g2658
  (
    n2703,
    n2687,
    n2685
  );


  and
  g2659
  (
    n2709,
    n1175,
    n2690
  );


  nand
  g2660
  (
    n2740,
    n2699,
    n1065,
    n2702,
    n2694
  );


  or
  g2661
  (
    n2711,
    n1065,
    n2701,
    n2706,
    n2418
  );


  nor
  g2662
  (
    n2741,
    n2424,
    n2423,
    n1065
  );


  or
  g2663
  (
    n2717,
    n2410,
    n2709,
    n2416,
    n2420
  );


  and
  g2664
  (
    n2728,
    n2410,
    n2417,
    n2432,
    n2705
  );


  xnor
  g2665
  (
    n2727,
    n2421,
    n1064,
    n2414,
    n2703
  );


  and
  g2666
  (
    n2725,
    n2429,
    n2419,
    n2413,
    n2415
  );


  nand
  g2667
  (
    n2738,
    n2426,
    n2698,
    n2411
  );


  nand
  g2668
  (
    n2732,
    n2425,
    n2421,
    n2704,
    n2411
  );


  and
  g2669
  (
    n2729,
    n2413,
    n2410,
    n2418,
    n2430
  );


  and
  g2670
  (
    n2745,
    n2427,
    n2413,
    n2707,
    n2431
  );


  xnor
  g2671
  (
    n2716,
    n2426,
    n2709,
    n2707,
    n2705
  );


  nor
  g2672
  (
    n2722,
    n2424,
    n2708,
    n2426
  );


  and
  g2673
  (
    n2718,
    n2428,
    n2431,
    n2703,
    n2416
  );


  and
  g2674
  (
    n2730,
    n2412,
    n2416,
    n2425,
    n1064
  );


  nor
  g2675
  (
    n2714,
    n2704,
    n2697,
    n2430,
    n2420
  );


  xnor
  g2676
  (
    n2712,
    n2412,
    n2427,
    n2415,
    n2431
  );


  or
  g2677
  (
    n2724,
    n2700,
    n2429,
    n2701
  );


  or
  g2678
  (
    n2723,
    n2432,
    n2703,
    n2419,
    n2706
  );


  and
  g2679
  (
    n2744,
    n2423,
    n2412,
    n2414,
    n2425
  );


  nand
  g2680
  (
    n2710,
    n2413,
    n2706,
    n2416,
    n2428
  );


  or
  g2681
  (
    n2731,
    n2424,
    n2708,
    n2414,
    n2420
  );


  xnor
  g2682
  (
    n2743,
    n2702,
    n2409,
    n2415
  );


  and
  g2683
  (
    n2736,
    n2419,
    n2709,
    n2704
  );


  nor
  g2684
  (
    n2726,
    n2707,
    n2703,
    n2422,
    n2417
  );


  and
  g2685
  (
    n2734,
    n2431,
    n2428,
    n2702,
    n2412
  );


  or
  g2686
  (
    n2713,
    n2701,
    n2709,
    n2708,
    n2705
  );


  nor
  g2687
  (
    n2720,
    n2708,
    n1065,
    n2422,
    n2414
  );


  nand
  g2688
  (
    n2739,
    n2430,
    n2422,
    n2419,
    n2705
  );


  or
  g2689
  (
    n2735,
    n2409,
    n2421,
    n2420,
    n2424
  );


  xnor
  g2690
  (
    n2733,
    n2696,
    n2425,
    n2410,
    n2421
  );


  nand
  g2691
  (
    n2715,
    n2702,
    n2415,
    n2417
  );


  nand
  g2692
  (
    n2719,
    n2418,
    n2428,
    n2423,
    n2422
  );


  nand
  g2693
  (
    n2742,
    n2430,
    n2706,
    n2418,
    n2429
  );


  xor
  g2694
  (
    n2737,
    n1064,
    n2409,
    n2427
  );


  xor
  g2695
  (
    n2721,
    n2707,
    n2701,
    n2411,
    n2695
  );


  xor
  g2696
  (
    n2748,
    n2735,
    n2485,
    n2441,
    n2719
  );


  nand
  g2697
  (
    n2783,
    n2435,
    n2493,
    n2728,
    n2717
  );


  xor
  g2698
  (
    n2889,
    n2434,
    n2461,
    n2506,
    n2721
  );


  nand
  g2699
  (
    n2764,
    n2499,
    n2466,
    n2491,
    n2740
  );


  nand
  g2700
  (
    n2749,
    n2494,
    n2713,
    n2501,
    n2727
  );


  nor
  g2701
  (
    n2780,
    n2436,
    n2457,
    n2451,
    n2710
  );


  xnor
  g2702
  (
    n2767,
    n2722,
    n2454,
    n2732,
    n2470
  );


  xnor
  g2703
  (
    n2791,
    n2490,
    n2498,
    n2724,
    n2723
  );


  and
  g2704
  (
    n2883,
    n2434,
    n2737,
    n2461
  );


  xor
  g2705
  (
    n2842,
    n2494,
    n2527,
    n2450,
    n2507
  );


  xor
  g2706
  (
    n2835,
    n2487,
    n2724,
    n2502,
    n2471
  );


  nor
  g2707
  (
    n2817,
    n2716,
    n2734,
    n2515,
    n2680
  );


  or
  g2708
  (
    n2875,
    n2452,
    n2515,
    n2510,
    n2502
  );


  and
  g2709
  (
    n2870,
    n2483,
    n2537,
    n2454,
    n2489
  );


  nor
  g2710
  (
    n2867,
    n2742,
    n2507,
    n2524,
    n2517
  );


  nand
  g2711
  (
    n2761,
    n2513,
    n2482,
    n2458,
    n2465
  );


  and
  g2712
  (
    n2855,
    n2451,
    n2721,
    n2446,
    n2717
  );


  nand
  g2713
  (
    n2811,
    n2505,
    n2730,
    n2448,
    n2442
  );


  or
  g2714
  (
    n2759,
    n2481,
    n2470,
    n2526,
    n2468
  );


  xor
  g2715
  (
    n2768,
    n2744,
    n2488,
    n2492,
    n2533
  );


  or
  g2716
  (
    n2886,
    n2711,
    n2460,
    n2735,
    n2714
  );


  xnor
  g2717
  (
    n2805,
    n2743,
    n2715,
    n2469,
    n2726
  );


  xnor
  g2718
  (
    n2873,
    n2526,
    n2460,
    n2506,
    n2505
  );


  and
  g2719
  (
    n2782,
    n2450,
    n2449,
    n2529,
    n2480
  );


  nor
  g2720
  (
    n2844,
    n2476,
    n2738,
    n2727,
    n2534
  );


  nor
  g2721
  (
    n2752,
    n2474,
    n2718,
    n2484,
    n2532
  );


  nor
  g2722
  (
    n2884,
    n2537,
    n2463,
    n2720,
    n2739
  );


  nand
  g2723
  (
    n2834,
    n2502,
    n2463,
    n2490
  );


  xnor
  g2724
  (
    n2874,
    n2719,
    n2446,
    n2466
  );


  xor
  g2725
  (
    n2830,
    n2465,
    n2489,
    n2722,
    n2443
  );


  nor
  g2726
  (
    n2845,
    n2451,
    n2724,
    n2459,
    n2463
  );


  nand
  g2727
  (
    n2813,
    n2480,
    n2727,
    n2712,
    n2452
  );


  xor
  g2728
  (
    n2779,
    n2514,
    n2734,
    n2455,
    n2537
  );


  xnor
  g2729
  (
    n2885,
    n2740,
    n2712,
    n2499,
    n2450
  );


  nor
  g2730
  (
    n2887,
    n2485,
    n2733,
    n2515,
    n2503
  );


  or
  g2731
  (
    n2824,
    n2435,
    n2490,
    n2535,
    n2519
  );


  nor
  g2732
  (
    n2831,
    n2457,
    n2744,
    n2497,
    n2451
  );


  nor
  g2733
  (
    n2786,
    n2729,
    n2743,
    n2513,
    n2467
  );


  nor
  g2734
  (
    n2800,
    n2736,
    n2530,
    n2501,
    n2718
  );


  or
  g2735
  (
    n2819,
    n2488,
    n2453,
    n2711,
    n2472
  );


  nor
  g2736
  (
    n2776,
    n2713,
    n2491,
    n2483,
    n2722
  );


  nor
  g2737
  (
    n2829,
    n2525,
    n2734,
    n2477,
    n2713
  );


  or
  g2738
  (
    n2861,
    n2720,
    n2714,
    n2445,
    n2512
  );


  or
  g2739
  (
    n2880,
    n2448,
    n2486,
    n2462,
    n2680
  );


  nor
  g2740
  (
    n2888,
    n2526,
    n2718,
    n2433,
    n2497
  );


  xor
  g2741
  (
    n2823,
    n2521,
    n2739,
    n2490,
    n2535
  );


  or
  g2742
  (
    n2878,
    n2486,
    n2452,
    n2519,
    n2710
  );


  xor
  g2743
  (
    n2832,
    n2437,
    n2441,
    n2442,
    n2450
  );


  and
  g2744
  (
    n2766,
    n2440,
    n2446,
    n2491,
    n2432
  );


  xor
  g2745
  (
    n2857,
    n2507,
    n2488,
    n2509,
    n2499
  );


  xor
  g2746
  (
    n2746,
    n2496,
    n2472,
    n2522,
    n2536
  );


  xor
  g2747
  (
    n2787,
    n2517,
    n2492,
    n2460,
    n2532
  );


  or
  g2748
  (
    n2772,
    n2731,
    n2533,
    n2498,
    n2723
  );


  and
  g2749
  (
    n2784,
    n2496,
    n2721,
    n2433,
    n2471
  );


  nor
  g2750
  (
    n2802,
    n2711,
    n2437,
    n2508,
    n2517
  );


  and
  g2751
  (
    n2762,
    n2460,
    n2469,
    n2472,
    n2532
  );


  xor
  g2752
  (
    n2753,
    n2474,
    n2725,
    n2462
  );


  xnor
  g2753
  (
    n2814,
    n2737,
    n2725,
    n2455,
    n2454
  );


  nor
  g2754
  (
    n2778,
    n2729,
    n2516,
    n2523,
    n2731
  );


  and
  g2755
  (
    n2879,
    n2715,
    n2742,
    n2745,
    n2442
  );


  xnor
  g2756
  (
    n2809,
    n2529,
    n2456,
    n2481,
    n2538
  );


  and
  g2757
  (
    n2852,
    n2466,
    n2519,
    n2493,
    n2445
  );


  nand
  g2758
  (
    n2825,
    n2717,
    n2504,
    n2464,
    n2480
  );


  nor
  g2759
  (
    n2803,
    n2444,
    n2532,
    n2739,
    n2504
  );


  nand
  g2760
  (
    n2765,
    n2738,
    n2475,
    n2433,
    n2534
  );


  nand
  g2761
  (
    n2858,
    n2518,
    n2448,
    n2512,
    n2443
  );


  nor
  g2762
  (
    n2843,
    n2444,
    n2524,
    n2434,
    n2461
  );


  xnor
  g2763
  (
    n2771,
    n2516,
    n2439,
    n2735,
    n2447
  );


  xnor
  g2764
  (
    KeyWire_0_34,
    n2494,
    n2474,
    n2723,
    n2711
  );


  nand
  g2765
  (
    n2785,
    n2508,
    n2473,
    n2455,
    n2459
  );


  and
  g2766
  (
    n2854,
    n2514,
    n2454,
    n2492,
    n2743
  );


  nor
  g2767
  (
    n2850,
    n2458,
    n2441,
    n2521,
    n2438
  );


  xor
  g2768
  (
    n2774,
    n2500,
    n2500,
    n2476,
    n2729
  );


  or
  g2769
  (
    n2763,
    n2742,
    n2478,
    n2712,
    n2524
  );


  xor
  g2770
  (
    n2820,
    n2457,
    n2503,
    n2717,
    n2453
  );


  or
  g2771
  (
    n2841,
    n2474,
    n2458,
    n2487,
    n2433
  );


  nor
  g2772
  (
    KeyWire_0_40,
    n2720,
    n2538,
    n2516,
    n2496
  );


  nand
  g2773
  (
    n2755,
    n2467,
    n2435,
    n2469,
    n2479
  );


  nand
  g2774
  (
    n2796,
    n2453,
    n2506,
    n2713,
    n2443
  );


  nand
  g2775
  (
    n2773,
    n2468,
    n2514,
    n2525,
    n2523
  );


  xor
  g2776
  (
    n2806,
    n2724,
    n2468,
    n2491,
    n2465
  );


  nor
  g2777
  (
    n2860,
    n2471,
    n2468,
    n2531,
    n2440
  );


  and
  g2778
  (
    n2797,
    n2529,
    n2528,
    n2715,
    n2511
  );


  xnor
  g2779
  (
    n2754,
    n2441,
    n2501,
    n2439,
    n2740
  );


  nor
  g2780
  (
    n2821,
    n2726,
    n2727,
    n2484,
    n2523
  );


  or
  g2781
  (
    n2836,
    n2745,
    n2477,
    n2509,
    n2495
  );


  or
  g2782
  (
    n2865,
    n2514,
    n2459,
    n2455,
    n2478
  );


  or
  g2783
  (
    n2839,
    n2457,
    n2447,
    n2459,
    n2475
  );


  xor
  g2784
  (
    n2827,
    n2741,
    n2730,
    n2493,
    n2508
  );


  xnor
  g2785
  (
    n2856,
    n2715,
    n2736,
    n2742,
    n2483
  );


  nor
  g2786
  (
    n2810,
    n2477,
    n2506,
    n2479,
    n2719
  );


  xnor
  g2787
  (
    n2822,
    n2469,
    n2745,
    n2533,
    n2440
  );


  or
  g2788
  (
    n2792,
    n2721,
    n2464,
    n2534,
    n2449
  );


  and
  g2789
  (
    n2794,
    n2481,
    n2732,
    n2443,
    n2479
  );


  nand
  g2790
  (
    n2849,
    n2710,
    n2733,
    n2538,
    n2511
  );


  or
  g2791
  (
    n2770,
    n2744,
    n2501,
    n2504,
    n2533
  );


  and
  g2792
  (
    n2760,
    n2462,
    n2467,
    n2508,
    n2442
  );


  nor
  g2793
  (
    n2747,
    n2448,
    n2513,
    n2444,
    n2480
  );


  and
  g2794
  (
    n2777,
    n2513,
    n2447,
    n2730,
    n2522
  );


  xor
  g2795
  (
    n2788,
    n2528,
    n2720,
    n2505,
    n2525
  );


  xor
  g2796
  (
    n2769,
    n2732,
    n2436,
    n2539
  );


  or
  g2797
  (
    n2807,
    n2488,
    n2729,
    n2518,
    n2516
  );


  nor
  g2798
  (
    KeyWire_0_38,
    n2740,
    n2528,
    n2511,
    n2539
  );


  xnor
  g2799
  (
    n2871,
    n2741,
    n2481,
    n2731,
    n2728
  );


  or
  g2800
  (
    n2838,
    n2486,
    n2725,
    n2728,
    n2517
  );


  or
  g2801
  (
    n2790,
    n2445,
    n2536,
    n2726,
    n2449
  );


  xnor
  g2802
  (
    n2866,
    n2495,
    n2723,
    n2436,
    n2498
  );


  or
  g2803
  (
    n2750,
    n2444,
    n2736,
    n2502,
    n2476
  );


  nor
  g2804
  (
    n2848,
    n2730,
    n2470,
    n2738,
    n2445
  );


  nor
  g2805
  (
    n2812,
    n2531,
    n2435,
    n2475,
    n2438
  );


  or
  g2806
  (
    n2756,
    n2473,
    n2712,
    n2522,
    n2466
  );


  or
  g2807
  (
    n2801,
    n2537,
    n2465,
    n2535,
    n2728
  );


  nor
  g2808
  (
    n2851,
    n2475,
    n2478,
    n2487,
    n2522
  );


  or
  g2809
  (
    n2781,
    n2741,
    n2710,
    n2539,
    n2432
  );


  xnor
  g2810
  (
    n2863,
    n2458,
    n2526,
    n2437,
    n2529
  );


  or
  g2811
  (
    n2799,
    n2484,
    n2510,
    n2527,
    n2520
  );


  or
  g2812
  (
    n2798,
    n2528,
    n2456,
    n2482,
    n2489
  );


  xnor
  g2813
  (
    n2815,
    n2521,
    n2470,
    n2484,
    n2482
  );


  or
  g2814
  (
    n2789,
    n2732,
    n2486,
    n2438,
    n2536
  );


  nor
  g2815
  (
    n2751,
    n2743,
    n2494,
    n2520,
    n2733
  );


  nor
  g2816
  (
    n2816,
    n2437,
    n2734,
    n2536,
    n2519
  );


  and
  g2817
  (
    n2775,
    n2487,
    n2714,
    n2511,
    n2483
  );


  xnor
  g2818
  (
    n2853,
    n2453,
    n2485,
    n2518,
    n2499
  );


  nor
  g2819
  (
    n2758,
    n2512,
    n2504,
    n2733,
    n2523
  );


  and
  g2820
  (
    n2862,
    n2449,
    n2530,
    n2745,
    n2489
  );


  nand
  g2821
  (
    n2846,
    n2527,
    n2521,
    n2456,
    n2493
  );


  nand
  g2822
  (
    n2837,
    n2510,
    n2716,
    n2479,
    n2737
  );


  xnor
  g2823
  (
    n2757,
    n2477,
    n2512,
    n2716,
    n2738
  );


  nor
  g2824
  (
    n2881,
    n2476,
    n2438,
    n2434,
    n2741
  );


  or
  g2825
  (
    n2859,
    n2518,
    n2485,
    n2739,
    n2440
  );


  and
  g2826
  (
    n2868,
    n2472,
    n2718,
    n2714,
    n2473
  );


  xor
  g2827
  (
    n2877,
    n2452,
    n2726,
    n2498,
    n2497
  );


  xor
  g2828
  (
    n2864,
    n2439,
    n2524,
    n2539,
    n2473
  );


  xor
  g2829
  (
    n2872,
    n2478,
    n2722,
    n2515,
    n2495
  );


  nor
  g2830
  (
    n2818,
    n2447,
    n2731,
    n2503
  );


  xor
  g2831
  (
    n2826,
    n2439,
    n2505,
    n2735,
    n2520
  );


  or
  g2832
  (
    n2808,
    n2462,
    n2500,
    n2530,
    n2497
  );


  or
  g2833
  (
    n2833,
    n2495,
    n2716,
    n2482,
    n2525
  );


  nand
  g2834
  (
    n2804,
    n2500,
    n2538,
    n2507,
    n2535
  );


  xnor
  g2835
  (
    n2882,
    n2471,
    n2736,
    n2534,
    n2464
  );


  nor
  g2836
  (
    n2793,
    n2531,
    n2510,
    n2520,
    n2496
  );


  and
  g2837
  (
    n2847,
    n2719,
    n2527,
    n2744,
    n2492
  );


  xnor
  g2838
  (
    n2828,
    n2530,
    n2461,
    n2464,
    n2531
  );


  xnor
  g2839
  (
    n2869,
    n2467,
    n2509,
    n2456
  );


  xnor
  g2840
  (
    n2938,
    n2781,
    n2859,
    n2819,
    n2812
  );


  nand
  g2841
  (
    n2931,
    n2835,
    n2877,
    n2796,
    n2827
  );


  xnor
  g2842
  (
    n2929,
    n2751,
    n2836,
    n2845,
    n2785
  );


  nand
  g2843
  (
    n2922,
    n2884,
    n2845,
    n2804,
    n2838
  );


  nor
  g2844
  (
    n2890,
    n2882,
    n2846,
    n2774,
    n2888
  );


  and
  g2845
  (
    n2948,
    n2828,
    n2802,
    n2860,
    n2883
  );


  nor
  g2846
  (
    KeyWire_0_8,
    n2867,
    n2772,
    n2862,
    n2881
  );


  or
  g2847
  (
    n2909,
    n2756,
    n2816,
    n2794,
    n2852
  );


  or
  g2848
  (
    n2925,
    n2780,
    n2884,
    n2788,
    n2770
  );


  nand
  g2849
  (
    n2895,
    n2878,
    n2857,
    n2876,
    n2820
  );


  nor
  g2850
  (
    n2939,
    n2870,
    n2811,
    n2837,
    n2832
  );


  xnor
  g2851
  (
    n2902,
    n2752,
    n2875,
    n2880,
    n2854
  );


  and
  g2852
  (
    n2913,
    n2838,
    n2881,
    n2849,
    n2753
  );


  nand
  g2853
  (
    n2899,
    n2811,
    n2866,
    n2874,
    n2807
  );


  nor
  g2854
  (
    n2911,
    n2746,
    n2880,
    n2862,
    n2800
  );


  xor
  g2855
  (
    n2950,
    n2826,
    n2876,
    n2802,
    n2869
  );


  or
  g2856
  (
    n2951,
    n2833,
    n2831,
    n2791,
    n2842
  );


  and
  g2857
  (
    n2944,
    n2856,
    n2867,
    n2760,
    n2836
  );


  xnor
  g2858
  (
    n2952,
    n2889,
    n2824,
    n2847,
    n2812
  );


  and
  g2859
  (
    n2907,
    n2866,
    n2776,
    n2834,
    n2886
  );


  and
  g2860
  (
    n2937,
    n2885,
    n2878,
    n2879,
    n2821
  );


  nor
  g2861
  (
    n2896,
    n2843,
    n2844,
    n2801,
    n2871
  );


  xor
  g2862
  (
    n2910,
    n2883,
    n2848,
    n2830
  );


  xor
  g2863
  (
    n2916,
    n2754,
    n2825,
    n2824,
    n2813
  );


  xnor
  g2864
  (
    n2892,
    n2854,
    n2793,
    n2840,
    n2883
  );


  nor
  g2865
  (
    n2940,
    n2840,
    n2810,
    n2881,
    n2879
  );


  nand
  g2866
  (
    n2914,
    n2880,
    n2805,
    n2848,
    n2809
  );


  nor
  g2867
  (
    n2915,
    n2822,
    n2889,
    n2818,
    n2750
  );


  and
  g2868
  (
    n2930,
    n2766,
    n2778,
    n2800,
    n2808
  );


  xor
  g2869
  (
    n2904,
    n2882,
    n2843,
    n2777,
    n2762
  );


  and
  g2870
  (
    n2918,
    n2860,
    n2779,
    n2771,
    n2853
  );


  nand
  g2871
  (
    n2933,
    n2821,
    n2768,
    n2801,
    n2856
  );


  xor
  g2872
  (
    n2923,
    n2884,
    n2826,
    n2846,
    n2858
  );


  or
  g2873
  (
    n2897,
    n2852,
    n2818,
    n2839,
    n2825
  );


  xnor
  g2874
  (
    n2932,
    n2815,
    n2808,
    n2881,
    n2885
  );


  and
  g2875
  (
    n2936,
    n2749,
    n2869,
    n2803,
    n2816
  );


  and
  g2876
  (
    n2903,
    n2829,
    n2865,
    n2831,
    n2786
  );


  xor
  g2877
  (
    n2921,
    n2763,
    n2877,
    n2813,
    n2828
  );


  nor
  g2878
  (
    n2891,
    n2787,
    n2775,
    n2874,
    n2764
  );


  xnor
  g2879
  (
    n2893,
    n2855,
    n2887,
    n2872,
    n2769
  );


  and
  g2880
  (
    n2945,
    n2817,
    n2841,
    n2773,
    n2820
  );


  xor
  g2881
  (
    n2949,
    n2759,
    n2757,
    n2814,
    n2868
  );


  xor
  g2882
  (
    n2941,
    n2809,
    n2803,
    n2886,
    n2807
  );


  nor
  g2883
  (
    n2906,
    n2853,
    n2832,
    n2873,
    n2839
  );


  nand
  g2884
  (
    n2946,
    n2810,
    n2789,
    n2761,
    n2790
  );


  nand
  g2885
  (
    n2917,
    n2850,
    n2823,
    n2849,
    n2782
  );


  or
  g2886
  (
    n2919,
    n2870,
    n2857,
    n2842,
    n2868
  );


  xnor
  g2887
  (
    n2926,
    n2887,
    n2880,
    n2882,
    n2872
  );


  xor
  g2888
  (
    n2901,
    n2806,
    n2829,
    n2835,
    n2863
  );


  and
  g2889
  (
    n2927,
    n2884,
    n2889,
    n2834,
    n2783
  );


  xor
  g2890
  (
    n2900,
    n2767,
    n2879,
    n2888,
    n2855
  );


  or
  g2891
  (
    n2905,
    n2864,
    n2889,
    n2863,
    n2850
  );


  xnor
  g2892
  (
    n2953,
    n2792,
    n2887,
    n2841,
    n2888
  );


  and
  g2893
  (
    n2920,
    n2879,
    n2755,
    n2819,
    n2864
  );


  nor
  g2894
  (
    n2894,
    n2865,
    n2837,
    n2888,
    n2822
  );


  or
  g2895
  (
    n2935,
    n2748,
    n2844,
    n2758,
    n2847
  );


  and
  g2896
  (
    n2942,
    n2861,
    n2882,
    n2804,
    n2823
  );


  xor
  g2897
  (
    n2908,
    n2797,
    n2833,
    n2859,
    n2806
  );


  or
  g2898
  (
    n2924,
    n2887,
    n2747,
    n2875,
    n2765
  );


  nand
  g2899
  (
    n2943,
    n2817,
    n2805,
    n2814,
    n2795
  );


  xor
  g2900
  (
    n2898,
    n2886,
    n2784,
    n2858,
    n2815
  );


  xnor
  g2901
  (
    n2912,
    n2827,
    n2851,
    n2883,
    n2885
  );


  xnor
  g2902
  (
    n2934,
    n2799,
    n2886,
    n2851,
    n2861
  );


  nor
  g2903
  (
    n2947,
    n2871,
    n2798,
    n2885,
    n2873
  );


  nor
  g2904
  (
    n2955,
    n2906,
    n2926,
    n2953,
    n2924
  );


  xor
  g2905
  (
    n2960,
    n2914,
    n2905,
    n2937,
    n2947
  );


  nor
  g2906
  (
    n2957,
    n2936,
    n2945,
    n2894,
    n2940
  );


  or
  g2907
  (
    n2967,
    n2917,
    n2913,
    n2948,
    n2898
  );


  nand
  g2908
  (
    n2958,
    n2939,
    n2949,
    n2900,
    n2922
  );


  nor
  g2909
  (
    n2954,
    n2938,
    n2941,
    n2891,
    n2946
  );


  nand
  g2910
  (
    n2959,
    n2943,
    n2950,
    n2942,
    n2920
  );


  or
  g2911
  (
    n2965,
    n2916,
    n2892,
    n2931,
    n2951
  );


  nand
  g2912
  (
    KeyWire_0_37,
    n2911,
    n2925,
    n2935,
    n2896
  );


  and
  g2913
  (
    n2962,
    n2912,
    n2930,
    n2923,
    n2910
  );


  and
  g2914
  (
    n2963,
    n2899,
    n2890,
    n2919,
    n2934
  );


  xor
  g2915
  (
    n2969,
    n2895,
    n2921,
    n2897,
    n2908
  );


  or
  g2916
  (
    n2956,
    n2927,
    n2933,
    n2918,
    n2944
  );


  nor
  g2917
  (
    n2964,
    n2928,
    n2903,
    n2902,
    n2915
  );


  or
  g2918
  (
    n2961,
    n2901,
    n2952,
    n2929,
    n2909
  );


  xor
  g2919
  (
    n2968,
    n2932,
    n2907,
    n2893,
    n2904
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n182,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1138,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n145,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n422,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1968,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1762,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n2593,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1315,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n2928,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n701,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1417,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1864,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n765,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n379,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n418,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1867,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1729,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n960,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n1780,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n611,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n2580,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n2255,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n410,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n779,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1492,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n2275,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n1012,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n626,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n2144,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n899,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n2242,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n750,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n2085,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n1524,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n2876,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n796,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1756,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n2966,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n2795,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n80,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n2840,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n2496,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n2595,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n1176,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n547,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n1569,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n2080,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n1161,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n922,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n2352,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n930,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n2664,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n677,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n610,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n2447,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n1613,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n2701,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n769,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n491,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n444,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n2062,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n1771,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n112,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n1565,
    KeyNOTWire_0_63
  );


endmodule

