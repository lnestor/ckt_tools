

module Stat_1430_17_9
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n208,
  n861,
  n984,
  n1220,
  n1334,
  n1441,
  n1439,
  n1447,
  n1449,
  n1437,
  n1440,
  n1438,
  n1445,
  n1453,
  n1442,
  n1454,
  n1452,
  n1436,
  n1444,
  n1434,
  n1448,
  n1443,
  n1435,
  n1451,
  n1450,
  n1446,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n208;
  output n861;
  output n984;
  output n1220;
  output n1334;
  output n1441;
  output n1439;
  output n1447;
  output n1449;
  output n1437;
  output n1440;
  output n1438;
  output n1445;
  output n1453;
  output n1442;
  output n1454;
  output n1452;
  output n1436;
  output n1444;
  output n1434;
  output n1448;
  output n1443;
  output n1435;
  output n1451;
  output n1450;
  output n1446;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    KeyWire_0_10,
    n1
  );


  buf
  g1
  (
    n36,
    n6
  );


  not
  g2
  (
    n37,
    n5
  );


  buf
  g3
  (
    n86,
    n16
  );


  not
  g4
  (
    n80,
    n21
  );


  not
  g5
  (
    n108,
    n14
  );


  buf
  g6
  (
    n100,
    n12
  );


  not
  g7
  (
    n53,
    n11
  );


  not
  g8
  (
    n90,
    n8
  );


  buf
  g9
  (
    n51,
    n4
  );


  buf
  g10
  (
    n89,
    n1
  );


  not
  g11
  (
    n30,
    n19
  );


  buf
  g12
  (
    n62,
    n21
  );


  buf
  g13
  (
    n63,
    n22
  );


  not
  g14
  (
    n87,
    n9
  );


  buf
  g15
  (
    n45,
    n18
  );


  not
  g16
  (
    n32,
    n3
  );


  not
  g17
  (
    n42,
    n9
  );


  buf
  g18
  (
    n48,
    n14
  );


  not
  g19
  (
    n75,
    n6
  );


  not
  g20
  (
    n102,
    n3
  );


  not
  g21
  (
    n84,
    n7
  );


  buf
  g22
  (
    n33,
    n19
  );


  buf
  g23
  (
    n112,
    n11
  );


  not
  g24
  (
    n41,
    n10
  );


  buf
  g25
  (
    n40,
    n4
  );


  not
  g26
  (
    n47,
    n13
  );


  not
  g27
  (
    n38,
    n16
  );


  buf
  g28
  (
    n106,
    n5
  );


  buf
  g29
  (
    n70,
    n17
  );


  not
  g30
  (
    n101,
    n10
  );


  buf
  g31
  (
    n88,
    n8
  );


  not
  g32
  (
    n52,
    n8
  );


  buf
  g33
  (
    n57,
    n13
  );


  not
  g34
  (
    n94,
    n8
  );


  not
  g35
  (
    n91,
    n12
  );


  buf
  g36
  (
    n69,
    n18
  );


  not
  g37
  (
    n93,
    n17
  );


  not
  g38
  (
    n39,
    n18
  );


  buf
  g39
  (
    n56,
    n2
  );


  buf
  g40
  (
    n76,
    n13
  );


  not
  g41
  (
    n67,
    n10
  );


  not
  g42
  (
    n65,
    n11
  );


  not
  g43
  (
    n109,
    n2
  );


  buf
  g44
  (
    n35,
    n3
  );


  not
  g45
  (
    n95,
    n15
  );


  buf
  g46
  (
    n92,
    n10
  );


  not
  g47
  (
    n54,
    n22
  );


  not
  g48
  (
    n98,
    n7
  );


  buf
  g49
  (
    KeyWire_0_29,
    n18
  );


  buf
  g50
  (
    n82,
    n1
  );


  not
  g51
  (
    n104,
    n19
  );


  buf
  g52
  (
    n72,
    n16
  );


  not
  g53
  (
    n68,
    n5
  );


  not
  g54
  (
    n58,
    n20
  );


  not
  g55
  (
    n46,
    n12
  );


  not
  g56
  (
    n105,
    n16
  );


  not
  g57
  (
    n111,
    n21
  );


  buf
  g58
  (
    n55,
    n14
  );


  buf
  g59
  (
    n59,
    n4
  );


  buf
  g60
  (
    n97,
    n15
  );


  not
  g61
  (
    n81,
    n20
  );


  not
  g62
  (
    n79,
    n6
  );


  not
  g63
  (
    n74,
    n22
  );


  buf
  g64
  (
    n29,
    n9
  );


  buf
  g65
  (
    n60,
    n14
  );


  not
  g66
  (
    n103,
    n7
  );


  not
  g67
  (
    n25,
    n3
  );


  buf
  g68
  (
    n44,
    n1
  );


  buf
  g69
  (
    n61,
    n20
  );


  not
  g70
  (
    n66,
    n7
  );


  buf
  g71
  (
    n31,
    n9
  );


  buf
  g72
  (
    n43,
    n17
  );


  not
  g73
  (
    n27,
    n22
  );


  not
  g74
  (
    n99,
    n5
  );


  buf
  g75
  (
    n73,
    n4
  );


  buf
  g76
  (
    n83,
    n6
  );


  not
  g77
  (
    n96,
    n13
  );


  buf
  g78
  (
    n49,
    n19
  );


  not
  g79
  (
    n26,
    n15
  );


  buf
  g80
  (
    n50,
    n2
  );


  buf
  g81
  (
    n71,
    n21
  );


  not
  g82
  (
    n34,
    n15
  );


  buf
  g83
  (
    n78,
    n17
  );


  not
  g84
  (
    n64,
    n2
  );


  not
  g85
  (
    n110,
    n12
  );


  not
  g86
  (
    n77,
    n11
  );


  buf
  g87
  (
    n85,
    n20
  );


  not
  g88
  (
    n321,
    n103
  );


  not
  g89
  (
    n215,
    n65
  );


  not
  g90
  (
    n384,
    n105
  );


  not
  g91
  (
    n154,
    n78
  );


  not
  g92
  (
    n223,
    n58
  );


  not
  g93
  (
    n364,
    n74
  );


  buf
  g94
  (
    n325,
    n51
  );


  buf
  g95
  (
    n291,
    n28
  );


  not
  g96
  (
    KeyWire_0_6,
    n58
  );


  buf
  g97
  (
    KeyWire_0_1,
    n40
  );


  not
  g98
  (
    n360,
    n85
  );


  buf
  g99
  (
    n126,
    n37
  );


  buf
  g100
  (
    n258,
    n75
  );


  buf
  g101
  (
    n337,
    n90
  );


  not
  g102
  (
    n310,
    n79
  );


  buf
  g103
  (
    n368,
    n61
  );


  not
  g104
  (
    n351,
    n82
  );


  not
  g105
  (
    n140,
    n74
  );


  buf
  g106
  (
    n281,
    n102
  );


  not
  g107
  (
    n228,
    n101
  );


  not
  g108
  (
    n221,
    n106
  );


  buf
  g109
  (
    n285,
    n67
  );


  buf
  g110
  (
    n218,
    n68
  );


  not
  g111
  (
    n194,
    n65
  );


  not
  g112
  (
    n252,
    n106
  );


  not
  g113
  (
    n333,
    n90
  );


  buf
  g114
  (
    n260,
    n67
  );


  not
  g115
  (
    n251,
    n52
  );


  not
  g116
  (
    n180,
    n96
  );


  not
  g117
  (
    n381,
    n56
  );


  not
  g118
  (
    n213,
    n99
  );


  buf
  g119
  (
    n244,
    n96
  );


  not
  g120
  (
    n214,
    n76
  );


  buf
  g121
  (
    n173,
    n36
  );


  buf
  g122
  (
    n365,
    n31
  );


  not
  g123
  (
    n168,
    n73
  );


  buf
  g124
  (
    n131,
    n104
  );


  buf
  g125
  (
    KeyWire_0_2,
    n92
  );


  not
  g126
  (
    n340,
    n99
  );


  buf
  g127
  (
    n141,
    n36
  );


  not
  g128
  (
    n170,
    n56
  );


  buf
  g129
  (
    n367,
    n75
  );


  buf
  g130
  (
    n302,
    n94
  );


  buf
  g131
  (
    n193,
    n109
  );


  not
  g132
  (
    n374,
    n109
  );


  buf
  g133
  (
    n243,
    n70
  );


  buf
  g134
  (
    n254,
    n80
  );


  not
  g135
  (
    n118,
    n48
  );


  not
  g136
  (
    n138,
    n89
  );


  buf
  g137
  (
    n220,
    n108
  );


  not
  g138
  (
    n253,
    n34
  );


  buf
  g139
  (
    n169,
    n80
  );


  not
  g140
  (
    n272,
    n86
  );


  buf
  g141
  (
    n265,
    n70
  );


  not
  g142
  (
    n235,
    n85
  );


  not
  g143
  (
    n342,
    n76
  );


  not
  g144
  (
    n239,
    n101
  );


  not
  g145
  (
    n356,
    n80
  );


  buf
  g146
  (
    n225,
    n37
  );


  buf
  g147
  (
    n149,
    n93
  );


  buf
  g148
  (
    n155,
    n104
  );


  buf
  g149
  (
    n159,
    n97
  );


  not
  g150
  (
    n307,
    n53
  );


  not
  g151
  (
    n232,
    n91
  );


  buf
  g152
  (
    n171,
    n107
  );


  buf
  g153
  (
    n276,
    n35
  );


  buf
  g154
  (
    n361,
    n26
  );


  buf
  g155
  (
    n280,
    n59
  );


  not
  g156
  (
    n116,
    n102
  );


  buf
  g157
  (
    n147,
    n105
  );


  not
  g158
  (
    n346,
    n66
  );


  not
  g159
  (
    n234,
    n105
  );


  not
  g160
  (
    n248,
    n42
  );


  not
  g161
  (
    n335,
    n43
  );


  not
  g162
  (
    n120,
    n69
  );


  not
  g163
  (
    n330,
    n54
  );


  not
  g164
  (
    n240,
    n92
  );


  not
  g165
  (
    n296,
    n46
  );


  buf
  g166
  (
    n275,
    n112
  );


  not
  g167
  (
    n370,
    n108
  );


  buf
  g168
  (
    n270,
    n43
  );


  buf
  g169
  (
    n249,
    n45
  );


  buf
  g170
  (
    n184,
    n25
  );


  not
  g171
  (
    n237,
    n76
  );


  buf
  g172
  (
    n202,
    n67
  );


  buf
  g173
  (
    n277,
    n94
  );


  buf
  g174
  (
    n231,
    n32
  );


  buf
  g175
  (
    n167,
    n81
  );


  buf
  g176
  (
    n255,
    n102
  );


  not
  g177
  (
    n306,
    n63
  );


  buf
  g178
  (
    n363,
    n95
  );


  not
  g179
  (
    n246,
    n45
  );


  not
  g180
  (
    n124,
    n68
  );


  not
  g181
  (
    n196,
    n84
  );


  not
  g182
  (
    n143,
    n101
  );


  not
  g183
  (
    n375,
    n42
  );


  not
  g184
  (
    n150,
    n30
  );


  not
  g185
  (
    n377,
    n111
  );


  not
  g186
  (
    n380,
    n112
  );


  not
  g187
  (
    n156,
    n28
  );


  buf
  g188
  (
    n129,
    n80
  );


  not
  g189
  (
    n348,
    n104
  );


  not
  g190
  (
    n279,
    n103
  );


  not
  g191
  (
    n316,
    n98
  );


  buf
  g192
  (
    n115,
    n88
  );


  not
  g193
  (
    n132,
    n46
  );


  buf
  g194
  (
    n192,
    n99
  );


  buf
  g195
  (
    n125,
    n44
  );


  buf
  g196
  (
    n226,
    n74
  );


  not
  g197
  (
    n323,
    n94
  );


  buf
  g198
  (
    n186,
    n41
  );


  buf
  g199
  (
    n336,
    n84
  );


  not
  g200
  (
    n345,
    n30
  );


  buf
  g201
  (
    n317,
    n57
  );


  buf
  g202
  (
    n241,
    n105
  );


  buf
  g203
  (
    n303,
    n74
  );


  not
  g204
  (
    n148,
    n87
  );


  not
  g205
  (
    n211,
    n96
  );


  not
  g206
  (
    n206,
    n107
  );


  buf
  g207
  (
    n114,
    n83
  );


  not
  g208
  (
    n344,
    n59
  );


  not
  g209
  (
    n127,
    n61
  );


  not
  g210
  (
    n201,
    n106
  );


  not
  g211
  (
    n359,
    n62
  );


  not
  g212
  (
    n136,
    n68
  );


  not
  g213
  (
    n178,
    n81
  );


  not
  g214
  (
    n174,
    n71
  );


  not
  g215
  (
    n290,
    n108
  );


  buf
  g216
  (
    n271,
    n98
  );


  not
  g217
  (
    n200,
    n107
  );


  not
  g218
  (
    n224,
    n35
  );


  not
  g219
  (
    n257,
    n29
  );


  not
  g220
  (
    n378,
    n68
  );


  buf
  g221
  (
    n299,
    n33
  );


  not
  g222
  (
    n287,
    n107
  );


  buf
  g223
  (
    n158,
    n62
  );


  not
  g224
  (
    n229,
    n55
  );


  buf
  g225
  (
    n349,
    n88
  );


  buf
  g226
  (
    n289,
    n110
  );


  buf
  g227
  (
    n236,
    n103
  );


  not
  g228
  (
    n183,
    n100
  );


  not
  g229
  (
    n165,
    n70
  );


  buf
  g230
  (
    n233,
    n79
  );


  buf
  g231
  (
    n305,
    n72
  );


  not
  g232
  (
    n372,
    n102
  );


  not
  g233
  (
    n146,
    n81
  );


  buf
  g234
  (
    n162,
    n100
  );


  not
  g235
  (
    n151,
    n39
  );


  buf
  g236
  (
    n217,
    n29
  );


  buf
  g237
  (
    n242,
    n77
  );


  not
  g238
  (
    KeyWire_0_23,
    n26
  );


  buf
  g239
  (
    n350,
    n63
  );


  buf
  g240
  (
    n163,
    n93
  );


  not
  g241
  (
    n179,
    n72
  );


  not
  g242
  (
    n308,
    n47
  );


  not
  g243
  (
    n119,
    n85
  );


  buf
  g244
  (
    n177,
    n76
  );


  buf
  g245
  (
    n259,
    n71
  );


  not
  g246
  (
    n369,
    n77
  );


  buf
  g247
  (
    n212,
    n34
  );


  not
  g248
  (
    n334,
    n88
  );


  not
  g249
  (
    n318,
    n44
  );


  buf
  g250
  (
    n264,
    n73
  );


  not
  g251
  (
    n332,
    n82
  );


  buf
  g252
  (
    n382,
    n79
  );


  not
  g253
  (
    n135,
    n66
  );


  buf
  g254
  (
    n230,
    n78
  );


  buf
  g255
  (
    n379,
    n39
  );


  not
  g256
  (
    n269,
    n90
  );


  not
  g257
  (
    n195,
    n25
  );


  not
  g258
  (
    n347,
    n64
  );


  buf
  g259
  (
    n210,
    n78
  );


  not
  g260
  (
    n256,
    n84
  );


  buf
  g261
  (
    n203,
    n112
  );


  not
  g262
  (
    n309,
    n54
  );


  not
  g263
  (
    n250,
    n87
  );


  buf
  g264
  (
    n198,
    n73
  );


  buf
  g265
  (
    n204,
    n88
  );


  buf
  g266
  (
    n142,
    n96
  );


  buf
  g267
  (
    n190,
    n57
  );


  buf
  g268
  (
    n268,
    n66
  );


  buf
  g269
  (
    n358,
    n75
  );


  buf
  g270
  (
    n331,
    n95
  );


  buf
  g271
  (
    n267,
    n85
  );


  buf
  g272
  (
    n304,
    n109
  );


  buf
  g273
  (
    n284,
    n101
  );


  not
  g274
  (
    n227,
    n31
  );


  buf
  g275
  (
    n145,
    n27
  );


  buf
  g276
  (
    n161,
    n47
  );


  not
  g277
  (
    n371,
    n94
  );


  buf
  g278
  (
    n117,
    n99
  );


  buf
  g279
  (
    n187,
    n83
  );


  not
  g280
  (
    n320,
    n100
  );


  not
  g281
  (
    n298,
    n72
  );


  buf
  g282
  (
    n383,
    n109
  );


  not
  g283
  (
    n362,
    n95
  );


  not
  g284
  (
    n355,
    n49
  );


  buf
  g285
  (
    n292,
    n97
  );


  buf
  g286
  (
    n128,
    n60
  );


  buf
  g287
  (
    n282,
    n27
  );


  buf
  g288
  (
    n133,
    n91
  );


  not
  g289
  (
    n274,
    n111
  );


  buf
  g290
  (
    n209,
    n89
  );


  not
  g291
  (
    n182,
    n53
  );


  buf
  g292
  (
    KeyWire_0_9,
    n100
  );


  not
  g293
  (
    n288,
    n70
  );


  not
  g294
  (
    n160,
    n87
  );


  not
  g295
  (
    n352,
    n33
  );


  buf
  g296
  (
    n315,
    n111
  );


  buf
  g297
  (
    n113,
    n91
  );


  not
  g298
  (
    n266,
    n75
  );


  buf
  g299
  (
    n122,
    n90
  );


  buf
  g300
  (
    n343,
    n52
  );


  buf
  g301
  (
    n294,
    n65
  );


  buf
  g302
  (
    n297,
    n112
  );


  not
  g303
  (
    n123,
    n97
  );


  not
  g304
  (
    n164,
    n51
  );


  buf
  g305
  (
    n262,
    n93
  );


  buf
  g306
  (
    n273,
    n78
  );


  buf
  g307
  (
    n172,
    n83
  );


  buf
  g308
  (
    n314,
    n60
  );


  buf
  g309
  (
    n181,
    n41
  );


  buf
  g310
  (
    n354,
    n65
  );


  buf
  g311
  (
    n189,
    n69
  );


  buf
  g312
  (
    n338,
    n86
  );


  not
  g313
  (
    n341,
    n81
  );


  buf
  g314
  (
    n139,
    n83
  );


  not
  g315
  (
    n311,
    n110
  );


  buf
  g316
  (
    n247,
    n97
  );


  not
  g317
  (
    n324,
    n50
  );


  buf
  g318
  (
    n322,
    n66
  );


  not
  g319
  (
    n153,
    n55
  );


  not
  g320
  (
    n137,
    n71
  );


  buf
  g321
  (
    n216,
    n95
  );


  buf
  g322
  (
    n199,
    n77
  );


  not
  g323
  (
    n144,
    n103
  );


  buf
  g324
  (
    n261,
    n92
  );


  buf
  g325
  (
    n222,
    n69
  );


  not
  g326
  (
    n238,
    n82
  );


  buf
  g327
  (
    n263,
    n73
  );


  not
  g328
  (
    n205,
    n40
  );


  not
  g329
  (
    n326,
    n86
  );


  not
  g330
  (
    n157,
    n77
  );


  buf
  g331
  (
    n283,
    n93
  );


  not
  g332
  (
    n197,
    n92
  );


  buf
  g333
  (
    n357,
    n71
  );


  buf
  g334
  (
    n312,
    n111
  );


  buf
  g335
  (
    n245,
    n72
  );


  buf
  g336
  (
    n166,
    n38
  );


  not
  g337
  (
    n219,
    n108
  );


  not
  g338
  (
    n300,
    n32
  );


  buf
  g339
  (
    n208,
    n38
  );


  not
  g340
  (
    n134,
    n84
  );


  not
  g341
  (
    n191,
    n87
  );


  not
  g342
  (
    n185,
    n89
  );


  not
  g343
  (
    n301,
    n110
  );


  buf
  g344
  (
    n313,
    n91
  );


  buf
  g345
  (
    n295,
    n79
  );


  not
  g346
  (
    n366,
    n104
  );


  buf
  g347
  (
    n339,
    n64
  );


  buf
  g348
  (
    n293,
    n110
  );


  buf
  g349
  (
    KeyWire_0_15,
    n49
  );


  buf
  g350
  (
    n327,
    n67
  );


  not
  g351
  (
    n376,
    n50
  );


  not
  g352
  (
    n329,
    n69
  );


  not
  g353
  (
    n207,
    n82
  );


  buf
  g354
  (
    n328,
    n86
  );


  buf
  g355
  (
    n176,
    n98
  );


  not
  g356
  (
    n373,
    n48
  );


  not
  g357
  (
    n286,
    n106
  );


  buf
  g358
  (
    n188,
    n89
  );


  buf
  g359
  (
    n319,
    n98
  );


  buf
  g360
  (
    n742,
    n273
  );


  buf
  g361
  (
    n630,
    n140
  );


  not
  g362
  (
    n414,
    n213
  );


  buf
  g363
  (
    n482,
    n142
  );


  buf
  g364
  (
    n514,
    n145
  );


  not
  g365
  (
    n573,
    n116
  );


  buf
  g366
  (
    n493,
    n284
  );


  buf
  g367
  (
    n732,
    n115
  );


  buf
  g368
  (
    n486,
    n132
  );


  not
  g369
  (
    n523,
    n276
  );


  not
  g370
  (
    n696,
    n235
  );


  buf
  g371
  (
    n483,
    n218
  );


  buf
  g372
  (
    KeyWire_0_4,
    n280
  );


  buf
  g373
  (
    n727,
    n140
  );


  buf
  g374
  (
    n413,
    n282
  );


  buf
  g375
  (
    n632,
    n188
  );


  not
  g376
  (
    n496,
    n161
  );


  not
  g377
  (
    n465,
    n155
  );


  buf
  g378
  (
    n565,
    n196
  );


  not
  g379
  (
    n724,
    n297
  );


  not
  g380
  (
    n693,
    n139
  );


  not
  g381
  (
    n598,
    n260
  );


  not
  g382
  (
    n478,
    n184
  );


  buf
  g383
  (
    n734,
    n153
  );


  not
  g384
  (
    n574,
    n297
  );


  buf
  g385
  (
    n544,
    n128
  );


  buf
  g386
  (
    n389,
    n162
  );


  not
  g387
  (
    n563,
    n171
  );


  buf
  g388
  (
    KeyWire_0_20,
    n174
  );


  not
  g389
  (
    n476,
    n227
  );


  buf
  g390
  (
    n641,
    n301
  );


  not
  g391
  (
    n456,
    n134
  );


  buf
  g392
  (
    n590,
    n223
  );


  not
  g393
  (
    n455,
    n187
  );


  buf
  g394
  (
    KeyWire_0_3,
    n284
  );


  not
  g395
  (
    n599,
    n124
  );


  buf
  g396
  (
    n485,
    n301
  );


  not
  g397
  (
    n705,
    n216
  );


  not
  g398
  (
    n568,
    n161
  );


  not
  g399
  (
    n664,
    n215
  );


  not
  g400
  (
    n488,
    n300
  );


  buf
  g401
  (
    n540,
    n141
  );


  not
  g402
  (
    n704,
    n230
  );


  buf
  g403
  (
    n521,
    n252
  );


  not
  g404
  (
    n614,
    n264
  );


  buf
  g405
  (
    n558,
    n139
  );


  not
  g406
  (
    n694,
    n228
  );


  not
  g407
  (
    n675,
    n265
  );


  buf
  g408
  (
    n718,
    n231
  );


  buf
  g409
  (
    n658,
    n118
  );


  not
  g410
  (
    n394,
    n191
  );


  not
  g411
  (
    n662,
    n248
  );


  not
  g412
  (
    n602,
    n243
  );


  buf
  g413
  (
    n690,
    n152
  );


  buf
  g414
  (
    n492,
    n201
  );


  not
  g415
  (
    n637,
    n284
  );


  buf
  g416
  (
    n562,
    n170
  );


  not
  g417
  (
    n513,
    n226
  );


  not
  g418
  (
    n583,
    n254
  );


  not
  g419
  (
    n719,
    n248
  );


  buf
  g420
  (
    n661,
    n282
  );


  buf
  g421
  (
    n612,
    n253
  );


  buf
  g422
  (
    n571,
    n271
  );


  not
  g423
  (
    n435,
    n245
  );


  not
  g424
  (
    n398,
    n278
  );


  not
  g425
  (
    n616,
    n299
  );


  buf
  g426
  (
    n386,
    n180
  );


  not
  g427
  (
    n495,
    n291
  );


  not
  g428
  (
    n452,
    n255
  );


  buf
  g429
  (
    n564,
    n204
  );


  not
  g430
  (
    n622,
    n175
  );


  buf
  g431
  (
    n406,
    n233
  );


  not
  g432
  (
    n680,
    n156
  );


  not
  g433
  (
    n607,
    n233
  );


  not
  g434
  (
    n667,
    n225
  );


  not
  g435
  (
    n735,
    n276
  );


  buf
  g436
  (
    n408,
    n286
  );


  not
  g437
  (
    n588,
    n220
  );


  not
  g438
  (
    n620,
    n180
  );


  not
  g439
  (
    n733,
    n302
  );


  not
  g440
  (
    n744,
    n244
  );


  not
  g441
  (
    n454,
    n169
  );


  buf
  g442
  (
    n451,
    n176
  );


  buf
  g443
  (
    n529,
    n177
  );


  not
  g444
  (
    n611,
    n234
  );


  not
  g445
  (
    n459,
    n174
  );


  not
  g446
  (
    n422,
    n219
  );


  not
  g447
  (
    n427,
    n286
  );


  buf
  g448
  (
    n619,
    n278
  );


  not
  g449
  (
    n432,
    n130
  );


  not
  g450
  (
    n655,
    n207
  );


  buf
  g451
  (
    n535,
    n278
  );


  not
  g452
  (
    n400,
    n269
  );


  buf
  g453
  (
    n541,
    n253
  );


  not
  g454
  (
    n751,
    n248
  );


  not
  g455
  (
    n566,
    n196
  );


  buf
  g456
  (
    n712,
    n301
  );


  buf
  g457
  (
    n431,
    n249
  );


  not
  g458
  (
    KeyWire_0_25,
    n265
  );


  not
  g459
  (
    n393,
    n142
  );


  buf
  g460
  (
    n403,
    n283
  );


  not
  g461
  (
    n700,
    n239
  );


  buf
  g462
  (
    n723,
    n119
  );


  buf
  g463
  (
    n683,
    n170
  );


  not
  g464
  (
    n746,
    n220
  );


  buf
  g465
  (
    n710,
    n164
  );


  not
  g466
  (
    n450,
    n298
  );


  buf
  g467
  (
    n551,
    n183
  );


  buf
  g468
  (
    n396,
    n136
  );


  buf
  g469
  (
    KeyWire_0_17,
    n245
  );


  buf
  g470
  (
    n511,
    n155
  );


  buf
  g471
  (
    n728,
    n126
  );


  not
  g472
  (
    n706,
    n255
  );


  buf
  g473
  (
    n678,
    n135
  );


  not
  g474
  (
    n392,
    n190
  );


  buf
  g475
  (
    n585,
    n279
  );


  not
  g476
  (
    n674,
    n207
  );


  buf
  g477
  (
    n397,
    n160
  );


  buf
  g478
  (
    n600,
    n197
  );


  buf
  g479
  (
    n460,
    n113
  );


  not
  g480
  (
    n685,
    n192
  );


  not
  g481
  (
    n587,
    n177
  );


  buf
  g482
  (
    n480,
    n225
  );


  not
  g483
  (
    n522,
    n241
  );


  buf
  g484
  (
    n660,
    n277
  );


  buf
  g485
  (
    n548,
    n166
  );


  not
  g486
  (
    n442,
    n133
  );


  buf
  g487
  (
    n748,
    n178
  );


  not
  g488
  (
    n472,
    n218
  );


  not
  g489
  (
    n552,
    n143
  );


  not
  g490
  (
    n645,
    n292
  );


  buf
  g491
  (
    n453,
    n190
  );


  buf
  g492
  (
    n575,
    n243
  );


  buf
  g493
  (
    n399,
    n181
  );


  buf
  g494
  (
    n416,
    n133
  );


  buf
  g495
  (
    n519,
    n242
  );


  buf
  g496
  (
    n640,
    n256
  );


  buf
  g497
  (
    n409,
    n289
  );


  buf
  g498
  (
    n639,
    n115
  );


  buf
  g499
  (
    n433,
    n257
  );


  not
  g500
  (
    n462,
    n129
  );


  not
  g501
  (
    n624,
    n246
  );


  buf
  g502
  (
    n385,
    n118
  );


  buf
  g503
  (
    n651,
    n213
  );


  not
  g504
  (
    n387,
    n234
  );


  not
  g505
  (
    n458,
    n216
  );


  not
  g506
  (
    n671,
    n222
  );


  buf
  g507
  (
    n609,
    n264
  );


  buf
  g508
  (
    n713,
    n240
  );


  not
  g509
  (
    n430,
    n216
  );


  buf
  g510
  (
    n688,
    n189
  );


  not
  g511
  (
    n569,
    n124
  );


  not
  g512
  (
    n621,
    n125
  );


  not
  g513
  (
    n729,
    n235
  );


  buf
  g514
  (
    n592,
    n199
  );


  not
  g515
  (
    n487,
    n292
  );


  buf
  g516
  (
    n554,
    n141
  );


  not
  g517
  (
    n536,
    n285
  );


  not
  g518
  (
    n401,
    n290
  );


  not
  g519
  (
    n510,
    n174
  );


  not
  g520
  (
    n533,
    n127
  );


  buf
  g521
  (
    n412,
    n230
  );


  not
  g522
  (
    n497,
    n134
  );


  not
  g523
  (
    n507,
    n238
  );


  not
  g524
  (
    n643,
    n262
  );


  not
  g525
  (
    n494,
    n165
  );


  buf
  g526
  (
    n550,
    n134
  );


  buf
  g527
  (
    n449,
    n258
  );


  buf
  g528
  (
    n601,
    n264
  );


  buf
  g529
  (
    n730,
    n200
  );


  buf
  g530
  (
    n539,
    n194
  );


  not
  g531
  (
    n512,
    n151
  );


  buf
  g532
  (
    n475,
    n146
  );


  not
  g533
  (
    n638,
    n251
  );


  buf
  g534
  (
    n448,
    n143
  );


  not
  g535
  (
    n752,
    n218
  );


  buf
  g536
  (
    n596,
    n132
  );


  not
  g537
  (
    n635,
    n276
  );


  buf
  g538
  (
    n720,
    n288
  );


  buf
  g539
  (
    n740,
    n172
  );


  not
  g540
  (
    n707,
    n153
  );


  buf
  g541
  (
    n423,
    n227
  );


  not
  g542
  (
    n697,
    n209
  );


  not
  g543
  (
    n518,
    n226
  );


  buf
  g544
  (
    n532,
    n229
  );


  buf
  g545
  (
    n468,
    n201
  );


  buf
  g546
  (
    n546,
    n240
  );


  buf
  g547
  (
    n747,
    n127
  );


  buf
  g548
  (
    n725,
    n274
  );


  buf
  g549
  (
    n466,
    n183
  );


  buf
  g550
  (
    n410,
    n210
  );


  buf
  g551
  (
    n745,
    n271
  );


  buf
  g552
  (
    n471,
    n224
  );


  buf
  g553
  (
    n434,
    n148
  );


  buf
  g554
  (
    n543,
    n198
  );


  not
  g555
  (
    n677,
    n261
  );


  buf
  g556
  (
    n576,
    n189
  );


  buf
  g557
  (
    n684,
    n135
  );


  buf
  g558
  (
    n666,
    n161
  );


  buf
  g559
  (
    n555,
    n170
  );


  buf
  g560
  (
    n516,
    n165
  );


  not
  g561
  (
    n402,
    n182
  );


  not
  g562
  (
    n542,
    n187
  );


  buf
  g563
  (
    n531,
    n261
  );


  buf
  g564
  (
    n443,
    n137
  );


  buf
  g565
  (
    n577,
    n287
  );


  buf
  g566
  (
    n686,
    n271
  );


  buf
  g567
  (
    n390,
    n293
  );


  buf
  g568
  (
    n418,
    n203
  );


  buf
  g569
  (
    n438,
    n136
  );


  not
  g570
  (
    n714,
    n200
  );


  buf
  g571
  (
    n663,
    n128
  );


  buf
  g572
  (
    n593,
    n229
  );


  buf
  g573
  (
    KeyWire_0_13,
    n290
  );


  not
  g574
  (
    KeyWire_0_22,
    n153
  );


  not
  g575
  (
    n654,
    n300
  );


  buf
  g576
  (
    n477,
    n208
  );


  buf
  g577
  (
    n428,
    n272
  );


  buf
  g578
  (
    n715,
    n159
  );


  not
  g579
  (
    n499,
    n155
  );


  buf
  g580
  (
    n673,
    n117
  );


  not
  g581
  (
    n594,
    n175
  );


  buf
  g582
  (
    n738,
    n294
  );


  not
  g583
  (
    KeyWire_0_12,
    n119
  );


  buf
  g584
  (
    n419,
    n217
  );


  not
  g585
  (
    n534,
    n217
  );


  not
  g586
  (
    KeyWire_0_8,
    n283
  );


  buf
  g587
  (
    n527,
    n113
  );


  buf
  g588
  (
    n470,
    n144
  );


  not
  g589
  (
    n464,
    n122
  );


  buf
  g590
  (
    n646,
    n251
  );


  not
  g591
  (
    n461,
    n247
  );


  buf
  g592
  (
    n549,
    n176
  );


  not
  g593
  (
    n629,
    n250
  );


  buf
  g594
  (
    n479,
    n237
  );


  buf
  g595
  (
    n623,
    n138
  );


  buf
  g596
  (
    n446,
    n244
  );


  buf
  g597
  (
    n515,
    n261
  );


  buf
  g598
  (
    n524,
    n168
  );


  not
  g599
  (
    n586,
    n259
  );


  nor
  g600
  (
    n502,
    n172,
    n156,
    n180,
    n136
  );


  xor
  g601
  (
    n625,
    n220,
    n163,
    n114,
    n136
  );


  nor
  g602
  (
    n404,
    n132,
    n280,
    n245,
    n238
  );


  xnor
  g603
  (
    n703,
    n205,
    n232,
    n169,
    n207
  );


  and
  g604
  (
    n561,
    n209,
    n147,
    n157,
    n203
  );


  nand
  g605
  (
    n580,
    n223,
    n290,
    n255,
    n186
  );


  and
  g606
  (
    n526,
    n158,
    n130,
    n243,
    n236
  );


  and
  g607
  (
    n695,
    n185,
    n206,
    n198,
    n128
  );


  nor
  g608
  (
    n420,
    n296,
    n195,
    n268,
    n184
  );


  or
  g609
  (
    n709,
    n297,
    n139,
    n127,
    n237
  );


  or
  g610
  (
    n652,
    n175,
    n295,
    n273,
    n293
  );


  xnor
  g611
  (
    n388,
    n221,
    n221,
    n167,
    n253
  );


  xor
  g612
  (
    n681,
    n125,
    n231,
    n204,
    n240
  );


  xnor
  g613
  (
    n642,
    n147,
    n285,
    n250,
    n277
  );


  xnor
  g614
  (
    n711,
    n200,
    n160,
    n208,
    n258
  );


  xor
  g615
  (
    n676,
    n273,
    n152,
    n212,
    n293
  );


  xnor
  g616
  (
    n572,
    n295,
    n241,
    n276,
    n160
  );


  or
  g617
  (
    n506,
    n141,
    n201,
    n190,
    n166
  );


  nor
  g618
  (
    n589,
    n117,
    n256,
    n254,
    n158
  );


  and
  g619
  (
    n659,
    n173,
    n127,
    n212,
    n118
  );


  xor
  g620
  (
    n440,
    n280,
    n179,
    n171,
    n123
  );


  nand
  g621
  (
    KeyWire_0_7,
    n227,
    n192,
    n137,
    n126
  );


  xor
  g622
  (
    n437,
    n148,
    n205,
    n125,
    n228
  );


  xnor
  g623
  (
    n741,
    n239,
    n124,
    n138,
    n150
  );


  xor
  g624
  (
    n649,
    n281,
    n118,
    n121,
    n244
  );


  or
  g625
  (
    n708,
    n157,
    n154,
    n194,
    n299
  );


  xnor
  g626
  (
    n417,
    n237,
    n201,
    n299,
    n283
  );


  nor
  g627
  (
    KeyWire_0_16,
    n258,
    n165,
    n209,
    n117
  );


  xnor
  g628
  (
    n606,
    n180,
    n149,
    n234,
    n166
  );


  nor
  g629
  (
    n636,
    n211,
    n177,
    n267,
    n302
  );


  xnor
  g630
  (
    n736,
    n250,
    n260,
    n132,
    n235
  );


  nor
  g631
  (
    n670,
    n235,
    n147,
    n269,
    n149
  );


  nor
  g632
  (
    n474,
    n267,
    n232,
    n139,
    n249
  );


  xnor
  g633
  (
    n457,
    n203,
    n258,
    n225,
    n250
  );


  and
  g634
  (
    n750,
    n122,
    n126,
    n171,
    n154
  );


  nor
  g635
  (
    n537,
    n164,
    n273,
    n285,
    n270
  );


  nand
  g636
  (
    n618,
    n248,
    n159,
    n197,
    n254
  );


  nor
  g637
  (
    n439,
    n267,
    n187,
    n275,
    n214
  );


  xor
  g638
  (
    n603,
    n162,
    n287,
    n300,
    n245
  );


  and
  g639
  (
    n610,
    n215,
    n207,
    n242,
    n266
  );


  xor
  g640
  (
    n578,
    n277,
    n269,
    n256,
    n206
  );


  or
  g641
  (
    n613,
    n268,
    n225,
    n215,
    n219
  );


  and
  g642
  (
    n567,
    n188,
    n210,
    n266,
    n256
  );


  or
  g643
  (
    KeyWire_0_11,
    n151,
    n236,
    n295,
    n217
  );


  nor
  g644
  (
    n668,
    n241,
    n221,
    n175,
    n145
  );


  nor
  g645
  (
    n749,
    n249,
    n202,
    n281,
    n292
  );


  nor
  g646
  (
    n581,
    n186,
    n224,
    n196,
    n198
  );


  xor
  g647
  (
    n669,
    n114,
    n287,
    n288,
    n268
  );


  or
  g648
  (
    n447,
    n209,
    n286,
    n252,
    n150
  );


  xnor
  g649
  (
    n722,
    n260,
    n189,
    n281,
    n116
  );


  nor
  g650
  (
    n411,
    n124,
    n216,
    n237,
    n272
  );


  or
  g651
  (
    n731,
    n133,
    n271,
    n131,
    n191
  );


  nor
  g652
  (
    n739,
    n229,
    n164,
    n224,
    n251
  );


  and
  g653
  (
    n591,
    n158,
    n277,
    n115,
    n119
  );


  xnor
  g654
  (
    n491,
    n213,
    n275,
    n157,
    n227
  );


  and
  g655
  (
    n445,
    n299,
    n228,
    n206,
    n223
  );


  nor
  g656
  (
    n545,
    n211,
    n223,
    n272,
    n228
  );


  xor
  g657
  (
    n415,
    n138,
    n128,
    n241,
    n213
  );


  nor
  g658
  (
    n557,
    n171,
    n170,
    n233,
    n145
  );


  or
  g659
  (
    n608,
    n150,
    n212,
    n145,
    n263
  );


  nand
  g660
  (
    n553,
    n202,
    n192,
    n298,
    n288
  );


  xor
  g661
  (
    n717,
    n161,
    n261,
    n120,
    n293
  );


  xnor
  g662
  (
    n650,
    n266,
    n135,
    n222,
    n279
  );


  and
  g663
  (
    n633,
    n148,
    n280,
    n275,
    n287
  );


  nor
  g664
  (
    n691,
    n249,
    n265,
    n160,
    n274
  );


  and
  g665
  (
    n626,
    n167,
    n291,
    n204,
    n144
  );


  or
  g666
  (
    n530,
    n152,
    n243,
    n162,
    n154
  );


  and
  g667
  (
    KeyWire_0_27,
    n177,
    n212,
    n238,
    n189
  );


  nand
  g668
  (
    n644,
    n137,
    n140,
    n178,
    n193
  );


  or
  g669
  (
    n498,
    n122,
    n281,
    n150,
    n156
  );


  xor
  g670
  (
    n504,
    n251,
    n211,
    n129,
    n115
  );


  xnor
  g671
  (
    n509,
    n205,
    n193,
    n172,
    n268
  );


  xnor
  g672
  (
    n716,
    n130,
    n144,
    n126,
    n176
  );


  xor
  g673
  (
    n682,
    n142,
    n240,
    n121,
    n179
  );


  nor
  g674
  (
    n500,
    n294,
    n259,
    n169,
    n174
  );


  nor
  g675
  (
    n605,
    n259,
    n195,
    n158,
    n186
  );


  nand
  g676
  (
    n665,
    n246,
    n230,
    n188,
    n129
  );


  nor
  g677
  (
    n520,
    n168,
    n208,
    n284,
    n120
  );


  xor
  g678
  (
    n634,
    n219,
    n226,
    n148,
    n236
  );


  nor
  g679
  (
    n426,
    n279,
    n289,
    n296,
    n143
  );


  nand
  g680
  (
    n672,
    n183,
    n146,
    n292,
    n246
  );


  nand
  g681
  (
    n441,
    n181,
    n294,
    n236,
    n221
  );


  xor
  g682
  (
    n559,
    n159,
    n185,
    n202,
    n272
  );


  and
  g683
  (
    n689,
    n263,
    n267,
    n257,
    n155
  );


  or
  g684
  (
    n692,
    n246,
    n247,
    n199
  );


  nor
  g685
  (
    n473,
    n185,
    n181,
    n290,
    n289
  );


  xor
  g686
  (
    n481,
    n198,
    n208,
    n291,
    n239
  );


  or
  g687
  (
    n582,
    n168,
    n131,
    n296,
    n257
  );


  xnor
  g688
  (
    n584,
    n239,
    n120,
    n296,
    n151
  );


  xnor
  g689
  (
    n657,
    n182,
    n191,
    n185,
    n173
  );


  xnor
  g690
  (
    n424,
    n188,
    n116,
    n131,
    n214
  );


  xor
  g691
  (
    n436,
    n242,
    n191,
    n123,
    n294
  );


  nor
  g692
  (
    n698,
    n283,
    n247,
    n178,
    n194
  );


  nand
  g693
  (
    n648,
    n194,
    n142,
    n144,
    n178
  );


  or
  g694
  (
    n538,
    n234,
    n156,
    n114
  );


  nand
  g695
  (
    n467,
    n263,
    n200,
    n117,
    n244
  );


  nand
  g696
  (
    n647,
    n206,
    n266,
    n229,
    n133
  );


  xor
  g697
  (
    n679,
    n152,
    n187,
    n129,
    n167
  );


  nor
  g698
  (
    n463,
    n173,
    n262,
    n242,
    n298
  );


  xor
  g699
  (
    n421,
    n270,
    n255,
    n184,
    n214
  );


  xnor
  g700
  (
    n503,
    n164,
    n210,
    n297,
    n186
  );


  nor
  g701
  (
    n405,
    n123,
    n196,
    n182,
    n226
  );


  xor
  g702
  (
    n444,
    n130,
    n222,
    n195,
    n269
  );


  xor
  g703
  (
    n604,
    n125,
    n120,
    n233,
    n137
  );


  xnor
  g704
  (
    n579,
    n173,
    n193,
    n262,
    n218
  );


  nand
  g705
  (
    n425,
    n278,
    n254,
    n238,
    n166
  );


  nand
  g706
  (
    n489,
    n279,
    n252,
    n197,
    n232
  );


  xor
  g707
  (
    n469,
    n147,
    n122,
    n182,
    n183
  );


  xnor
  g708
  (
    n627,
    n217,
    n190,
    n264,
    n146
  );


  nand
  g709
  (
    n628,
    n270,
    n169,
    n289,
    n203
  );


  xnor
  g710
  (
    n597,
    n222,
    n119,
    n211,
    n193
  );


  xnor
  g711
  (
    n484,
    n172,
    n205,
    n138,
    n257
  );


  nor
  g712
  (
    n743,
    n159,
    n168,
    n252,
    n298
  );


  or
  g713
  (
    n528,
    n195,
    n274,
    n262,
    n179
  );


  or
  g714
  (
    n501,
    n140,
    n295,
    n224,
    n288
  );


  nand
  g715
  (
    n617,
    n300,
    n253,
    n149,
    n270
  );


  or
  g716
  (
    n490,
    n231,
    n260,
    n141,
    n181
  );


  or
  g717
  (
    n687,
    n210,
    n121,
    n143,
    n259
  );


  xor
  g718
  (
    n505,
    n202,
    n274,
    n123,
    n192
  );


  nor
  g719
  (
    n391,
    n214,
    n265,
    n282
  );


  or
  g720
  (
    n556,
    n153,
    n263,
    n204,
    n285
  );


  xor
  g721
  (
    n560,
    n199,
    n163,
    n167,
    n286
  );


  nand
  g722
  (
    n656,
    n149,
    n220,
    n176,
    n163
  );


  or
  g723
  (
    n395,
    n165,
    n131,
    n184,
    n231
  );


  nand
  g724
  (
    n429,
    n154,
    n162,
    n135,
    n134
  );


  and
  g725
  (
    n570,
    n121,
    n157,
    n230,
    n219
  );


  nor
  g726
  (
    n653,
    n275,
    n232,
    n163,
    n291
  );


  and
  g727
  (
    n737,
    n116,
    n215,
    n179,
    n197
  );


  xnor
  g728
  (
    n753,
    n151,
    n146,
    n199,
    n301
  );


  buf
  g729
  (
    n817,
    n508
  );


  not
  g730
  (
    n840,
    n463
  );


  buf
  g731
  (
    n841,
    n480
  );


  buf
  g732
  (
    n779,
    n533
  );


  not
  g733
  (
    n836,
    n450
  );


  buf
  g734
  (
    n784,
    n457
  );


  buf
  g735
  (
    n776,
    n433
  );


  buf
  g736
  (
    n760,
    n439
  );


  not
  g737
  (
    n849,
    n410
  );


  buf
  g738
  (
    n765,
    n486
  );


  buf
  g739
  (
    n801,
    n522
  );


  buf
  g740
  (
    n772,
    n504
  );


  not
  g741
  (
    n835,
    n432
  );


  not
  g742
  (
    n834,
    n407
  );


  buf
  g743
  (
    n791,
    n471
  );


  buf
  g744
  (
    n788,
    n420
  );


  not
  g745
  (
    n783,
    n387
  );


  not
  g746
  (
    n810,
    n512
  );


  buf
  g747
  (
    n755,
    n435
  );


  buf
  g748
  (
    n821,
    n481
  );


  not
  g749
  (
    n759,
    n507
  );


  buf
  g750
  (
    n820,
    n494
  );


  buf
  g751
  (
    n837,
    n430
  );


  buf
  g752
  (
    n781,
    n456
  );


  not
  g753
  (
    n832,
    n479
  );


  not
  g754
  (
    n819,
    n538
  );


  buf
  g755
  (
    n825,
    n501
  );


  not
  g756
  (
    n764,
    n506
  );


  buf
  g757
  (
    n770,
    n510
  );


  not
  g758
  (
    n774,
    n514
  );


  not
  g759
  (
    n806,
    n518
  );


  buf
  g760
  (
    n846,
    n467
  );


  buf
  g761
  (
    n793,
    n515
  );


  buf
  g762
  (
    n850,
    n444
  );


  not
  g763
  (
    n811,
    n483
  );


  buf
  g764
  (
    n826,
    n452
  );


  buf
  g765
  (
    n844,
    n423
  );


  buf
  g766
  (
    n795,
    n519
  );


  buf
  g767
  (
    n786,
    n438
  );


  buf
  g768
  (
    n813,
    n528
  );


  buf
  g769
  (
    n767,
    n442
  );


  buf
  g770
  (
    n773,
    n498
  );


  buf
  g771
  (
    n782,
    n530
  );


  buf
  g772
  (
    n787,
    n509
  );


  not
  g773
  (
    n798,
    n446
  );


  buf
  g774
  (
    n828,
    n393
  );


  not
  g775
  (
    n799,
    n451
  );


  not
  g776
  (
    n839,
    n389
  );


  not
  g777
  (
    n808,
    n476
  );


  not
  g778
  (
    n831,
    n517
  );


  not
  g779
  (
    n775,
    n443
  );


  buf
  g780
  (
    n756,
    n412
  );


  buf
  g781
  (
    n792,
    n391
  );


  not
  g782
  (
    n824,
    n497
  );


  not
  g783
  (
    n790,
    n500
  );


  not
  g784
  (
    n807,
    n395
  );


  buf
  g785
  (
    n766,
    n426
  );


  buf
  g786
  (
    n816,
    n474
  );


  buf
  g787
  (
    n803,
    n468
  );


  buf
  g788
  (
    n796,
    n492
  );


  buf
  g789
  (
    n778,
    n539
  );


  not
  g790
  (
    n827,
    n511
  );


  buf
  g791
  (
    n818,
    n529
  );


  buf
  g792
  (
    n842,
    n427
  );


  not
  g793
  (
    n815,
    n513
  );


  not
  g794
  (
    n794,
    n470
  );


  buf
  g795
  (
    n809,
    n472
  );


  buf
  g796
  (
    n852,
    n464
  );


  not
  g797
  (
    n780,
    n535
  );


  not
  g798
  (
    n797,
    n449
  );


  buf
  g799
  (
    n829,
    n390
  );


  buf
  g800
  (
    n838,
    n408
  );


  not
  g801
  (
    n769,
    n396
  );


  not
  g802
  (
    n763,
    n437
  );


  not
  g803
  (
    n771,
    n489
  );


  buf
  g804
  (
    n785,
    n392
  );


  buf
  g805
  (
    n812,
    n417
  );


  buf
  g806
  (
    n800,
    n455
  );


  buf
  g807
  (
    n777,
    n540
  );


  buf
  g808
  (
    n758,
    n490
  );


  and
  g809
  (
    n802,
    n459,
    n536,
    n413,
    n425
  );


  xor
  g810
  (
    n804,
    n441,
    n405,
    n429,
    n406
  );


  nand
  g811
  (
    n768,
    n484,
    n394,
    n385,
    n487
  );


  nand
  g812
  (
    n762,
    n465,
    n414,
    n503,
    n482
  );


  xor
  g813
  (
    n848,
    n462,
    n527,
    n523,
    n516
  );


  xor
  g814
  (
    n843,
    n404,
    n421,
    n409,
    n502
  );


  xor
  g815
  (
    n830,
    n521,
    n499,
    n478,
    n399
  );


  or
  g816
  (
    n814,
    n469,
    n520,
    n488,
    n422
  );


  nand
  g817
  (
    n845,
    n526,
    n397,
    n491,
    n505
  );


  nand
  g818
  (
    n757,
    n440,
    n411,
    n403,
    n419
  );


  and
  g819
  (
    n822,
    n466,
    n447,
    n461,
    n460
  );


  nand
  g820
  (
    n761,
    n402,
    n398,
    n485,
    n458
  );


  xor
  g821
  (
    n833,
    n534,
    n428,
    n496,
    n448
  );


  and
  g822
  (
    n789,
    n495,
    n445,
    n431,
    n418
  );


  nand
  g823
  (
    n823,
    n401,
    n473,
    n416,
    n475
  );


  and
  g824
  (
    n805,
    n531,
    n477,
    n388,
    n434
  );


  nand
  g825
  (
    n847,
    n524,
    n493,
    n436,
    n454
  );


  xor
  g826
  (
    n851,
    n424,
    n537,
    n415,
    n400
  );


  xnor
  g827
  (
    n754,
    n532,
    n525,
    n453,
    n386
  );


  not
  g828
  (
    n860,
    n759
  );


  buf
  g829
  (
    n853,
    n754
  );


  buf
  g830
  (
    n859,
    n756
  );


  not
  g831
  (
    n856,
    n755
  );


  buf
  g832
  (
    n861,
    n757
  );


  not
  g833
  (
    n855,
    n755
  );


  not
  g834
  (
    n854,
    n758
  );


  buf
  g835
  (
    n862,
    n758
  );


  not
  g836
  (
    n857,
    n759
  );


  not
  g837
  (
    n863,
    n756
  );


  not
  g838
  (
    n858,
    n757
  );


  or
  g839
  (
    n869,
    n542,
    n862,
    n565,
    n541
  );


  and
  g840
  (
    n865,
    n543,
    n551,
    n858,
    n567
  );


  and
  g841
  (
    n866,
    n549,
    n857,
    n553,
    n855
  );


  xor
  g842
  (
    n872,
    n859,
    n544,
    n566,
    n548
  );


  and
  g843
  (
    n870,
    n559,
    n550,
    n547,
    n562
  );


  or
  g844
  (
    n864,
    n557,
    n558,
    n860,
    n856
  );


  xor
  g845
  (
    n867,
    n569,
    n554,
    n560,
    n861
  );


  xnor
  g846
  (
    n868,
    n564,
    n568,
    n863,
    n546
  );


  nand
  g847
  (
    n873,
    n552,
    n556,
    n555,
    n561
  );


  or
  g848
  (
    n871,
    n863,
    n545,
    n563,
    n570
  );


  buf
  g849
  (
    n886,
    n871
  );


  not
  g850
  (
    n881,
    n867
  );


  nand
  g851
  (
    n879,
    n588,
    n596,
    n873,
    n577
  );


  nor
  g852
  (
    n889,
    n864,
    n869,
    n870,
    n592
  );


  nand
  g853
  (
    n893,
    n868,
    n760,
    n23,
    n591
  );


  xnor
  g854
  (
    n883,
    n583,
    n576,
    n580,
    n761
  );


  nand
  g855
  (
    n884,
    n586,
    n869,
    n871,
    n584
  );


  nand
  g856
  (
    n878,
    n872,
    n760,
    n870,
    n871
  );


  nand
  g857
  (
    n888,
    n865,
    n872,
    n868,
    n867
  );


  nor
  g858
  (
    n885,
    n579,
    n581,
    n868,
    n590
  );


  xnor
  g859
  (
    n882,
    n597,
    n865,
    n593,
    n864
  );


  or
  g860
  (
    n891,
    n582,
    n867,
    n866
  );


  nor
  g861
  (
    n890,
    n868,
    n869,
    n864,
    n599
  );


  xnor
  g862
  (
    n892,
    n595,
    n572,
    n866,
    n871
  );


  xnor
  g863
  (
    n877,
    n870,
    n573,
    n761,
    n864
  );


  xnor
  g864
  (
    n875,
    n873,
    n873,
    n867,
    n870
  );


  or
  g865
  (
    n876,
    n873,
    n872,
    n574,
    n587
  );


  or
  g866
  (
    n887,
    n869,
    n575,
    n865,
    n589
  );


  or
  g867
  (
    n874,
    n578,
    n865,
    n872,
    n585
  );


  xnor
  g868
  (
    n880,
    n866,
    n598,
    n571,
    n594
  );


  not
  g869
  (
    n930,
    n767
  );


  not
  g870
  (
    n908,
    n821
  );


  buf
  g871
  (
    n918,
    n802
  );


  buf
  g872
  (
    n950,
    n817
  );


  not
  g873
  (
    n957,
    n23
  );


  not
  g874
  (
    n903,
    n887
  );


  not
  g875
  (
    n916,
    n24
  );


  buf
  g876
  (
    n942,
    n771
  );


  buf
  g877
  (
    n947,
    n791
  );


  not
  g878
  (
    n948,
    n770
  );


  not
  g879
  (
    n964,
    n813
  );


  not
  g880
  (
    n954,
    n885
  );


  not
  g881
  (
    n936,
    n775
  );


  not
  g882
  (
    n926,
    n893
  );


  buf
  g883
  (
    n965,
    n606
  );


  not
  g884
  (
    n911,
    n887
  );


  buf
  g885
  (
    n935,
    n790
  );


  not
  g886
  (
    n939,
    n806
  );


  buf
  g887
  (
    n902,
    n805
  );


  buf
  g888
  (
    n955,
    n780
  );


  buf
  g889
  (
    n919,
    n23
  );


  buf
  g890
  (
    n894,
    n792
  );


  buf
  g891
  (
    n967,
    n881
  );


  buf
  g892
  (
    n959,
    n876
  );


  xnor
  g893
  (
    n949,
    n776,
    n886
  );


  xnor
  g894
  (
    n920,
    n610,
    n795,
    n778,
    n788
  );


  nand
  g895
  (
    n932,
    n772,
    n789,
    n24,
    n811
  );


  or
  g896
  (
    n915,
    n881,
    n615,
    n877,
    n883
  );


  nor
  g897
  (
    n951,
    n786,
    n879,
    n889,
    n791
  );


  nor
  g898
  (
    n958,
    n789,
    n884,
    n877,
    n883
  );


  or
  g899
  (
    n928,
    n800,
    n883,
    n875,
    n765
  );


  and
  g900
  (
    n961,
    n809,
    n602,
    n818,
    n783
  );


  and
  g901
  (
    n901,
    n787,
    n303,
    n771,
    n890
  );


  nand
  g902
  (
    n909,
    n763,
    n880,
    n879,
    n782
  );


  nand
  g903
  (
    n905,
    n818,
    n814,
    n801,
    n875
  );


  nor
  g904
  (
    n956,
    n882,
    n779,
    n879,
    n820
  );


  nand
  g905
  (
    n946,
    n885,
    n801,
    n803,
    n802
  );


  nor
  g906
  (
    n923,
    n797,
    n878,
    n815,
    n303
  );


  nand
  g907
  (
    n944,
    n884,
    n604,
    n603,
    n796
  );


  xor
  g908
  (
    n962,
    n773,
    n806,
    n874,
    n800
  );


  and
  g909
  (
    n933,
    n890,
    n23,
    n804,
    n886
  );


  xor
  g910
  (
    n929,
    n816,
    n784,
    n611,
    n889
  );


  xor
  g911
  (
    n906,
    n793,
    n881,
    n885,
    n810
  );


  or
  g912
  (
    n963,
    n803,
    n766,
    n884,
    n614
  );


  and
  g913
  (
    n897,
    n892,
    n882,
    n805,
    n891
  );


  or
  g914
  (
    n960,
    n819,
    n607,
    n817,
    n888
  );


  nor
  g915
  (
    n941,
    n797,
    n795,
    n891,
    n878
  );


  or
  g916
  (
    n904,
    n820,
    n892,
    n814,
    n762
  );


  xor
  g917
  (
    n914,
    n787,
    n886,
    n780,
    n302
  );


  nor
  g918
  (
    n899,
    n891,
    n785,
    n769,
    n790
  );


  or
  g919
  (
    n922,
    n778,
    n893,
    n880,
    n601
  );


  xor
  g920
  (
    n945,
    n788,
    n878,
    n890,
    n879
  );


  nor
  g921
  (
    n934,
    n812,
    n882,
    n772,
    n819
  );


  nor
  g922
  (
    n912,
    n762,
    n807,
    n808,
    n893
  );


  xnor
  g923
  (
    n966,
    n765,
    n776,
    n883,
    n887
  );


  xnor
  g924
  (
    n953,
    n608,
    n769,
    n893,
    n605
  );


  and
  g925
  (
    n940,
    n809,
    n768,
    n785,
    n796
  );


  nand
  g926
  (
    n900,
    n799,
    n773,
    n813,
    n891
  );


  or
  g927
  (
    n910,
    n810,
    n799,
    n600,
    n777
  );


  xnor
  g928
  (
    n931,
    n792,
    n815,
    n880,
    n768
  );


  and
  g929
  (
    n952,
    n612,
    n886,
    n782,
    n874
  );


  xnor
  g930
  (
    n898,
    n786,
    n764,
    n816,
    n774
  );


  nand
  g931
  (
    n921,
    n767,
    n770,
    n303,
    n808
  );


  xnor
  g932
  (
    n938,
    n302,
    n888,
    n794
  );


  nand
  g933
  (
    n927,
    n877,
    n889,
    n783,
    n798
  );


  or
  g934
  (
    n925,
    n763,
    n892,
    n798,
    n811
  );


  and
  g935
  (
    n907,
    n781,
    n880,
    n764,
    n609
  );


  nor
  g936
  (
    n924,
    n807,
    n303,
    n876,
    n24
  );


  xnor
  g937
  (
    n913,
    n812,
    n890,
    n781,
    n882
  );


  and
  g938
  (
    n917,
    n775,
    n774,
    n884,
    n887
  );


  and
  g939
  (
    n943,
    n766,
    n878,
    n885,
    n892
  );


  nand
  g940
  (
    n895,
    n804,
    n881,
    n24,
    n779
  );


  or
  g941
  (
    n937,
    n888,
    n613,
    n794,
    n777
  );


  xnor
  g942
  (
    n896,
    n877,
    n793,
    n784,
    n889
  );


  nand
  g943
  (
    n982,
    n937,
    n934,
    n915,
    n930
  );


  or
  g944
  (
    n975,
    n909,
    n898,
    n904,
    n953
  );


  xor
  g945
  (
    n968,
    n905,
    n941,
    n924,
    n942
  );


  nor
  g946
  (
    n974,
    n950,
    n929,
    n943,
    n933
  );


  xnor
  g947
  (
    n980,
    n907,
    n948,
    n917,
    n927
  );


  and
  g948
  (
    n972,
    n919,
    n899,
    n916,
    n900
  );


  xor
  g949
  (
    n978,
    n938,
    n903,
    n931,
    n951
  );


  and
  g950
  (
    n976,
    n928,
    n952,
    n901,
    n925
  );


  nor
  g951
  (
    n970,
    n897,
    n947,
    n918,
    n939
  );


  xnor
  g952
  (
    KeyWire_0_24,
    n902,
    n896,
    n935,
    n944
  );


  and
  g953
  (
    n973,
    n946,
    n945,
    n949,
    n926
  );


  or
  g954
  (
    n979,
    n923,
    n914,
    n894,
    n908
  );


  nand
  g955
  (
    n977,
    n911,
    n906,
    n910,
    n932
  );


  xnor
  g956
  (
    n981,
    n921,
    n920,
    n936,
    n912
  );


  xor
  g957
  (
    n971,
    n940,
    n922,
    n913,
    n895
  );


  not
  g958
  (
    n991,
    n971
  );


  not
  g959
  (
    n985,
    n970
  );


  buf
  g960
  (
    n990,
    n982
  );


  buf
  g961
  (
    n987,
    n982
  );


  not
  g962
  (
    n995,
    n972
  );


  not
  g963
  (
    n992,
    n974
  );


  not
  g964
  (
    n986,
    n980
  );


  buf
  g965
  (
    n993,
    n981
  );


  not
  g966
  (
    n984,
    n976
  );


  buf
  g967
  (
    n997,
    n968
  );


  buf
  g968
  (
    n983,
    n973
  );


  not
  g969
  (
    n994,
    n975
  );


  not
  g970
  (
    n996,
    n977
  );


  not
  g971
  (
    n989,
    n978
  );


  buf
  g972
  (
    n998,
    n979
  );


  not
  g973
  (
    n988,
    n969
  );


  buf
  g974
  (
    KeyWire_0_14,
    n983
  );


  buf
  g975
  (
    n1005,
    n988
  );


  not
  g976
  (
    n1007,
    n989
  );


  not
  g977
  (
    n1009,
    n987
  );


  buf
  g978
  (
    n1015,
    n986
  );


  not
  g979
  (
    n1006,
    n987
  );


  buf
  g980
  (
    n1022,
    n989
  );


  not
  g981
  (
    n1014,
    n985
  );


  not
  g982
  (
    n1008,
    n988
  );


  not
  g983
  (
    n1019,
    n986
  );


  buf
  g984
  (
    n1020,
    n989
  );


  not
  g985
  (
    n1012,
    n986
  );


  not
  g986
  (
    n1021,
    n985
  );


  not
  g987
  (
    n1011,
    n988
  );


  buf
  g988
  (
    n1017,
    n983
  );


  not
  g989
  (
    n999,
    n987
  );


  buf
  g990
  (
    n1001,
    n984
  );


  buf
  g991
  (
    n1000,
    n986
  );


  not
  g992
  (
    n1010,
    n987
  );


  not
  g993
  (
    n1002,
    n989
  );


  buf
  g994
  (
    n1018,
    n984
  );


  not
  g995
  (
    n1004,
    n985
  );


  not
  g996
  (
    n1003,
    n988
  );


  not
  g997
  (
    n1013,
    n985
  );


  xor
  g998
  (
    n1071,
    n348,
    n349,
    n321,
    n1015
  );


  nor
  g999
  (
    n1103,
    n638,
    n340,
    n352,
    n327
  );


  nand
  g1000
  (
    n1043,
    n312,
    n314,
    n307,
    n309
  );


  nor
  g1001
  (
    n1090,
    n345,
    n350,
    n327,
    n331
  );


  nand
  g1002
  (
    n1044,
    n345,
    n1004,
    n362,
    n305
  );


  nor
  g1003
  (
    n1099,
    n356,
    n316,
    n1001,
    n633
  );


  nand
  g1004
  (
    n1064,
    n353,
    n1012,
    n308,
    n316
  );


  or
  g1005
  (
    n1107,
    n351,
    n1014,
    n1008,
    n334
  );


  and
  g1006
  (
    n1075,
    n326,
    n1015,
    n328,
    n337
  );


  xor
  g1007
  (
    n1034,
    n353,
    n304,
    n334,
    n315
  );


  xor
  g1008
  (
    n1048,
    n357,
    n618,
    n649,
    n309
  );


  xnor
  g1009
  (
    n1085,
    n644,
    n341,
    n628,
    n328
  );


  xnor
  g1010
  (
    n1038,
    n1018,
    n630,
    n647,
    n629
  );


  xor
  g1011
  (
    n1106,
    n321,
    n1002,
    n1020,
    n347
  );


  nor
  g1012
  (
    n1116,
    n1020,
    n335,
    n334,
    n311
  );


  xor
  g1013
  (
    n1058,
    n327,
    n1005,
    n616,
    n619
  );


  nand
  g1014
  (
    n1028,
    n1007,
    n1016,
    n335,
    n322
  );


  or
  g1015
  (
    n1053,
    n1018,
    n333,
    n1021,
    n1017
  );


  xnor
  g1016
  (
    n1050,
    n1009,
    n309,
    n1016,
    n623
  );


  nand
  g1017
  (
    n1055,
    n360,
    n315,
    n325,
    n1000
  );


  xor
  g1018
  (
    n1080,
    n333,
    n329,
    n364,
    n352
  );


  xor
  g1019
  (
    n1114,
    n338,
    n363,
    n361,
    n640
  );


  nand
  g1020
  (
    n1083,
    n1008,
    n332,
    n1011,
    n364
  );


  and
  g1021
  (
    n1036,
    n339,
    n1000,
    n359,
    n306
  );


  nor
  g1022
  (
    n1061,
    n1001,
    n346,
    n315,
    n322
  );


  and
  g1023
  (
    n1027,
    n360,
    n1013,
    n343,
    n325
  );


  xnor
  g1024
  (
    n1066,
    n353,
    n364,
    n348,
    n338
  );


  nand
  g1025
  (
    n1098,
    n1010,
    n336,
    n331,
    n1005
  );


  xor
  g1026
  (
    n1087,
    n344,
    n1011,
    n341,
    n363
  );


  nand
  g1027
  (
    n1041,
    n1000,
    n361,
    n1002,
    n1004
  );


  xor
  g1028
  (
    n1029,
    n330,
    n632,
    n1017,
    n329
  );


  or
  g1029
  (
    n1035,
    n1008,
    n339,
    n1000,
    n347
  );


  nand
  g1030
  (
    n1100,
    n318,
    n345,
    n324,
    n1009
  );


  nor
  g1031
  (
    n1024,
    n323,
    n349,
    n362,
    n361
  );


  nor
  g1032
  (
    n1072,
    n319,
    n320,
    n327,
    n341
  );


  xor
  g1033
  (
    n1088,
    n318,
    n1002,
    n326,
    n359
  );


  or
  g1034
  (
    n1054,
    n1010,
    n1006,
    n361,
    n357
  );


  xnor
  g1035
  (
    n1076,
    n353,
    n349,
    n1014,
    n626
  );


  nand
  g1036
  (
    n1065,
    n641,
    n342,
    n346
  );


  and
  g1037
  (
    n1091,
    n310,
    n1019,
    n338,
    n342
  );


  nor
  g1038
  (
    n1060,
    n355,
    n329,
    n348,
    n314
  );


  and
  g1039
  (
    n1069,
    n304,
    n326,
    n311,
    n1001
  );


  nand
  g1040
  (
    n1084,
    n346,
    n310,
    n305,
    n333
  );


  and
  g1041
  (
    n1057,
    n340,
    n1019,
    n624,
    n332
  );


  xnor
  g1042
  (
    n1023,
    n358,
    n1007,
    n312,
    n1003
  );


  nand
  g1043
  (
    n1089,
    n324,
    n639,
    n321,
    n305
  );


  nand
  g1044
  (
    n1073,
    n1009,
    n651,
    n637,
    n1006
  );


  and
  g1045
  (
    n1109,
    n645,
    n337,
    n310,
    n341
  );


  and
  g1046
  (
    n1067,
    n1007,
    n318,
    n627,
    n343
  );


  nor
  g1047
  (
    n1105,
    n1017,
    n650,
    n322,
    n324
  );


  nor
  g1048
  (
    n1082,
    n308,
    n1011,
    n651,
    n1022
  );


  nor
  g1049
  (
    n1101,
    n335,
    n634,
    n1014,
    n339
  );


  nand
  g1050
  (
    n1115,
    n323,
    n362,
    n1009,
    n307
  );


  nand
  g1051
  (
    n1102,
    n338,
    n317,
    n363,
    n1019
  );


  and
  g1052
  (
    n1110,
    n337,
    n357,
    n1007,
    n1006
  );


  nor
  g1053
  (
    n1045,
    n1021,
    n1021,
    n1015,
    n1013
  );


  nand
  g1054
  (
    n1031,
    n356,
    n306,
    n362,
    n316
  );


  or
  g1055
  (
    n1112,
    n329,
    n336,
    n310,
    n335
  );


  and
  g1056
  (
    n1093,
    n1008,
    n337,
    n355,
    n314
  );


  or
  g1057
  (
    n1079,
    n351,
    n348,
    n1018,
    n1022
  );


  and
  g1058
  (
    n1026,
    n325,
    n307,
    n324,
    n345
  );


  and
  g1059
  (
    KeyWire_0_21,
    n317,
    n354,
    n316,
    n999
  );


  nand
  g1060
  (
    n1033,
    n347,
    n351,
    n356,
    n1016
  );


  nor
  g1061
  (
    n1030,
    n330,
    n308,
    n350,
    n1002
  );


  nand
  g1062
  (
    n1068,
    n1010,
    n317,
    n1015,
    n643
  );


  xnor
  g1063
  (
    n1111,
    n1022,
    n1018,
    n312,
    n319
  );


  xnor
  g1064
  (
    n1078,
    n1019,
    n352,
    n313,
    n1016
  );


  xnor
  g1065
  (
    n1097,
    n1011,
    n321,
    n309,
    n631
  );


  xnor
  g1066
  (
    n1063,
    n360,
    n306,
    n326,
    n363
  );


  nand
  g1067
  (
    n1056,
    n305,
    n328,
    n330
  );


  and
  g1068
  (
    n1039,
    n340,
    n1003,
    n360,
    n356
  );


  nor
  g1069
  (
    n1094,
    n617,
    n358,
    n1012,
    n311
  );


  nand
  g1070
  (
    n1051,
    n313,
    n635,
    n1021,
    n342
  );


  xor
  g1071
  (
    n1062,
    n349,
    n319,
    n312,
    n320
  );


  xnor
  g1072
  (
    n1040,
    n320,
    n307,
    n336,
    n646
  );


  xor
  g1073
  (
    n1077,
    n642,
    n1004,
    n1010,
    n1020
  );


  and
  g1074
  (
    n1025,
    n317,
    n320,
    n331,
    n358
  );


  nor
  g1075
  (
    n1081,
    n350,
    n323,
    n622,
    n365
  );


  nor
  g1076
  (
    n1092,
    n344,
    n621,
    n1003
  );


  or
  g1077
  (
    n1113,
    n1020,
    n306,
    n1017,
    n636
  );


  and
  g1078
  (
    n1047,
    n333,
    n358,
    n1022,
    n1012
  );


  xor
  g1079
  (
    n1059,
    n354,
    n322,
    n339,
    n350
  );


  or
  g1080
  (
    n1086,
    n620,
    n332,
    n364,
    n999
  );


  xor
  g1081
  (
    n1070,
    n1005,
    n314,
    n331,
    n355
  );


  xnor
  g1082
  (
    n1096,
    n355,
    n1013,
    n1014,
    n1006
  );


  or
  g1083
  (
    n1104,
    n313,
    n325,
    n332,
    n625
  );


  nor
  g1084
  (
    n1042,
    n359,
    n351,
    n1012,
    n304
  );


  nand
  g1085
  (
    n1046,
    n346,
    n1013,
    n304,
    n340
  );


  nor
  g1086
  (
    n1037,
    n1001,
    n313,
    n343,
    n347
  );


  or
  g1087
  (
    n1074,
    n330,
    n343,
    n344,
    n357
  );


  xor
  g1088
  (
    n1108,
    n344,
    n1005,
    n352,
    n318
  );


  nor
  g1089
  (
    n1049,
    n319,
    n308,
    n336,
    n311
  );


  and
  g1090
  (
    n1052,
    n354,
    n1004,
    n323,
    n315
  );


  and
  g1091
  (
    n1032,
    n334,
    n359,
    n648,
    n354
  );


  not
  g1092
  (
    n1118,
    n1044
  );


  buf
  g1093
  (
    n1154,
    n1055
  );


  not
  g1094
  (
    n1155,
    n1045
  );


  buf
  g1095
  (
    n1133,
    n1048
  );


  buf
  g1096
  (
    n1137,
    n1051
  );


  not
  g1097
  (
    n1148,
    n1039
  );


  buf
  g1098
  (
    n1117,
    n1049
  );


  buf
  g1099
  (
    n1129,
    n1028
  );


  buf
  g1100
  (
    n1122,
    n1031
  );


  not
  g1101
  (
    n1125,
    n1037
  );


  not
  g1102
  (
    n1152,
    n1056
  );


  not
  g1103
  (
    n1153,
    n1046
  );


  not
  g1104
  (
    n1149,
    n1047
  );


  buf
  g1105
  (
    n1146,
    n1052
  );


  not
  g1106
  (
    n1143,
    n1026
  );


  not
  g1107
  (
    n1130,
    n1050
  );


  not
  g1108
  (
    n1136,
    n1061
  );


  not
  g1109
  (
    n1147,
    n1023
  );


  buf
  g1110
  (
    KeyWire_0_28,
    n1062
  );


  buf
  g1111
  (
    n1156,
    n1042
  );


  not
  g1112
  (
    n1132,
    n1038
  );


  not
  g1113
  (
    n1151,
    n1035
  );


  not
  g1114
  (
    n1142,
    n1034
  );


  buf
  g1115
  (
    n1131,
    n1032
  );


  buf
  g1116
  (
    n1120,
    n1054
  );


  buf
  g1117
  (
    n1150,
    n1057
  );


  not
  g1118
  (
    n1140,
    n1024
  );


  not
  g1119
  (
    n1141,
    n1040
  );


  buf
  g1120
  (
    n1134,
    n1027
  );


  buf
  g1121
  (
    n1139,
    n1059
  );


  not
  g1122
  (
    n1138,
    n1036
  );


  buf
  g1123
  (
    n1128,
    n1025
  );


  not
  g1124
  (
    n1127,
    n1030
  );


  buf
  g1125
  (
    n1119,
    n1029
  );


  buf
  g1126
  (
    n1121,
    n1058
  );


  not
  g1127
  (
    n1126,
    n1033
  );


  not
  g1128
  (
    n1124,
    n1043
  );


  buf
  g1129
  (
    n1144,
    n1060
  );


  buf
  g1130
  (
    n1145,
    n1053
  );


  buf
  g1131
  (
    n1123,
    n1041
  );


  nand
  g1132
  (
    n1161,
    n1142,
    n1145,
    n1137
  );


  nand
  g1133
  (
    n1190,
    n1132,
    n1150,
    n994,
    n368
  );


  xnor
  g1134
  (
    n1197,
    n1135,
    n847,
    n1143,
    n844
  );


  or
  g1135
  (
    n1169,
    n1119,
    n1119,
    n369,
    n380
  );


  and
  g1136
  (
    n1211,
    n1065,
    n1128,
    n1123,
    n849
  );


  xor
  g1137
  (
    n1226,
    n846,
    n846,
    n1156,
    n1127
  );


  and
  g1138
  (
    n1198,
    n997,
    n995,
    n841,
    n1082
  );


  and
  g1139
  (
    n1162,
    n1138,
    n1147,
    n1153,
    n1071
  );


  xnor
  g1140
  (
    n1225,
    n847,
    n1068,
    n374,
    n375
  );


  and
  g1141
  (
    n1187,
    n366,
    n843,
    n372,
    n1129
  );


  or
  g1142
  (
    n1224,
    n368,
    n851,
    n1067,
    n997
  );


  nand
  g1143
  (
    n1244,
    n1148,
    n1134,
    n375,
    n848
  );


  xor
  g1144
  (
    n1246,
    n825,
    n365,
    n370,
    n996
  );


  xnor
  g1145
  (
    n1191,
    n843,
    n1066,
    n1081,
    n1121
  );


  nand
  g1146
  (
    n1204,
    n366,
    n841,
    n1149,
    n998
  );


  or
  g1147
  (
    n1201,
    n1120,
    n840,
    n1070,
    n822
  );


  or
  g1148
  (
    n1184,
    n1137,
    n828,
    n1072,
    n1152
  );


  nand
  g1149
  (
    n1239,
    n1118,
    n1140,
    n1131,
    n1119
  );


  nand
  g1150
  (
    n1180,
    n383,
    n997,
    n1133,
    n1123
  );


  and
  g1151
  (
    n1241,
    n1146,
    n993,
    n1142,
    n1144
  );


  nand
  g1152
  (
    n1221,
    n1117,
    n842,
    n1127,
    n1142
  );


  or
  g1153
  (
    n1194,
    n1124,
    n1154,
    n1130,
    n1129
  );


  xnor
  g1154
  (
    n1216,
    n371,
    n848,
    n1138,
    n1131
  );


  nand
  g1155
  (
    n1218,
    n1140,
    n1143,
    n837
  );


  xnor
  g1156
  (
    n1167,
    n1118,
    n369,
    n990,
    n1133
  );


  xor
  g1157
  (
    n1196,
    n1132,
    n1150,
    n1141,
    n1133
  );


  xnor
  g1158
  (
    n1163,
    n372,
    n827,
    n835,
    n1123
  );


  xor
  g1159
  (
    n1250,
    n1152,
    n992,
    n379,
    n376
  );


  nor
  g1160
  (
    n1193,
    n990,
    n852,
    n842,
    n844
  );


  and
  g1161
  (
    n1240,
    n365,
    n1126,
    n1147,
    n1128
  );


  or
  g1162
  (
    KeyWire_0_30,
    n368,
    n1145,
    n1139,
    n1124
  );


  or
  g1163
  (
    n1249,
    n367,
    n991,
    n1126,
    n1144
  );


  and
  g1164
  (
    n1248,
    n1148,
    n369,
    n821,
    n1127
  );


  or
  g1165
  (
    n1189,
    n373,
    n852,
    n1151,
    n848
  );


  and
  g1166
  (
    n1220,
    n845,
    n823,
    n1118,
    n1128
  );


  or
  g1167
  (
    n1251,
    n1136,
    n1122,
    n1146,
    n830
  );


  and
  g1168
  (
    n1206,
    n844,
    n1129,
    n1076,
    n1145
  );


  or
  g1169
  (
    n1179,
    n1081,
    n367,
    n372,
    n996
  );


  or
  g1170
  (
    n1202,
    n384,
    n380,
    n832,
    n996
  );


  and
  g1171
  (
    n1181,
    n850,
    n833,
    n1079,
    n1124
  );


  or
  g1172
  (
    n1200,
    n991,
    n377,
    n366,
    n1122
  );


  or
  g1173
  (
    n1186,
    n998,
    n373,
    n1150,
    n378
  );


  nor
  g1174
  (
    n1212,
    n380,
    n383,
    n833,
    n1130
  );


  nor
  g1175
  (
    n1233,
    n838,
    n1134,
    n1121,
    n376
  );


  xnor
  g1176
  (
    n1217,
    n845,
    n1080,
    n825,
    n368
  );


  xnor
  g1177
  (
    n1231,
    n374,
    n851,
    n1135,
    n1154
  );


  nor
  g1178
  (
    n1219,
    n1117,
    n1149,
    n843,
    n378
  );


  xor
  g1179
  (
    n1242,
    n1082,
    n1156,
    n1155,
    n823
  );


  or
  g1180
  (
    n1174,
    n838,
    n847,
    n365,
    n1122
  );


  nand
  g1181
  (
    n1247,
    n381,
    n1140,
    n842,
    n1149
  );


  or
  g1182
  (
    n1223,
    n998,
    n996,
    n836,
    n1126
  );


  or
  g1183
  (
    n1209,
    n846,
    n1138,
    n1139,
    n836
  );


  and
  g1184
  (
    n1173,
    n851,
    n832,
    n378,
    n1134
  );


  and
  g1185
  (
    n1253,
    n850,
    n995,
    n831,
    n372
  );


  xor
  g1186
  (
    n1213,
    n991,
    n1147,
    n370,
    n1148
  );


  xor
  g1187
  (
    n1199,
    n824,
    n375,
    n1140,
    n1135
  );


  and
  g1188
  (
    n1188,
    n1125,
    n845,
    n829,
    n1146
  );


  nand
  g1189
  (
    n1165,
    n840,
    n835,
    n828,
    n1075
  );


  xnor
  g1190
  (
    n1168,
    n380,
    n826,
    n993,
    n379
  );


  nor
  g1191
  (
    n1183,
    n1120,
    n1138,
    n1117,
    n1126
  );


  or
  g1192
  (
    n1208,
    n1123,
    n382,
    n1150,
    n377
  );


  and
  g1193
  (
    n1175,
    n382,
    n849,
    n1151
  );


  and
  g1194
  (
    n1230,
    n998,
    n1121,
    n1155,
    n383
  );


  or
  g1195
  (
    n1210,
    n1124,
    n849,
    n994,
    n1154
  );


  nor
  g1196
  (
    n1195,
    n1129,
    n1079,
    n827,
    n1144
  );


  and
  g1197
  (
    n1178,
    n1083,
    n841,
    n1135,
    n1136
  );


  nor
  g1198
  (
    n1172,
    n826,
    n1078,
    n377,
    n1120
  );


  nand
  g1199
  (
    n1177,
    n374,
    n379,
    n1146,
    n381
  );


  nor
  g1200
  (
    n1185,
    n1064,
    n1152,
    n1127,
    n824
  );


  nor
  g1201
  (
    n1157,
    n1148,
    n851,
    n1153,
    n378
  );


  and
  g1202
  (
    n1171,
    n1154,
    n1132,
    n834,
    n377
  );


  nand
  g1203
  (
    n1182,
    n1142,
    n995,
    n1134,
    n382
  );


  nand
  g1204
  (
    n1235,
    n1144,
    n990,
    n1125,
    n1121
  );


  nand
  g1205
  (
    n1214,
    n1119,
    n995,
    n1149,
    n383
  );


  and
  g1206
  (
    n1237,
    n1063,
    n1077,
    n831,
    n839
  );


  xnor
  g1207
  (
    n1238,
    n841,
    n1143,
    n993,
    n1147
  );


  or
  g1208
  (
    n1245,
    n381,
    n370,
    n844,
    n367
  );


  xor
  g1209
  (
    n1158,
    n384,
    n1156,
    n1141
  );


  xnor
  g1210
  (
    n1192,
    n1128,
    n1074,
    n852,
    n384
  );


  and
  g1211
  (
    n1205,
    n847,
    n990,
    n992
  );


  xnor
  g1212
  (
    n1160,
    n371,
    n1136,
    n1141
  );


  nor
  g1213
  (
    n1170,
    n846,
    n1131,
    n1139,
    n369
  );


  nor
  g1214
  (
    n1166,
    n371,
    n1125,
    n1137,
    n830
  );


  nor
  g1215
  (
    n1164,
    n1137,
    n373,
    n370,
    n850
  );


  xor
  g1216
  (
    n1203,
    n843,
    n1155,
    n371,
    n373
  );


  or
  g1217
  (
    n1252,
    n992,
    n1117,
    n1152,
    n839
  );


  nor
  g1218
  (
    n1228,
    n822,
    n848,
    n1122,
    n367
  );


  xnor
  g1219
  (
    n1236,
    n1125,
    n1145,
    n1156,
    n1143
  );


  xor
  g1220
  (
    n1243,
    n1080,
    n376,
    n1151
  );


  xnor
  g1221
  (
    n1176,
    n993,
    n994,
    n1130,
    n375
  );


  xor
  g1222
  (
    n1232,
    n850,
    n1069,
    n997,
    n379
  );


  nor
  g1223
  (
    n1229,
    n842,
    n1153,
    n1133,
    n845
  );


  nand
  g1224
  (
    n1207,
    n1118,
    n834,
    n829,
    n991
  );


  nor
  g1225
  (
    n1215,
    n382,
    n852,
    n384,
    n381
  );


  and
  g1226
  (
    n1234,
    n1155,
    n1153,
    n994,
    n1131
  );


  xnor
  g1227
  (
    n1159,
    n1120,
    n366,
    n1130,
    n1132
  );


  nor
  g1228
  (
    n1227,
    n1073,
    n1139,
    n1151,
    n374
  );


  nand
  g1229
  (
    n1275,
    n720,
    n1227,
    n1173,
    n741
  );


  or
  g1230
  (
    n1342,
    n1201,
    n693,
    n1087,
    n1086
  );


  or
  g1231
  (
    n1297,
    n654,
    n683,
    n699,
    n749
  );


  or
  g1232
  (
    n1293,
    n1100,
    n725,
    n751,
    n685
  );


  and
  g1233
  (
    n1263,
    n1102,
    n742,
    n1105,
    n1219
  );


  and
  g1234
  (
    n1269,
    n734,
    n1178,
    n736
  );


  xnor
  g1235
  (
    n1296,
    n653,
    n1212,
    n963,
    n721
  );


  xnor
  g1236
  (
    n1330,
    n724,
    n730,
    n1215,
    n722
  );


  nand
  g1237
  (
    n1254,
    n707,
    n672,
    n961,
    n1229
  );


  or
  g1238
  (
    n1345,
    n745,
    n740,
    n1096,
    n1213
  );


  xnor
  g1239
  (
    n1295,
    n749,
    n690,
    n1251,
    n1099
  );


  xnor
  g1240
  (
    n1258,
    n962,
    n1084,
    n682,
    n1109
  );


  nor
  g1241
  (
    n1306,
    n689,
    n682,
    n1203,
    n1112
  );


  xnor
  g1242
  (
    n1262,
    n1102,
    n670,
    n1165,
    n674
  );


  nand
  g1243
  (
    n1294,
    n717,
    n721,
    n1084,
    n1237
  );


  nand
  g1244
  (
    n1267,
    n693,
    n679,
    n717,
    n738
  );


  nand
  g1245
  (
    n1325,
    n1191,
    n734,
    n713,
    n694
  );


  and
  g1246
  (
    KeyWire_0_18,
    n1189,
    n1221,
    n671,
    n957
  );


  or
  g1247
  (
    n1333,
    n718,
    n1192,
    n1232,
    n695
  );


  xnor
  g1248
  (
    n1282,
    n1185,
    n960,
    n716,
    n1244
  );


  and
  g1249
  (
    n1304,
    n733,
    n675,
    n700,
    n660
  );


  and
  g1250
  (
    n1312,
    n1095,
    n702,
    n1195,
    n1111
  );


  xor
  g1251
  (
    n1316,
    n658,
    n724,
    n1222,
    n664
  );


  nor
  g1252
  (
    n1303,
    n669,
    n656,
    n728,
    n1085
  );


  xnor
  g1253
  (
    n1319,
    n1115,
    n1083,
    n685,
    n667
  );


  nand
  g1254
  (
    n1311,
    n1233,
    n1096,
    n1163,
    n719
  );


  xor
  g1255
  (
    n1309,
    n1247,
    n715,
    n714,
    n1248
  );


  and
  g1256
  (
    n1308,
    n711,
    n1089,
    n1107,
    n1180
  );


  and
  g1257
  (
    n1313,
    n657,
    n696,
    n701,
    n684
  );


  and
  g1258
  (
    n1341,
    n695,
    n688,
    n677,
    n1114
  );


  nor
  g1259
  (
    n1332,
    n705,
    n710,
    n1239,
    n704
  );


  or
  g1260
  (
    n1317,
    n690,
    n672,
    n1181,
    n709
  );


  and
  g1261
  (
    n1302,
    n1169,
    n1115,
    n656,
    n698
  );


  xor
  g1262
  (
    n1335,
    n1087,
    n687,
    n726,
    n1182
  );


  nor
  g1263
  (
    n1277,
    n1093,
    n747,
    n707,
    n1176
  );


  nor
  g1264
  (
    n1291,
    n664,
    n673,
    n1242,
    n1160
  );


  xnor
  g1265
  (
    n1327,
    n1231,
    n1101,
    n701
  );


  xnor
  g1266
  (
    n1270,
    n1177,
    n1197,
    n731,
    n1091
  );


  nor
  g1267
  (
    n1322,
    n718,
    n1085,
    n1250,
    n657
  );


  nor
  g1268
  (
    n1307,
    n1190,
    n1100,
    n1217,
    n1194
  );


  xor
  g1269
  (
    n1346,
    n745,
    n727,
    n744,
    n668
  );


  xnor
  g1270
  (
    n1257,
    n748,
    n1164,
    n1179,
    n1094
  );


  nand
  g1271
  (
    n1310,
    n700,
    n716,
    n697,
    n967
  );


  and
  g1272
  (
    n1260,
    n1112,
    n681,
    n733,
    n753
  );


  nand
  g1273
  (
    n1271,
    n653,
    n1226,
    n1089,
    n738
  );


  xnor
  g1274
  (
    n1347,
    n688,
    n1090,
    n739,
    n1116
  );


  nand
  g1275
  (
    n1318,
    n663,
    n699,
    n1104,
    n1223
  );


  nor
  g1276
  (
    n1256,
    n966,
    n661,
    n1092,
    n735
  );


  or
  g1277
  (
    n1315,
    n1208,
    n1116,
    n1110,
    n1224
  );


  xnor
  g1278
  (
    n1290,
    n1162,
    n1111,
    n740,
    n964
  );


  and
  g1279
  (
    n1261,
    n729,
    n696,
    n692,
    n666
  );


  or
  g1280
  (
    n1328,
    n723,
    n1186,
    n1193,
    n1109
  );


  and
  g1281
  (
    n1334,
    n747,
    n1252,
    n719,
    n1113
  );


  xnor
  g1282
  (
    n1323,
    n742,
    n710,
    n1098,
    n712
  );


  or
  g1283
  (
    n1320,
    n1108,
    n679,
    n751,
    n705
  );


  nand
  g1284
  (
    n1259,
    n730,
    n680,
    n752,
    n729
  );


  nand
  g1285
  (
    n1279,
    n965,
    n741,
    n708,
    n1241
  );


  and
  g1286
  (
    n1283,
    n731,
    n708,
    n692,
    n743
  );


  nand
  g1287
  (
    n1305,
    n675,
    n1110,
    n659,
    n750
  );


  nand
  g1288
  (
    n1339,
    n722,
    n691,
    n1092,
    n686
  );


  nand
  g1289
  (
    n1278,
    n686,
    n1243,
    n1105,
    n1236
  );


  nand
  g1290
  (
    n1329,
    n1206,
    n956,
    n665,
    n666
  );


  or
  g1291
  (
    n1289,
    n659,
    n1218,
    n677,
    n683
  );


  nand
  g1292
  (
    KeyWire_0_31,
    n711,
    n1108,
    n1113,
    n1199
  );


  nor
  g1293
  (
    n1292,
    n655,
    n1106,
    n665
  );


  nand
  g1294
  (
    n1337,
    n663,
    n715,
    n655,
    n669
  );


  nand
  g1295
  (
    n1286,
    n1183,
    n966,
    n726,
    n732
  );


  and
  g1296
  (
    n1348,
    n1114,
    n1086,
    n703,
    n1166
  );


  xor
  g1297
  (
    KeyWire_0_19,
    n955,
    n661,
    n1225,
    n732
  );


  and
  g1298
  (
    n1326,
    n1175,
    n1235,
    n668,
    n703
  );


  xor
  g1299
  (
    n1265,
    n1204,
    n1099,
    n1187,
    n1094
  );


  nor
  g1300
  (
    n1344,
    n746,
    n1172,
    n684,
    n723
  );


  xor
  g1301
  (
    n1274,
    n1103,
    n1220,
    n1249,
    n652
  );


  xor
  g1302
  (
    n1284,
    n1097,
    n697,
    n673,
    n670
  );


  or
  g1303
  (
    n1276,
    n746,
    n680,
    n712,
    n1174
  );


  and
  g1304
  (
    n1314,
    n1200,
    n1196,
    n725,
    n1184
  );


  nand
  g1305
  (
    n1287,
    n654,
    n1245,
    n1188,
    n1161
  );


  xnor
  g1306
  (
    n1264,
    n728,
    n1170,
    n676,
    n1167
  );


  xnor
  g1307
  (
    n1336,
    n1240,
    n737,
    n1098,
    n662
  );


  xnor
  g1308
  (
    n1321,
    n667,
    n698,
    n706,
    n720
  );


  nor
  g1309
  (
    n1298,
    n694,
    n967,
    n1216,
    n706
  );


  xor
  g1310
  (
    n1255,
    n714,
    n744,
    n1091,
    n1171
  );


  xnor
  g1311
  (
    n1343,
    n1090,
    n1158,
    n735,
    n737
  );


  xnor
  g1312
  (
    n1349,
    n1107,
    n1238,
    n1088,
    n652
  );


  xnor
  g1313
  (
    n1281,
    n1103,
    n743,
    n1207,
    n660
  );


  xor
  g1314
  (
    n1268,
    n750,
    n671,
    n691,
    n1234
  );


  nor
  g1315
  (
    n1299,
    n681,
    n958,
    n1210,
    n674
  );


  and
  g1316
  (
    n1301,
    n748,
    n1246,
    n689,
    n678
  );


  nand
  g1317
  (
    n1280,
    n702,
    n1228,
    n1097,
    n704
  );


  xnor
  g1318
  (
    KeyWire_0_26,
    n687,
    n752,
    n1168,
    n1211
  );


  xor
  g1319
  (
    n1331,
    n1088,
    n1104,
    n713,
    n1253
  );


  xnor
  g1320
  (
    n1272,
    n739,
    n753,
    n1095,
    n959
  );


  nor
  g1321
  (
    n1288,
    n1093,
    n965,
    n1159,
    n1209
  );


  or
  g1322
  (
    n1300,
    n954,
    n727,
    n678,
    n709
  );


  nand
  g1323
  (
    n1338,
    n658,
    n1214,
    n676,
    n662
  );


  nor
  g1324
  (
    n1266,
    n1230,
    n1202,
    n1198,
    n1205
  );


  xor
  g1325
  (
    n1396,
    n1309,
    n1345,
    n1299,
    n1304
  );


  nand
  g1326
  (
    n1378,
    n1324,
    n1272,
    n1285,
    n1298
  );


  xnor
  g1327
  (
    n1413,
    n1323,
    n1303,
    n1307,
    n1267
  );


  and
  g1328
  (
    n1376,
    n1289,
    n1292,
    n1283,
    n1282
  );


  or
  g1329
  (
    n1410,
    n1263,
    n1287,
    n1277,
    n1318
  );


  nand
  g1330
  (
    n1428,
    n1322,
    n1312,
    n1327,
    n1266
  );


  xor
  g1331
  (
    n1398,
    n1344,
    n1326,
    n1283,
    n1337
  );


  and
  g1332
  (
    n1374,
    n1309,
    n1281,
    n1254
  );


  xor
  g1333
  (
    n1367,
    n1304,
    n1329,
    n1288,
    n1258
  );


  xnor
  g1334
  (
    n1356,
    n1291,
    n1294,
    n1256
  );


  xor
  g1335
  (
    n1364,
    n1301,
    n1259,
    n1290,
    n1317
  );


  xor
  g1336
  (
    n1393,
    n1297,
    n1305,
    n1340,
    n1341
  );


  and
  g1337
  (
    n1425,
    n1286,
    n1341,
    n1326,
    n1315
  );


  xnor
  g1338
  (
    n1414,
    n1261,
    n1314,
    n1331,
    n1279
  );


  nand
  g1339
  (
    n1427,
    n1329,
    n1320,
    n1293,
    n1340
  );


  and
  g1340
  (
    n1368,
    n1339,
    n1278,
    n1307,
    n1326
  );


  or
  g1341
  (
    n1400,
    n1286,
    n1276,
    n1324,
    n1296
  );


  or
  g1342
  (
    n1429,
    n1349,
    n1324,
    n1284,
    n1311
  );


  and
  g1343
  (
    n1417,
    n1322,
    n1309,
    n1339,
    n1265
  );


  and
  g1344
  (
    n1397,
    n1302,
    n1312,
    n1268,
    n1328
  );


  and
  g1345
  (
    n1401,
    n1345,
    n1346,
    n1343,
    n1336
  );


  nand
  g1346
  (
    n1424,
    n1318,
    n1318,
    n1295,
    n1290
  );


  or
  g1347
  (
    n1420,
    n1316,
    n1280,
    n1277,
    n1337
  );


  xor
  g1348
  (
    n1419,
    n1271,
    n1313,
    n1299,
    n1323
  );


  xor
  g1349
  (
    KeyWire_0_5,
    n1327,
    n1288,
    n1349,
    n1283
  );


  nor
  g1350
  (
    n1377,
    n1311,
    n1257,
    n1335,
    n1310
  );


  nor
  g1351
  (
    n1383,
    n1344,
    n1304,
    n1341,
    n1349
  );


  xor
  g1352
  (
    n1379,
    n1271,
    n1342,
    n1257,
    n1287
  );


  nand
  g1353
  (
    n1359,
    n1284,
    n1279,
    n1343,
    n1308
  );


  xor
  g1354
  (
    n1380,
    n1330,
    n1330,
    n1319,
    n1255
  );


  xor
  g1355
  (
    n1363,
    n1275,
    n1339,
    n1320,
    n1329
  );


  nor
  g1356
  (
    n1402,
    n1315,
    n1298,
    n1338,
    n1285
  );


  or
  g1357
  (
    n1362,
    n1306,
    n1258,
    n1278,
    n1307
  );


  nand
  g1358
  (
    n1421,
    n1288,
    n1284,
    n1292,
    n1327
  );


  nor
  g1359
  (
    n1423,
    n1343,
    n1308,
    n1281,
    n1319
  );


  and
  g1360
  (
    n1418,
    n1332,
    n1287,
    n1331,
    n1274
  );


  nor
  g1361
  (
    n1384,
    n1334,
    n1308,
    n1342,
    n1317
  );


  and
  g1362
  (
    n1354,
    n1311,
    n1265,
    n1317,
    n1322
  );


  nor
  g1363
  (
    n1355,
    n1336,
    n1331,
    n1297,
    n1270
  );


  and
  g1364
  (
    n1352,
    n1330,
    n1319,
    n1345,
    n1290
  );


  nor
  g1365
  (
    n1381,
    n1286,
    n1334,
    n1283,
    n1264
  );


  nor
  g1366
  (
    n1350,
    n1346,
    n1305,
    n1278,
    n1296
  );


  nor
  g1367
  (
    n1370,
    n1301,
    n1290,
    n1255,
    n1280
  );


  and
  g1368
  (
    n1416,
    n1325,
    n1260,
    n1270,
    n1289
  );


  nor
  g1369
  (
    n1399,
    n1295,
    n1312,
    n1313,
    n1343
  );


  or
  g1370
  (
    n1422,
    n1264,
    n1314,
    n1348,
    n1282
  );


  xnor
  g1371
  (
    n1372,
    n1299,
    n1254,
    n1260,
    n1315
  );


  xnor
  g1372
  (
    n1409,
    n1335,
    n1289,
    n1316,
    n1337
  );


  nand
  g1373
  (
    n1387,
    n1295,
    n1306,
    n1327,
    n1279
  );


  nand
  g1374
  (
    n1433,
    n1319,
    n1262,
    n1303,
    n1259
  );


  and
  g1375
  (
    n1408,
    n1268,
    n1347,
    n1325,
    n1284
  );


  nor
  g1376
  (
    n1431,
    n1295,
    n1338,
    n1293,
    n1298
  );


  or
  g1377
  (
    n1373,
    n1294,
    n1348,
    n1309,
    n1310
  );


  or
  g1378
  (
    n1395,
    n1289,
    n1313,
    n1310,
    n1336
  );


  nand
  g1379
  (
    n1353,
    n1296,
    n1276,
    n1321,
    n1285
  );


  xnor
  g1380
  (
    KeyWire_0_0,
    n1312,
    n1282,
    n1291,
    n1337
  );


  and
  g1381
  (
    n1403,
    n1313,
    n1302,
    n1340,
    n1342
  );


  xnor
  g1382
  (
    n1389,
    n1347,
    n1332,
    n1267,
    n1298
  );


  nor
  g1383
  (
    n1358,
    n1310,
    n1307,
    n1263,
    n1300
  );


  nand
  g1384
  (
    n1388,
    n1314,
    n1274,
    n1344,
    n1293
  );


  and
  g1385
  (
    n1412,
    n1262,
    n1335,
    n1332,
    n1300
  );


  nor
  g1386
  (
    n1371,
    n1348,
    n1303,
    n1326,
    n1304
  );


  or
  g1387
  (
    n1369,
    n1272,
    n1302,
    n1336,
    n1282
  );


  xor
  g1388
  (
    n1394,
    n1338,
    n1288,
    n1349,
    n1346
  );


  or
  g1389
  (
    n1406,
    n1305,
    n1320,
    n1300,
    n1342
  );


  nor
  g1390
  (
    n1382,
    n1275,
    n1279,
    n1301,
    n1292
  );


  nor
  g1391
  (
    n1375,
    n1339,
    n1347,
    n1314,
    n1340
  );


  xnor
  g1392
  (
    n1385,
    n1333,
    n1321,
    n1324
  );


  nand
  g1393
  (
    n1386,
    n1328,
    n1317,
    n1305,
    n1301
  );


  nor
  g1394
  (
    n1426,
    n1296,
    n1329,
    n1338,
    n1334
  );


  or
  g1395
  (
    n1391,
    n1303,
    n1333,
    n1297,
    n1293
  );


  and
  g1396
  (
    n1366,
    n1316,
    n1328,
    n1333,
    n1285
  );


  nor
  g1397
  (
    n1361,
    n1331,
    n1332,
    n1261,
    n1315
  );


  xnor
  g1398
  (
    n1360,
    n1280,
    n1302,
    n1300,
    n1294
  );


  and
  g1399
  (
    n1432,
    n1330,
    n1321,
    n1328,
    n1318
  );


  nand
  g1400
  (
    n1415,
    n1287,
    n1316,
    n1323,
    n1299
  );


  xnor
  g1401
  (
    n1392,
    n1322,
    n1341,
    n1269
  );


  xnor
  g1402
  (
    n1390,
    n1320,
    n1256,
    n1306,
    n1308
  );


  xnor
  g1403
  (
    n1357,
    n1291,
    n1291,
    n1347,
    n1345
  );


  nor
  g1404
  (
    n1430,
    n1266,
    n1273,
    n1325,
    n1344
  );


  xnor
  g1405
  (
    n1365,
    n1306,
    n1278,
    n1348,
    n1325
  );


  xnor
  g1406
  (
    n1404,
    n1333,
    n1334,
    n1323,
    n1280
  );


  nand
  g1407
  (
    n1405,
    n1335,
    n1311,
    n1273,
    n1281
  );


  xor
  g1408
  (
    n1407,
    n1292,
    n1286,
    n1297,
    n1346
  );


  nand
  g1409
  (
    n1445,
    n1389,
    n1365,
    n1384,
    n1425
  );


  or
  g1410
  (
    n1439,
    n1370,
    n1361,
    n1382,
    n1426
  );


  nor
  g1411
  (
    n1436,
    n1350,
    n1364,
    n1383,
    n1391
  );


  nor
  g1412
  (
    n1452,
    n1394,
    n1373,
    n1418,
    n1352
  );


  xor
  g1413
  (
    n1443,
    n1400,
    n1379,
    n1398,
    n1399
  );


  nand
  g1414
  (
    n1434,
    n1408,
    n1406,
    n1362,
    n1431
  );


  or
  g1415
  (
    n1444,
    n1351,
    n1377,
    n1416,
    n1386
  );


  xnor
  g1416
  (
    n1441,
    n1414,
    n1422,
    n1415,
    n1413
  );


  nand
  g1417
  (
    n1446,
    n1409,
    n1353,
    n1411,
    n1407
  );


  nand
  g1418
  (
    n1447,
    n1424,
    n1363,
    n1360,
    n1369
  );


  or
  g1419
  (
    n1450,
    n1354,
    n1378,
    n1387,
    n1420
  );


  or
  g1420
  (
    n1440,
    n1355,
    n1419,
    n1402,
    n1404
  );


  nor
  g1421
  (
    n1435,
    n1396,
    n1393,
    n1356,
    n1417
  );


  nor
  g1422
  (
    n1448,
    n1428,
    n1371,
    n1430,
    n1397
  );


  nor
  g1423
  (
    n1449,
    n1429,
    n1368,
    n1390,
    n1401
  );


  xor
  g1424
  (
    n1437,
    n1423,
    n1376,
    n1367,
    n1410
  );


  nand
  g1425
  (
    n1451,
    n1381,
    n1366,
    n1392,
    n1433
  );


  xnor
  g1426
  (
    n1454,
    n1357,
    n1405,
    n1375,
    n1359
  );


  xnor
  g1427
  (
    n1438,
    n1358,
    n1372,
    n1395,
    n1427
  );


  nor
  g1428
  (
    n1453,
    n1385,
    n1374,
    n1421,
    n1412
  );


  xor
  g1429
  (
    n1442,
    n1403,
    n1380,
    n1432,
    n1388
  );


  xnor
  KeyGate_0_0
  (
    n1411,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n121,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n152,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n726,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n702,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n1351,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n175,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n615,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n631,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n130,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n107,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n508,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n701,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n525,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1016,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n353,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n699,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n547,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n1324,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n1273,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n517,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1095,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n595,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n278,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n969,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n407,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1340,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n721,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1135,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n28,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1222,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1285,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

