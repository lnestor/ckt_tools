

module Stat_1000_201
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n871,
  n847,
  n863,
  n850,
  n858,
  n841,
  n854,
  n852,
  n955,
  n966,
  n943,
  n965,
  n957,
  n956,
  n952,
  n958,
  n954,
  n961,
  n968,
  n946,
  n950,
  n970,
  n976,
  n973,
  n1021,
  n1025,
  n1023,
  n1028,
  n1031,
  n1030,
  n1032,
  n1029,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n871;
  output n847;
  output n863;
  output n850;
  output n858;
  output n841;
  output n854;
  output n852;
  output n955;
  output n966;
  output n943;
  output n965;
  output n957;
  output n956;
  output n952;
  output n958;
  output n954;
  output n961;
  output n968;
  output n946;
  output n950;
  output n970;
  output n976;
  output n973;
  output n1021;
  output n1025;
  output n1023;
  output n1028;
  output n1031;
  output n1030;
  output n1032;
  output n1029;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n848;
  wire n849;
  wire n851;
  wire n853;
  wire n855;
  wire n856;
  wire n857;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n944;
  wire n945;
  wire n947;
  wire n948;
  wire n949;
  wire n951;
  wire n953;
  wire n959;
  wire n960;
  wire n962;
  wire n963;
  wire n964;
  wire n967;
  wire n969;
  wire n971;
  wire n972;
  wire n974;
  wire n975;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1022;
  wire n1024;
  wire n1026;
  wire n1027;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n51,
    n6
  );


  not
  g1
  (
    n70,
    n31
  );


  buf
  g2
  (
    n131,
    n12
  );


  not
  g3
  (
    n154,
    n1
  );


  buf
  g4
  (
    n110,
    n7
  );


  not
  g5
  (
    n113,
    n3
  );


  not
  g6
  (
    n77,
    n31
  );


  not
  g7
  (
    n105,
    n17
  );


  not
  g8
  (
    n145,
    n7
  );


  not
  g9
  (
    n78,
    n15
  );


  not
  g10
  (
    n148,
    n18
  );


  buf
  g11
  (
    n129,
    n26
  );


  buf
  g12
  (
    n33,
    n11
  );


  not
  g13
  (
    n128,
    n21
  );


  not
  g14
  (
    n104,
    n3
  );


  buf
  g15
  (
    n119,
    n31
  );


  not
  g16
  (
    n97,
    n2
  );


  buf
  g17
  (
    n120,
    n17
  );


  buf
  g18
  (
    n138,
    n29
  );


  buf
  g19
  (
    n48,
    n6
  );


  buf
  g20
  (
    n90,
    n26
  );


  not
  g21
  (
    n92,
    n24
  );


  not
  g22
  (
    n144,
    n8
  );


  buf
  g23
  (
    n80,
    n22
  );


  not
  g24
  (
    n137,
    n25
  );


  buf
  g25
  (
    n108,
    n8
  );


  not
  g26
  (
    n151,
    n18
  );


  buf
  g27
  (
    n107,
    n8
  );


  buf
  g28
  (
    n50,
    n22
  );


  not
  g29
  (
    n63,
    n9
  );


  not
  g30
  (
    n62,
    n27
  );


  not
  g31
  (
    n140,
    n13
  );


  not
  g32
  (
    n123,
    n19
  );


  buf
  g33
  (
    n85,
    n19
  );


  buf
  g34
  (
    n156,
    n25
  );


  not
  g35
  (
    n44,
    n18
  );


  not
  g36
  (
    n114,
    n12
  );


  buf
  g37
  (
    n112,
    n22
  );


  not
  g38
  (
    n117,
    n5
  );


  not
  g39
  (
    n57,
    n28
  );


  buf
  g40
  (
    n139,
    n23
  );


  buf
  g41
  (
    n155,
    n11
  );


  buf
  g42
  (
    n126,
    n23
  );


  not
  g43
  (
    n40,
    n13
  );


  buf
  g44
  (
    n74,
    n5
  );


  buf
  g45
  (
    n106,
    n16
  );


  buf
  g46
  (
    n135,
    n1
  );


  buf
  g47
  (
    n149,
    n25
  );


  not
  g48
  (
    KeyWire_0_15,
    n7
  );


  buf
  g49
  (
    n86,
    n11
  );


  buf
  g50
  (
    n45,
    n10
  );


  buf
  g51
  (
    n143,
    n3
  );


  buf
  g52
  (
    n41,
    n18
  );


  not
  g53
  (
    n71,
    n29
  );


  buf
  g54
  (
    n73,
    n10
  );


  buf
  g55
  (
    n141,
    n4
  );


  buf
  g56
  (
    n121,
    n5
  );


  not
  g57
  (
    n58,
    n23
  );


  not
  g58
  (
    n94,
    n24
  );


  not
  g59
  (
    n47,
    n9
  );


  buf
  g60
  (
    n118,
    n19
  );


  not
  g61
  (
    n66,
    n28
  );


  buf
  g62
  (
    n95,
    n27
  );


  not
  g63
  (
    n87,
    n20
  );


  buf
  g64
  (
    n133,
    n28
  );


  not
  g65
  (
    n52,
    n29
  );


  buf
  g66
  (
    n124,
    n21
  );


  not
  g67
  (
    n98,
    n19
  );


  not
  g68
  (
    n43,
    n17
  );


  buf
  g69
  (
    n103,
    n22
  );


  buf
  g70
  (
    n56,
    n26
  );


  buf
  g71
  (
    n82,
    n12
  );


  buf
  g72
  (
    n38,
    n14
  );


  not
  g73
  (
    n81,
    n2
  );


  buf
  g74
  (
    n134,
    n17
  );


  buf
  g75
  (
    n147,
    n30
  );


  buf
  g76
  (
    n67,
    n15
  );


  buf
  g77
  (
    n35,
    n29
  );


  not
  g78
  (
    n152,
    n27
  );


  not
  g79
  (
    n64,
    n25
  );


  not
  g80
  (
    n96,
    n4
  );


  not
  g81
  (
    n91,
    n7
  );


  buf
  g82
  (
    n142,
    n24
  );


  not
  g83
  (
    n36,
    n21
  );


  buf
  g84
  (
    n61,
    n23
  );


  buf
  g85
  (
    n54,
    n10
  );


  buf
  g86
  (
    n39,
    n16
  );


  not
  g87
  (
    n65,
    n10
  );


  not
  g88
  (
    n59,
    n32
  );


  not
  g89
  (
    n122,
    n28
  );


  not
  g90
  (
    n132,
    n14
  );


  buf
  g91
  (
    n88,
    n4
  );


  not
  g92
  (
    n102,
    n20
  );


  buf
  g93
  (
    n109,
    n15
  );


  not
  g94
  (
    n76,
    n30
  );


  not
  g95
  (
    n72,
    n5
  );


  buf
  g96
  (
    n84,
    n15
  );


  not
  g97
  (
    n69,
    n30
  );


  buf
  g98
  (
    n127,
    n9
  );


  not
  g99
  (
    n55,
    n31
  );


  buf
  g100
  (
    n116,
    n12
  );


  not
  g101
  (
    n111,
    n6
  );


  not
  g102
  (
    n146,
    n13
  );


  not
  g103
  (
    n34,
    n21
  );


  buf
  g104
  (
    n89,
    n20
  );


  buf
  g105
  (
    n93,
    n9
  );


  not
  g106
  (
    n100,
    n11
  );


  buf
  g107
  (
    n53,
    n4
  );


  not
  g108
  (
    n60,
    n20
  );


  not
  g109
  (
    n153,
    n1
  );


  buf
  g110
  (
    n79,
    n13
  );


  buf
  g111
  (
    n42,
    n2
  );


  not
  g112
  (
    n125,
    n24
  );


  buf
  g113
  (
    n46,
    n16
  );


  not
  g114
  (
    n83,
    n6
  );


  not
  g115
  (
    n101,
    n30
  );


  buf
  g116
  (
    n136,
    n14
  );


  buf
  g117
  (
    n37,
    n3
  );


  not
  g118
  (
    n75,
    n16
  );


  not
  g119
  (
    n115,
    n14
  );


  not
  g120
  (
    n99,
    n26
  );


  not
  g121
  (
    n130,
    n27
  );


  not
  g122
  (
    n150,
    n8
  );


  buf
  g123
  (
    n68,
    n2
  );


  buf
  g124
  (
    n236,
    n89
  );


  not
  g125
  (
    n399,
    n81
  );


  buf
  g126
  (
    n410,
    n117
  );


  buf
  g127
  (
    n374,
    n52
  );


  buf
  g128
  (
    n322,
    n154
  );


  buf
  g129
  (
    n407,
    n39
  );


  not
  g130
  (
    KeyWire_0_10,
    n121
  );


  not
  g131
  (
    n288,
    n85
  );


  not
  g132
  (
    n245,
    n49
  );


  not
  g133
  (
    n224,
    n126
  );


  not
  g134
  (
    n257,
    n58
  );


  not
  g135
  (
    n246,
    n66
  );


  not
  g136
  (
    n300,
    n110
  );


  not
  g137
  (
    n433,
    n41
  );


  buf
  g138
  (
    n427,
    n135
  );


  not
  g139
  (
    n392,
    n36
  );


  not
  g140
  (
    n178,
    n35
  );


  buf
  g141
  (
    n317,
    n40
  );


  buf
  g142
  (
    n183,
    n106
  );


  buf
  g143
  (
    n185,
    n151
  );


  not
  g144
  (
    n434,
    n102
  );


  not
  g145
  (
    n237,
    n126
  );


  not
  g146
  (
    n174,
    n108
  );


  buf
  g147
  (
    n309,
    n143
  );


  buf
  g148
  (
    n318,
    n61
  );


  buf
  g149
  (
    n342,
    n44
  );


  buf
  g150
  (
    n331,
    n50
  );


  not
  g151
  (
    KeyWire_0_14,
    n150
  );


  buf
  g152
  (
    n321,
    n128
  );


  not
  g153
  (
    n217,
    n34
  );


  buf
  g154
  (
    n296,
    n80
  );


  buf
  g155
  (
    n388,
    n97
  );


  not
  g156
  (
    n378,
    n152
  );


  not
  g157
  (
    n219,
    n141
  );


  not
  g158
  (
    n370,
    n145
  );


  buf
  g159
  (
    n250,
    n39
  );


  not
  g160
  (
    n394,
    n128
  );


  buf
  g161
  (
    n170,
    n109
  );


  not
  g162
  (
    n166,
    n114
  );


  not
  g163
  (
    n382,
    n142
  );


  buf
  g164
  (
    n179,
    n83
  );


  not
  g165
  (
    n232,
    n50
  );


  not
  g166
  (
    n403,
    n81
  );


  buf
  g167
  (
    n228,
    n51
  );


  not
  g168
  (
    n314,
    n115
  );


  not
  g169
  (
    n262,
    n116
  );


  not
  g170
  (
    n160,
    n149
  );


  buf
  g171
  (
    n171,
    n74
  );


  not
  g172
  (
    n371,
    n55
  );


  buf
  g173
  (
    n240,
    n94
  );


  not
  g174
  (
    n199,
    n84
  );


  not
  g175
  (
    n249,
    n111
  );


  buf
  g176
  (
    n325,
    n114
  );


  buf
  g177
  (
    n337,
    n39
  );


  buf
  g178
  (
    n426,
    n98
  );


  not
  g179
  (
    n428,
    n33
  );


  not
  g180
  (
    n406,
    n38
  );


  not
  g181
  (
    n276,
    n104
  );


  buf
  g182
  (
    n226,
    n121
  );


  not
  g183
  (
    n292,
    n47
  );


  buf
  g184
  (
    n443,
    n56
  );


  not
  g185
  (
    n369,
    n57
  );


  buf
  g186
  (
    n400,
    n36
  );


  not
  g187
  (
    n347,
    n38
  );


  buf
  g188
  (
    n281,
    n67
  );


  buf
  g189
  (
    n381,
    n76
  );


  not
  g190
  (
    n188,
    n99
  );


  buf
  g191
  (
    n377,
    n147
  );


  not
  g192
  (
    n293,
    n141
  );


  buf
  g193
  (
    n405,
    n113
  );


  buf
  g194
  (
    n176,
    n103
  );


  not
  g195
  (
    n303,
    n75
  );


  buf
  g196
  (
    n338,
    n55
  );


  not
  g197
  (
    n316,
    n34
  );


  buf
  g198
  (
    n420,
    n136
  );


  not
  g199
  (
    n366,
    n134
  );


  buf
  g200
  (
    n215,
    n95
  );


  buf
  g201
  (
    n299,
    n115
  );


  not
  g202
  (
    n329,
    n33
  );


  not
  g203
  (
    n326,
    n127
  );


  not
  g204
  (
    n286,
    n144
  );


  buf
  g205
  (
    n421,
    n154
  );


  buf
  g206
  (
    n398,
    n122
  );


  buf
  g207
  (
    n157,
    n73
  );


  buf
  g208
  (
    n423,
    n49
  );


  buf
  g209
  (
    n206,
    n60
  );


  not
  g210
  (
    n162,
    n130
  );


  buf
  g211
  (
    n290,
    n75
  );


  not
  g212
  (
    n247,
    n130
  );


  buf
  g213
  (
    n213,
    n82
  );


  not
  g214
  (
    n356,
    n50
  );


  buf
  g215
  (
    KeyWire_0_0,
    n51
  );


  not
  g216
  (
    n279,
    n153
  );


  buf
  g217
  (
    n256,
    n139
  );


  not
  g218
  (
    n163,
    n82
  );


  not
  g219
  (
    n354,
    n71
  );


  not
  g220
  (
    n208,
    n83
  );


  buf
  g221
  (
    n308,
    n153
  );


  not
  g222
  (
    n263,
    n104
  );


  not
  g223
  (
    n319,
    n69
  );


  buf
  g224
  (
    n415,
    n138
  );


  buf
  g225
  (
    n436,
    n37
  );


  not
  g226
  (
    n203,
    n102
  );


  not
  g227
  (
    n209,
    n95
  );


  not
  g228
  (
    n181,
    n47
  );


  buf
  g229
  (
    n343,
    n53
  );


  not
  g230
  (
    n190,
    n118
  );


  buf
  g231
  (
    n417,
    n100
  );


  buf
  g232
  (
    n275,
    n70
  );


  not
  g233
  (
    n442,
    n111
  );


  buf
  g234
  (
    n412,
    n41
  );


  buf
  g235
  (
    n386,
    n83
  );


  not
  g236
  (
    n207,
    n135
  );


  buf
  g237
  (
    n327,
    n72
  );


  buf
  g238
  (
    n201,
    n127
  );


  not
  g239
  (
    n419,
    n142
  );


  buf
  g240
  (
    n324,
    n153
  );


  buf
  g241
  (
    n254,
    n57
  );


  buf
  g242
  (
    n367,
    n148
  );


  buf
  g243
  (
    n175,
    n62
  );


  buf
  g244
  (
    n159,
    n68
  );


  buf
  g245
  (
    n169,
    n54
  );


  not
  g246
  (
    n221,
    n145
  );


  buf
  g247
  (
    n204,
    n95
  );


  not
  g248
  (
    n306,
    n72
  );


  not
  g249
  (
    n233,
    n97
  );


  buf
  g250
  (
    n211,
    n147
  );


  not
  g251
  (
    n383,
    n35
  );


  not
  g252
  (
    n258,
    n152
  );


  not
  g253
  (
    n198,
    n66
  );


  buf
  g254
  (
    n333,
    n46
  );


  buf
  g255
  (
    n271,
    n71
  );


  not
  g256
  (
    n267,
    n131
  );


  not
  g257
  (
    KeyWire_0_3,
    n94
  );


  buf
  g258
  (
    n395,
    n151
  );


  not
  g259
  (
    n380,
    n140
  );


  not
  g260
  (
    n350,
    n48
  );


  not
  g261
  (
    n283,
    n137
  );


  not
  g262
  (
    KeyWire_0_11,
    n143
  );


  buf
  g263
  (
    n205,
    n93
  );


  not
  g264
  (
    n251,
    n133
  );


  buf
  g265
  (
    n365,
    n92
  );


  not
  g266
  (
    n411,
    n147
  );


  buf
  g267
  (
    n304,
    n52
  );


  not
  g268
  (
    n172,
    n48
  );


  buf
  g269
  (
    n298,
    n72
  );


  buf
  g270
  (
    n429,
    n101
  );


  buf
  g271
  (
    n297,
    n67
  );


  buf
  g272
  (
    n241,
    n149
  );


  not
  g273
  (
    n424,
    n129
  );


  buf
  g274
  (
    n362,
    n146
  );


  not
  g275
  (
    n242,
    n63
  );


  not
  g276
  (
    n387,
    n122
  );


  not
  g277
  (
    n282,
    n148
  );


  not
  g278
  (
    n401,
    n68
  );


  buf
  g279
  (
    n334,
    n129
  );


  not
  g280
  (
    n260,
    n94
  );


  buf
  g281
  (
    n345,
    n44
  );


  not
  g282
  (
    n189,
    n140
  );


  buf
  g283
  (
    n220,
    n86
  );


  buf
  g284
  (
    n408,
    n52
  );


  buf
  g285
  (
    n359,
    n105
  );


  buf
  g286
  (
    n344,
    n132
  );


  not
  g287
  (
    n280,
    n51
  );


  not
  g288
  (
    n285,
    n55
  );


  not
  g289
  (
    n200,
    n69
  );


  not
  g290
  (
    n210,
    n42
  );


  not
  g291
  (
    n158,
    n91
  );


  buf
  g292
  (
    n268,
    n116
  );


  not
  g293
  (
    n384,
    n133
  );


  not
  g294
  (
    n244,
    n109
  );


  buf
  g295
  (
    n368,
    n135
  );


  not
  g296
  (
    n379,
    n128
  );


  buf
  g297
  (
    n441,
    n107
  );


  not
  g298
  (
    n252,
    n107
  );


  buf
  g299
  (
    n349,
    n132
  );


  not
  g300
  (
    n414,
    n113
  );


  buf
  g301
  (
    n375,
    n96
  );


  buf
  g302
  (
    n230,
    n146
  );


  buf
  g303
  (
    n389,
    n108
  );


  not
  g304
  (
    n278,
    n100
  );


  not
  g305
  (
    n165,
    n42
  );


  not
  g306
  (
    n358,
    n85
  );


  not
  g307
  (
    KeyWire_0_1,
    n149
  );


  buf
  g308
  (
    n302,
    n34
  );


  buf
  g309
  (
    n255,
    n119
  );


  not
  g310
  (
    n301,
    n151
  );


  buf
  g311
  (
    n216,
    n37
  );


  buf
  g312
  (
    n161,
    n125
  );


  not
  g313
  (
    n231,
    n87
  );


  buf
  g314
  (
    n191,
    n86
  );


  buf
  g315
  (
    n335,
    n59
  );


  buf
  g316
  (
    n167,
    n58
  );


  not
  g317
  (
    n346,
    n124
  );


  buf
  g318
  (
    n432,
    n140
  );


  not
  g319
  (
    n248,
    n40
  );


  buf
  g320
  (
    n376,
    n88
  );


  not
  g321
  (
    n409,
    n108
  );


  buf
  g322
  (
    n364,
    n59
  );


  buf
  g323
  (
    n438,
    n131
  );


  not
  g324
  (
    n194,
    n117
  );


  not
  g325
  (
    n284,
    n65
  );


  not
  g326
  (
    n265,
    n56
  );


  buf
  g327
  (
    n440,
    n61
  );


  buf
  g328
  (
    n312,
    n38
  );


  not
  g329
  (
    n402,
    n110
  );


  buf
  g330
  (
    n239,
    n106
  );


  buf
  g331
  (
    n273,
    n111
  );


  not
  g332
  (
    n332,
    n154
  );


  buf
  g333
  (
    n192,
    n133
  );


  buf
  g334
  (
    n348,
    n124
  );


  buf
  g335
  (
    n393,
    n91
  );


  buf
  g336
  (
    n289,
    n112
  );


  not
  g337
  (
    n307,
    n115
  );


  not
  g338
  (
    n397,
    n35
  );


  buf
  g339
  (
    n272,
    n91
  );


  not
  g340
  (
    n270,
    n130
  );


  not
  g341
  (
    n391,
    n137
  );


  not
  g342
  (
    n363,
    n139
  );


  buf
  g343
  (
    n404,
    n123
  );


  buf
  g344
  (
    n339,
    n87
  );


  buf
  g345
  (
    n336,
    n54
  );


  buf
  g346
  (
    n385,
    n90
  );


  buf
  g347
  (
    n253,
    n112
  );


  not
  g348
  (
    n195,
    n126
  );


  buf
  g349
  (
    n187,
    n141
  );


  buf
  g350
  (
    n355,
    n88
  );


  not
  g351
  (
    n291,
    n42
  );


  buf
  g352
  (
    n164,
    n79
  );


  not
  g353
  (
    n182,
    n86
  );


  buf
  g354
  (
    n340,
    n106
  );


  not
  g355
  (
    n277,
    n93
  );


  buf
  g356
  (
    n180,
    n144
  );


  not
  g357
  (
    n227,
    n74
  );


  buf
  g358
  (
    n274,
    n110
  );


  buf
  g359
  (
    n416,
    n58
  );


  not
  g360
  (
    n444,
    n76
  );


  not
  g361
  (
    n222,
    n81
  );


  buf
  g362
  (
    n294,
    n129
  );


  not
  g363
  (
    n218,
    n134
  );


  not
  g364
  (
    n430,
    n87
  );


  not
  g365
  (
    n320,
    n75
  );


  not
  g366
  (
    n177,
    n98
  );


  not
  g367
  (
    n431,
    n99
  );


  buf
  g368
  (
    n184,
    n125
  );


  not
  g369
  (
    n261,
    n103
  );


  not
  g370
  (
    n341,
    n114
  );


  not
  g371
  (
    n225,
    n132
  );


  not
  g372
  (
    n305,
    n37
  );


  not
  g373
  (
    n295,
    n48
  );


  buf
  g374
  (
    n197,
    n136
  );


  buf
  g375
  (
    n223,
    n155
  );


  buf
  g376
  (
    n310,
    n80
  );


  buf
  g377
  (
    n196,
    n46
  );


  buf
  g378
  (
    n425,
    n57
  );


  buf
  g379
  (
    n357,
    n134
  );


  not
  g380
  (
    n259,
    n118
  );


  buf
  g381
  (
    n396,
    n93
  );


  buf
  g382
  (
    n373,
    n90
  );


  buf
  g383
  (
    n243,
    n60
  );


  buf
  g384
  (
    n186,
    n78
  );


  xor
  g385
  (
    n353,
    n41,
    n60
  );


  xnor
  g386
  (
    n437,
    n117,
    n33,
    n77,
    n113
  );


  nand
  g387
  (
    n229,
    n98,
    n45,
    n138,
    n85
  );


  xor
  g388
  (
    n193,
    n150,
    n36,
    n146,
    n88
  );


  xnor
  g389
  (
    n323,
    n70,
    n67,
    n62,
    n79
  );


  xnor
  g390
  (
    n435,
    n53,
    n64,
    n145,
    n70
  );


  or
  g391
  (
    n264,
    n121,
    n90,
    n79,
    n120
  );


  nor
  g392
  (
    n330,
    n77,
    n53,
    n54,
    n62
  );


  nand
  g393
  (
    n372,
    n74,
    n49,
    n66,
    n143
  );


  nand
  g394
  (
    n168,
    n112,
    n82,
    n123,
    n89
  );


  xnor
  g395
  (
    n238,
    n102,
    n43,
    n122,
    n107
  );


  xnor
  g396
  (
    n287,
    n116,
    n65,
    n105,
    n43
  );


  or
  g397
  (
    n361,
    n68,
    n119,
    n127,
    n64
  );


  nand
  g398
  (
    n352,
    n101,
    n44,
    n45
  );


  or
  g399
  (
    n234,
    n46,
    n59,
    n73,
    n84
  );


  xor
  g400
  (
    n422,
    n92,
    n96,
    n100
  );


  xor
  g401
  (
    n311,
    n152,
    n63,
    n43,
    n65
  );


  nand
  g402
  (
    n390,
    n71,
    n137,
    n47,
    n123
  );


  nand
  g403
  (
    n173,
    n89,
    n78,
    n109
  );


  and
  g404
  (
    n214,
    n99,
    n73,
    n142,
    n77
  );


  nand
  g405
  (
    n266,
    n101,
    n148,
    n63,
    n80
  );


  or
  g406
  (
    n439,
    n131,
    n76,
    n92,
    n105
  );


  or
  g407
  (
    n315,
    n64,
    n104,
    n120,
    n97
  );


  xor
  g408
  (
    n269,
    n118,
    n150,
    n136,
    n69
  );


  xnor
  g409
  (
    n360,
    n120,
    n84,
    n103,
    n144
  );


  xnor
  g410
  (
    n418,
    n56,
    n124,
    n139,
    n61
  );


  nand
  g411
  (
    n328,
    n40,
    n125,
    n119,
    n138
  );


  xor
  g412
  (
    n553,
    n274,
    n365,
    n330,
    n288
  );


  nor
  g413
  (
    n509,
    n390,
    n184,
    n320,
    n346
  );


  xor
  g414
  (
    n554,
    n272,
    n191,
    n179,
    n366
  );


  nor
  g415
  (
    n450,
    n322,
    n361,
    n365,
    n168
  );


  and
  g416
  (
    n447,
    n283,
    n197,
    n316,
    n311
  );


  or
  g417
  (
    n490,
    n278,
    n292,
    n386,
    n260
  );


  xnor
  g418
  (
    n488,
    n165,
    n232,
    n213,
    n247
  );


  or
  g419
  (
    n558,
    n262,
    n299,
    n234,
    n386
  );


  or
  g420
  (
    n599,
    n229,
    n354,
    n230,
    n351
  );


  nand
  g421
  (
    n526,
    n263,
    n362,
    n270,
    n230
  );


  xor
  g422
  (
    n583,
    n335,
    n394,
    n244,
    n393
  );


  xnor
  g423
  (
    n592,
    n374,
    n178,
    n275,
    n285
  );


  or
  g424
  (
    n533,
    n254,
    n232,
    n332,
    n290
  );


  or
  g425
  (
    n454,
    n385,
    n212,
    n215,
    n331
  );


  and
  g426
  (
    n517,
    n382,
    n308,
    n276,
    n252
  );


  xnor
  g427
  (
    n467,
    n392,
    n372,
    n274,
    n316
  );


  xor
  g428
  (
    n458,
    n202,
    n291,
    n282,
    n381
  );


  nand
  g429
  (
    n564,
    n334,
    n306,
    n293,
    n195
  );


  xor
  g430
  (
    n565,
    n312,
    n289,
    n320,
    n261
  );


  nand
  g431
  (
    n576,
    n201,
    n393,
    n333,
    n377
  );


  nand
  g432
  (
    n487,
    n182,
    n357,
    n342,
    n372
  );


  nor
  g433
  (
    n544,
    n199,
    n301,
    n277,
    n276
  );


  nand
  g434
  (
    n597,
    n249,
    n236,
    n318,
    n182
  );


  nand
  g435
  (
    n469,
    n396,
    n396,
    n283,
    n180
  );


  xor
  g436
  (
    n477,
    n171,
    n248,
    n395,
    n169
  );


  or
  g437
  (
    n507,
    n368,
    n255,
    n277,
    n328
  );


  nand
  g438
  (
    n545,
    n217,
    n372,
    n315,
    n392
  );


  nor
  g439
  (
    n522,
    n161,
    n288,
    n257,
    n211
  );


  nand
  g440
  (
    n459,
    n284,
    n395,
    n292,
    n307
  );


  nor
  g441
  (
    n465,
    n300,
    n302,
    n364,
    n309
  );


  and
  g442
  (
    n537,
    n259,
    n241,
    n173,
    n308
  );


  nand
  g443
  (
    n571,
    n352,
    n199,
    n190,
    n254
  );


  nand
  g444
  (
    n481,
    n363,
    n183,
    n394,
    n373
  );


  and
  g445
  (
    n499,
    n345,
    n366,
    n390,
    n175
  );


  xnor
  g446
  (
    n505,
    n298,
    n253,
    n387,
    n187
  );


  nor
  g447
  (
    n491,
    n297,
    n332,
    n388,
    n357
  );


  xor
  g448
  (
    n542,
    n386,
    n267,
    n172,
    n266
  );


  xnor
  g449
  (
    n562,
    n231,
    n387,
    n296,
    n345
  );


  nand
  g450
  (
    n575,
    n279,
    n158,
    n185,
    n253
  );


  and
  g451
  (
    n478,
    n242,
    n302,
    n387,
    n158
  );


  or
  g452
  (
    n574,
    n157,
    n212,
    n368,
    n381
  );


  xnor
  g453
  (
    n483,
    n318,
    n286,
    n364,
    n383
  );


  xor
  g454
  (
    n588,
    n258,
    n172,
    n162,
    n242
  );


  nand
  g455
  (
    n559,
    n338,
    n169,
    n240,
    n207
  );


  and
  g456
  (
    n600,
    n220,
    n319,
    n163,
    n346
  );


  xor
  g457
  (
    n446,
    n265,
    n175,
    n285,
    n223
  );


  and
  g458
  (
    n540,
    n316,
    n350,
    n297,
    n166
  );


  and
  g459
  (
    n535,
    n181,
    n185,
    n180,
    n384
  );


  or
  g460
  (
    n510,
    n243,
    n270,
    n351,
    n353
  );


  xnor
  g461
  (
    n550,
    n167,
    n215,
    n268,
    n304
  );


  nand
  g462
  (
    n474,
    n289,
    n375,
    n234,
    n296
  );


  or
  g463
  (
    n548,
    n360,
    n341,
    n373,
    n259
  );


  xnor
  g464
  (
    n513,
    n282,
    n334,
    n317,
    n319
  );


  or
  g465
  (
    n561,
    n221,
    n251,
    n218,
    n241
  );


  and
  g466
  (
    n568,
    n326,
    n318,
    n299,
    n164
  );


  xnor
  g467
  (
    n578,
    n320,
    n183,
    n225,
    n160
  );


  and
  g468
  (
    n515,
    n378,
    n356,
    n210,
    n396
  );


  and
  g469
  (
    n518,
    n330,
    n257,
    n173,
    n290
  );


  nor
  g470
  (
    n536,
    n233,
    n379,
    n323
  );


  xnor
  g471
  (
    n464,
    n262,
    n359,
    n354,
    n310
  );


  nor
  g472
  (
    n572,
    n267,
    n312,
    n245,
    n382
  );


  nand
  g473
  (
    n496,
    n343,
    n348,
    n222,
    n336
  );


  and
  g474
  (
    n506,
    n192,
    n305,
    n166,
    n304
  );


  and
  g475
  (
    n475,
    n355,
    n361,
    n250,
    n176
  );


  xor
  g476
  (
    n557,
    n192,
    n293,
    n252,
    n321
  );


  or
  g477
  (
    n460,
    n284,
    n294,
    n340,
    n303
  );


  or
  g478
  (
    n586,
    n314,
    n236,
    n174,
    n258
  );


  xor
  g479
  (
    n479,
    n295,
    n374,
    n174,
    n287
  );


  nand
  g480
  (
    n591,
    n378,
    n189,
    n295,
    n280
  );


  xnor
  g481
  (
    n589,
    n214,
    n296,
    n325,
    n339
  );


  and
  g482
  (
    n525,
    n306,
    n397,
    n377,
    n328
  );


  and
  g483
  (
    n551,
    n159,
    n321,
    n195,
    n293
  );


  nand
  g484
  (
    n449,
    n272,
    n206,
    n382,
    n246
  );


  and
  g485
  (
    n529,
    n177,
    n339,
    n371,
    n163
  );


  xnor
  g486
  (
    n451,
    n209,
    n340,
    n251,
    n356
  );


  xnor
  g487
  (
    n471,
    n333,
    n268,
    n353,
    n346
  );


  nand
  g488
  (
    n470,
    n395,
    n184,
    n349,
    n295
  );


  nor
  g489
  (
    n511,
    n325,
    n196,
    n377,
    n216
  );


  nand
  g490
  (
    n452,
    n304,
    n365,
    n221,
    n193
  );


  nand
  g491
  (
    n569,
    n392,
    n256,
    n362,
    n194
  );


  xnor
  g492
  (
    n566,
    n383,
    n275,
    n385,
    n343
  );


  nand
  g493
  (
    n555,
    n191,
    n312,
    n309,
    n314
  );


  xnor
  g494
  (
    n567,
    n351,
    n347,
    n266,
    n373
  );


  nor
  g495
  (
    n519,
    n343,
    n287,
    n326,
    n194
  );


  nor
  g496
  (
    n539,
    n264,
    n219,
    n335,
    n348
  );


  or
  g497
  (
    n585,
    n269,
    n285,
    n203,
    n176
  );


  or
  g498
  (
    n560,
    n235,
    n208,
    n266,
    n267
  );


  xor
  g499
  (
    n579,
    n201,
    n376,
    n352,
    n247
  );


  xnor
  g500
  (
    n455,
    n281,
    n324,
    n352,
    n338
  );


  and
  g501
  (
    KeyWire_0_4,
    n347,
    n301,
    n336,
    n292
  );


  xnor
  g502
  (
    n527,
    n282,
    n389,
    n278,
    n193
  );


  nor
  g503
  (
    n573,
    n273,
    n257,
    n186,
    n376
  );


  or
  g504
  (
    n472,
    n181,
    n294,
    n337,
    n210
  );


  nand
  g505
  (
    n570,
    n367,
    n385,
    n324,
    n391
  );


  and
  g506
  (
    n486,
    n313,
    n283,
    n381,
    n272
  );


  and
  g507
  (
    n530,
    n256,
    n379,
    n190,
    n289
  );


  xor
  g508
  (
    n594,
    n311,
    n356,
    n202,
    n238
  );


  xnor
  g509
  (
    n508,
    n237,
    n305,
    n342,
    n229
  );


  nand
  g510
  (
    n497,
    n369,
    n198,
    n349,
    n239
  );


  nor
  g511
  (
    n514,
    n261,
    n369,
    n329,
    n393
  );


  nor
  g512
  (
    n590,
    n275,
    n235,
    n279,
    n348
  );


  nand
  g513
  (
    n524,
    n265,
    n220,
    n269,
    n188
  );


  nand
  g514
  (
    n453,
    n265,
    n273,
    n164,
    n177
  );


  and
  g515
  (
    n448,
    n228,
    n213,
    n286,
    n340
  );


  or
  g516
  (
    n456,
    n345,
    n358,
    n363,
    n357
  );


  xor
  g517
  (
    n543,
    n354,
    n313,
    n189,
    n226
  );


  and
  g518
  (
    n484,
    n157,
    n271,
    n314,
    n281
  );


  or
  g519
  (
    n556,
    n211,
    n350,
    n233,
    n256
  );


  xor
  g520
  (
    n523,
    n170,
    n205,
    n206,
    n200
  );


  nand
  g521
  (
    n457,
    n380,
    n264,
    n227,
    n310
  );


  xnor
  g522
  (
    n463,
    n279,
    n325,
    n198,
    n291
  );


  xnor
  g523
  (
    n462,
    n287,
    n260,
    n331,
    n171
  );


  nor
  g524
  (
    KeyWire_0_5,
    n162,
    n226,
    n246,
    n294
  );


  xor
  g525
  (
    n532,
    n336,
    n208,
    n355,
    n260
  );


  xnor
  g526
  (
    n587,
    n219,
    n204,
    n390,
    n239
  );


  or
  g527
  (
    n503,
    n341,
    n300,
    n360,
    n259
  );


  or
  g528
  (
    n445,
    n324,
    n248,
    n380,
    n326
  );


  nand
  g529
  (
    n521,
    n355,
    n167,
    n353,
    n306
  );


  xor
  g530
  (
    n563,
    n187,
    n327,
    n376,
    n159
  );


  xnor
  g531
  (
    n528,
    n317,
    n337,
    n397,
    n244
  );


  xnor
  g532
  (
    n476,
    n261,
    n371,
    n209,
    n301
  );


  xor
  g533
  (
    n495,
    n371,
    n364,
    n280,
    n310
  );


  nand
  g534
  (
    n500,
    n263,
    n268,
    n350,
    n224
  );


  and
  g535
  (
    n582,
    n305,
    n297,
    n178,
    n307
  );


  xnor
  g536
  (
    n595,
    n245,
    n271,
    n224,
    n363
  );


  nor
  g537
  (
    n498,
    n338,
    n335,
    n264,
    n391
  );


  or
  g538
  (
    n473,
    n302,
    n327,
    n331,
    n328
  );


  xnor
  g539
  (
    n547,
    n160,
    n308,
    n231,
    n367
  );


  xnor
  g540
  (
    n502,
    n311,
    n374,
    n227,
    n378
  );


  nor
  g541
  (
    n492,
    n339,
    n280,
    n360,
    n271
  );


  xnor
  g542
  (
    n512,
    n222,
    n298,
    n367
  );


  and
  g543
  (
    n461,
    n375,
    n262,
    n223,
    n361
  );


  and
  g544
  (
    n493,
    n362,
    n228,
    n379,
    n315
  );


  or
  g545
  (
    n546,
    n237,
    n388,
    n359,
    n384
  );


  xnor
  g546
  (
    n549,
    n288,
    n214,
    n369,
    n286
  );


  nand
  g547
  (
    n552,
    n217,
    n258,
    n330,
    n225
  );


  nor
  g548
  (
    n468,
    n370,
    n276,
    n329,
    n344
  );


  xor
  g549
  (
    n501,
    n307,
    n165,
    n216,
    n290
  );


  and
  g550
  (
    n494,
    n309,
    n315,
    n359,
    n334
  );


  xnor
  g551
  (
    n485,
    n196,
    n341,
    n300,
    n332
  );


  nand
  g552
  (
    n593,
    n263,
    n329,
    n388,
    n273
  );


  xor
  g553
  (
    n489,
    n218,
    n370,
    n270,
    n333
  );


  and
  g554
  (
    n482,
    n322,
    n358,
    n284,
    n375
  );


  xnor
  g555
  (
    n534,
    n368,
    n319,
    n383,
    n322
  );


  and
  g556
  (
    n516,
    n207,
    n278,
    n274,
    n337
  );


  xnor
  g557
  (
    n577,
    n303,
    n281,
    n179,
    n391
  );


  and
  g558
  (
    n466,
    n323,
    n317,
    n349,
    n389
  );


  nand
  g559
  (
    n480,
    n291,
    n250,
    n170,
    n168
  );


  xor
  g560
  (
    n580,
    n321,
    n204,
    n370,
    n389
  );


  or
  g561
  (
    n520,
    n344,
    n186,
    n238,
    n161
  );


  nand
  g562
  (
    n504,
    n240,
    n313,
    n344,
    n205
  );


  and
  g563
  (
    n581,
    n200,
    n255,
    n384,
    n188
  );


  nor
  g564
  (
    n538,
    n397,
    n394,
    n380,
    n327
  );


  and
  g565
  (
    n598,
    n347,
    n358,
    n249,
    n269
  );


  or
  g566
  (
    n584,
    n277,
    n203,
    n303,
    n342
  );


  or
  g567
  (
    n541,
    n243,
    n366,
    n299,
    n197
  );


  buf
  g568
  (
    n614,
    n480
  );


  buf
  g569
  (
    n676,
    n471
  );


  not
  g570
  (
    n632,
    n483
  );


  not
  g571
  (
    n699,
    n577
  );


  buf
  g572
  (
    n675,
    n531
  );


  buf
  g573
  (
    n666,
    n530
  );


  not
  g574
  (
    n636,
    n569
  );


  not
  g575
  (
    n628,
    n551
  );


  buf
  g576
  (
    n645,
    n524
  );


  buf
  g577
  (
    n672,
    n523
  );


  buf
  g578
  (
    n634,
    n596
  );


  not
  g579
  (
    n613,
    n595
  );


  not
  g580
  (
    n706,
    n487
  );


  buf
  g581
  (
    n629,
    n538
  );


  not
  g582
  (
    n667,
    n546
  );


  not
  g583
  (
    n647,
    n591
  );


  not
  g584
  (
    n607,
    n567
  );


  not
  g585
  (
    n609,
    n518
  );


  buf
  g586
  (
    n704,
    n495
  );


  buf
  g587
  (
    n601,
    n593
  );


  buf
  g588
  (
    n688,
    n453
  );


  buf
  g589
  (
    n610,
    n552
  );


  buf
  g590
  (
    n650,
    n579
  );


  not
  g591
  (
    n651,
    n562
  );


  not
  g592
  (
    n661,
    n535
  );


  buf
  g593
  (
    n640,
    n541
  );


  buf
  g594
  (
    n653,
    n593
  );


  buf
  g595
  (
    n631,
    n595
  );


  not
  g596
  (
    n633,
    n560
  );


  not
  g597
  (
    n641,
    n555
  );


  buf
  g598
  (
    n689,
    n527
  );


  not
  g599
  (
    n649,
    n554
  );


  not
  g600
  (
    n627,
    n546
  );


  not
  g601
  (
    n707,
    n505
  );


  buf
  g602
  (
    n696,
    n504
  );


  buf
  g603
  (
    n700,
    n600
  );


  buf
  g604
  (
    n665,
    n581
  );


  not
  g605
  (
    KeyWire_0_6,
    n597
  );


  buf
  g606
  (
    n659,
    n538
  );


  buf
  g607
  (
    n652,
    n577
  );


  buf
  g608
  (
    n695,
    n525
  );


  buf
  g609
  (
    n677,
    n581
  );


  buf
  g610
  (
    n639,
    n510
  );


  buf
  g611
  (
    n658,
    n584
  );


  not
  g612
  (
    n657,
    n594
  );


  buf
  g613
  (
    n617,
    n463
  );


  buf
  g614
  (
    n680,
    n587
  );


  not
  g615
  (
    n693,
    n502
  );


  not
  g616
  (
    n626,
    n481
  );


  buf
  g617
  (
    n606,
    n456
  );


  not
  g618
  (
    n608,
    n490
  );


  buf
  g619
  (
    n669,
    n455
  );


  buf
  g620
  (
    n654,
    n573
  );


  not
  g621
  (
    n690,
    n469
  );


  buf
  g622
  (
    n674,
    n528
  );


  not
  g623
  (
    n604,
    n568
  );


  not
  g624
  (
    n670,
    n559
  );


  buf
  g625
  (
    n687,
    n493
  );


  not
  g626
  (
    n681,
    n494
  );


  not
  g627
  (
    n698,
    n470
  );


  not
  g628
  (
    n630,
    n547
  );


  buf
  g629
  (
    n637,
    n497
  );


  buf
  g630
  (
    n644,
    n592
  );


  buf
  g631
  (
    n621,
    n457
  );


  buf
  g632
  (
    n703,
    n565
  );


  not
  g633
  (
    n622,
    n539
  );


  buf
  g634
  (
    n663,
    n503
  );


  not
  g635
  (
    n664,
    n561
  );


  not
  g636
  (
    n710,
    n534
  );


  buf
  g637
  (
    n643,
    n492
  );


  not
  g638
  (
    n602,
    n553
  );


  nor
  g639
  (
    n697,
    n563,
    n576,
    n543,
    n552
  );


  xor
  g640
  (
    n611,
    n536,
    n600,
    n526,
    n554
  );


  xnor
  g641
  (
    n625,
    n501,
    n446,
    n474,
    n589
  );


  or
  g642
  (
    n702,
    n567,
    n450,
    n566,
    n475
  );


  nand
  g643
  (
    n655,
    n516,
    n467,
    n485,
    n568
  );


  nor
  g644
  (
    n671,
    n536,
    n520,
    n556,
    n569
  );


  and
  g645
  (
    n684,
    n539,
    n541,
    n461,
    n599
  );


  and
  g646
  (
    n692,
    n570,
    n556,
    n550,
    n540
  );


  or
  g647
  (
    n642,
    n584,
    n543,
    n557,
    n445
  );


  nor
  g648
  (
    n708,
    n589,
    n573,
    n590,
    n558
  );


  nor
  g649
  (
    n660,
    n496,
    n508,
    n553,
    n537
  );


  nor
  g650
  (
    n662,
    n563,
    n564,
    n557,
    n521
  );


  or
  g651
  (
    n678,
    n533,
    n571,
    n580,
    n489
  );


  xor
  g652
  (
    n615,
    n533,
    n507,
    n544,
    n560
  );


  nor
  g653
  (
    n605,
    n500,
    n572,
    n545,
    n486
  );


  or
  g654
  (
    n682,
    n462,
    n562,
    n561,
    n513
  );


  or
  g655
  (
    n668,
    n534,
    n515,
    n590,
    n537
  );


  nor
  g656
  (
    n691,
    n473,
    n449,
    n558,
    n571
  );


  xnor
  g657
  (
    KeyWire_0_8,
    n594,
    n522,
    n548,
    n596
  );


  and
  g658
  (
    n686,
    n532,
    n578,
    n452,
    n545
  );


  nor
  g659
  (
    n701,
    n597,
    n551,
    n570,
    n565
  );


  or
  g660
  (
    n673,
    n509,
    n465,
    n459,
    n550
  );


  nor
  g661
  (
    n618,
    n466,
    n519,
    n476,
    n511
  );


  nor
  g662
  (
    n635,
    n512,
    n542,
    n598,
    n549
  );


  and
  g663
  (
    n603,
    n529,
    n588,
    n506,
    n464
  );


  or
  g664
  (
    n612,
    n586,
    n532,
    n591,
    n542
  );


  or
  g665
  (
    n679,
    n599,
    n549,
    n488,
    n448
  );


  xnor
  g666
  (
    n624,
    n559,
    n451,
    n530,
    n454
  );


  xor
  g667
  (
    n620,
    n572,
    n583,
    n544,
    n535
  );


  or
  g668
  (
    n694,
    n479,
    n585,
    n499,
    n468
  );


  nand
  g669
  (
    n646,
    n578,
    n472,
    n547,
    n484
  );


  xnor
  g670
  (
    n619,
    n566,
    n548,
    n517,
    n498
  );


  or
  g671
  (
    n709,
    n586,
    n585,
    n582,
    n477
  );


  or
  g672
  (
    n623,
    n576,
    n575,
    n540,
    n580
  );


  and
  g673
  (
    n638,
    n514,
    n579,
    n598,
    n575
  );


  and
  g674
  (
    n656,
    n460,
    n583,
    n491,
    n478
  );


  or
  g675
  (
    n683,
    n587,
    n588,
    n458,
    n555
  );


  or
  g676
  (
    n705,
    n582,
    n592,
    n574
  );


  and
  g677
  (
    n685,
    n564,
    n482,
    n447,
    n531
  );


  xnor
  g678
  (
    n714,
    n613,
    n603,
    n610
  );


  xnor
  g679
  (
    n717,
    n616,
    n604,
    n607,
    n615
  );


  xnor
  g680
  (
    n715,
    n606,
    n613,
    n614,
    n608
  );


  xnor
  g681
  (
    n712,
    n617,
    n605,
    n613,
    n611
  );


  nor
  g682
  (
    n716,
    n607,
    n612,
    n615,
    n602
  );


  xnor
  g683
  (
    n719,
    n603,
    n609,
    n605,
    n615
  );


  or
  g684
  (
    n711,
    n602,
    n616,
    n612,
    n608
  );


  nand
  g685
  (
    n718,
    n602,
    n610,
    n604,
    n616
  );


  xnor
  g686
  (
    KeyWire_0_7,
    n608,
    n611,
    n605,
    n609
  );


  nand
  g687
  (
    n713,
    n614,
    n606,
    n601,
    n611
  );


  or
  g688
  (
    n722,
    n610,
    n614,
    n609,
    n601
  );


  xor
  g689
  (
    n721,
    n612,
    n606,
    n607,
    n604
  );


  not
  g690
  (
    n743,
    n716
  );


  buf
  g691
  (
    n734,
    n716
  );


  not
  g692
  (
    n730,
    n711
  );


  not
  g693
  (
    n744,
    n714
  );


  not
  g694
  (
    n729,
    n713
  );


  not
  g695
  (
    n732,
    n719
  );


  not
  g696
  (
    n727,
    n712
  );


  not
  g697
  (
    n731,
    n717
  );


  buf
  g698
  (
    n723,
    n713
  );


  not
  g699
  (
    n726,
    n715
  );


  not
  g700
  (
    n725,
    n717
  );


  not
  g701
  (
    n735,
    n711
  );


  not
  g702
  (
    n738,
    n718
  );


  not
  g703
  (
    n737,
    n715
  );


  buf
  g704
  (
    n733,
    n714
  );


  buf
  g705
  (
    n742,
    n718
  );


  not
  g706
  (
    n728,
    n714
  );


  buf
  g707
  (
    n736,
    n716
  );


  not
  g708
  (
    n741,
    n712
  );


  not
  g709
  (
    n724,
    n718
  );


  buf
  g710
  (
    n739,
    n715
  );


  buf
  g711
  (
    n740,
    n717
  );


  xnor
  g712
  (
    n794,
    n742,
    n645,
    n681,
    n740
  );


  or
  g713
  (
    n797,
    n631,
    n653,
    n744,
    n618
  );


  or
  g714
  (
    n771,
    n650,
    n741,
    n623,
    n672
  );


  nor
  g715
  (
    n747,
    n738,
    n734,
    n742,
    n732
  );


  xnor
  g716
  (
    n792,
    n634,
    n739,
    n665,
    n740
  );


  xor
  g717
  (
    n767,
    n743,
    n636,
    n682,
    n639
  );


  xor
  g718
  (
    n803,
    n737,
    n740,
    n617,
    n666
  );


  and
  g719
  (
    n785,
    n644,
    n648,
    n637,
    n732
  );


  nor
  g720
  (
    n796,
    n743,
    n653,
    n644,
    n737
  );


  nand
  g721
  (
    n802,
    n670,
    n739,
    n654,
    n678
  );


  xor
  g722
  (
    n759,
    n677,
    n618,
    n647,
    n739
  );


  nor
  g723
  (
    n775,
    n678,
    n641,
    n728,
    n741
  );


  xnor
  g724
  (
    n750,
    n736,
    n744,
    n652,
    n673
  );


  nand
  g725
  (
    n812,
    n729,
    n736,
    n656,
    n676
  );


  xor
  g726
  (
    n799,
    n678,
    n617,
    n649,
    n645
  );


  nand
  g727
  (
    n774,
    n653,
    n732,
    n677,
    n734
  );


  nand
  g728
  (
    n795,
    n621,
    n650,
    n676,
    n636
  );


  or
  g729
  (
    n763,
    n643,
    n657,
    n728,
    n641
  );


  nor
  g730
  (
    n784,
    n655,
    n669,
    n640,
    n635
  );


  or
  g731
  (
    n778,
    n736,
    n671,
    n723,
    n662
  );


  or
  g732
  (
    n772,
    n668,
    n724,
    n674,
    n682
  );


  nand
  g733
  (
    n814,
    n657,
    n680,
    n740,
    n682
  );


  nor
  g734
  (
    n748,
    n628,
    n621,
    n663,
    n726
  );


  nor
  g735
  (
    n761,
    n735,
    n732,
    n658,
    n662
  );


  xnor
  g736
  (
    n758,
    n619,
    n731,
    n663,
    n659
  );


  nor
  g737
  (
    n813,
    n643,
    n738,
    n648,
    n673
  );


  nor
  g738
  (
    n782,
    n658,
    n628,
    n624,
    n672
  );


  xor
  g739
  (
    n764,
    n661,
    n629,
    n664,
    n739
  );


  nor
  g740
  (
    n769,
    n625,
    n629,
    n642,
    n622
  );


  nor
  g741
  (
    n777,
    n731,
    n631,
    n671,
    n665
  );


  or
  g742
  (
    n805,
    n727,
    n624,
    n652,
    n656
  );


  or
  g743
  (
    n765,
    n730,
    n730,
    n669,
    n633
  );


  nor
  g744
  (
    n745,
    n724,
    n656,
    n735,
    n727
  );


  nand
  g745
  (
    n756,
    n622,
    n681,
    n620,
    n632
  );


  and
  g746
  (
    n789,
    n625,
    n658,
    n679,
    n743
  );


  and
  g747
  (
    n800,
    n636,
    n730,
    n742,
    n735
  );


  and
  g748
  (
    n760,
    n726,
    n651,
    n649,
    n741
  );


  xor
  g749
  (
    n753,
    n670,
    n633,
    n651,
    n664
  );


  or
  g750
  (
    n807,
    n637,
    n675,
    n627,
    n726
  );


  and
  g751
  (
    n773,
    n667,
    n647,
    n729,
    n666
  );


  xor
  g752
  (
    n801,
    n628,
    n632,
    n619,
    n625
  );


  or
  g753
  (
    n798,
    n627,
    n660,
    n725,
    n646
  );


  and
  g754
  (
    n762,
    n676,
    n669,
    n622,
    n634
  );


  nor
  g755
  (
    n776,
    n677,
    n741,
    n734,
    n727
  );


  or
  g756
  (
    n811,
    n723,
    n674,
    n635,
    n727
  );


  and
  g757
  (
    n806,
    n674,
    n627,
    n743,
    n638
  );


  and
  g758
  (
    n746,
    n733,
    n633,
    n623,
    n632
  );


  xor
  g759
  (
    n752,
    n733,
    n725,
    n728,
    n626
  );


  xnor
  g760
  (
    n770,
    n737,
    n726,
    n629,
    n725
  );


  nand
  g761
  (
    n783,
    n670,
    n665,
    n639,
    n646
  );


  or
  g762
  (
    n755,
    n634,
    n659,
    n650,
    n639
  );


  xnor
  g763
  (
    KeyWire_0_12,
    n649,
    n654,
    n624,
    n734
  );


  or
  g764
  (
    n768,
    n662,
    n642,
    n637,
    n652
  );


  or
  g765
  (
    n780,
    n663,
    n666,
    n744,
    n630
  );


  nor
  g766
  (
    n791,
    n661,
    n724,
    n644,
    n681
  );


  nand
  g767
  (
    n815,
    n630,
    n744,
    n672,
    n671
  );


  and
  g768
  (
    n790,
    n731,
    n655,
    n646,
    n647
  );


  nor
  g769
  (
    n779,
    n679,
    n648,
    n730,
    n620
  );


  xor
  g770
  (
    n804,
    n651,
    n724,
    n728,
    n638
  );


  nor
  g771
  (
    n793,
    n619,
    n738,
    n668,
    n729
  );


  nor
  g772
  (
    n781,
    n630,
    n725,
    n723,
    n742
  );


  xnor
  g773
  (
    n749,
    n731,
    n660,
    n621,
    n733
  );


  and
  g774
  (
    n754,
    n675,
    n664,
    n680,
    n642
  );


  and
  g775
  (
    n810,
    n655,
    n626,
    n640,
    n673
  );


  xor
  g776
  (
    n788,
    n631,
    n679,
    n729,
    n657
  );


  nor
  g777
  (
    n809,
    n661,
    n626,
    n640,
    n735
  );


  and
  g778
  (
    n751,
    n638,
    n618,
    n680,
    n635
  );


  xor
  g779
  (
    n787,
    n623,
    n620,
    n737,
    n641
  );


  nor
  g780
  (
    n757,
    n645,
    n667,
    n675
  );


  xor
  g781
  (
    n808,
    n659,
    n733,
    n654,
    n660
  );


  xnor
  g782
  (
    n786,
    n738,
    n668,
    n736,
    n643
  );


  nor
  g783
  (
    n823,
    n756,
    n748,
    n754,
    n745
  );


  nor
  g784
  (
    n827,
    n757,
    n769,
    n760,
    n755
  );


  xor
  g785
  (
    n820,
    n752,
    n775,
    n782,
    n767
  );


  xor
  g786
  (
    n832,
    n766,
    n768,
    n767,
    n751
  );


  or
  g787
  (
    n825,
    n776,
    n780,
    n781,
    n750
  );


  nand
  g788
  (
    n828,
    n779,
    n753,
    n764,
    n777
  );


  nand
  g789
  (
    n836,
    n758,
    n759,
    n753,
    n765
  );


  and
  g790
  (
    n824,
    n773,
    n785,
    n745,
    n757
  );


  or
  g791
  (
    n826,
    n754,
    n784,
    n749,
    n772
  );


  xor
  g792
  (
    n822,
    n786,
    n747,
    n780,
    n768
  );


  and
  g793
  (
    n821,
    n765,
    n762,
    n752,
    n774
  );


  and
  g794
  (
    n817,
    n770,
    n784,
    n773,
    n772
  );


  nand
  g795
  (
    n829,
    n774,
    n776,
    n746,
    n781
  );


  nand
  g796
  (
    n816,
    n778,
    n783,
    n777,
    n747
  );


  or
  g797
  (
    n834,
    n785,
    n760,
    n763,
    n746
  );


  nand
  g798
  (
    n819,
    n761,
    n759,
    n770,
    n766
  );


  or
  g799
  (
    n830,
    n786,
    n762,
    n756,
    n771
  );


  or
  g800
  (
    n831,
    n778,
    n750,
    n764,
    n763
  );


  nor
  g801
  (
    n835,
    n783,
    n761,
    n771,
    n751
  );


  xnor
  g802
  (
    n818,
    n782,
    n748,
    n769,
    n755
  );


  or
  g803
  (
    n833,
    n758,
    n779,
    n749,
    n775
  );


  xnor
  g804
  (
    n873,
    n816,
    n400
  );


  xnor
  g805
  (
    n862,
    n404,
    n835,
    n428,
    n414
  );


  nor
  g806
  (
    n851,
    n685,
    n685,
    n823,
    n427
  );


  and
  g807
  (
    n855,
    n424,
    n833,
    n421
  );


  xor
  g808
  (
    n848,
    n401,
    n422,
    n410,
    n423
  );


  nand
  g809
  (
    n857,
    n410,
    n683,
    n828,
    n418
  );


  nor
  g810
  (
    n838,
    n684,
    n402,
    n686,
    n407
  );


  xnor
  g811
  (
    n868,
    n427,
    n421,
    n823,
    n831
  );


  and
  g812
  (
    n866,
    n400,
    n406,
    n420,
    n403
  );


  nand
  g813
  (
    n842,
    n818,
    n415,
    n422,
    n408
  );


  and
  g814
  (
    n846,
    n420,
    n820,
    n422,
    n426
  );


  nand
  g815
  (
    n852,
    n820,
    n401,
    n417,
    n834
  );


  nor
  g816
  (
    n840,
    n399,
    n412,
    n418,
    n684
  );


  nor
  g817
  (
    n860,
    n414,
    n416,
    n817
  );


  nand
  g818
  (
    n853,
    n836,
    n822,
    n404,
    n423
  );


  xnor
  g819
  (
    n856,
    n419,
    n399,
    n428,
    n827
  );


  nand
  g820
  (
    n861,
    n411,
    n819,
    n818,
    n821
  );


  or
  g821
  (
    n871,
    n825,
    n398,
    n417,
    n420
  );


  or
  g822
  (
    n847,
    n414,
    n426,
    n835,
    n824
  );


  xnor
  g823
  (
    n843,
    n409,
    n819,
    n685,
    n418
  );


  xor
  g824
  (
    n849,
    n413,
    n412,
    n683,
    n408
  );


  xor
  g825
  (
    n869,
    n406,
    n424,
    n425
  );


  or
  g826
  (
    n839,
    n417,
    n826,
    n425,
    n825
  );


  nand
  g827
  (
    n864,
    n832,
    n408,
    n683,
    n403
  );


  and
  g828
  (
    n867,
    n426,
    n398,
    n830,
    n419
  );


  and
  g829
  (
    n845,
    n415,
    n416,
    n413,
    n411
  );


  and
  g830
  (
    n870,
    n427,
    n419,
    n826,
    n816
  );


  nor
  g831
  (
    n837,
    n827,
    n684,
    n829,
    n410
  );


  xor
  g832
  (
    n863,
    n404,
    n409,
    n424,
    n834
  );


  nor
  g833
  (
    n850,
    n411,
    n405,
    n829,
    n407
  );


  xor
  g834
  (
    n872,
    n406,
    n409,
    n423,
    n407
  );


  nor
  g835
  (
    n844,
    n831,
    n399,
    n415,
    n402
  );


  xor
  g836
  (
    n854,
    n821,
    n817,
    n830,
    n824
  );


  and
  g837
  (
    n858,
    n828,
    n428,
    n833,
    n405
  );


  xor
  g838
  (
    n859,
    n405,
    n403,
    n402,
    n398
  );


  or
  g839
  (
    n865,
    n412,
    n413,
    n400,
    n401
  );


  nand
  g840
  (
    n841,
    n822,
    n836,
    n832,
    n429
  );


  and
  g841
  (
    n894,
    n790,
    n433,
    n795,
    n793
  );


  xnor
  g842
  (
    n899,
    n802,
    n869,
    n859,
    n812
  );


  or
  g843
  (
    n884,
    n800,
    n430,
    n796,
    n810
  );


  nand
  g844
  (
    n901,
    n795,
    n849,
    n845,
    n815
  );


  nand
  g845
  (
    n881,
    n806,
    n815,
    n804
  );


  nor
  g846
  (
    n882,
    n811,
    n686,
    n793,
    n864
  );


  and
  g847
  (
    n885,
    n852,
    n815,
    n814,
    n431
  );


  or
  g848
  (
    n900,
    n796,
    n687,
    n871,
    n798
  );


  nor
  g849
  (
    n878,
    n432,
    n690,
    n809,
    n807
  );


  nand
  g850
  (
    n886,
    n789,
    n431,
    n794,
    n867
  );


  xnor
  g851
  (
    n896,
    n813,
    n863,
    n799,
    n868
  );


  or
  g852
  (
    KeyWire_0_2,
    n792,
    n801,
    n787,
    n788
  );


  or
  g853
  (
    n892,
    n431,
    n789,
    n794,
    n791
  );


  xor
  g854
  (
    n897,
    n429,
    n851,
    n799,
    n858
  );


  xor
  g855
  (
    n877,
    n432,
    n813,
    n429,
    n688
  );


  nor
  g856
  (
    n888,
    n686,
    n687,
    n800,
    n432
  );


  or
  g857
  (
    n880,
    n870,
    n802,
    n866,
    n808
  );


  nor
  g858
  (
    n874,
    n814,
    n862,
    n801,
    n689
  );


  or
  g859
  (
    n889,
    n814,
    n854,
    n810,
    n806
  );


  nand
  g860
  (
    n879,
    n812,
    n687,
    n847,
    n853
  );


  xor
  g861
  (
    n891,
    n803,
    n811,
    n797,
    n430
  );


  nor
  g862
  (
    n898,
    n788,
    n813,
    n787,
    n846
  );


  xnor
  g863
  (
    n875,
    n808,
    n803,
    n872,
    n850
  );


  and
  g864
  (
    n895,
    n873,
    n855,
    n809,
    n688
  );


  nor
  g865
  (
    n890,
    n812,
    n805,
    n861,
    n865
  );


  xor
  g866
  (
    n887,
    n792,
    n805,
    n791,
    n798
  );


  and
  g867
  (
    n883,
    n430,
    n857,
    n811,
    n860
  );


  nor
  g868
  (
    n893,
    n807,
    n856,
    n689,
    n848
  );


  or
  g869
  (
    n902,
    n689,
    n790,
    n797,
    n688
  );


  nor
  g870
  (
    KeyWire_0_9,
    n434,
    n702,
    n691,
    n899
  );


  nand
  g871
  (
    n904,
    n696,
    n882,
    n895,
    n700
  );


  and
  g872
  (
    n916,
    n888,
    n876,
    n896,
    n900
  );


  and
  g873
  (
    n915,
    n894,
    n875,
    n892,
    n886
  );


  or
  g874
  (
    n937,
    n898,
    n891,
    n896,
    n893
  );


  xor
  g875
  (
    n938,
    n698,
    n893,
    n693,
    n894
  );


  xor
  g876
  (
    n914,
    n896,
    n695,
    n887,
    n155
  );


  or
  g877
  (
    n936,
    n898,
    n891,
    n878,
    n889
  );


  xor
  g878
  (
    n934,
    n884,
    n696,
    n435
  );


  xor
  g879
  (
    n920,
    n892,
    n891,
    n32,
    n875
  );


  and
  g880
  (
    n906,
    n691,
    n895,
    n719,
    n704
  );


  nand
  g881
  (
    n909,
    n693,
    n902,
    n880,
    n697
  );


  xor
  g882
  (
    n940,
    n900,
    n880,
    n897,
    n888
  );


  xor
  g883
  (
    n917,
    n895,
    n876,
    n890,
    n692
  );


  xnor
  g884
  (
    n913,
    n881,
    n879,
    n898,
    n874
  );


  or
  g885
  (
    n935,
    n877,
    n701,
    n899,
    n875
  );


  and
  g886
  (
    n933,
    n901,
    n882,
    n879,
    n435
  );


  xnor
  g887
  (
    n921,
    n902,
    n876,
    n698,
    n898
  );


  xnor
  g888
  (
    n942,
    n433,
    n435,
    n880,
    n702
  );


  or
  g889
  (
    n912,
    n890,
    n720,
    n703,
    n694
  );


  xor
  g890
  (
    n918,
    n878,
    n889,
    n697,
    n720
  );


  and
  g891
  (
    n910,
    n721,
    n32,
    n894,
    n701
  );


  xor
  g892
  (
    n930,
    n698,
    n889,
    n899,
    n878
  );


  xor
  g893
  (
    n926,
    n883,
    n693,
    n884,
    n720
  );


  xor
  g894
  (
    n919,
    n888,
    n702,
    n886,
    n883
  );


  or
  g895
  (
    n908,
    n881,
    n704,
    n874,
    n691
  );


  nor
  g896
  (
    n923,
    n692,
    n877,
    n884,
    n885
  );


  xor
  g897
  (
    n925,
    n900,
    n694,
    n433,
    n877
  );


  xor
  g898
  (
    n932,
    n897,
    n695,
    n700,
    n887
  );


  or
  g899
  (
    n941,
    n902,
    n719,
    n882,
    n155
  );


  nand
  g900
  (
    n905,
    n879,
    n899,
    n156,
    n874
  );


  and
  g901
  (
    KeyWire_0_13,
    n900,
    n703,
    n901,
    n885
  );


  xor
  g902
  (
    n928,
    n699,
    n902,
    n893,
    n897
  );


  or
  g903
  (
    n924,
    n700,
    n434,
    n890,
    n692
  );


  and
  g904
  (
    n929,
    n699,
    n32,
    n896,
    n721
  );


  xor
  g905
  (
    n931,
    n434,
    n901,
    n697
  );


  xor
  g906
  (
    n922,
    n721,
    n703,
    n881,
    n886
  );


  nor
  g907
  (
    n903,
    n690,
    n885,
    n699,
    n887
  );


  xnor
  g908
  (
    n939,
    n897,
    n892,
    n694,
    n883
  );


  nor
  g909
  (
    n927,
    n690,
    n701,
    n722,
    n695
  );


  xor
  g910
  (
    n962,
    n921,
    n936,
    n928,
    n934
  );


  nand
  g911
  (
    n959,
    n923,
    n938,
    n937,
    n942
  );


  nor
  g912
  (
    n952,
    n933,
    n919,
    n914,
    n930
  );


  nand
  g913
  (
    n943,
    n905,
    n922,
    n929,
    n927
  );


  and
  g914
  (
    n960,
    n941,
    n926,
    n905,
    n939
  );


  nor
  g915
  (
    n945,
    n924,
    n910,
    n937
  );


  xor
  g916
  (
    n951,
    n926,
    n934,
    n925,
    n922
  );


  nor
  g917
  (
    n967,
    n941,
    n908,
    n932
  );


  nand
  g918
  (
    n946,
    n939,
    n920,
    n942,
    n940
  );


  xor
  g919
  (
    n958,
    n923,
    n935,
    n924,
    n939
  );


  or
  g920
  (
    n957,
    n920,
    n935,
    n917,
    n922
  );


  nand
  g921
  (
    n956,
    n906,
    n912,
    n928,
    n909
  );


  xor
  g922
  (
    n949,
    n929,
    n940,
    n436
  );


  or
  g923
  (
    n964,
    n907,
    n936,
    n921,
    n931
  );


  or
  g924
  (
    n969,
    n916,
    n935,
    n934,
    n156
  );


  nand
  g925
  (
    n953,
    n912,
    n929,
    n924,
    n903
  );


  and
  g926
  (
    n961,
    n436,
    n936,
    n437,
    n909
  );


  or
  g927
  (
    n944,
    n941,
    n916,
    n906,
    n921
  );


  nor
  g928
  (
    n963,
    n914,
    n903,
    n931,
    n938
  );


  xor
  g929
  (
    n947,
    n942,
    n931,
    n913,
    n938
  );


  xor
  g930
  (
    n968,
    n911,
    n940,
    n933
  );


  xor
  g931
  (
    n966,
    n918,
    n927,
    n913,
    n926
  );


  or
  g932
  (
    n948,
    n919,
    n932,
    n911,
    n915
  );


  or
  g933
  (
    n954,
    n937,
    n923,
    n930,
    n918
  );


  nand
  g934
  (
    n965,
    n928,
    n917,
    n908,
    n925
  );


  and
  g935
  (
    n955,
    n904,
    n927,
    n907,
    n437
  );


  or
  g936
  (
    n950,
    n930,
    n904,
    n915,
    n925
  );


  not
  g937
  (
    n973,
    n959
  );


  not
  g938
  (
    n972,
    n960
  );


  buf
  g939
  (
    n976,
    n967
  );


  not
  g940
  (
    n975,
    n966
  );


  buf
  g941
  (
    n977,
    n965
  );


  buf
  g942
  (
    n970,
    n962
  );


  nand
  g943
  (
    n974,
    n964,
    n956
  );


  nand
  g944
  (
    n971,
    n961,
    n963,
    n958,
    n957
  );


  not
  g945
  (
    n978,
    n973
  );


  buf
  g946
  (
    n981,
    n976
  );


  not
  g947
  (
    n980,
    n974
  );


  not
  g948
  (
    n979,
    n975
  );


  not
  g949
  (
    n988,
    n980
  );


  buf
  g950
  (
    n985,
    n980
  );


  buf
  g951
  (
    n986,
    n978
  );


  not
  g952
  (
    n983,
    n978
  );


  buf
  g953
  (
    n984,
    n979
  );


  not
  g954
  (
    n987,
    n981
  );


  and
  g955
  (
    n982,
    n981,
    n979
  );


  buf
  g956
  (
    n993,
    n441
  );


  not
  g957
  (
    n990,
    n987
  );


  not
  g958
  (
    n991,
    n986
  );


  buf
  g959
  (
    n989,
    n438
  );


  not
  g960
  (
    n992,
    n986
  );


  buf
  g961
  (
    n1007,
    n983
  );


  buf
  g962
  (
    n996,
    n437
  );


  buf
  g963
  (
    n999,
    n982
  );


  not
  g964
  (
    n1002,
    n441
  );


  buf
  g965
  (
    n1000,
    n988
  );


  buf
  g966
  (
    n1008,
    n983
  );


  buf
  g967
  (
    n997,
    n984
  );


  not
  g968
  (
    n1005,
    n977
  );


  or
  g969
  (
    n1003,
    n438,
    n984,
    n440
  );


  nor
  g970
  (
    n998,
    n442,
    n439,
    n984,
    n982
  );


  nor
  g971
  (
    n995,
    n988,
    n441,
    n439,
    n985
  );


  xnor
  g972
  (
    n994,
    n440,
    n987,
    n985,
    n443
  );


  nand
  g973
  (
    n1004,
    n987,
    n442,
    n985,
    n988
  );


  xnor
  g974
  (
    n1001,
    n440,
    n986,
    n443,
    n438
  );


  xnor
  g975
  (
    n1006,
    n442,
    n983,
    n439,
    n443
  );


  xnor
  g976
  (
    n1015,
    n1007,
    n1000,
    n991,
    n1008
  );


  nor
  g977
  (
    n1016,
    n1006,
    n1006,
    n995,
    n969
  );


  or
  g978
  (
    n1014,
    n1001,
    n1003,
    n1004,
    n1002
  );


  and
  g979
  (
    n1013,
    n998,
    n999,
    n1005,
    n989
  );


  nor
  g980
  (
    n1009,
    n1008,
    n981,
    n994,
    n990
  );


  or
  g981
  (
    n1012,
    n1004,
    n968,
    n1002,
    n1005
  );


  nand
  g982
  (
    n1017,
    n1007,
    n997,
    n993,
    n1003
  );


  and
  g983
  (
    n1010,
    n1001,
    n998,
    n999,
    n1000
  );


  or
  g984
  (
    n1011,
    n997,
    n156,
    n992,
    n996
  );


  buf
  g985
  (
    n1019,
    n1009
  );


  not
  g986
  (
    n1018,
    n1010
  );


  xor
  g987
  (
    n1024,
    n1012,
    n1018,
    n1015
  );


  xor
  g988
  (
    n1025,
    n1011,
    n1014,
    n1019
  );


  nor
  g989
  (
    n1026,
    n1018,
    n707,
    n1010
  );


  xnor
  g990
  (
    n1021,
    n706,
    n722,
    n1018,
    n705
  );


  and
  g991
  (
    n1020,
    n706,
    n722,
    n1015,
    n1013
  );


  nor
  g992
  (
    n1023,
    n706,
    n1011,
    n1016,
    n707
  );


  and
  g993
  (
    n1022,
    n704,
    n1012,
    n705,
    n1019
  );


  nor
  g994
  (
    n1027,
    n1013,
    n1014,
    n705,
    n1019
  );


  xor
  g995
  (
    n1028,
    n709,
    n708,
    n1017
  );


  nand
  g996
  (
    n1032,
    n1024,
    n444,
    n1025,
    n1016
  );


  or
  g997
  (
    n1030,
    n710,
    n1027,
    n709,
    n1017
  );


  xnor
  g998
  (
    n1031,
    n1023,
    n444,
    n1026
  );


  or
  g999
  (
    n1029,
    n708,
    n709,
    n710
  );


  xor
  KeyGate_0_0
  (
    n235,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n413,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n876,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n202,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n531,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n596,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n616,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n720,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n648,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n907,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n212,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n313,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n766,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n911,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n351,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n49,
    KeyNOTWire_0_15
  );


endmodule

