

module Stat_786_1023
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n807,
  n799,
  n801,
  n809,
  n811,
  n797,
  n813,
  n800,
  n796,
  n805,
  n806,
  n812,
  n804,
  n802,
  n808,
  n810,
  n803,
  n798
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n807;output n799;output n801;output n809;output n811;output n797;output n813;output n800;output n796;output n805;output n806;output n812;output n804;output n802;output n808;output n810;output n803;output n798;
  wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  not
  g0
  (
    n56,
    n9
  );


  not
  g1
  (
    n74,
    n11
  );


  not
  g2
  (
    n89,
    n13
  );


  not
  g3
  (
    n102,
    n13
  );


  buf
  g4
  (
    n93,
    n2
  );


  buf
  g5
  (
    n47,
    n10
  );


  buf
  g6
  (
    n126,
    n24
  );


  buf
  g7
  (
    n67,
    n13
  );


  not
  g8
  (
    n101,
    n18
  );


  buf
  g9
  (
    n120,
    n12
  );


  buf
  g10
  (
    n62,
    n20
  );


  buf
  g11
  (
    n52,
    n24
  );


  buf
  g12
  (
    n61,
    n25
  );


  not
  g13
  (
    n91,
    n1
  );


  buf
  g14
  (
    n68,
    n23
  );


  buf
  g15
  (
    n64,
    n14
  );


  buf
  g16
  (
    n42,
    n11
  );


  not
  g17
  (
    n78,
    n15
  );


  buf
  g18
  (
    n96,
    n4
  );


  not
  g19
  (
    n48,
    n20
  );


  not
  g20
  (
    n29,
    n16
  );


  not
  g21
  (
    n123,
    n24
  );


  buf
  g22
  (
    n109,
    n2
  );


  buf
  g23
  (
    n79,
    n18
  );


  buf
  g24
  (
    n41,
    n19
  );


  not
  g25
  (
    n57,
    n12
  );


  buf
  g26
  (
    n46,
    n17
  );


  not
  g27
  (
    n75,
    n12
  );


  not
  g28
  (
    n28,
    n9
  );


  not
  g29
  (
    n50,
    n16
  );


  buf
  g30
  (
    KeyWire_0_48,
    n3
  );


  buf
  g31
  (
    n94,
    n21
  );


  not
  g32
  (
    n100,
    n7
  );


  not
  g33
  (
    n39,
    n25
  );


  buf
  g34
  (
    n105,
    n15
  );


  not
  g35
  (
    n113,
    n13
  );


  not
  g36
  (
    n119,
    n21
  );


  not
  g37
  (
    n124,
    n25
  );


  not
  g38
  (
    KeyWire_0_12,
    n8
  );


  buf
  g39
  (
    n36,
    n7
  );


  not
  g40
  (
    n122,
    n8
  );


  not
  g41
  (
    n81,
    n19
  );


  not
  g42
  (
    n65,
    n1
  );


  buf
  g43
  (
    KeyWire_0_11,
    n18
  );


  buf
  g44
  (
    n92,
    n7
  );


  buf
  g45
  (
    n58,
    n10
  );


  buf
  g46
  (
    n35,
    n17
  );


  not
  g47
  (
    KeyWire_0_30,
    n23
  );


  not
  g48
  (
    n107,
    n3
  );


  buf
  g49
  (
    n103,
    n20
  );


  not
  g50
  (
    n71,
    n4
  );


  buf
  g51
  (
    n70,
    n10
  );


  buf
  g52
  (
    KeyWire_0_6,
    n4
  );


  not
  g53
  (
    n90,
    n21
  );


  not
  g54
  (
    n125,
    n1
  );


  buf
  g55
  (
    n106,
    n22
  );


  not
  g56
  (
    n33,
    n10
  );


  not
  g57
  (
    n77,
    n14
  );


  not
  g58
  (
    n45,
    n6
  );


  buf
  g59
  (
    n121,
    n1
  );


  not
  g60
  (
    n82,
    n17
  );


  not
  g61
  (
    n73,
    n23
  );


  buf
  g62
  (
    n87,
    n15
  );


  not
  g63
  (
    n110,
    n16
  );


  not
  g64
  (
    n98,
    n9
  );


  buf
  g65
  (
    n31,
    n8
  );


  not
  g66
  (
    n32,
    n3
  );


  not
  g67
  (
    n95,
    n14
  );


  buf
  g68
  (
    n69,
    n24
  );


  buf
  g69
  (
    n111,
    n23
  );


  not
  g70
  (
    n84,
    n22
  );


  buf
  g71
  (
    n117,
    n8
  );


  not
  g72
  (
    n85,
    n6
  );


  not
  g73
  (
    n115,
    n11
  );


  not
  g74
  (
    n88,
    n19
  );


  not
  g75
  (
    n97,
    n2
  );


  not
  g76
  (
    n60,
    n19
  );


  not
  g77
  (
    n108,
    n17
  );


  buf
  g78
  (
    n34,
    n5
  );


  buf
  g79
  (
    KeyWire_0_40,
    n6
  );


  buf
  g80
  (
    n38,
    n2
  );


  buf
  g81
  (
    n118,
    n22
  );


  not
  g82
  (
    KeyWire_0_47,
    n5
  );


  not
  g83
  (
    n104,
    n22
  );


  not
  g84
  (
    KeyWire_0_50,
    n4
  );


  not
  g85
  (
    n59,
    n7
  );


  buf
  g86
  (
    n63,
    n21
  );


  not
  g87
  (
    n40,
    n5
  );


  buf
  g88
  (
    n43,
    n12
  );


  buf
  g89
  (
    n66,
    n6
  );


  buf
  g90
  (
    n54,
    n18
  );


  not
  g91
  (
    n114,
    n14
  );


  not
  g92
  (
    n83,
    n15
  );


  not
  g93
  (
    n51,
    n3
  );


  buf
  g94
  (
    n37,
    n5
  );


  buf
  g95
  (
    n53,
    n20
  );


  buf
  g96
  (
    n86,
    n11
  );


  not
  g97
  (
    n44,
    n16
  );


  buf
  g98
  (
    n99,
    n9
  );


  not
  g99
  (
    n340,
    n81
  );


  not
  g100
  (
    n153,
    n66
  );


  not
  g101
  (
    n211,
    n61
  );


  not
  g102
  (
    KeyWire_0_52,
    n28
  );


  not
  g103
  (
    n140,
    n65
  );


  not
  g104
  (
    n166,
    n36
  );


  not
  g105
  (
    n315,
    n79
  );


  not
  g106
  (
    KeyWire_0_44,
    n76
  );


  buf
  g107
  (
    n306,
    n49
  );


  buf
  g108
  (
    n348,
    n36
  );


  not
  g109
  (
    n148,
    n68
  );


  not
  g110
  (
    n197,
    n64
  );


  not
  g111
  (
    n238,
    n84
  );


  buf
  g112
  (
    n325,
    n80
  );


  buf
  g113
  (
    n225,
    n73
  );


  buf
  g114
  (
    n203,
    n51
  );


  not
  g115
  (
    n233,
    n66
  );


  buf
  g116
  (
    n175,
    n29
  );


  buf
  g117
  (
    n324,
    n40
  );


  not
  g118
  (
    n156,
    n61
  );


  not
  g119
  (
    n209,
    n33
  );


  buf
  g120
  (
    n162,
    n70
  );


  buf
  g121
  (
    n163,
    n38
  );


  not
  g122
  (
    n249,
    n46
  );


  not
  g123
  (
    n292,
    n49
  );


  buf
  g124
  (
    n307,
    n44
  );


  buf
  g125
  (
    n174,
    n35
  );


  not
  g126
  (
    n178,
    n55
  );


  not
  g127
  (
    n154,
    n51
  );


  not
  g128
  (
    n239,
    n43
  );


  not
  g129
  (
    n221,
    n82
  );


  not
  g130
  (
    n206,
    n46
  );


  not
  g131
  (
    n346,
    n81
  );


  buf
  g132
  (
    n226,
    n61
  );


  buf
  g133
  (
    n349,
    n61
  );


  buf
  g134
  (
    n339,
    n60
  );


  not
  g135
  (
    n223,
    n44
  );


  buf
  g136
  (
    n183,
    n41
  );


  buf
  g137
  (
    n286,
    n75
  );


  buf
  g138
  (
    n257,
    n64
  );


  not
  g139
  (
    n334,
    n83
  );


  not
  g140
  (
    n289,
    n47
  );


  not
  g141
  (
    n318,
    n29
  );


  not
  g142
  (
    n130,
    n76
  );


  buf
  g143
  (
    n181,
    n70
  );


  buf
  g144
  (
    n290,
    n39
  );


  not
  g145
  (
    n227,
    n68
  );


  buf
  g146
  (
    n259,
    n38
  );


  buf
  g147
  (
    n232,
    n71
  );


  not
  g148
  (
    n144,
    n60
  );


  buf
  g149
  (
    n260,
    n34
  );


  not
  g150
  (
    n247,
    n37
  );


  buf
  g151
  (
    n344,
    n74
  );


  buf
  g152
  (
    n273,
    n53
  );


  not
  g153
  (
    n228,
    n68
  );


  buf
  g154
  (
    n245,
    n71
  );


  buf
  g155
  (
    n316,
    n77
  );


  buf
  g156
  (
    n244,
    n32
  );


  buf
  g157
  (
    n293,
    n69
  );


  not
  g158
  (
    n200,
    n54
  );


  not
  g159
  (
    n214,
    n69
  );


  buf
  g160
  (
    n150,
    n67
  );


  buf
  g161
  (
    n215,
    n51
  );


  not
  g162
  (
    n288,
    n77
  );


  buf
  g163
  (
    n275,
    n58
  );


  not
  g164
  (
    n177,
    n37
  );


  not
  g165
  (
    n345,
    n72
  );


  buf
  g166
  (
    n182,
    n34
  );


  buf
  g167
  (
    n313,
    n42
  );


  buf
  g168
  (
    KeyWire_0_25,
    n42
  );


  buf
  g169
  (
    n171,
    n55
  );


  not
  g170
  (
    n164,
    n77
  );


  not
  g171
  (
    n243,
    n67
  );


  not
  g172
  (
    KeyWire_0_21,
    n53
  );


  not
  g173
  (
    n139,
    n49
  );


  not
  g174
  (
    n263,
    n51
  );


  buf
  g175
  (
    n237,
    n76
  );


  not
  g176
  (
    n173,
    n60
  );


  not
  g177
  (
    n220,
    n34
  );


  buf
  g178
  (
    n311,
    n71
  );


  buf
  g179
  (
    KeyWire_0_41,
    n31
  );


  not
  g180
  (
    n354,
    n31
  );


  buf
  g181
  (
    KeyWire_0_15,
    n54
  );


  not
  g182
  (
    n287,
    n40
  );


  buf
  g183
  (
    n199,
    n80
  );


  buf
  g184
  (
    KeyWire_0_14,
    n59
  );


  buf
  g185
  (
    n256,
    n82
  );


  not
  g186
  (
    n276,
    n34
  );


  buf
  g187
  (
    n242,
    n69
  );


  buf
  g188
  (
    n176,
    n68
  );


  buf
  g189
  (
    n132,
    n75
  );


  not
  g190
  (
    n133,
    n65
  );


  buf
  g191
  (
    n342,
    n79
  );


  buf
  g192
  (
    n246,
    n54
  );


  buf
  g193
  (
    n184,
    n57
  );


  not
  g194
  (
    n157,
    n45
  );


  buf
  g195
  (
    KeyWire_0_26,
    n78
  );


  not
  g196
  (
    n278,
    n62
  );


  buf
  g197
  (
    n187,
    n45
  );


  not
  g198
  (
    n323,
    n43
  );


  not
  g199
  (
    KeyWire_0_62,
    n70
  );


  not
  g200
  (
    n169,
    n53
  );


  not
  g201
  (
    n317,
    n77
  );


  not
  g202
  (
    KeyWire_0_33,
    n28
  );


  buf
  g203
  (
    n322,
    n52
  );


  not
  g204
  (
    n250,
    n56
  );


  buf
  g205
  (
    n294,
    n80
  );


  not
  g206
  (
    n265,
    n33
  );


  buf
  g207
  (
    n192,
    n50
  );


  not
  g208
  (
    n219,
    n83
  );


  not
  g209
  (
    n191,
    n32
  );


  buf
  g210
  (
    n303,
    n57
  );


  buf
  g211
  (
    n305,
    n73
  );


  buf
  g212
  (
    n321,
    n47
  );


  not
  g213
  (
    n285,
    n41
  );


  not
  g214
  (
    n161,
    n74
  );


  buf
  g215
  (
    n281,
    n48
  );


  buf
  g216
  (
    n198,
    n47
  );


  buf
  g217
  (
    n134,
    n70
  );


  buf
  g218
  (
    n146,
    n62
  );


  buf
  g219
  (
    n296,
    n81
  );


  not
  g220
  (
    n241,
    n35
  );


  buf
  g221
  (
    n205,
    n33
  );


  not
  g222
  (
    n135,
    n59
  );


  not
  g223
  (
    n196,
    n56
  );


  not
  g224
  (
    n301,
    n47
  );


  not
  g225
  (
    n230,
    n54
  );


  not
  g226
  (
    n272,
    n78
  );


  buf
  g227
  (
    n213,
    n69
  );


  not
  g228
  (
    n353,
    n71
  );


  buf
  g229
  (
    n299,
    n72
  );


  buf
  g230
  (
    n319,
    n28
  );


  buf
  g231
  (
    n335,
    n40
  );


  buf
  g232
  (
    n158,
    n72
  );


  not
  g233
  (
    KeyWire_0_28,
    n48
  );


  buf
  g234
  (
    n222,
    n59
  );


  buf
  g235
  (
    n179,
    n37
  );


  not
  g236
  (
    n218,
    n50
  );


  not
  g237
  (
    n308,
    n57
  );


  buf
  g238
  (
    n152,
    n42
  );


  not
  g239
  (
    n337,
    n84
  );


  buf
  g240
  (
    n267,
    n42
  );


  not
  g241
  (
    n145,
    n37
  );


  buf
  g242
  (
    KeyWire_0_13,
    n76
  );


  not
  g243
  (
    n168,
    n73
  );


  not
  g244
  (
    n160,
    n84
  );


  not
  g245
  (
    n347,
    n31
  );


  not
  g246
  (
    KeyWire_0_45,
    n67
  );


  not
  g247
  (
    KeyWire_0_31,
    n30
  );


  not
  g248
  (
    n327,
    n63
  );


  not
  g249
  (
    n341,
    n40
  );


  buf
  g250
  (
    n258,
    n46
  );


  buf
  g251
  (
    n338,
    n43
  );


  not
  g252
  (
    n304,
    n38
  );


  not
  g253
  (
    n279,
    n33
  );


  not
  g254
  (
    n210,
    n74
  );


  not
  g255
  (
    n149,
    n65
  );


  buf
  g256
  (
    n255,
    n60
  );


  not
  g257
  (
    n131,
    n72
  );


  not
  g258
  (
    n207,
    n39
  );


  not
  g259
  (
    KeyWire_0_49,
    n29
  );


  not
  g260
  (
    n235,
    n53
  );


  buf
  g261
  (
    n180,
    n81
  );


  not
  g262
  (
    n329,
    n56
  );


  not
  g263
  (
    n234,
    n41
  );


  not
  g264
  (
    n282,
    n55
  );


  buf
  g265
  (
    n332,
    n82
  );


  buf
  g266
  (
    n253,
    n82
  );


  not
  g267
  (
    KeyWire_0_39,
    n80
  );


  buf
  g268
  (
    n283,
    n44
  );


  not
  g269
  (
    n350,
    n67
  );


  buf
  g270
  (
    n224,
    n52
  );


  buf
  g271
  (
    n127,
    n78
  );


  buf
  g272
  (
    n284,
    n64
  );


  not
  g273
  (
    n298,
    n32
  );


  buf
  g274
  (
    n254,
    n65
  );


  not
  g275
  (
    n185,
    n30
  );


  not
  g276
  (
    n136,
    n31
  );


  buf
  g277
  (
    n231,
    n66
  );


  not
  g278
  (
    n252,
    n83
  );


  buf
  g279
  (
    n295,
    n73
  );


  not
  g280
  (
    n195,
    n49
  );


  buf
  g281
  (
    n188,
    n35
  );


  buf
  g282
  (
    KeyWire_0_3,
    n43
  );


  not
  g283
  (
    n212,
    n39
  );


  buf
  g284
  (
    n343,
    n75
  );


  not
  g285
  (
    n248,
    n79
  );


  buf
  g286
  (
    n167,
    n59
  );


  not
  g287
  (
    n142,
    n74
  );


  not
  g288
  (
    KeyWire_0_61,
    n36
  );


  not
  g289
  (
    n236,
    n50
  );


  not
  g290
  (
    n217,
    n83
  );


  not
  g291
  (
    n309,
    n30
  );


  buf
  g292
  (
    n328,
    n78
  );


  not
  g293
  (
    n297,
    n35
  );


  buf
  g294
  (
    KeyWire_0_16,
    n39
  );


  buf
  g295
  (
    n194,
    n66
  );


  buf
  g296
  (
    n314,
    n36
  );


  buf
  g297
  (
    n159,
    n48
  );


  not
  g298
  (
    n270,
    n63
  );


  not
  g299
  (
    n170,
    n63
  );


  not
  g300
  (
    n138,
    n84
  );


  buf
  g301
  (
    n189,
    n45
  );


  not
  g302
  (
    n302,
    n41
  );


  not
  g303
  (
    n208,
    n56
  );


  not
  g304
  (
    n193,
    n58
  );


  not
  g305
  (
    n352,
    n62
  );


  buf
  g306
  (
    n312,
    n28
  );


  buf
  g307
  (
    n277,
    n48
  );


  buf
  g308
  (
    n251,
    n75
  );


  not
  g309
  (
    n268,
    n52
  );


  buf
  g310
  (
    n274,
    n79
  );


  not
  g311
  (
    n271,
    n45
  );


  not
  g312
  (
    n216,
    n30
  );


  buf
  g313
  (
    n165,
    n52
  );


  not
  g314
  (
    n143,
    n29
  );


  not
  g315
  (
    n240,
    n55
  );


  buf
  g316
  (
    n326,
    n58
  );


  buf
  g317
  (
    n320,
    n38
  );


  buf
  g318
  (
    n351,
    n44
  );


  buf
  g319
  (
    KeyWire_0_24,
    n64
  );


  buf
  g320
  (
    n262,
    n32
  );


  buf
  g321
  (
    n147,
    n62
  );


  not
  g322
  (
    n280,
    n63
  );


  buf
  g323
  (
    n172,
    n57
  );


  buf
  g324
  (
    n333,
    n58
  );


  not
  g325
  (
    n137,
    n50
  );


  not
  g326
  (
    n310,
    n46
  );


  not
  g327
  (
    n361,
    n146
  );


  buf
  g328
  (
    n377,
    n133
  );


  not
  g329
  (
    KeyWire_0_51,
    n135
  );


  not
  g330
  (
    n372,
    n145
  );


  not
  g331
  (
    n358,
    n127
  );


  buf
  g332
  (
    n363,
    n131
  );


  not
  g333
  (
    n365,
    n130
  );


  not
  g334
  (
    n364,
    n138
  );


  buf
  g335
  (
    n378,
    n142
  );


  not
  g336
  (
    n373,
    n129
  );


  buf
  g337
  (
    KeyWire_0_58,
    n136
  );


  buf
  g338
  (
    n375,
    n143
  );


  buf
  g339
  (
    KeyWire_0_22,
    n141
  );


  not
  g340
  (
    n371,
    n151
  );


  not
  g341
  (
    n374,
    n148
  );


  not
  g342
  (
    n369,
    n150
  );


  buf
  g343
  (
    n360,
    n149
  );


  buf
  g344
  (
    n379,
    n137
  );


  buf
  g345
  (
    n376,
    n152
  );


  not
  g346
  (
    n359,
    n147
  );


  not
  g347
  (
    n366,
    n134
  );


  not
  g348
  (
    n362,
    n144
  );


  buf
  g349
  (
    n357,
    n132
  );


  buf
  g350
  (
    n356,
    n128
  );


  not
  g351
  (
    n368,
    n140
  );


  not
  g352
  (
    KeyWire_0_18,
    n139
  );


  xnor
  g353
  (
    n427,
    n223,
    n241,
    n224,
    n173
  );


  or
  g354
  (
    n466,
    n361,
    n379,
    n374,
    n253
  );


  xnor
  g355
  (
    n454,
    n181,
    n356,
    n232,
    n168
  );


  xnor
  g356
  (
    n395,
    n206,
    n257,
    n367,
    n247
  );


  xor
  g357
  (
    n477,
    n221,
    n260,
    n193,
    n377
  );


  xnor
  g358
  (
    n385,
    n367,
    n254,
    n192,
    n205
  );


  or
  g359
  (
    n431,
    n230,
    n254,
    n365,
    n241
  );


  and
  g360
  (
    n425,
    n375,
    n162,
    n371,
    n182
  );


  or
  g361
  (
    n401,
    n201,
    n198,
    n256,
    n185
  );


  xnor
  g362
  (
    n390,
    n250,
    n376,
    n211,
    n160
  );


  xnor
  g363
  (
    n475,
    n218,
    n246,
    n224,
    n155
  );


  or
  g364
  (
    n430,
    n248,
    n229,
    n176,
    n223
  );


  xor
  g365
  (
    n406,
    n170,
    n360,
    n233,
    n176
  );


  and
  g366
  (
    KeyWire_0_60,
    n257,
    n364,
    n362,
    n157
  );


  nand
  g367
  (
    n472,
    n368,
    n358,
    n205,
    n202
  );


  xor
  g368
  (
    n479,
    n371,
    n190,
    n239,
    n153
  );


  xnor
  g369
  (
    n415,
    n222,
    n363,
    n183,
    n237
  );


  xor
  g370
  (
    n404,
    n251,
    n196,
    n226
  );


  xnor
  g371
  (
    n419,
    n204,
    n197,
    n164,
    n364
  );


  nor
  g372
  (
    n394,
    n251,
    n219,
    n261,
    n255
  );


  and
  g373
  (
    n468,
    n247,
    n235,
    n361,
    n369
  );


  or
  g374
  (
    n460,
    n212,
    n373,
    n232,
    n368
  );


  and
  g375
  (
    n450,
    n207,
    n218,
    n165,
    n256
  );


  or
  g376
  (
    KeyWire_0_36,
    n363,
    n240,
    n212,
    n195
  );


  nor
  g377
  (
    n384,
    n214,
    n194,
    n243,
    n366
  );


  xor
  g378
  (
    n478,
    n225,
    n231,
    n248,
    n154
  );


  xnor
  g379
  (
    n422,
    n204,
    n244,
    n245,
    n225
  );


  xor
  g380
  (
    n398,
    n367,
    n247,
    n187,
    n375
  );


  or
  g381
  (
    n474,
    n374,
    n227,
    n192,
    n379
  );


  xor
  g382
  (
    n391,
    n189,
    n213,
    n255,
    n235
  );


  nor
  g383
  (
    n418,
    n191,
    n214,
    n178,
    n355
  );


  xor
  g384
  (
    n435,
    n183,
    n214,
    n374,
    n217
  );


  xor
  g385
  (
    n464,
    n190,
    n366,
    n174,
    n178
  );


  and
  g386
  (
    n446,
    n229,
    n193,
    n228,
    n360
  );


  xnor
  g387
  (
    n423,
    n216,
    n378,
    n246,
    n225
  );


  xnor
  g388
  (
    n480,
    n236,
    n184,
    n165
  );


  nand
  g389
  (
    n449,
    n215,
    n164,
    n180,
    n209
  );


  or
  g390
  (
    n393,
    n192,
    n370,
    n372,
    n378
  );


  nor
  g391
  (
    n420,
    n251,
    n262,
    n230,
    n227
  );


  xor
  g392
  (
    n445,
    n242,
    n170,
    n362,
    n361
  );


  or
  g393
  (
    n483,
    n373,
    n177,
    n244,
    n210
  );


  xnor
  g394
  (
    n426,
    n209,
    n203,
    n177,
    n161
  );


  nand
  g395
  (
    n444,
    n175,
    n363,
    n185,
    n357
  );


  nor
  g396
  (
    n438,
    n379,
    n186,
    n198,
    n240
  );


  and
  g397
  (
    KeyWire_0_27,
    n212,
    n179,
    n256,
    n372
  );


  xor
  g398
  (
    n407,
    n252,
    n356,
    n210,
    n360
  );


  nor
  g399
  (
    KeyWire_0_20,
    n191,
    n187,
    n223,
    n184
  );


  xnor
  g400
  (
    n441,
    n372,
    n176,
    n201,
    n168
  );


  nor
  g401
  (
    n482,
    n235,
    n188,
    n239,
    n222
  );


  nand
  g402
  (
    n413,
    n180,
    n166,
    n356,
    n358
  );


  nor
  g403
  (
    n470,
    n187,
    n369,
    n238,
    n215
  );


  xnor
  g404
  (
    n443,
    n365,
    n178,
    n207,
    n215
  );


  or
  g405
  (
    n408,
    n355,
    n174,
    n167,
    n358
  );


  nand
  g406
  (
    n402,
    n373,
    n357,
    n359,
    n370
  );


  or
  g407
  (
    n424,
    n175,
    n199,
    n171,
    n226
  );


  nor
  g408
  (
    n457,
    n218,
    n380,
    n188,
    n233
  );


  and
  g409
  (
    n400,
    n364,
    n374,
    n179
  );


  and
  g410
  (
    n386,
    n246,
    n233,
    n193,
    n174
  );


  and
  g411
  (
    n452,
    n210,
    n222,
    n362,
    n167
  );


  xor
  g412
  (
    n455,
    n248,
    n379,
    n357,
    n368
  );


  or
  g413
  (
    n459,
    n360,
    n241,
    n258,
    n250
  );


  nand
  g414
  (
    n429,
    n211,
    n189,
    n205,
    n172
  );


  nand
  g415
  (
    n389,
    n158,
    n173,
    n166,
    n359
  );


  nand
  g416
  (
    n381,
    n234,
    n377,
    n195,
    n359
  );


  or
  g417
  (
    n382,
    n194,
    n249,
    n259,
    n209
  );


  nand
  g418
  (
    n396,
    n378,
    n258,
    n262,
    n259
  );


  nor
  g419
  (
    n388,
    n170,
    n377,
    n355,
    n213
  );


  xor
  g420
  (
    n463,
    n172,
    n200,
    n165,
    n240
  );


  xor
  g421
  (
    n458,
    n177,
    n188,
    n182,
    n208
  );


  nand
  g422
  (
    n410,
    n186,
    n221,
    n249,
    n197
  );


  or
  g423
  (
    n465,
    n227,
    n207,
    n228,
    n253
  );


  and
  g424
  (
    n411,
    n185,
    n186,
    n380,
    n220
  );


  xor
  g425
  (
    KeyWire_0_57,
    n234,
    n182,
    n263
  );


  or
  g426
  (
    n461,
    n236,
    n202,
    n380,
    n257
  );


  and
  g427
  (
    n448,
    n171,
    n372,
    n361,
    n375
  );


  nand
  g428
  (
    n383,
    n366,
    n169,
    n172,
    n211
  );


  xnor
  g429
  (
    n437,
    n163,
    n260,
    n365,
    n261
  );


  nor
  g430
  (
    n434,
    n357,
    n244,
    n191,
    n376
  );


  nand
  g431
  (
    n416,
    n245,
    n355,
    n368,
    n375
  );


  nand
  g432
  (
    n481,
    n380,
    n204,
    n359,
    n199
  );


  and
  g433
  (
    n409,
    n237,
    n231,
    n376,
    n252
  );


  xor
  g434
  (
    KeyWire_0_8,
    n181,
    n232,
    n169,
    n242
  );


  and
  g435
  (
    n439,
    n363,
    n231,
    n198,
    n371
  );


  xor
  g436
  (
    n417,
    n259,
    n228,
    n377,
    n216
  );


  nor
  g437
  (
    n436,
    n369,
    n189,
    n263,
    n183
  );


  xnor
  g438
  (
    n405,
    n243,
    n199,
    n195,
    n168
  );


  xnor
  g439
  (
    n433,
    n166,
    n221,
    n250,
    n261
  );


  and
  g440
  (
    n447,
    n262,
    n156,
    n203,
    n366
  );


  nor
  g441
  (
    n412,
    n229,
    n255,
    n365,
    n378
  );


  or
  g442
  (
    n476,
    n260,
    n258,
    n226,
    n216
  );


  xor
  g443
  (
    n399,
    n362,
    n203,
    n200,
    n220
  );


  nor
  g444
  (
    n392,
    n219,
    n237,
    n252,
    n230
  );


  or
  g445
  (
    n473,
    n249,
    n208,
    n190,
    n194
  );


  and
  g446
  (
    n428,
    n173,
    n196,
    n356,
    n175
  );


  and
  g447
  (
    n442,
    n376,
    n242,
    n169,
    n253
  );


  or
  g448
  (
    n456,
    n167,
    n243,
    n201,
    n371
  );


  xnor
  g449
  (
    n387,
    n200,
    n373,
    n234,
    n180
  );


  xor
  g450
  (
    n397,
    n370,
    n208,
    n217,
    n220
  );


  nand
  g451
  (
    n414,
    n202,
    n159,
    n264,
    n197
  );


  nor
  g452
  (
    n484,
    n171,
    n239,
    n181,
    n206
  );


  xor
  g453
  (
    KeyWire_0_10,
    n238,
    n236,
    n206,
    n245
  );


  nand
  g454
  (
    KeyWire_0_0,
    n364,
    n367,
    n217,
    n254
  );


  xnor
  g455
  (
    n462,
    n358,
    n219,
    n164,
    n224
  );


  or
  g456
  (
    n432,
    n370,
    n213,
    n369,
    n238
  );


  xor
  g457
  (
    n524,
    n385,
    n289,
    n337,
    n384
  );


  and
  g458
  (
    n556,
    n27,
    n340,
    n88,
    n344
  );


  and
  g459
  (
    n512,
    n400,
    n27,
    n417,
    n330
  );


  or
  g460
  (
    n543,
    n271,
    n413,
    n273,
    n390
  );


  nor
  g461
  (
    n497,
    n423,
    n335,
    n344,
    n403
  );


  or
  g462
  (
    n553,
    n422,
    n316,
    n290,
    n265
  );


  xor
  g463
  (
    n538,
    n299,
    n396,
    n392,
    n99
  );


  xor
  g464
  (
    KeyWire_0_5,
    n390,
    n287,
    n396,
    n418
  );


  xnor
  g465
  (
    KeyWire_0_56,
    n330,
    n409,
    n325,
    n289
  );


  and
  g466
  (
    n591,
    n288,
    n397,
    n402,
    n323
  );


  nor
  g467
  (
    KeyWire_0_59,
    n266,
    n306,
    n308,
    n320
  );


  nor
  g468
  (
    n494,
    n292,
    n338,
    n91,
    n422
  );


  nand
  g469
  (
    n568,
    n398,
    n314,
    n313,
    n26
  );


  xnor
  g470
  (
    n586,
    n382,
    n87,
    n267,
    n391
  );


  xnor
  g471
  (
    n507,
    n411,
    n391,
    n295,
    n322
  );


  nor
  g472
  (
    n585,
    n421,
    n271,
    n294
  );


  xor
  g473
  (
    n570,
    n412,
    n303,
    n98,
    n324
  );


  or
  g474
  (
    n516,
    n323,
    n291,
    n311,
    n334
  );


  xor
  g475
  (
    n565,
    n296,
    n267,
    n91,
    n316
  );


  and
  g476
  (
    n566,
    n92,
    n393,
    n415,
    n25
  );


  nand
  g477
  (
    n552,
    n342,
    n318,
    n274,
    n416
  );


  or
  g478
  (
    n536,
    n281,
    n312,
    n275,
    n406
  );


  nand
  g479
  (
    n559,
    n309,
    n97,
    n86,
    n89
  );


  nor
  g480
  (
    n519,
    n411,
    n266,
    n272,
    n331
  );


  and
  g481
  (
    n502,
    n328,
    n395,
    n85,
    n333
  );


  or
  g482
  (
    n540,
    n345,
    n383,
    n328,
    n96
  );


  nand
  g483
  (
    n555,
    n269,
    n389,
    n280,
    n402
  );


  nand
  g484
  (
    n593,
    n90,
    n343,
    n398
  );


  or
  g485
  (
    n492,
    n93,
    n27,
    n92,
    n303
  );


  nand
  g486
  (
    n589,
    n405,
    n325,
    n286,
    n324
  );


  or
  g487
  (
    n564,
    n273,
    n420,
    n400,
    n399
  );


  and
  g488
  (
    n493,
    n401,
    n399,
    n316,
    n315
  );


  xor
  g489
  (
    n557,
    n308,
    n405,
    n300,
    n336
  );


  xnor
  g490
  (
    n546,
    n387,
    n312,
    n404,
    n87
  );


  nor
  g491
  (
    n515,
    n294,
    n297,
    n27,
    n287
  );


  and
  g492
  (
    n594,
    n412,
    n272,
    n296,
    n298
  );


  xnor
  g493
  (
    n541,
    n418,
    n94,
    n97,
    n385
  );


  nand
  g494
  (
    n573,
    n422,
    n26,
    n339,
    n338
  );


  or
  g495
  (
    KeyWire_0_55,
    n315,
    n396,
    n412,
    n309
  );


  and
  g496
  (
    n579,
    n280,
    n312,
    n329,
    n272
  );


  xnor
  g497
  (
    n534,
    n318,
    n410,
    n279,
    n418
  );


  or
  g498
  (
    n578,
    n330,
    n282,
    n421,
    n335
  );


  nor
  g499
  (
    n574,
    n281,
    n89,
    n93,
    n265
  );


  and
  g500
  (
    n500,
    n303,
    n322,
    n343,
    n329
  );


  or
  g501
  (
    KeyWire_0_7,
    n270,
    n305,
    n398,
    n340
  );


  or
  g502
  (
    n503,
    n304,
    n390,
    n98,
    n317
  );


  nand
  g503
  (
    n537,
    n288,
    n286,
    n285,
    n325
  );


  xor
  g504
  (
    n517,
    n93,
    n331,
    n305,
    n394
  );


  xnor
  g505
  (
    n560,
    n94,
    n283,
    n320,
    n299
  );


  or
  g506
  (
    n505,
    n406,
    n293,
    n324,
    n414
  );


  and
  g507
  (
    n531,
    n90,
    n392,
    n298,
    n393
  );


  xor
  g508
  (
    n580,
    n295,
    n326,
    n268,
    n293
  );


  xor
  g509
  (
    n582,
    n419,
    n300,
    n279,
    n86
  );


  nand
  g510
  (
    n504,
    n332,
    n395,
    n342,
    n327
  );


  nor
  g511
  (
    n513,
    n97,
    n410,
    n284,
    n332
  );


  xnor
  g512
  (
    n498,
    n281,
    n397,
    n403,
    n399
  );


  or
  g513
  (
    n518,
    n284,
    n382,
    n98,
    n310
  );


  or
  g514
  (
    n532,
    n346,
    n388,
    n334,
    n264
  );


  xor
  g515
  (
    n525,
    n97,
    n333,
    n300,
    n323
  );


  or
  g516
  (
    n567,
    n394,
    n283,
    n387,
    n96
  );


  xor
  g517
  (
    n545,
    n320,
    n311,
    n381,
    n90
  );


  nor
  g518
  (
    n506,
    n410,
    n95,
    n341,
    n269
  );


  nand
  g519
  (
    n533,
    n385,
    n88,
    n383,
    n90
  );


  nand
  g520
  (
    n495,
    n99,
    n285,
    n301,
    n341
  );


  nor
  g521
  (
    n569,
    n291,
    n403,
    n405,
    n87
  );


  xor
  g522
  (
    n499,
    n423,
    n415,
    n292,
    n294
  );


  nor
  g523
  (
    n496,
    n290,
    n327,
    n339,
    n413
  );


  and
  g524
  (
    n544,
    n95,
    n397,
    n301,
    n319
  );


  nand
  g525
  (
    n563,
    n298,
    n393,
    n394,
    n409
  );


  nand
  g526
  (
    n530,
    n319,
    n89,
    n401,
    n278
  );


  nor
  g527
  (
    n520,
    n419,
    n411,
    n277,
    n305
  );


  xnor
  g528
  (
    n572,
    n286,
    n419,
    n282,
    n313
  );


  and
  g529
  (
    n554,
    n404,
    n384,
    n389,
    n94
  );


  xor
  g530
  (
    n523,
    n288,
    n284,
    n296,
    n273
  );


  nand
  g531
  (
    n583,
    n391,
    n292,
    n309,
    n388
  );


  nand
  g532
  (
    n571,
    n98,
    n310,
    n317,
    n416
  );


  nand
  g533
  (
    n527,
    n321,
    n297,
    n306,
    n409
  );


  xor
  g534
  (
    n562,
    n307,
    n88,
    n406,
    n413
  );


  xor
  g535
  (
    n510,
    n88,
    n314,
    n386,
    n297
  );


  or
  g536
  (
    KeyWire_0_46,
    n26,
    n337,
    n392
  );


  nand
  g537
  (
    n548,
    n387,
    n290,
    n302,
    n283
  );


  xor
  g538
  (
    n522,
    n91,
    n415,
    n96,
    n314
  );


  xor
  g539
  (
    n488,
    n277,
    n424,
    n95,
    n275
  );


  xor
  g540
  (
    n561,
    n386,
    n420,
    n287,
    n423
  );


  xor
  g541
  (
    n535,
    n99,
    n317,
    n96,
    n381
  );


  nor
  g542
  (
    n489,
    n322,
    n275,
    n270,
    n401
  );


  xnor
  g543
  (
    n485,
    n282,
    n291,
    n321,
    n384
  );


  nand
  g544
  (
    n550,
    n321,
    n414,
    n295,
    n417
  );


  nor
  g545
  (
    n529,
    n274,
    n345,
    n276
  );


  nor
  g546
  (
    n514,
    n408,
    n407,
    n92,
    n386
  );


  xnor
  g547
  (
    n590,
    n382,
    n334,
    n313,
    n274
  );


  nor
  g548
  (
    n490,
    n404,
    n26,
    n278,
    n407
  );


  or
  g549
  (
    n549,
    n92,
    n264,
    n416,
    n307
  );


  nor
  g550
  (
    KeyWire_0_1,
    n402,
    n335,
    n339,
    n94
  );


  xor
  g551
  (
    n587,
    n408,
    n86,
    n383,
    n333
  );


  xnor
  g552
  (
    n528,
    n420,
    n311,
    n326,
    n332
  );


  xnor
  g553
  (
    n558,
    n270,
    n267,
    n265,
    n266
  );


  nand
  g554
  (
    n576,
    n341,
    n268,
    n93,
    n276
  );


  xnor
  g555
  (
    n575,
    n268,
    n285,
    n408,
    n336
  );


  nand
  g556
  (
    n509,
    n85,
    n345,
    n302,
    n417
  );


  nand
  g557
  (
    n491,
    n421,
    n89,
    n85,
    n304
  );


  or
  g558
  (
    n501,
    n318,
    n304,
    n293,
    n277
  );


  nor
  g559
  (
    KeyWire_0_53,
    n344,
    n269,
    n328,
    n407
  );


  xor
  g560
  (
    n542,
    n331,
    n327,
    n306,
    n278
  );


  or
  g561
  (
    n521,
    n302,
    n336,
    n279,
    n85
  );


  xnor
  g562
  (
    n581,
    n315,
    n95,
    n414,
    n400
  );


  or
  g563
  (
    n487,
    n388,
    n308,
    n340,
    n342
  );


  and
  g564
  (
    n526,
    n301,
    n381,
    n307,
    n319
  );


  xnor
  g565
  (
    n539,
    n326,
    n86,
    n299,
    n91
  );


  nor
  g566
  (
    n547,
    n389,
    n310,
    n289,
    n280
  );


  xor
  g567
  (
    n551,
    n338,
    n329,
    n395,
    n87
  );


  xnor
  g568
  (
    n619,
    n429,
    n455,
    n447,
    n476
  );


  xor
  g569
  (
    n674,
    n559,
    n555,
    n508,
    n465
  );


  or
  g570
  (
    n607,
    n512,
    n465,
    n479,
    n500
  );


  nand
  g571
  (
    n655,
    n444,
    n560,
    n432,
    n442
  );


  xor
  g572
  (
    n601,
    n457,
    n505,
    n449,
    n545
  );


  xnor
  g573
  (
    n645,
    n426,
    n439,
    n438,
    n532
  );


  xor
  g574
  (
    KeyWire_0_43,
    n473,
    n472,
    n449,
    n429
  );


  xnor
  g575
  (
    n651,
    n550,
    n436,
    n470,
    n461
  );


  or
  g576
  (
    KeyWire_0_23,
    n106,
    n469,
    n547,
    n521
  );


  nand
  g577
  (
    n631,
    n463,
    n452,
    n425,
    n466
  );


  and
  g578
  (
    n602,
    n433,
    n518,
    n473,
    n502
  );


  or
  g579
  (
    n611,
    n549,
    n441,
    n103
  );


  nand
  g580
  (
    KeyWire_0_4,
    n427,
    n462,
    n444,
    n527
  );


  nand
  g581
  (
    n604,
    n437,
    n542,
    n456,
    n426
  );


  nor
  g582
  (
    n679,
    n443,
    n470,
    n432,
    n483
  );


  nor
  g583
  (
    n647,
    n493,
    n546,
    n482,
    n540
  );


  xor
  g584
  (
    n640,
    n437,
    n103,
    n104,
    n529
  );


  or
  g585
  (
    n618,
    n530,
    n543,
    n475,
    n471
  );


  or
  g586
  (
    n670,
    n106,
    n106,
    n454,
    n449
  );


  nor
  g587
  (
    n643,
    n472,
    n443,
    n486,
    n562
  );


  or
  g588
  (
    n634,
    n104,
    n455,
    n531,
    n446
  );


  xor
  g589
  (
    n676,
    n464,
    n474,
    n568,
    n434
  );


  nand
  g590
  (
    n678,
    n507,
    n503,
    n446,
    n445
  );


  nor
  g591
  (
    n616,
    n435,
    n453,
    n440,
    n460
  );


  xnor
  g592
  (
    n644,
    n102,
    n516,
    n432,
    n436
  );


  or
  g593
  (
    n597,
    n457,
    n475,
    n105,
    n484
  );


  or
  g594
  (
    n669,
    n484,
    n448,
    n517,
    n99
  );


  xnor
  g595
  (
    n660,
    n428,
    n455,
    n480,
    n434
  );


  xnor
  g596
  (
    n646,
    n438,
    n491,
    n468,
    n536
  );


  or
  g597
  (
    n621,
    n465,
    n451,
    n458,
    n431
  );


  xnor
  g598
  (
    n617,
    n101,
    n461,
    n557,
    n564
  );


  xnor
  g599
  (
    KeyWire_0_38,
    n447,
    n435,
    n563,
    n519
  );


  xor
  g600
  (
    n641,
    n475,
    n479,
    n448,
    n438
  );


  nand
  g601
  (
    n630,
    n489,
    n107,
    n470,
    n556
  );


  or
  g602
  (
    n605,
    n439,
    n477,
    n476,
    n473
  );


  or
  g603
  (
    n653,
    n425,
    n484,
    n428,
    n446
  );


  xor
  g604
  (
    n608,
    n466,
    n520,
    n472,
    n480
  );


  xnor
  g605
  (
    n612,
    n469,
    n522,
    n477,
    n447
  );


  xor
  g606
  (
    n635,
    n470,
    n444,
    n454,
    n453
  );


  and
  g607
  (
    n610,
    n440,
    n526,
    n101,
    n498
  );


  xnor
  g608
  (
    n652,
    n100,
    n487,
    n442,
    n459
  );


  nor
  g609
  (
    n680,
    n544,
    n460,
    n450,
    n485
  );


  or
  g610
  (
    n661,
    n482,
    n424,
    n461,
    n454
  );


  nor
  g611
  (
    n659,
    n465,
    n431,
    n453,
    n450
  );


  xnor
  g612
  (
    n628,
    n467,
    n471,
    n436,
    n431
  );


  nand
  g613
  (
    n598,
    n479,
    n456,
    n477,
    n482
  );


  and
  g614
  (
    n657,
    n570,
    n103,
    n496,
    n102
  );


  nand
  g615
  (
    n675,
    n440,
    n426,
    n441,
    n455
  );


  xor
  g616
  (
    n648,
    n449,
    n481,
    n442,
    n447
  );


  xor
  g617
  (
    n658,
    n100,
    n459,
    n424,
    n482
  );


  xnor
  g618
  (
    n609,
    n494,
    n471,
    n458,
    n561
  );


  or
  g619
  (
    n615,
    n433,
    n102,
    n483,
    n515
  );


  nor
  g620
  (
    n599,
    n525,
    n471,
    n475,
    n433
  );


  nor
  g621
  (
    n625,
    n483,
    n554,
    n504,
    n528
  );


  nor
  g622
  (
    n620,
    n483,
    n514,
    n467,
    n492
  );


  and
  g623
  (
    n603,
    n481,
    n100,
    n429,
    n104
  );


  nor
  g624
  (
    n629,
    n444,
    n523,
    n468,
    n448
  );


  nand
  g625
  (
    n665,
    n480,
    n506,
    n435,
    n477
  );


  xnor
  g626
  (
    n633,
    n464,
    n459,
    n100,
    n104
  );


  nand
  g627
  (
    n600,
    n472,
    n452,
    n105,
    n467
  );


  and
  g628
  (
    n626,
    n456,
    n551,
    n453,
    n458
  );


  nor
  g629
  (
    n668,
    n476,
    n480,
    n497,
    n464
  );


  and
  g630
  (
    n614,
    n460,
    n448,
    n481,
    n466
  );


  xor
  g631
  (
    n637,
    n430,
    n478,
    n437,
    n510
  );


  nor
  g632
  (
    n681,
    n442,
    n452,
    n462,
    n439
  );


  nand
  g633
  (
    n650,
    n509,
    n459,
    n479,
    n445
  );


  xor
  g634
  (
    n667,
    n524,
    n478,
    n107,
    n450
  );


  xnor
  g635
  (
    n639,
    n457,
    n463,
    n469,
    n103
  );


  or
  g636
  (
    n624,
    n101,
    n458,
    n476,
    n553
  );


  xnor
  g637
  (
    n638,
    n539,
    n481,
    n474,
    n105
  );


  xnor
  g638
  (
    KeyWire_0_63,
    n452,
    n513,
    n501,
    n495
  );


  and
  g639
  (
    n654,
    n430,
    n430,
    n460,
    n445
  );


  or
  g640
  (
    n606,
    n566,
    n101,
    n461,
    n534
  );


  nor
  g641
  (
    n622,
    n538,
    n468,
    n427,
    n451
  );


  and
  g642
  (
    n613,
    n474,
    n467,
    n463,
    n441
  );


  and
  g643
  (
    KeyWire_0_35,
    n450,
    n464,
    n443,
    n473
  );


  and
  g644
  (
    n662,
    n533,
    n106,
    n552,
    n558
  );


  or
  g645
  (
    n642,
    n102,
    n548,
    n457,
    n466
  );


  nor
  g646
  (
    n673,
    n462,
    n456,
    n478,
    n425
  );


  nor
  g647
  (
    n664,
    n488,
    n478,
    n565,
    n434
  );


  nor
  g648
  (
    n656,
    n454,
    n468,
    n490,
    n484
  );


  or
  g649
  (
    n632,
    n474,
    n499,
    n535,
    n427
  );


  nand
  g650
  (
    n627,
    n541,
    n451,
    n462,
    n469
  );


  xnor
  g651
  (
    n636,
    n446,
    n511,
    n443,
    n463
  );


  or
  g652
  (
    n677,
    n105,
    n445,
    n428,
    n567
  );


  xnor
  g653
  (
    n649,
    n451,
    n569,
    n440,
    n537
  );


  buf
  g654
  (
    n684,
    n592
  );


  not
  g655
  (
    n688,
    n610
  );


  buf
  g656
  (
    n702,
    n351
  );


  not
  g657
  (
    n685,
    n350
  );


  xnor
  g658
  (
    n694,
    n576,
    n583
  );


  nand
  g659
  (
    n692,
    n347,
    n354,
    n350,
    n615
  );


  and
  g660
  (
    n703,
    n353,
    n354,
    n579,
    n581
  );


  xor
  g661
  (
    n699,
    n601,
    n573,
    n353,
    n606
  );


  nand
  g662
  (
    n682,
    n591,
    n575,
    n572,
    n346
  );


  xor
  g663
  (
    n697,
    n590,
    n587,
    n350,
    n348
  );


  nand
  g664
  (
    n701,
    n349,
    n595,
    n354,
    n353
  );


  nand
  g665
  (
    n686,
    n351,
    n612,
    n615,
    n348
  );


  or
  g666
  (
    KeyWire_0_9,
    n574,
    n593,
    n349,
    n600
  );


  xor
  g667
  (
    n696,
    n614,
    n347,
    n605,
    n582
  );


  nand
  g668
  (
    n687,
    n351,
    n604,
    n602,
    n578
  );


  nor
  g669
  (
    n683,
    n594,
    n577,
    n346,
    n608
  );


  xor
  g670
  (
    n689,
    n615,
    n586,
    n597,
    n607
  );


  nand
  g671
  (
    KeyWire_0_29,
    n585,
    n354,
    n599,
    n352
  );


  and
  g672
  (
    n695,
    n609,
    n349,
    n596,
    n352
  );


  or
  g673
  (
    n698,
    n347,
    n603,
    n598,
    n352
  );


  xnor
  g674
  (
    n700,
    n588,
    n348,
    n571,
    n589
  );


  or
  g675
  (
    n691,
    n584,
    n613,
    n611,
    n580
  );


  or
  g676
  (
    n752,
    n110,
    n641,
    n701,
    n669
  );


  nor
  g677
  (
    n762,
    n638,
    n660,
    n644,
    n654
  );


  xor
  g678
  (
    n753,
    n624,
    n683,
    n628,
    n109
  );


  xnor
  g679
  (
    n750,
    n679,
    n696,
    n109,
    n701
  );


  nand
  g680
  (
    n749,
    n702,
    n681,
    n110,
    n660
  );


  xnor
  g681
  (
    n767,
    n627,
    n678,
    n682
  );


  and
  g682
  (
    n725,
    n663,
    n111,
    n648,
    n622
  );


  nand
  g683
  (
    n724,
    n109,
    n687,
    n700
  );


  nor
  g684
  (
    n737,
    n670,
    n681,
    n627,
    n649
  );


  or
  g685
  (
    n765,
    n702,
    n634,
    n695
  );


  nor
  g686
  (
    n718,
    n666,
    n628,
    n697,
    n685
  );


  xor
  g687
  (
    n722,
    n694,
    n698,
    n703,
    n629
  );


  and
  g688
  (
    n732,
    n663,
    n674,
    n677,
    n670
  );


  nor
  g689
  (
    n766,
    n672,
    n633,
    n668,
    n639
  );


  or
  g690
  (
    n771,
    n631,
    n690,
    n636,
    n111
  );


  and
  g691
  (
    n741,
    n698,
    n658,
    n690,
    n672
  );


  and
  g692
  (
    n734,
    n650,
    n640,
    n636,
    n679
  );


  nand
  g693
  (
    KeyWire_0_42,
    n639,
    n623,
    n649,
    n673
  );


  nand
  g694
  (
    n731,
    n624,
    n684,
    n617,
    n638
  );


  nor
  g695
  (
    n726,
    n619,
    n669,
    n659,
    n625
  );


  nand
  g696
  (
    n761,
    n632,
    n657,
    n635,
    n691
  );


  and
  g697
  (
    n739,
    n647,
    n655,
    n650,
    n621
  );


  xor
  g698
  (
    n759,
    n661,
    n676,
    n626,
    n668
  );


  nand
  g699
  (
    n720,
    n678,
    n665,
    n634,
    n632
  );


  nor
  g700
  (
    n706,
    n656,
    n622,
    n674,
    n693
  );


  nor
  g701
  (
    n758,
    n686,
    n636,
    n620,
    n651
  );


  or
  g702
  (
    n713,
    n686,
    n672,
    n688
  );


  xnor
  g703
  (
    n774,
    n655,
    n655,
    n701,
    n684
  );


  xor
  g704
  (
    n719,
    n617,
    n659,
    n671,
    n676
  );


  nor
  g705
  (
    n733,
    n630,
    n620,
    n702,
    n652
  );


  xnor
  g706
  (
    n714,
    n671,
    n662,
    n630,
    n107
  );


  xor
  g707
  (
    n730,
    n691,
    n616,
    n617,
    n698
  );


  xor
  g708
  (
    KeyWire_0_34,
    n661,
    n623,
    n685,
    n616
  );


  xor
  g709
  (
    n751,
    n618,
    n676,
    n656,
    n642
  );


  and
  g710
  (
    n772,
    n651,
    n699,
    n621,
    n695
  );


  and
  g711
  (
    n738,
    n662,
    n664,
    n665,
    n688
  );


  nand
  g712
  (
    n747,
    n649,
    n647,
    n624,
    n646
  );


  or
  g713
  (
    n712,
    n626,
    n658,
    n628,
    n700
  );


  xnor
  g714
  (
    n763,
    n673,
    n664,
    n686,
    n679
  );


  nor
  g715
  (
    n704,
    n653,
    n641,
    n644,
    n684
  );


  or
  g716
  (
    n716,
    n640,
    n638,
    n674,
    n678
  );


  xor
  g717
  (
    n743,
    n675,
    n622,
    n692,
    n694
  );


  nor
  g718
  (
    n756,
    n652,
    n677,
    n702,
    n668
  );


  nand
  g719
  (
    n740,
    n619,
    n642,
    n108,
    n648
  );


  or
  g720
  (
    n769,
    n696,
    n699,
    n620,
    n625
  );


  xnor
  g721
  (
    n717,
    n662,
    n698,
    n657,
    n697
  );


  and
  g722
  (
    n711,
    n646,
    n632,
    n696,
    n107
  );


  and
  g723
  (
    n775,
    n700,
    n671,
    n111,
    n659
  );


  nand
  g724
  (
    n715,
    n657,
    n660,
    n629,
    n631
  );


  or
  g725
  (
    n748,
    n639,
    n637,
    n689,
    n626
  );


  xor
  g726
  (
    n735,
    n703,
    n647,
    n680,
    n653
  );


  nor
  g727
  (
    KeyWire_0_19,
    n680,
    n637,
    n645,
    n667
  );


  xor
  g728
  (
    n723,
    n664,
    n642,
    n693,
    n643
  );


  nand
  g729
  (
    n728,
    n665,
    n619,
    n634,
    n691
  );


  nor
  g730
  (
    n727,
    n646,
    n633,
    n110
  );


  xor
  g731
  (
    n757,
    n693,
    n627,
    n651,
    n683
  );


  or
  g732
  (
    n754,
    n689,
    n683,
    n687,
    n650
  );


  and
  g733
  (
    n770,
    n680,
    n616,
    n108,
    n621
  );


  xor
  g734
  (
    n744,
    n701,
    n666,
    n673,
    n703
  );


  nor
  g735
  (
    n729,
    n637,
    n652,
    n677,
    n625
  );


  xor
  g736
  (
    KeyWire_0_37,
    n675,
    n685,
    n667,
    n700
  );


  xnor
  g737
  (
    n708,
    n631,
    n635,
    n644,
    n661
  );


  xnor
  g738
  (
    n746,
    n697,
    n643,
    n675,
    n653
  );


  or
  g739
  (
    KeyWire_0_32,
    n643,
    n645,
    n623,
    n641
  );


  xor
  g740
  (
    n705,
    n690,
    n663,
    n667,
    n654
  );


  and
  g741
  (
    n760,
    n658,
    n703,
    n670,
    n654
  );


  or
  g742
  (
    n707,
    n108,
    n669,
    n656,
    n629
  );


  xnor
  g743
  (
    n721,
    n699,
    n645,
    n689,
    n682
  );


  and
  g744
  (
    n773,
    n618,
    n630,
    n635,
    n699
  );


  nor
  g745
  (
    n710,
    n633,
    n681,
    n618,
    n692
  );


  or
  g746
  (
    KeyWire_0_54,
    n648,
    n108,
    n109,
    n694
  );


  or
  g747
  (
    n764,
    n692,
    n640,
    n111,
    n666
  );


  xnor
  g748
  (
    n781,
    n718,
    n723,
    n121,
    n123
  );


  xnor
  g749
  (
    n793,
    n715,
    n125,
    n124
  );


  xor
  g750
  (
    n779,
    n707,
    n116,
    n122,
    n117
  );


  xnor
  g751
  (
    n784,
    n710,
    n115,
    n118,
    n123
  );


  nor
  g752
  (
    n787,
    n122,
    n120,
    n125,
    n722
  );


  nor
  g753
  (
    n788,
    n125,
    n121,
    n115,
    n119
  );


  nand
  g754
  (
    n776,
    n712,
    n711,
    n121,
    n120
  );


  xor
  g755
  (
    KeyWire_0_2,
    n113,
    n113,
    n126,
    n120
  );


  and
  g756
  (
    n786,
    n116,
    n116,
    n115,
    n120
  );


  or
  g757
  (
    n791,
    n112,
    n716,
    n119,
    n124
  );


  xor
  g758
  (
    n789,
    n117,
    n720,
    n115,
    n713
  );


  and
  g759
  (
    n790,
    n116,
    n119,
    n126,
    n114
  );


  nor
  g760
  (
    n780,
    n719,
    n124,
    n717
  );


  xnor
  g761
  (
    n792,
    n704,
    n112,
    n117,
    n709
  );


  nor
  g762
  (
    n795,
    n114,
    n112
  );


  xnor
  g763
  (
    n783,
    n714,
    n118,
    n123
  );


  nand
  g764
  (
    n785,
    n118,
    n126,
    n117,
    n122
  );


  xnor
  g765
  (
    KeyWire_0_17,
    n708,
    n123,
    n126,
    n113
  );


  and
  g766
  (
    n778,
    n121,
    n705,
    n122,
    n706
  );


  xnor
  g767
  (
    n794,
    n114,
    n721,
    n119,
    n113
  );


  and
  g768
  (
    n796,
    n759,
    n740,
    n783,
    n792
  );


  xnor
  g769
  (
    n799,
    n755,
    n725,
    n788,
    n747
  );


  nand
  g770
  (
    n806,
    n777,
    n746,
    n734,
    n763
  );


  and
  g771
  (
    n810,
    n794,
    n795,
    n771,
    n738
  );


  nor
  g772
  (
    n807,
    n781,
    n766,
    n752,
    n769
  );


  or
  g773
  (
    n802,
    n737,
    n782,
    n750,
    n784
  );


  and
  g774
  (
    n805,
    n735,
    n741,
    n727,
    n758
  );


  or
  g775
  (
    n797,
    n754,
    n751,
    n785,
    n791
  );


  or
  g776
  (
    n804,
    n739,
    n743,
    n745,
    n731
  );


  xor
  g777
  (
    n800,
    n770,
    n730,
    n768,
    n761
  );


  nor
  g778
  (
    n803,
    n765,
    n729,
    n772,
    n724
  );


  xnor
  g779
  (
    n811,
    n728,
    n780,
    n776,
    n744
  );


  nand
  g780
  (
    n798,
    n749,
    n764,
    n774,
    n767
  );


  nand
  g781
  (
    n801,
    n760,
    n789,
    n756,
    n742
  );


  xnor
  g782
  (
    n808,
    n748,
    n786,
    n787,
    n732
  );


  and
  g783
  (
    n813,
    n779,
    n790,
    n736,
    n753
  );


  xnor
  g784
  (
    n809,
    n733,
    n726,
    n762,
    n778
  );


  and
  g785
  (
    n812,
    n773,
    n757,
    n775,
    n793
  );


  xnor
  KeyGate_0_0
  (
    n471,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n508,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n782,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n186,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n671,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n577,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n30,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n584,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n403,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n693,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n451,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n49,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n80,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n129,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n336,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n202,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n151,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n777,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n355,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n736,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n469,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n128,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n367,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n623,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n141,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n269,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n155,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n421,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n331,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n690,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n55,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n201,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n709,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n229,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n745,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n663,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n440,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n742,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n666,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n261,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n116,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n190,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n755,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n672,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n330,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n204,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n486,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n112,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n72,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n266,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n76,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n380,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n300,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n588,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n768,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n595,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n592,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n453,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n370,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n511,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n467,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n291,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n264,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n596,
    KeyNOTWire_0_63
  );


endmodule


