

module Stat_1000_151
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n767,
  n1008,
  n1011,
  n1021,
  n1027,
  n1025,
  n1032,
  n1006,
  n1017,
  n1031,
  n1010,
  n1012,
  n1013,
  n1014,
  n1003,
  n1026,
  n1028,
  n1005,
  n1020,
  n1029,
  n1030,
  n1019,
  n1018,
  n1022,
  n1002,
  n1015,
  n1023,
  n1024,
  n1016,
  n1004,
  n1009,
  n1007
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n767;output n1008;output n1011;output n1021;output n1027;output n1025;output n1032;output n1006;output n1017;output n1031;output n1010;output n1012;output n1013;output n1014;output n1003;output n1026;output n1028;output n1005;output n1020;output n1029;output n1030;output n1019;output n1018;output n1022;output n1002;output n1015;output n1023;output n1024;output n1016;output n1004;output n1009;output n1007;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n54,
    n13
  );


  not
  g1
  (
    n116,
    n2
  );


  buf
  g2
  (
    n69,
    n22
  );


  not
  g3
  (
    n42,
    n26
  );


  buf
  g4
  (
    n130,
    n24
  );


  not
  g5
  (
    n129,
    n12
  );


  buf
  g6
  (
    KeyWire_0_12,
    n7
  );


  not
  g7
  (
    n47,
    n8
  );


  buf
  g8
  (
    n127,
    n5
  );


  buf
  g9
  (
    n92,
    n17
  );


  not
  g10
  (
    KeyWire_0_4,
    n22
  );


  buf
  g11
  (
    n132,
    n27
  );


  buf
  g12
  (
    n86,
    n11
  );


  buf
  g13
  (
    n142,
    n17
  );


  buf
  g14
  (
    n89,
    n11
  );


  buf
  g15
  (
    KeyWire_0_16,
    n29
  );


  not
  g16
  (
    n78,
    n16
  );


  buf
  g17
  (
    n147,
    n11
  );


  buf
  g18
  (
    KeyWire_0_2,
    n4
  );


  buf
  g19
  (
    n96,
    n17
  );


  not
  g20
  (
    n114,
    n22
  );


  not
  g21
  (
    n57,
    n30
  );


  buf
  g22
  (
    n94,
    n9
  );


  buf
  g23
  (
    n103,
    n10
  );


  not
  g24
  (
    n75,
    n28
  );


  buf
  g25
  (
    n124,
    n22
  );


  not
  g26
  (
    n146,
    n18
  );


  buf
  g27
  (
    n49,
    n12
  );


  buf
  g28
  (
    n115,
    n29
  );


  buf
  g29
  (
    n95,
    n10
  );


  not
  g30
  (
    n133,
    n29
  );


  not
  g31
  (
    n38,
    n30
  );


  buf
  g32
  (
    n126,
    n6
  );


  buf
  g33
  (
    n98,
    n11
  );


  buf
  g34
  (
    n79,
    n28
  );


  buf
  g35
  (
    n36,
    n3
  );


  buf
  g36
  (
    n145,
    n25
  );


  not
  g37
  (
    n80,
    n23
  );


  buf
  g38
  (
    n149,
    n15
  );


  not
  g39
  (
    n134,
    n26
  );


  buf
  g40
  (
    n43,
    n25
  );


  not
  g41
  (
    n77,
    n26
  );


  not
  g42
  (
    n152,
    n27
  );


  buf
  g43
  (
    n55,
    n25
  );


  not
  g44
  (
    n143,
    n28
  );


  buf
  g45
  (
    n131,
    n21
  );


  not
  g46
  (
    n108,
    n21
  );


  not
  g47
  (
    n150,
    n23
  );


  buf
  g48
  (
    n70,
    n4
  );


  not
  g49
  (
    n53,
    n14
  );


  buf
  g50
  (
    n59,
    n23
  );


  not
  g51
  (
    n64,
    n14
  );


  buf
  g52
  (
    n72,
    n20
  );


  buf
  g53
  (
    n120,
    n17
  );


  buf
  g54
  (
    n119,
    n31
  );


  not
  g55
  (
    n37,
    n18
  );


  buf
  g56
  (
    n123,
    n30
  );


  not
  g57
  (
    n68,
    n7
  );


  buf
  g58
  (
    KeyWire_0_21,
    n1
  );


  buf
  g59
  (
    n140,
    n19
  );


  not
  g60
  (
    KeyWire_0_15,
    n20
  );


  buf
  g61
  (
    n88,
    n13
  );


  buf
  g62
  (
    n60,
    n18
  );


  buf
  g63
  (
    KeyWire_0_3,
    n10
  );


  buf
  g64
  (
    n46,
    n31
  );


  not
  g65
  (
    n35,
    n27
  );


  buf
  g66
  (
    n107,
    n15
  );


  not
  g67
  (
    n73,
    n29
  );


  buf
  g68
  (
    n121,
    n10
  );


  buf
  g69
  (
    n93,
    n7
  );


  not
  g70
  (
    n136,
    n12
  );


  buf
  g71
  (
    n97,
    n6
  );


  buf
  g72
  (
    n40,
    n32
  );


  buf
  g73
  (
    n139,
    n21
  );


  not
  g74
  (
    n51,
    n13
  );


  not
  g75
  (
    n122,
    n14
  );


  not
  g76
  (
    n81,
    n15
  );


  buf
  g77
  (
    n118,
    n7
  );


  not
  g78
  (
    n65,
    n9
  );


  not
  g79
  (
    n135,
    n15
  );


  not
  g80
  (
    n101,
    n25
  );


  not
  g81
  (
    n52,
    n5
  );


  buf
  g82
  (
    n137,
    n12
  );


  buf
  g83
  (
    n117,
    n8
  );


  not
  g84
  (
    n91,
    n24
  );


  not
  g85
  (
    n63,
    n23
  );


  buf
  g86
  (
    n100,
    n26
  );


  not
  g87
  (
    n110,
    n32
  );


  not
  g88
  (
    n125,
    n16
  );


  buf
  g89
  (
    n39,
    n27
  );


  buf
  g90
  (
    n148,
    n18
  );


  buf
  g91
  (
    n33,
    n13
  );


  not
  g92
  (
    n111,
    n20
  );


  not
  g93
  (
    n62,
    n5
  );


  buf
  g94
  (
    n105,
    n31
  );


  not
  g95
  (
    n109,
    n32
  );


  buf
  g96
  (
    n106,
    n4
  );


  buf
  g97
  (
    n102,
    n3
  );


  not
  g98
  (
    n44,
    n5
  );


  not
  g99
  (
    n34,
    n30
  );


  not
  g100
  (
    n50,
    n9
  );


  not
  g101
  (
    n144,
    n8
  );


  buf
  g102
  (
    n71,
    n19
  );


  buf
  g103
  (
    n61,
    n16
  );


  not
  g104
  (
    n90,
    n32
  );


  not
  g105
  (
    n85,
    n21
  );


  buf
  g106
  (
    n151,
    n28
  );


  buf
  g107
  (
    n41,
    n19
  );


  buf
  g108
  (
    n113,
    n16
  );


  not
  g109
  (
    n58,
    n6
  );


  buf
  g110
  (
    n104,
    n9
  );


  not
  g111
  (
    n128,
    n24
  );


  not
  g112
  (
    n83,
    n8
  );


  buf
  g113
  (
    n66,
    n20
  );


  not
  g114
  (
    n112,
    n31
  );


  buf
  g115
  (
    n82,
    n14
  );


  not
  g116
  (
    n99,
    n24
  );


  buf
  g117
  (
    n48,
    n19
  );


  not
  g118
  (
    n87,
    n6
  );


  not
  g119
  (
    n76,
    n4
  );


  not
  g120
  (
    n179,
    n89
  );


  not
  g121
  (
    n260,
    n95
  );


  not
  g122
  (
    n383,
    n73
  );


  not
  g123
  (
    n164,
    n112
  );


  not
  g124
  (
    n173,
    n62
  );


  not
  g125
  (
    n344,
    n102
  );


  not
  g126
  (
    n219,
    n101
  );


  buf
  g127
  (
    n284,
    n62
  );


  buf
  g128
  (
    n285,
    n74
  );


  buf
  g129
  (
    n154,
    n110
  );


  buf
  g130
  (
    n255,
    n146
  );


  buf
  g131
  (
    n238,
    n113
  );


  buf
  g132
  (
    n340,
    n123
  );


  not
  g133
  (
    n155,
    n51
  );


  not
  g134
  (
    n321,
    n94
  );


  buf
  g135
  (
    n312,
    n108
  );


  not
  g136
  (
    n362,
    n56
  );


  buf
  g137
  (
    n210,
    n64
  );


  buf
  g138
  (
    n246,
    n89
  );


  buf
  g139
  (
    n262,
    n76
  );


  not
  g140
  (
    n264,
    n107
  );


  not
  g141
  (
    n370,
    n58
  );


  not
  g142
  (
    n190,
    n59
  );


  buf
  g143
  (
    n395,
    n33
  );


  nand
  g144
  (
    n266,
    n59,
    n111
  );


  nor
  g145
  (
    n314,
    n101,
    n66
  );


  or
  g146
  (
    n298,
    n67,
    n88
  );


  and
  g147
  (
    n328,
    n143,
    n148
  );


  or
  g148
  (
    n365,
    n37,
    n45
  );


  xnor
  g149
  (
    n191,
    n121,
    n72
  );


  xnor
  g150
  (
    n270,
    n48,
    n121
  );


  or
  g151
  (
    n300,
    n60,
    n120
  );


  xor
  g152
  (
    n239,
    n47,
    n121
  );


  nand
  g153
  (
    n189,
    n122,
    n86
  );


  or
  g154
  (
    n243,
    n135,
    n110
  );


  or
  g155
  (
    n261,
    n128,
    n132
  );


  xnor
  g156
  (
    n332,
    n72,
    n51
  );


  or
  g157
  (
    n160,
    n76,
    n115
  );


  nor
  g158
  (
    n311,
    n66,
    n74
  );


  and
  g159
  (
    n318,
    n130,
    n143
  );


  xnor
  g160
  (
    n221,
    n49,
    n129
  );


  nand
  g161
  (
    n323,
    n97,
    n55
  );


  or
  g162
  (
    KeyWire_0_17,
    n34,
    n112
  );


  or
  g163
  (
    n306,
    n56,
    n35
  );


  or
  g164
  (
    n237,
    n90,
    n92
  );


  nand
  g165
  (
    n315,
    n82,
    n41
  );


  xor
  g166
  (
    n329,
    n34,
    n96
  );


  nand
  g167
  (
    n186,
    n43,
    n94
  );


  xor
  g168
  (
    n276,
    n62,
    n143
  );


  or
  g169
  (
    n334,
    n71,
    n108
  );


  xor
  g170
  (
    n265,
    n88,
    n147
  );


  nand
  g171
  (
    n220,
    n136,
    n67
  );


  and
  g172
  (
    n163,
    n87,
    n146
  );


  or
  g173
  (
    n387,
    n61,
    n68
  );


  or
  g174
  (
    n172,
    n78,
    n142
  );


  xnor
  g175
  (
    n282,
    n40,
    n65
  );


  nor
  g176
  (
    n162,
    n58,
    n122
  );


  or
  g177
  (
    n401,
    n52,
    n114
  );


  xnor
  g178
  (
    n380,
    n71,
    n136
  );


  xnor
  g179
  (
    n386,
    n59,
    n50
  );


  nor
  g180
  (
    n388,
    n69,
    n80
  );


  and
  g181
  (
    n215,
    n55,
    n111
  );


  or
  g182
  (
    n229,
    n106,
    n45
  );


  nand
  g183
  (
    n242,
    n130,
    n53
  );


  or
  g184
  (
    n302,
    n68,
    n111
  );


  xnor
  g185
  (
    n212,
    n59,
    n66
  );


  nor
  g186
  (
    n377,
    n70,
    n97
  );


  nand
  g187
  (
    n288,
    n91,
    n102
  );


  and
  g188
  (
    n356,
    n149,
    n132
  );


  and
  g189
  (
    n308,
    n41,
    n123
  );


  xor
  g190
  (
    n222,
    n106,
    n91
  );


  or
  g191
  (
    n198,
    n83,
    n58
  );


  and
  g192
  (
    n252,
    n127,
    n114
  );


  or
  g193
  (
    n287,
    n37,
    n75
  );


  or
  g194
  (
    n345,
    n116,
    n151
  );


  and
  g195
  (
    n274,
    n77,
    n36
  );


  nor
  g196
  (
    n398,
    n80,
    n108
  );


  nor
  g197
  (
    n223,
    n125,
    n110
  );


  nor
  g198
  (
    n165,
    n105,
    n45
  );


  nand
  g199
  (
    n289,
    n103,
    n50
  );


  xnor
  g200
  (
    n317,
    n131,
    n79
  );


  nand
  g201
  (
    n389,
    n139,
    n83
  );


  or
  g202
  (
    n382,
    n65,
    n78
  );


  xnor
  g203
  (
    n159,
    n57,
    n98
  );


  nor
  g204
  (
    n211,
    n109,
    n81
  );


  xnor
  g205
  (
    n241,
    n85,
    n52
  );


  and
  g206
  (
    n180,
    n105,
    n92
  );


  nor
  g207
  (
    n218,
    n126,
    n137
  );


  xnor
  g208
  (
    n374,
    n145,
    n134
  );


  and
  g209
  (
    n158,
    n116,
    n44
  );


  xor
  g210
  (
    n205,
    n100,
    n144
  );


  not
  g211
  (
    n203,
    n93
  );


  nor
  g212
  (
    n326,
    n88,
    n130
  );


  nand
  g213
  (
    n225,
    n63,
    n141
  );


  nand
  g214
  (
    n336,
    n90,
    n82
  );


  xor
  g215
  (
    n235,
    n131,
    n40
  );


  or
  g216
  (
    n337,
    n112,
    n101
  );


  nand
  g217
  (
    n299,
    n99,
    n55
  );


  and
  g218
  (
    n293,
    n36,
    n77
  );


  nand
  g219
  (
    n197,
    n73,
    n135
  );


  and
  g220
  (
    n355,
    n117,
    n124
  );


  nand
  g221
  (
    n316,
    n115,
    n127
  );


  nand
  g222
  (
    n335,
    n70,
    n60
  );


  xor
  g223
  (
    n240,
    n150,
    n86
  );


  and
  g224
  (
    n324,
    n142,
    n102
  );


  and
  g225
  (
    n319,
    n146,
    n42
  );


  nand
  g226
  (
    n368,
    n80,
    n120
  );


  or
  g227
  (
    n167,
    n151,
    n115
  );


  and
  g228
  (
    n204,
    n66,
    n63
  );


  xor
  g229
  (
    n250,
    n144,
    n94
  );


  nor
  g230
  (
    n343,
    n133,
    n37
  );


  nor
  g231
  (
    n402,
    n133,
    n87
  );


  xnor
  g232
  (
    n350,
    n63,
    n126
  );


  nor
  g233
  (
    n193,
    n88,
    n137
  );


  xor
  g234
  (
    n292,
    n57,
    n95
  );


  or
  g235
  (
    n322,
    n84,
    n141
  );


  xor
  g236
  (
    n258,
    n49,
    n103
  );


  nand
  g237
  (
    n283,
    n75,
    n45
  );


  and
  g238
  (
    n202,
    n57,
    n52
  );


  or
  g239
  (
    KeyWire_0_10,
    n81,
    n86
  );


  xnor
  g240
  (
    n177,
    n85,
    n99
  );


  nor
  g241
  (
    n303,
    n106,
    n128
  );


  nor
  g242
  (
    n233,
    n43,
    n56
  );


  xnor
  g243
  (
    n245,
    n94,
    n69
  );


  and
  g244
  (
    n174,
    n140,
    n50
  );


  or
  g245
  (
    n267,
    n62,
    n64
  );


  and
  g246
  (
    n347,
    n122,
    n150
  );


  and
  g247
  (
    n339,
    n102,
    n104
  );


  nor
  g248
  (
    n330,
    n68,
    n125
  );


  and
  g249
  (
    n175,
    n70,
    n101
  );


  or
  g250
  (
    n301,
    n107,
    n91
  );


  xor
  g251
  (
    n206,
    n141,
    n119
  );


  xor
  g252
  (
    n279,
    n53,
    n71
  );


  nor
  g253
  (
    n184,
    n97,
    n36
  );


  xor
  g254
  (
    n397,
    n49,
    n64
  );


  or
  g255
  (
    n178,
    n98,
    n119
  );


  and
  g256
  (
    n181,
    n149,
    n93
  );


  nand
  g257
  (
    n351,
    n37,
    n46
  );


  or
  g258
  (
    n170,
    n131,
    n68
  );


  nand
  g259
  (
    n269,
    n65,
    n44
  );


  xnor
  g260
  (
    n183,
    n141,
    n70
  );


  xor
  g261
  (
    n304,
    n137,
    n114
  );


  xor
  g262
  (
    n227,
    n96,
    n69
  );


  xor
  g263
  (
    n349,
    n138,
    n150
  );


  xnor
  g264
  (
    n320,
    n149,
    n33
  );


  xor
  g265
  (
    n358,
    n125,
    n111
  );


  xnor
  g266
  (
    n352,
    n95,
    n118
  );


  nor
  g267
  (
    KeyWire_0_27,
    n71,
    n73
  );


  nor
  g268
  (
    n157,
    n124,
    n82
  );


  xnor
  g269
  (
    n376,
    n130,
    n43
  );


  nor
  g270
  (
    n259,
    n44,
    n80
  );


  nor
  g271
  (
    n373,
    n108,
    n72
  );


  xnor
  g272
  (
    n272,
    n110,
    n41
  );


  and
  g273
  (
    n313,
    n51,
    n46
  );


  nand
  g274
  (
    n232,
    n61,
    n40
  );


  or
  g275
  (
    n153,
    n82,
    n92
  );


  nand
  g276
  (
    n369,
    n135,
    n63
  );


  nand
  g277
  (
    n213,
    n134,
    n119
  );


  xnor
  g278
  (
    n208,
    n148,
    n136
  );


  xor
  g279
  (
    n224,
    n87,
    n81
  );


  and
  g280
  (
    n278,
    n90,
    n120
  );


  nor
  g281
  (
    n400,
    n127,
    n128
  );


  or
  g282
  (
    n357,
    n128,
    n73
  );


  nor
  g283
  (
    n348,
    n96,
    n142
  );


  or
  g284
  (
    n294,
    n91,
    n76
  );


  nand
  g285
  (
    n384,
    n61,
    n142
  );


  or
  g286
  (
    n214,
    n147,
    n145
  );


  xnor
  g287
  (
    n161,
    n123,
    n38
  );


  xnor
  g288
  (
    n359,
    n84,
    n116
  );


  and
  g289
  (
    n360,
    n54,
    n139
  );


  xnor
  g290
  (
    n354,
    n61,
    n47
  );


  nand
  g291
  (
    n333,
    n67,
    n75
  );


  xnor
  g292
  (
    n363,
    n85,
    n78
  );


  nand
  g293
  (
    n200,
    n72,
    n109
  );


  xnor
  g294
  (
    n196,
    n127,
    n104
  );


  xnor
  g295
  (
    n207,
    n124,
    n58
  );


  and
  g296
  (
    KeyWire_0_9,
    n107,
    n99
  );


  xnor
  g297
  (
    n361,
    n148,
    n123
  );


  or
  g298
  (
    n367,
    n129,
    n47
  );


  and
  g299
  (
    n230,
    n126,
    n55
  );


  xnor
  g300
  (
    n234,
    n122,
    n50
  );


  and
  g301
  (
    n166,
    n99,
    n98
  );


  xor
  g302
  (
    n277,
    n115,
    n51
  );


  xor
  g303
  (
    n257,
    n118,
    n147
  );


  nand
  g304
  (
    n309,
    n98,
    n34
  );


  or
  g305
  (
    n256,
    n83,
    n42
  );


  and
  g306
  (
    n216,
    n57,
    n95
  );


  and
  g307
  (
    n201,
    n133,
    n126
  );


  xor
  g308
  (
    KeyWire_0_1,
    n151,
    n138
  );


  xnor
  g309
  (
    n271,
    n42,
    n75
  );


  and
  g310
  (
    n192,
    n100,
    n77
  );


  xnor
  g311
  (
    n195,
    n39,
    n113
  );


  xnor
  g312
  (
    n226,
    n105,
    n76
  );


  nor
  g313
  (
    n194,
    n109,
    n52
  );


  nor
  g314
  (
    n391,
    n113,
    n140
  );


  and
  g315
  (
    n372,
    n41,
    n103
  );


  xnor
  g316
  (
    n392,
    n48,
    n113
  );


  nand
  g317
  (
    n378,
    n140,
    n134
  );


  nand
  g318
  (
    n342,
    n43,
    n38
  );


  nand
  g319
  (
    n156,
    n129,
    n100
  );


  nand
  g320
  (
    n251,
    n105,
    n118
  );


  nor
  g321
  (
    n393,
    n145,
    n60
  );


  and
  g322
  (
    n281,
    n106,
    n53
  );


  nand
  g323
  (
    n366,
    n146,
    n84
  );


  nor
  g324
  (
    n396,
    n46,
    n74
  );


  xnor
  g325
  (
    n295,
    n116,
    n87
  );


  nand
  g326
  (
    n254,
    n65,
    n33
  );


  nand
  g327
  (
    n297,
    n89,
    n56
  );


  and
  g328
  (
    n280,
    n84,
    n107
  );


  or
  g329
  (
    n346,
    n39,
    n133
  );


  and
  g330
  (
    n390,
    n46,
    n93
  );


  xnor
  g331
  (
    n249,
    n34,
    n143
  );


  nand
  g332
  (
    n375,
    n54,
    n35
  );


  xor
  g333
  (
    n244,
    n54,
    n42
  );


  or
  g334
  (
    n247,
    n117,
    n145
  );


  or
  g335
  (
    n185,
    n38,
    n35
  );


  nand
  g336
  (
    n291,
    n147,
    n83
  );


  nor
  g337
  (
    n381,
    n124,
    n119
  );


  or
  g338
  (
    n379,
    n79,
    n104
  );


  or
  g339
  (
    n305,
    n92,
    n137
  );


  xnor
  g340
  (
    n325,
    n139,
    n39
  );


  or
  g341
  (
    n385,
    n117,
    n33
  );


  xor
  g342
  (
    n327,
    n79,
    n74
  );


  xnor
  g343
  (
    n307,
    n49,
    n148
  );


  nor
  g344
  (
    n187,
    n103,
    n90
  );


  xnor
  g345
  (
    n399,
    n138,
    n79
  );


  nand
  g346
  (
    n171,
    n38,
    n89
  );


  nor
  g347
  (
    n253,
    n81,
    n64
  );


  xor
  g348
  (
    n394,
    n53,
    n60
  );


  and
  g349
  (
    n248,
    n132,
    n96
  );


  nand
  g350
  (
    n209,
    n44,
    n135
  );


  xor
  g351
  (
    KeyWire_0_26,
    n85,
    n131
  );


  xor
  g352
  (
    n182,
    n39,
    n97
  );


  xnor
  g353
  (
    n275,
    n77,
    n112
  );


  and
  g354
  (
    n217,
    n36,
    n48
  );


  xnor
  g355
  (
    KeyWire_0_0,
    n78,
    n140
  );


  nand
  g356
  (
    n310,
    n136,
    n86
  );


  xor
  g357
  (
    n199,
    n139,
    n48
  );


  xor
  g358
  (
    n188,
    n129,
    n132
  );


  xor
  g359
  (
    n290,
    n117,
    n149
  );


  xor
  g360
  (
    n236,
    n104,
    n144
  );


  nor
  g361
  (
    n231,
    n47,
    n118
  );


  xor
  g362
  (
    n168,
    n150,
    n69
  );


  xnor
  g363
  (
    n364,
    n54,
    n109
  );


  nor
  g364
  (
    n341,
    n114,
    n100
  );


  nand
  g365
  (
    n228,
    n138,
    n67
  );


  xnor
  g366
  (
    n371,
    n35,
    n125
  );


  xnor
  g367
  (
    n338,
    n144,
    n40
  );


  nand
  g368
  (
    n331,
    n151,
    n120
  );


  nand
  g369
  (
    n268,
    n121,
    n134
  );


  not
  g370
  (
    n451,
    n221
  );


  buf
  g371
  (
    n438,
    n160
  );


  buf
  g372
  (
    n413,
    n197
  );


  buf
  g373
  (
    n426,
    n198
  );


  not
  g374
  (
    n425,
    n204
  );


  not
  g375
  (
    n414,
    n225
  );


  buf
  g376
  (
    n422,
    n153
  );


  not
  g377
  (
    n431,
    n170
  );


  not
  g378
  (
    n472,
    n173
  );


  not
  g379
  (
    n416,
    n213
  );


  buf
  g380
  (
    n474,
    n186
  );


  buf
  g381
  (
    n418,
    n176
  );


  buf
  g382
  (
    n454,
    n214
  );


  not
  g383
  (
    n432,
    n169
  );


  not
  g384
  (
    n444,
    n187
  );


  not
  g385
  (
    n427,
    n162
  );


  buf
  g386
  (
    n450,
    n167
  );


  buf
  g387
  (
    KeyWire_0_5,
    n201
  );


  buf
  g388
  (
    n421,
    n179
  );


  not
  g389
  (
    n423,
    n157
  );


  buf
  g390
  (
    n436,
    n181
  );


  buf
  g391
  (
    n405,
    n164
  );


  not
  g392
  (
    n437,
    n180
  );


  not
  g393
  (
    n419,
    n163
  );


  not
  g394
  (
    n466,
    n191
  );


  buf
  g395
  (
    n430,
    n206
  );


  buf
  g396
  (
    n448,
    n215
  );


  buf
  g397
  (
    n462,
    n210
  );


  not
  g398
  (
    n420,
    n168
  );


  buf
  g399
  (
    n409,
    n158
  );


  buf
  g400
  (
    n441,
    n183
  );


  not
  g401
  (
    n467,
    n207
  );


  not
  g402
  (
    n445,
    n203
  );


  buf
  g403
  (
    n424,
    n175
  );


  not
  g404
  (
    n461,
    n217
  );


  not
  g405
  (
    n407,
    n216
  );


  buf
  g406
  (
    n410,
    n202
  );


  not
  g407
  (
    n458,
    n205
  );


  buf
  g408
  (
    n452,
    n209
  );


  buf
  g409
  (
    n459,
    n190
  );


  buf
  g410
  (
    n456,
    n196
  );


  not
  g411
  (
    n417,
    n159
  );


  buf
  g412
  (
    n428,
    n154
  );


  buf
  g413
  (
    n476,
    n165
  );


  not
  g414
  (
    n475,
    n184
  );


  not
  g415
  (
    n457,
    n219
  );


  not
  g416
  (
    n435,
    n194
  );


  not
  g417
  (
    n442,
    n223
  );


  buf
  g418
  (
    n411,
    n222
  );


  not
  g419
  (
    n465,
    n182
  );


  not
  g420
  (
    n446,
    n193
  );


  not
  g421
  (
    n455,
    n166
  );


  buf
  g422
  (
    n447,
    n174
  );


  buf
  g423
  (
    n406,
    n200
  );


  not
  g424
  (
    n433,
    n226
  );


  buf
  g425
  (
    n440,
    n171
  );


  not
  g426
  (
    n412,
    n155
  );


  not
  g427
  (
    n471,
    n185
  );


  buf
  g428
  (
    n429,
    n211
  );


  not
  g429
  (
    n460,
    n177
  );


  buf
  g430
  (
    n408,
    n172
  );


  not
  g431
  (
    n464,
    n195
  );


  not
  g432
  (
    n473,
    n192
  );


  not
  g433
  (
    n434,
    n188
  );


  not
  g434
  (
    n415,
    n220
  );


  not
  g435
  (
    KeyWire_0_20,
    n212
  );


  buf
  g436
  (
    n404,
    n189
  );


  not
  g437
  (
    n453,
    n178
  );


  not
  g438
  (
    n449,
    n161
  );


  buf
  g439
  (
    n468,
    n208
  );


  buf
  g440
  (
    n463,
    n156
  );


  buf
  g441
  (
    n470,
    n224
  );


  buf
  g442
  (
    n469,
    n218
  );


  not
  g443
  (
    n443,
    n199
  );


  not
  g444
  (
    n483,
    n407
  );


  buf
  g445
  (
    n486,
    n411
  );


  buf
  g446
  (
    n478,
    n405
  );


  not
  g447
  (
    n487,
    n406
  );


  not
  g448
  (
    n489,
    n408
  );


  buf
  g449
  (
    n477,
    n406
  );


  not
  g450
  (
    n485,
    n408
  );


  not
  g451
  (
    n480,
    n407
  );


  xor
  g452
  (
    n484,
    n407,
    n409,
    n411,
    n410
  );


  or
  g453
  (
    n479,
    n410,
    n410,
    n406,
    n412
  );


  nor
  g454
  (
    n488,
    n407,
    n404,
    n411,
    n406
  );


  xor
  g455
  (
    n482,
    n410,
    n408,
    n409
  );


  and
  g456
  (
    n481,
    n408,
    n403,
    n411,
    n409
  );


  buf
  g457
  (
    n507,
    n412
  );


  buf
  g458
  (
    n517,
    n486
  );


  not
  g459
  (
    n516,
    n421
  );


  buf
  g460
  (
    n513,
    n413
  );


  not
  g461
  (
    n529,
    n480
  );


  buf
  g462
  (
    n537,
    n426
  );


  xnor
  g463
  (
    n505,
    n238,
    n417,
    n237,
    n419
  );


  xor
  g464
  (
    n522,
    n481,
    n423,
    n436,
    n418
  );


  xor
  g465
  (
    n526,
    n482,
    n419,
    n415,
    n424
  );


  or
  g466
  (
    n532,
    n412,
    n487,
    n488
  );


  xor
  g467
  (
    n515,
    n421,
    n433,
    n479,
    n480
  );


  xnor
  g468
  (
    n512,
    n432,
    n489,
    n416
  );


  or
  g469
  (
    n509,
    n424,
    n486,
    n484,
    n436
  );


  xnor
  g470
  (
    n500,
    n485,
    n485,
    n420,
    n486
  );


  xor
  g471
  (
    n496,
    n426,
    n248,
    n425,
    n483
  );


  and
  g472
  (
    n534,
    n414,
    n429,
    n427,
    n477
  );


  and
  g473
  (
    n504,
    n481,
    n152,
    n229,
    n484
  );


  nand
  g474
  (
    n535,
    n489,
    n488,
    n228,
    n425
  );


  nand
  g475
  (
    n511,
    n489,
    n414,
    n484,
    n428
  );


  xnor
  g476
  (
    n521,
    n245,
    n431,
    n428,
    n417
  );


  and
  g477
  (
    n519,
    n435,
    n435,
    n233,
    n420
  );


  nor
  g478
  (
    KeyWire_0_18,
    n414,
    n421,
    n422,
    n435
  );


  xor
  g479
  (
    n530,
    n488,
    n422,
    n478,
    n427
  );


  xor
  g480
  (
    n523,
    n418,
    n486,
    n428,
    n480
  );


  and
  g481
  (
    n518,
    n425,
    n434,
    n485,
    n423
  );


  nor
  g482
  (
    n527,
    n244,
    n426,
    n412,
    n418
  );


  xor
  g483
  (
    n502,
    n247,
    n433,
    n485
  );


  nand
  g484
  (
    n498,
    n246,
    n413,
    n487,
    n436
  );


  xnor
  g485
  (
    n495,
    n249,
    n251,
    n428,
    n423
  );


  nand
  g486
  (
    n531,
    n418,
    n416,
    n227,
    n417
  );


  nand
  g487
  (
    n490,
    n416,
    n419,
    n488,
    n480
  );


  and
  g488
  (
    n533,
    n419,
    n427,
    n478,
    n482
  );


  or
  g489
  (
    n528,
    n234,
    n422,
    n243,
    n430
  );


  and
  g490
  (
    n525,
    n414,
    n252,
    n417,
    n482
  );


  nand
  g491
  (
    n499,
    n477,
    n483,
    n429
  );


  or
  g492
  (
    n508,
    n427,
    n432,
    n424,
    n434
  );


  or
  g493
  (
    n506,
    n432,
    n483,
    n230,
    n433
  );


  or
  g494
  (
    n493,
    n239,
    n436,
    n434,
    n240
  );


  xor
  g495
  (
    KeyWire_0_22,
    n479,
    n421,
    n484,
    n481
  );


  nor
  g496
  (
    n497,
    n434,
    n241,
    n425,
    n242
  );


  xor
  g497
  (
    n503,
    n250,
    n431,
    n432,
    n435
  );


  nor
  g498
  (
    n514,
    n420,
    n430,
    n232,
    n415
  );


  xnor
  g499
  (
    n501,
    n415,
    n426,
    n431
  );


  and
  g500
  (
    n510,
    n235,
    n479,
    n482,
    n422
  );


  nor
  g501
  (
    n492,
    n424,
    n231,
    n416,
    n236
  );


  and
  g502
  (
    n536,
    n430,
    n481,
    n429,
    n413
  );


  and
  g503
  (
    n524,
    n430,
    n429,
    n413,
    n415
  );


  xnor
  g504
  (
    n491,
    n423,
    n479,
    n487,
    n420
  );


  buf
  g505
  (
    n722,
    n504
  );


  not
  g506
  (
    n574,
    n491
  );


  not
  g507
  (
    n668,
    n501
  );


  buf
  g508
  (
    n554,
    n527
  );


  buf
  g509
  (
    KeyWire_0_23,
    n506
  );


  not
  g510
  (
    n569,
    n529
  );


  buf
  g511
  (
    n548,
    n532
  );


  buf
  g512
  (
    n589,
    n503
  );


  not
  g513
  (
    n539,
    n523
  );


  not
  g514
  (
    n547,
    n493
  );


  not
  g515
  (
    n670,
    n508
  );


  not
  g516
  (
    n540,
    n493
  );


  buf
  g517
  (
    n665,
    n496
  );


  not
  g518
  (
    n584,
    n509
  );


  buf
  g519
  (
    n612,
    n520
  );


  not
  g520
  (
    n549,
    n507
  );


  buf
  g521
  (
    n608,
    n532
  );


  not
  g522
  (
    n557,
    n505
  );


  buf
  g523
  (
    n633,
    n530
  );


  not
  g524
  (
    n568,
    n490
  );


  not
  g525
  (
    n630,
    n528
  );


  not
  g526
  (
    n685,
    n523
  );


  not
  g527
  (
    n694,
    n507
  );


  buf
  g528
  (
    n626,
    n508
  );


  buf
  g529
  (
    n690,
    n280
  );


  buf
  g530
  (
    n669,
    n520
  );


  buf
  g531
  (
    n648,
    n511
  );


  buf
  g532
  (
    n708,
    n279
  );


  not
  g533
  (
    n662,
    n271
  );


  not
  g534
  (
    n651,
    n536
  );


  buf
  g535
  (
    n622,
    n510
  );


  buf
  g536
  (
    n700,
    n506
  );


  not
  g537
  (
    n678,
    n518
  );


  not
  g538
  (
    n611,
    n491
  );


  buf
  g539
  (
    n601,
    n520
  );


  buf
  g540
  (
    n570,
    n268
  );


  buf
  g541
  (
    n596,
    n522
  );


  not
  g542
  (
    n564,
    n535
  );


  buf
  g543
  (
    n663,
    n272
  );


  buf
  g544
  (
    n684,
    n508
  );


  not
  g545
  (
    n620,
    n533
  );


  not
  g546
  (
    n543,
    n535
  );


  buf
  g547
  (
    n573,
    n517
  );


  buf
  g548
  (
    n604,
    n524
  );


  buf
  g549
  (
    n562,
    n498
  );


  buf
  g550
  (
    n621,
    n495
  );


  buf
  g551
  (
    n666,
    n497
  );


  buf
  g552
  (
    n565,
    n257
  );


  buf
  g553
  (
    n591,
    n529
  );


  not
  g554
  (
    n642,
    n269
  );


  not
  g555
  (
    n718,
    n531
  );


  buf
  g556
  (
    n671,
    n502
  );


  buf
  g557
  (
    n649,
    n529
  );


  buf
  g558
  (
    n687,
    n513
  );


  not
  g559
  (
    n638,
    n511
  );


  buf
  g560
  (
    n542,
    n260
  );


  buf
  g561
  (
    n639,
    n267
  );


  not
  g562
  (
    n624,
    n496
  );


  buf
  g563
  (
    n587,
    n516
  );


  not
  g564
  (
    n593,
    n505
  );


  buf
  g565
  (
    n640,
    n526
  );


  buf
  g566
  (
    n681,
    n521
  );


  buf
  g567
  (
    n585,
    n492
  );


  not
  g568
  (
    n616,
    n491
  );


  buf
  g569
  (
    n652,
    n531
  );


  not
  g570
  (
    n724,
    n516
  );


  buf
  g571
  (
    n541,
    n497
  );


  buf
  g572
  (
    n650,
    n518
  );


  buf
  g573
  (
    n660,
    n494
  );


  buf
  g574
  (
    n689,
    n492
  );


  not
  g575
  (
    n546,
    n528
  );


  not
  g576
  (
    n698,
    n490
  );


  buf
  g577
  (
    n688,
    n525
  );


  buf
  g578
  (
    n628,
    n528
  );


  buf
  g579
  (
    n632,
    n518
  );


  buf
  g580
  (
    n701,
    n502
  );


  not
  g581
  (
    n605,
    n513
  );


  not
  g582
  (
    n590,
    n522
  );


  not
  g583
  (
    n713,
    n255
  );


  buf
  g584
  (
    n682,
    n525
  );


  buf
  g585
  (
    n706,
    n521
  );


  buf
  g586
  (
    n653,
    n525
  );


  buf
  g587
  (
    n710,
    n262
  );


  not
  g588
  (
    n545,
    n273
  );


  not
  g589
  (
    n641,
    n498
  );


  buf
  g590
  (
    n577,
    n504
  );


  not
  g591
  (
    n544,
    n265
  );


  buf
  g592
  (
    n625,
    n512
  );


  buf
  g593
  (
    n606,
    n518
  );


  buf
  g594
  (
    n656,
    n501
  );


  not
  g595
  (
    n563,
    n496
  );


  buf
  g596
  (
    n686,
    n499
  );


  not
  g597
  (
    n692,
    n278
  );


  buf
  g598
  (
    n711,
    n259
  );


  not
  g599
  (
    n594,
    n515
  );


  not
  g600
  (
    n643,
    n517
  );


  not
  g601
  (
    KeyWire_0_24,
    n514
  );


  buf
  g602
  (
    n646,
    n531
  );


  not
  g603
  (
    n552,
    n514
  );


  buf
  g604
  (
    n629,
    n515
  );


  not
  g605
  (
    n696,
    n508
  );


  not
  g606
  (
    KeyWire_0_19,
    n525
  );


  not
  g607
  (
    n721,
    n496
  );


  not
  g608
  (
    n615,
    n497
  );


  not
  g609
  (
    n558,
    n504
  );


  buf
  g610
  (
    n592,
    n515
  );


  buf
  g611
  (
    n725,
    n534
  );


  not
  g612
  (
    n726,
    n519
  );


  buf
  g613
  (
    n683,
    n522
  );


  not
  g614
  (
    n635,
    n254
  );


  not
  g615
  (
    n614,
    n516
  );


  buf
  g616
  (
    n575,
    n512
  );


  buf
  g617
  (
    n645,
    n261
  );


  not
  g618
  (
    n598,
    n494
  );


  buf
  g619
  (
    n695,
    n500
  );


  buf
  g620
  (
    n623,
    n524
  );


  buf
  g621
  (
    n659,
    n497
  );


  not
  g622
  (
    n561,
    n537
  );


  buf
  g623
  (
    n572,
    n274
  );


  not
  g624
  (
    n559,
    n523
  );


  not
  g625
  (
    n664,
    n530
  );


  not
  g626
  (
    n609,
    n506
  );


  buf
  g627
  (
    n667,
    n499
  );


  buf
  g628
  (
    n709,
    n534
  );


  not
  g629
  (
    n538,
    n510
  );


  not
  g630
  (
    n704,
    n490
  );


  buf
  g631
  (
    n673,
    n513
  );


  not
  g632
  (
    n567,
    n500
  );


  not
  g633
  (
    n550,
    n519
  );


  buf
  g634
  (
    n617,
    n529
  );


  not
  g635
  (
    n636,
    n526
  );


  buf
  g636
  (
    n714,
    n516
  );


  buf
  g637
  (
    n693,
    n513
  );


  buf
  g638
  (
    n716,
    n493
  );


  not
  g639
  (
    n644,
    n499
  );


  buf
  g640
  (
    n619,
    n498
  );


  buf
  g641
  (
    n566,
    n505
  );


  buf
  g642
  (
    n603,
    n534
  );


  buf
  g643
  (
    n560,
    n495
  );


  buf
  g644
  (
    n661,
    n491
  );


  not
  g645
  (
    n707,
    n527
  );


  buf
  g646
  (
    n679,
    n535
  );


  not
  g647
  (
    n719,
    n501
  );


  buf
  g648
  (
    n571,
    n498
  );


  not
  g649
  (
    n676,
    n517
  );


  buf
  g650
  (
    KeyWire_0_11,
    n521
  );


  buf
  g651
  (
    n600,
    n264
  );


  buf
  g652
  (
    n597,
    n532
  );


  not
  g653
  (
    n627,
    n519
  );


  not
  g654
  (
    n647,
    n505
  );


  buf
  g655
  (
    n578,
    n512
  );


  buf
  g656
  (
    n551,
    n536
  );


  not
  g657
  (
    n555,
    n503
  );


  buf
  g658
  (
    n580,
    n507
  );


  not
  g659
  (
    n631,
    n530
  );


  buf
  g660
  (
    n723,
    n526
  );


  not
  g661
  (
    n607,
    n500
  );


  buf
  g662
  (
    n715,
    n510
  );


  buf
  g663
  (
    n705,
    n507
  );


  not
  g664
  (
    n675,
    n526
  );


  not
  g665
  (
    n576,
    n256
  );


  not
  g666
  (
    n699,
    n276
  );


  buf
  g667
  (
    n720,
    n524
  );


  buf
  g668
  (
    n634,
    n506
  );


  buf
  g669
  (
    KeyWire_0_8,
    n537
  );


  not
  g670
  (
    n677,
    n527
  );


  buf
  g671
  (
    n702,
    n275
  );


  buf
  g672
  (
    n658,
    n532
  );


  not
  g673
  (
    n697,
    n501
  );


  buf
  g674
  (
    n581,
    n533
  );


  not
  g675
  (
    n637,
    n495
  );


  not
  g676
  (
    KeyWire_0_29,
    n509
  );


  buf
  g677
  (
    n618,
    n510
  );


  not
  g678
  (
    n672,
    n502
  );


  buf
  g679
  (
    n595,
    n492
  );


  not
  g680
  (
    n680,
    n490
  );


  buf
  g681
  (
    n613,
    n521
  );


  buf
  g682
  (
    n599,
    n527
  );


  not
  g683
  (
    n674,
    n509
  );


  buf
  g684
  (
    n717,
    n270
  );


  and
  g685
  (
    n582,
    n535,
    n533,
    n494,
    n523
  );


  and
  g686
  (
    n579,
    n536,
    n503,
    n504,
    n502
  );


  nand
  g687
  (
    n588,
    n277,
    n509,
    n524,
    n531
  );


  xnor
  g688
  (
    n657,
    n512,
    n537,
    n517,
    n495
  );


  nor
  g689
  (
    n610,
    n503,
    n514,
    n500,
    n253
  );


  xnor
  g690
  (
    n712,
    n492,
    n522,
    n494,
    n515
  );


  and
  g691
  (
    n691,
    n499,
    n534,
    n266,
    n530
  );


  or
  g692
  (
    n553,
    n511,
    n533,
    n493,
    n519
  );


  and
  g693
  (
    n727,
    n258,
    n514,
    n536,
    n263
  );


  and
  g694
  (
    n583,
    n537,
    n511,
    n528,
    n520
  );


  not
  g695
  (
    n729,
    n549
  );


  buf
  g696
  (
    n732,
    n552
  );


  buf
  g697
  (
    n736,
    n556
  );


  not
  g698
  (
    n733,
    n538
  );


  not
  g699
  (
    n737,
    n541
  );


  not
  g700
  (
    n734,
    n543
  );


  nor
  g701
  (
    n735,
    n544,
    n551
  );


  nand
  g702
  (
    n730,
    n554,
    n539,
    n545,
    n540
  );


  or
  g703
  (
    n728,
    n557,
    n548,
    n550,
    n546
  );


  or
  g704
  (
    n731,
    n547,
    n553,
    n555,
    n542
  );


  or
  g705
  (
    n765,
    n332,
    n737,
    n286,
    n307
  );


  or
  g706
  (
    n750,
    n350,
    n349,
    n354,
    n735
  );


  xnor
  g707
  (
    n761,
    n728,
    n734,
    n287
  );


  nor
  g708
  (
    n740,
    n734,
    n304,
    n320,
    n371
  );


  nor
  g709
  (
    n744,
    n361,
    n347,
    n336,
    n348
  );


  and
  g710
  (
    n749,
    n300,
    n322,
    n736,
    n297
  );


  nand
  g711
  (
    n746,
    n324,
    n352,
    n299,
    n306
  );


  xor
  g712
  (
    n755,
    n362,
    n729,
    n737,
    n334
  );


  or
  g713
  (
    n766,
    n285,
    n333,
    n335,
    n735
  );


  xor
  g714
  (
    n757,
    n732,
    n344,
    n338,
    n735
  );


  nor
  g715
  (
    n738,
    n730,
    n327,
    n311,
    n329
  );


  xnor
  g716
  (
    n764,
    n356,
    n302,
    n359,
    n736
  );


  nor
  g717
  (
    n751,
    n298,
    n737,
    n731,
    n357
  );


  xnor
  g718
  (
    n762,
    n340,
    n325,
    n305,
    n370
  );


  nand
  g719
  (
    n763,
    n345,
    n353,
    n737,
    n326
  );


  or
  g720
  (
    n754,
    n369,
    n346,
    n315,
    n317
  );


  nand
  g721
  (
    n760,
    n292,
    n343,
    n288,
    n731
  );


  nand
  g722
  (
    n753,
    n296,
    n732,
    n736
  );


  xnor
  g723
  (
    n758,
    n733,
    n733,
    n313,
    n365
  );


  nor
  g724
  (
    n739,
    n283,
    n337,
    n308,
    n293
  );


  nand
  g725
  (
    n767,
    n729,
    n323,
    n368,
    n316
  );


  and
  g726
  (
    n741,
    n331,
    n330,
    n366,
    n281
  );


  or
  g727
  (
    n768,
    n321,
    n314,
    n291,
    n733
  );


  nor
  g728
  (
    n759,
    n373,
    n355,
    n351,
    n310
  );


  or
  g729
  (
    n743,
    n364,
    n295,
    n318,
    n363
  );


  or
  g730
  (
    n747,
    n360,
    n358,
    n328,
    n309
  );


  xor
  g731
  (
    n756,
    n367,
    n736,
    n284,
    n303
  );


  nor
  g732
  (
    n745,
    n733,
    n290,
    n312,
    n339
  );


  nor
  g733
  (
    n742,
    n341,
    n735,
    n319,
    n301
  );


  xor
  g734
  (
    n748,
    n732,
    n282,
    n342,
    n289
  );


  nand
  g735
  (
    n752,
    n294,
    n730,
    n734,
    n372
  );


  or
  g736
  (
    n772,
    n446,
    n453,
    n377,
    n745
  );


  or
  g737
  (
    KeyWire_0_28,
    n452,
    n438,
    n448,
    n739
  );


  or
  g738
  (
    n784,
    n446,
    n449,
    n440,
    n445
  );


  nand
  g739
  (
    n792,
    n448,
    n743,
    n447,
    n378
  );


  or
  g740
  (
    n795,
    n437,
    n454,
    n739,
    n452
  );


  xnor
  g741
  (
    n770,
    n744,
    n376,
    n449,
    n444
  );


  nand
  g742
  (
    n791,
    n374,
    n441,
    n438,
    n739
  );


  nor
  g743
  (
    n783,
    n452,
    n438,
    n453,
    n441
  );


  nand
  g744
  (
    n771,
    n742,
    n450,
    n448,
    n440
  );


  xor
  g745
  (
    n779,
    n444,
    n447,
    n453,
    n742
  );


  xnor
  g746
  (
    n769,
    n437,
    n450,
    n740
  );


  nor
  g747
  (
    n776,
    n738,
    n437,
    n440
  );


  xnor
  g748
  (
    n782,
    n451,
    n449,
    n447,
    n443
  );


  and
  g749
  (
    n785,
    n741,
    n447,
    n445,
    n443
  );


  or
  g750
  (
    n793,
    n441,
    n385,
    n443,
    n375
  );


  and
  g751
  (
    n788,
    n740,
    n444,
    n446,
    n382
  );


  and
  g752
  (
    n774,
    n742,
    n450,
    n380,
    n744
  );


  or
  g753
  (
    n777,
    n741,
    n743
  );


  xnor
  g754
  (
    n786,
    n453,
    n448,
    n451,
    n438
  );


  nor
  g755
  (
    n787,
    n441,
    n744,
    n738,
    n379
  );


  xor
  g756
  (
    n778,
    n446,
    n442,
    n445
  );


  nand
  g757
  (
    n794,
    n449,
    n742,
    n443,
    n439
  );


  and
  g758
  (
    n790,
    n451,
    n451,
    n442,
    n439
  );


  nand
  g759
  (
    n773,
    n444,
    n383,
    n439,
    n381
  );


  xor
  g760
  (
    n789,
    n437,
    n744,
    n741,
    n450
  );


  xnor
  g761
  (
    n780,
    n740,
    n741,
    n442,
    n739
  );


  xor
  g762
  (
    n775,
    n384,
    n445,
    n452,
    n439
  );


  nand
  g763
  (
    n810,
    n458,
    n468,
    n466
  );


  and
  g764
  (
    n798,
    n785,
    n473,
    n787,
    n464
  );


  or
  g765
  (
    n818,
    n788,
    n459,
    n465,
    n457
  );


  and
  g766
  (
    n801,
    n779,
    n466,
    n467,
    n464
  );


  xor
  g767
  (
    n814,
    n463,
    n778,
    n771,
    n791
  );


  xor
  g768
  (
    n796,
    n471,
    n469,
    n472
  );


  xnor
  g769
  (
    n804,
    n465,
    n463,
    n795,
    n460
  );


  and
  g770
  (
    n817,
    n777,
    n792,
    n795,
    n774
  );


  nand
  g771
  (
    n816,
    n454,
    n468,
    n786,
    n461
  );


  and
  g772
  (
    n800,
    n456,
    n455,
    n458,
    n470
  );


  xnor
  g773
  (
    n797,
    n469,
    n454,
    n783,
    n471
  );


  or
  g774
  (
    n809,
    n457,
    n465,
    n784,
    n461
  );


  nor
  g775
  (
    n808,
    n462,
    n463,
    n459,
    n789
  );


  nand
  g776
  (
    n819,
    n459,
    n775,
    n474,
    n472
  );


  xor
  g777
  (
    n807,
    n473,
    n456,
    n455
  );


  or
  g778
  (
    n806,
    n460,
    n464,
    n472,
    n466
  );


  nand
  g779
  (
    n813,
    n776,
    n474,
    n458,
    n462
  );


  nor
  g780
  (
    n815,
    n464,
    n780,
    n456,
    n465
  );


  nand
  g781
  (
    n822,
    n458,
    n460,
    n461,
    n472
  );


  nand
  g782
  (
    n812,
    n454,
    n462,
    n794,
    n471
  );


  and
  g783
  (
    n803,
    n457,
    n460,
    n770,
    n470
  );


  xor
  g784
  (
    KeyWire_0_13,
    n456,
    n473,
    n463,
    n769
  );


  nand
  g785
  (
    n820,
    n474,
    n461,
    n470,
    n475
  );


  nor
  g786
  (
    n823,
    n467,
    n782,
    n790,
    n457
  );


  nor
  g787
  (
    n802,
    n471,
    n470,
    n459,
    n793
  );


  or
  g788
  (
    n805,
    n772,
    n468,
    n473,
    n462
  );


  nand
  g789
  (
    n799,
    n455,
    n469,
    n773,
    n466
  );


  xor
  g790
  (
    n821,
    n781,
    n467,
    n474
  );


  or
  g791
  (
    n860,
    n616,
    n823,
    n819,
    n797
  );


  nor
  g792
  (
    n850,
    n803,
    n640,
    n799,
    n587
  );


  xor
  g793
  (
    n854,
    n395,
    n397,
    n816,
    n613
  );


  and
  g794
  (
    n845,
    n819,
    n799,
    n572,
    n805
  );


  nand
  g795
  (
    n858,
    n589,
    n596,
    n391,
    n820
  );


  or
  g796
  (
    n855,
    n562,
    n625,
    n806,
    n624
  );


  xnor
  g797
  (
    n824,
    n558,
    n817,
    n626
  );


  and
  g798
  (
    n864,
    n817,
    n582,
    n563,
    n801
  );


  xnor
  g799
  (
    n867,
    n810,
    n817,
    n390,
    n623
  );


  xor
  g800
  (
    n829,
    n809,
    n819,
    n152,
    n642
  );


  nand
  g801
  (
    KeyWire_0_25,
    n588,
    n638,
    n636,
    n814
  );


  nand
  g802
  (
    n861,
    n823,
    n152,
    n811,
    n584
  );


  xor
  g803
  (
    n825,
    n823,
    n394,
    n821,
    n592
  );


  nand
  g804
  (
    n832,
    n614,
    n618,
    n807,
    n565
  );


  nand
  g805
  (
    n839,
    n561,
    n813,
    n602,
    n615
  );


  xnor
  g806
  (
    n843,
    n822,
    n822,
    n805,
    n601
  );


  nand
  g807
  (
    n848,
    n816,
    n804,
    n802,
    n396
  );


  or
  g808
  (
    n842,
    n617,
    n822,
    n569,
    n575
  );


  or
  g809
  (
    n833,
    n607,
    n566,
    n612,
    n632
  );


  and
  g810
  (
    n849,
    n392,
    n796,
    n627,
    n611
  );


  nand
  g811
  (
    n847,
    n637,
    n798,
    n593,
    n574
  );


  nor
  g812
  (
    n844,
    n567,
    n571,
    n821,
    n807
  );


  xor
  g813
  (
    n862,
    n585,
    n633,
    n820,
    n634
  );


  and
  g814
  (
    n840,
    n818,
    n819,
    n595,
    n578
  );


  nor
  g815
  (
    n827,
    n389,
    n604,
    n573,
    n619
  );


  or
  g816
  (
    n836,
    n641,
    n399,
    n622,
    n629
  );


  nor
  g817
  (
    n826,
    n610,
    n797,
    n631,
    n401
  );


  and
  g818
  (
    n834,
    n820,
    n796,
    n811,
    n598
  );


  and
  g819
  (
    n835,
    n815,
    n603,
    n818,
    n808
  );


  nor
  g820
  (
    n863,
    n398,
    n570,
    n630,
    n606
  );


  xor
  g821
  (
    n853,
    n798,
    n639,
    n560,
    n608
  );


  xnor
  g822
  (
    n841,
    n815,
    n821,
    n813,
    n393
  );


  or
  g823
  (
    n852,
    n152,
    n816,
    n820,
    n628
  );


  and
  g824
  (
    n851,
    n810,
    n590,
    n600,
    n581
  );


  nand
  g825
  (
    n830,
    n580,
    n801,
    n400,
    n591
  );


  or
  g826
  (
    n857,
    n559,
    n594,
    n586,
    n806
  );


  xor
  g827
  (
    n846,
    n800,
    n621,
    n568,
    n577
  );


  and
  g828
  (
    n866,
    n818,
    n386,
    n821,
    n803
  );


  nor
  g829
  (
    n837,
    n564,
    n814,
    n800,
    n597
  );


  or
  g830
  (
    n828,
    n605,
    n388,
    n808,
    n620
  );


  nor
  g831
  (
    n859,
    n579,
    n609,
    n809,
    n802
  );


  xnor
  g832
  (
    n865,
    n804,
    n823,
    n387,
    n635
  );


  or
  g833
  (
    n831,
    n599,
    n822,
    n816,
    n576
  );


  or
  g834
  (
    n838,
    n812,
    n812,
    n583,
    n818
  );


  nand
  g835
  (
    n881,
    n657,
    n662,
    n862,
    n824
  );


  xor
  g836
  (
    n879,
    n836,
    n643,
    n847,
    n645
  );


  xor
  g837
  (
    n875,
    n651,
    n835,
    n656,
    n664
  );


  xnor
  g838
  (
    n868,
    n666,
    n661,
    n828,
    n648
  );


  and
  g839
  (
    n877,
    n653,
    n867,
    n854,
    n826
  );


  xnor
  g840
  (
    n882,
    n860,
    n848,
    n866,
    n838
  );


  xor
  g841
  (
    n880,
    n840,
    n863,
    n861,
    n853
  );


  xor
  g842
  (
    n878,
    n659,
    n856,
    n844,
    n647
  );


  and
  g843
  (
    n876,
    n649,
    n845,
    n846,
    n834
  );


  xnor
  g844
  (
    n873,
    n850,
    n831,
    n829,
    n652
  );


  and
  g845
  (
    n874,
    n663,
    n833,
    n660,
    n841
  );


  nand
  g846
  (
    n871,
    n864,
    n855,
    n830,
    n832
  );


  or
  g847
  (
    n872,
    n858,
    n843,
    n655,
    n842
  );


  or
  g848
  (
    n870,
    n865,
    n644,
    n654,
    n825
  );


  xnor
  g849
  (
    n883,
    n857,
    n839,
    n837,
    n665
  );


  xor
  g850
  (
    n884,
    n658,
    n851,
    n859,
    n827
  );


  nand
  g851
  (
    n869,
    n650,
    n646,
    n849,
    n852
  );


  not
  g852
  (
    n919,
    n701
  );


  not
  g853
  (
    n888,
    n879
  );


  not
  g854
  (
    n917,
    n710
  );


  buf
  g855
  (
    n902,
    n869
  );


  buf
  g856
  (
    n885,
    n672
  );


  not
  g857
  (
    n901,
    n876
  );


  not
  g858
  (
    n892,
    n714
  );


  not
  g859
  (
    n886,
    n713
  );


  buf
  g860
  (
    n910,
    n693
  );


  not
  g861
  (
    n893,
    n667
  );


  not
  g862
  (
    n904,
    n880
  );


  buf
  g863
  (
    n908,
    n709
  );


  buf
  g864
  (
    n906,
    n871
  );


  buf
  g865
  (
    n891,
    n671
  );


  buf
  g866
  (
    n914,
    n706
  );


  buf
  g867
  (
    n918,
    n694
  );


  buf
  g868
  (
    n907,
    n712
  );


  not
  g869
  (
    n921,
    n687
  );


  not
  g870
  (
    n916,
    n689
  );


  nor
  g871
  (
    n915,
    n675,
    n878,
    n677
  );


  nand
  g872
  (
    n911,
    n875,
    n673,
    n871,
    n874
  );


  xor
  g873
  (
    n895,
    n692,
    n878,
    n880,
    n708
  );


  xnor
  g874
  (
    n896,
    n668,
    n877,
    n676,
    n881
  );


  nor
  g875
  (
    n890,
    n684,
    n707,
    n872,
    n711
  );


  nor
  g876
  (
    n912,
    n685,
    n884,
    n882
  );


  xor
  g877
  (
    n887,
    n703,
    n678,
    n682,
    n700
  );


  xnor
  g878
  (
    n898,
    n877,
    n870,
    n670,
    n884
  );


  and
  g879
  (
    n899,
    n475,
    n702,
    n882,
    n874
  );


  or
  g880
  (
    n903,
    n475,
    n686,
    n690,
    n683
  );


  xnor
  g881
  (
    n920,
    n669,
    n881,
    n873,
    n882
  );


  or
  g882
  (
    n905,
    n883,
    n679,
    n873,
    n476
  );


  nand
  g883
  (
    n909,
    n879,
    n695,
    n882,
    n883
  );


  or
  g884
  (
    n900,
    n884,
    n697,
    n698,
    n681
  );


  nand
  g885
  (
    n913,
    n704,
    n875,
    n883,
    n699
  );


  nor
  g886
  (
    n897,
    n705,
    n876,
    n674,
    n872
  );


  nand
  g887
  (
    n889,
    n680,
    n883,
    n696,
    n868
  );


  or
  g888
  (
    n894,
    n691,
    n475,
    n688,
    n476
  );


  not
  g889
  (
    n996,
    n909
  );


  not
  g890
  (
    KeyWire_0_6,
    n897
  );


  buf
  g891
  (
    n930,
    n752
  );


  buf
  g892
  (
    n968,
    n720
  );


  not
  g893
  (
    n998,
    n755
  );


  not
  g894
  (
    n926,
    n746
  );


  buf
  g895
  (
    n941,
    n763
  );


  buf
  g896
  (
    n984,
    n763
  );


  not
  g897
  (
    n972,
    n749
  );


  buf
  g898
  (
    n924,
    n919
  );


  not
  g899
  (
    n931,
    n909
  );


  not
  g900
  (
    n980,
    n765
  );


  buf
  g901
  (
    n994,
    n886
  );


  buf
  g902
  (
    n957,
    n921
  );


  buf
  g903
  (
    n934,
    n756
  );


  not
  g904
  (
    n970,
    n750
  );


  buf
  g905
  (
    n938,
    n759
  );


  not
  g906
  (
    n942,
    n716
  );


  buf
  g907
  (
    n964,
    n920
  );


  not
  g908
  (
    KeyWire_0_31,
    n910
  );


  buf
  g909
  (
    n954,
    n893
  );


  not
  g910
  (
    n956,
    n914
  );


  not
  g911
  (
    n991,
    n756
  );


  not
  g912
  (
    n962,
    n726
  );


  not
  g913
  (
    n932,
    n758
  );


  buf
  g914
  (
    KeyWire_0_7,
    n907
  );


  buf
  g915
  (
    n981,
    n726
  );


  buf
  g916
  (
    n946,
    n749
  );


  not
  g917
  (
    n989,
    n752
  );


  not
  g918
  (
    n979,
    n914
  );


  buf
  g919
  (
    n978,
    n717
  );


  not
  g920
  (
    n971,
    n889
  );


  not
  g921
  (
    n948,
    n908
  );


  buf
  g922
  (
    n929,
    n748
  );


  buf
  g923
  (
    n927,
    n911
  );


  buf
  g924
  (
    n966,
    n745
  );


  not
  g925
  (
    n939,
    n759
  );


  buf
  g926
  (
    n953,
    n909
  );


  buf
  g927
  (
    n1000,
    n721
  );


  buf
  g928
  (
    n999,
    n890
  );


  buf
  g929
  (
    KeyWire_0_14,
    n920
  );


  xor
  g930
  (
    n949,
    n758,
    n725
  );


  nand
  g931
  (
    n985,
    n911,
    n920
  );


  xnor
  g932
  (
    n977,
    n766,
    n768,
    n753,
    n726
  );


  nor
  g933
  (
    n937,
    n910,
    n754,
    n895,
    n919
  );


  and
  g934
  (
    n943,
    n719,
    n888,
    n748,
    n761
  );


  or
  g935
  (
    n963,
    n916,
    n756,
    n903,
    n768
  );


  nor
  g936
  (
    n983,
    n749,
    n754,
    n892,
    n905
  );


  xor
  g937
  (
    n923,
    n914,
    n746,
    n906,
    n912
  );


  xor
  g938
  (
    n995,
    n753,
    n908,
    n766,
    n476
  );


  nand
  g939
  (
    n1001,
    n767,
    n755,
    n921,
    n751
  );


  nand
  g940
  (
    n951,
    n917,
    n891,
    n915,
    n754
  );


  or
  g941
  (
    n990,
    n752,
    n747,
    n722,
    n760
  );


  nor
  g942
  (
    n992,
    n908,
    n764,
    n745
  );


  xor
  g943
  (
    n935,
    n907,
    n751,
    n918,
    n902
  );


  xor
  g944
  (
    n960,
    n913,
    n913,
    n908,
    n753
  );


  and
  g945
  (
    n993,
    n759,
    n918,
    n757,
    n767
  );


  nand
  g946
  (
    n928,
    n751,
    n476,
    n750,
    n904
  );


  xnor
  g947
  (
    n936,
    n746,
    n762,
    n885,
    n755
  );


  nand
  g948
  (
    n958,
    n760,
    n916,
    n767,
    n913
  );


  xnor
  g949
  (
    n986,
    n761,
    n754,
    n915,
    n911
  );


  or
  g950
  (
    n965,
    n760,
    n915,
    n767,
    n916
  );


  nand
  g951
  (
    n982,
    n763,
    n750,
    n910,
    n757
  );


  nand
  g952
  (
    n988,
    n766,
    n899,
    n749,
    n750
  );


  or
  g953
  (
    n967,
    n747,
    n762,
    n887,
    n748
  );


  nor
  g954
  (
    n940,
    n765,
    n757,
    n909,
    n766
  );


  nand
  g955
  (
    n976,
    n762,
    n725,
    n914,
    n715
  );


  and
  g956
  (
    n955,
    n918,
    n912,
    n753,
    n919
  );


  and
  g957
  (
    n944,
    n759,
    n760,
    n768,
    n745
  );


  nand
  g958
  (
    n969,
    n917,
    n764,
    n751,
    n901
  );


  nand
  g959
  (
    n947,
    n911,
    n758,
    n917,
    n761
  );


  nor
  g960
  (
    n952,
    n755,
    n894,
    n748,
    n763
  );


  nor
  g961
  (
    n945,
    n912,
    n896,
    n916,
    n758
  );


  nand
  g962
  (
    n987,
    n919,
    n724,
    n765,
    n756
  );


  xnor
  g963
  (
    n925,
    n761,
    n920,
    n723,
    n718
  );


  and
  g964
  (
    n997,
    n747,
    n746,
    n913,
    n764
  );


  or
  g965
  (
    n974,
    n917,
    n898,
    n910,
    n921
  );


  xor
  g966
  (
    n950,
    n768,
    n918,
    n752,
    n747
  );


  nor
  g967
  (
    n961,
    n765,
    n757,
    n915,
    n912
  );


  nor
  g968
  (
    n922,
    n921,
    n762,
    n726,
    n900
  );


  nand
  g969
  (
    n1003,
    n990,
    n936,
    n938,
    n402
  );


  and
  g970
  (
    n1026,
    n727,
    n926,
    n928,
    n989
  );


  xor
  g971
  (
    n1025,
    n967,
    n1001,
    n944,
    n989
  );


  and
  g972
  (
    n1016,
    n995,
    n962,
    n990,
    n956
  );


  nor
  g973
  (
    KeyWire_0_30,
    n954,
    n984,
    n998,
    n974
  );


  xnor
  g974
  (
    n1011,
    n971,
    n1000,
    n999,
    n922
  );


  nand
  g975
  (
    n1014,
    n994,
    n959,
    n953,
    n955
  );


  and
  g976
  (
    n1028,
    n932,
    n993,
    n998,
    n981
  );


  or
  g977
  (
    n1032,
    n1001,
    n949,
    n994
  );


  xor
  g978
  (
    n1015,
    n972,
    n940,
    n973,
    n992
  );


  or
  g979
  (
    n1004,
    n994,
    n996,
    n995,
    n930
  );


  xor
  g980
  (
    n1012,
    n997,
    n946,
    n995,
    n996
  );


  nand
  g981
  (
    n1002,
    n982,
    n934,
    n988,
    n998
  );


  xnor
  g982
  (
    n1019,
    n978,
    n976,
    n990,
    n997
  );


  xnor
  g983
  (
    n1017,
    n998,
    n991,
    n980
  );


  nor
  g984
  (
    n1021,
    n999,
    n999,
    n996,
    n992
  );


  xor
  g985
  (
    n1010,
    n924,
    n987,
    n950,
    n935
  );


  nand
  g986
  (
    n1023,
    n958,
    n999,
    n979,
    n992
  );


  nand
  g987
  (
    n1008,
    n931,
    n966,
    n727,
    n951
  );


  or
  g988
  (
    n1013,
    n1000,
    n969,
    n961,
    n933
  );


  nand
  g989
  (
    n1020,
    n727,
    n947,
    n975,
    n991
  );


  nand
  g990
  (
    n1024,
    n942,
    n996,
    n989,
    n952
  );


  xnor
  g991
  (
    n1030,
    n1001,
    n983,
    n992,
    n986
  );


  nand
  g992
  (
    n1029,
    n948,
    n989,
    n727,
    n941
  );


  xnor
  g993
  (
    n1031,
    n993,
    n964,
    n927,
    n965
  );


  and
  g994
  (
    n1009,
    n960,
    n943,
    n993
  );


  xor
  g995
  (
    n1005,
    n925,
    n1000,
    n991,
    n997
  );


  nand
  g996
  (
    n1007,
    n963,
    n957,
    n970,
    n977
  );


  nor
  g997
  (
    n1018,
    n968,
    n997,
    n945,
    n923
  );


  nand
  g998
  (
    n1006,
    n995,
    n1001,
    n937,
    n939
  );


  xnor
  g999
  (
    n1027,
    n1000,
    n985,
    n929,
    n990
  );


  xnor
  KeyGate_0_0
  (
    n263,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n273,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n138,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n74,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n67,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n403,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n959,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n973,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n655,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n296,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n353,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n703,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n45,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n811,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n975,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n56,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n141,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n176,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n494,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n602,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n439,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n84,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n520,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n586,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n556,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n856,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n286,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n169,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n781,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n654,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1022,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n933,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


