

module Stat_1000_157
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n638,
  n733,
  n759,
  n753,
  n778,
  n775,
  n768,
  n748,
  n758,
  n779,
  n754,
  n750,
  n734,
  n751,
  n745,
  n762,
  n771,
  n767,
  n776,
  n747,
  n740,
  n756,
  n798,
  n1032,
  n1027,
  n1024,
  n1025,
  n1030,
  n1026,
  n1028,
  n1029,
  n1031
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n638;output n733;output n759;output n753;output n778;output n775;output n768;output n748;output n758;output n779;output n754;output n750;output n734;output n751;output n745;output n762;output n771;output n767;output n776;output n747;output n740;output n756;output n798;output n1032;output n1027;output n1024;output n1025;output n1030;output n1026;output n1028;output n1029;output n1031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n735;wire n736;wire n737;wire n738;wire n739;wire n741;wire n742;wire n743;wire n744;wire n746;wire n749;wire n752;wire n755;wire n757;wire n760;wire n761;wire n763;wire n764;wire n765;wire n766;wire n769;wire n770;wire n772;wire n773;wire n774;wire n777;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  not
  g0
  (
    n50,
    n13
  );


  buf
  g1
  (
    n69,
    n11
  );


  not
  g2
  (
    n86,
    n20
  );


  buf
  g3
  (
    n84,
    n17
  );


  not
  g4
  (
    n37,
    n21
  );


  buf
  g5
  (
    n43,
    n4
  );


  not
  g6
  (
    n115,
    n7
  );


  not
  g7
  (
    n49,
    n14
  );


  not
  g8
  (
    n88,
    n17
  );


  buf
  g9
  (
    n100,
    n16
  );


  buf
  g10
  (
    n98,
    n19
  );


  buf
  g11
  (
    n44,
    n10
  );


  buf
  g12
  (
    n63,
    n4
  );


  buf
  g13
  (
    n87,
    n16
  );


  buf
  g14
  (
    n108,
    n7
  );


  buf
  g15
  (
    n111,
    n7
  );


  not
  g16
  (
    n104,
    n16
  );


  not
  g17
  (
    n67,
    n13
  );


  buf
  g18
  (
    n113,
    n22
  );


  not
  g19
  (
    n70,
    n2
  );


  buf
  g20
  (
    n106,
    n3
  );


  not
  g21
  (
    n81,
    n12
  );


  not
  g22
  (
    n38,
    n9
  );


  buf
  g23
  (
    n91,
    n6
  );


  buf
  g24
  (
    n55,
    n18
  );


  not
  g25
  (
    n33,
    n8
  );


  buf
  g26
  (
    n90,
    n5
  );


  not
  g27
  (
    n85,
    n9
  );


  not
  g28
  (
    n116,
    n20
  );


  buf
  g29
  (
    n41,
    n21
  );


  buf
  g30
  (
    n114,
    n3
  );


  buf
  g31
  (
    n34,
    n12
  );


  buf
  g32
  (
    n53,
    n2
  );


  buf
  g33
  (
    n93,
    n10
  );


  not
  g34
  (
    n71,
    n6
  );


  buf
  g35
  (
    n51,
    n10
  );


  buf
  g36
  (
    n79,
    n14
  );


  buf
  g37
  (
    n110,
    n7
  );


  not
  g38
  (
    n74,
    n1
  );


  buf
  g39
  (
    n54,
    n21
  );


  not
  g40
  (
    n95,
    n14
  );


  buf
  g41
  (
    n82,
    n18
  );


  buf
  g42
  (
    n105,
    n3
  );


  not
  g43
  (
    n39,
    n13
  );


  not
  g44
  (
    n59,
    n1
  );


  buf
  g45
  (
    n47,
    n15
  );


  buf
  g46
  (
    n76,
    n1
  );


  buf
  g47
  (
    n60,
    n19
  );


  buf
  g48
  (
    KeyWire_0_12,
    n20
  );


  buf
  g49
  (
    n64,
    n18
  );


  not
  g50
  (
    n102,
    n17
  );


  not
  g51
  (
    n89,
    n12
  );


  buf
  g52
  (
    n118,
    n19
  );


  buf
  g53
  (
    n48,
    n11
  );


  buf
  g54
  (
    n40,
    n8
  );


  buf
  g55
  (
    n107,
    n22
  );


  buf
  g56
  (
    n112,
    n6
  );


  buf
  g57
  (
    n78,
    n9
  );


  not
  g58
  (
    n72,
    n11
  );


  not
  g59
  (
    n36,
    n12
  );


  not
  g60
  (
    n97,
    n5
  );


  not
  g61
  (
    n80,
    n8
  );


  not
  g62
  (
    n109,
    n1
  );


  not
  g63
  (
    n57,
    n2
  );


  buf
  g64
  (
    n52,
    n3
  );


  buf
  g65
  (
    n73,
    n18
  );


  buf
  g66
  (
    n68,
    n14
  );


  not
  g67
  (
    n42,
    n5
  );


  buf
  g68
  (
    n46,
    n20
  );


  not
  g69
  (
    n83,
    n8
  );


  buf
  g70
  (
    n56,
    n2
  );


  not
  g71
  (
    n94,
    n6
  );


  not
  g72
  (
    n45,
    n4
  );


  buf
  g73
  (
    n66,
    n16
  );


  buf
  g74
  (
    n101,
    n15
  );


  not
  g75
  (
    n58,
    n15
  );


  buf
  g76
  (
    n35,
    n5
  );


  not
  g77
  (
    n62,
    n9
  );


  buf
  g78
  (
    n61,
    n19
  );


  buf
  g79
  (
    n77,
    n15
  );


  buf
  g80
  (
    n99,
    n21
  );


  not
  g81
  (
    n65,
    n4
  );


  buf
  g82
  (
    n92,
    n11
  );


  buf
  g83
  (
    n96,
    n13
  );


  not
  g84
  (
    n117,
    n17
  );


  not
  g85
  (
    n103,
    n10
  );


  not
  g86
  (
    n163,
    n72
  );


  not
  g87
  (
    n172,
    n49
  );


  buf
  g88
  (
    n150,
    n70
  );


  not
  g89
  (
    n209,
    n39
  );


  not
  g90
  (
    n169,
    n46
  );


  buf
  g91
  (
    n242,
    n48
  );


  not
  g92
  (
    n282,
    n46
  );


  not
  g93
  (
    n141,
    n34
  );


  not
  g94
  (
    n243,
    n62
  );


  not
  g95
  (
    KeyWire_0_11,
    n68
  );


  not
  g96
  (
    n232,
    n35
  );


  not
  g97
  (
    n143,
    n63
  );


  buf
  g98
  (
    n193,
    n57
  );


  not
  g99
  (
    n170,
    n62
  );


  not
  g100
  (
    n192,
    n55
  );


  buf
  g101
  (
    n124,
    n55
  );


  not
  g102
  (
    n203,
    n43
  );


  buf
  g103
  (
    n182,
    n36
  );


  not
  g104
  (
    n119,
    n47
  );


  buf
  g105
  (
    n228,
    n40
  );


  not
  g106
  (
    n259,
    n73
  );


  buf
  g107
  (
    n175,
    n63
  );


  buf
  g108
  (
    n186,
    n53
  );


  buf
  g109
  (
    n146,
    n50
  );


  buf
  g110
  (
    n256,
    n74
  );


  not
  g111
  (
    n204,
    n41
  );


  buf
  g112
  (
    n248,
    n48
  );


  buf
  g113
  (
    n247,
    n64
  );


  not
  g114
  (
    n158,
    n69
  );


  buf
  g115
  (
    n178,
    n74
  );


  not
  g116
  (
    n221,
    n71
  );


  buf
  g117
  (
    n196,
    n74
  );


  buf
  g118
  (
    n128,
    n57
  );


  buf
  g119
  (
    n260,
    n59
  );


  not
  g120
  (
    n273,
    n66
  );


  buf
  g121
  (
    n162,
    n45
  );


  not
  g122
  (
    n250,
    n43
  );


  buf
  g123
  (
    n263,
    n75
  );


  not
  g124
  (
    n153,
    n67
  );


  not
  g125
  (
    n202,
    n75
  );


  buf
  g126
  (
    n223,
    n35
  );


  not
  g127
  (
    n244,
    n38
  );


  not
  g128
  (
    n293,
    n42
  );


  buf
  g129
  (
    n218,
    n56
  );


  not
  g130
  (
    n165,
    n37
  );


  not
  g131
  (
    n206,
    n34
  );


  not
  g132
  (
    n281,
    n40
  );


  buf
  g133
  (
    n227,
    n44
  );


  not
  g134
  (
    n230,
    n36
  );


  buf
  g135
  (
    n171,
    n53
  );


  buf
  g136
  (
    n144,
    n77
  );


  not
  g137
  (
    n274,
    n42
  );


  not
  g138
  (
    n145,
    n71
  );


  not
  g139
  (
    n164,
    n63
  );


  not
  g140
  (
    n131,
    n39
  );


  not
  g141
  (
    n139,
    n72
  );


  not
  g142
  (
    n138,
    n65
  );


  buf
  g143
  (
    n199,
    n72
  );


  not
  g144
  (
    n268,
    n45
  );


  not
  g145
  (
    n147,
    n48
  );


  not
  g146
  (
    n253,
    n46
  );


  buf
  g147
  (
    n200,
    n47
  );


  not
  g148
  (
    n127,
    n36
  );


  buf
  g149
  (
    n246,
    n49
  );


  buf
  g150
  (
    n217,
    n69
  );


  buf
  g151
  (
    n135,
    n69
  );


  not
  g152
  (
    n180,
    n38
  );


  buf
  g153
  (
    n160,
    n52
  );


  buf
  g154
  (
    n213,
    n47
  );


  buf
  g155
  (
    n215,
    n54
  );


  buf
  g156
  (
    n264,
    n65
  );


  not
  g157
  (
    n185,
    n53
  );


  buf
  g158
  (
    n262,
    n33
  );


  not
  g159
  (
    n129,
    n68
  );


  buf
  g160
  (
    n208,
    n61
  );


  not
  g161
  (
    n212,
    n58
  );


  buf
  g162
  (
    n149,
    n38
  );


  not
  g163
  (
    n234,
    n45
  );


  buf
  g164
  (
    n177,
    n50
  );


  not
  g165
  (
    n214,
    n57
  );


  not
  g166
  (
    n152,
    n46
  );


  not
  g167
  (
    n132,
    n73
  );


  buf
  g168
  (
    n181,
    n34
  );


  not
  g169
  (
    n183,
    n74
  );


  buf
  g170
  (
    n220,
    n34
  );


  buf
  g171
  (
    n276,
    n40
  );


  buf
  g172
  (
    KeyWire_0_8,
    n63
  );


  buf
  g173
  (
    n222,
    n49
  );


  buf
  g174
  (
    n151,
    n33
  );


  buf
  g175
  (
    n252,
    n56
  );


  not
  g176
  (
    n195,
    n70
  );


  not
  g177
  (
    n184,
    n76
  );


  buf
  g178
  (
    n142,
    n60
  );


  buf
  g179
  (
    n155,
    n61
  );


  not
  g180
  (
    n122,
    n54
  );


  buf
  g181
  (
    n271,
    n41
  );


  not
  g182
  (
    n156,
    n65
  );


  buf
  g183
  (
    n189,
    n39
  );


  buf
  g184
  (
    n159,
    n72
  );


  not
  g185
  (
    n279,
    n53
  );


  not
  g186
  (
    n236,
    n44
  );


  buf
  g187
  (
    n261,
    n51
  );


  buf
  g188
  (
    n266,
    n44
  );


  not
  g189
  (
    n201,
    n52
  );


  buf
  g190
  (
    n205,
    n76
  );


  not
  g191
  (
    n283,
    n66
  );


  buf
  g192
  (
    KeyWire_0_1,
    n37
  );


  buf
  g193
  (
    n297,
    n50
  );


  not
  g194
  (
    n290,
    n62
  );


  not
  g195
  (
    n207,
    n71
  );


  buf
  g196
  (
    n120,
    n35
  );


  not
  g197
  (
    n284,
    n70
  );


  buf
  g198
  (
    n148,
    n42
  );


  buf
  g199
  (
    n157,
    n70
  );


  not
  g200
  (
    n133,
    n51
  );


  not
  g201
  (
    n278,
    n65
  );


  not
  g202
  (
    n167,
    n60
  );


  not
  g203
  (
    n211,
    n61
  );


  not
  g204
  (
    n254,
    n66
  );


  not
  g205
  (
    n225,
    n71
  );


  buf
  g206
  (
    n123,
    n59
  );


  buf
  g207
  (
    n229,
    n58
  );


  buf
  g208
  (
    n237,
    n76
  );


  not
  g209
  (
    n191,
    n66
  );


  not
  g210
  (
    n251,
    n56
  );


  buf
  g211
  (
    n277,
    n52
  );


  not
  g212
  (
    n289,
    n77
  );


  not
  g213
  (
    n187,
    n33
  );


  not
  g214
  (
    n291,
    n55
  );


  buf
  g215
  (
    n296,
    n36
  );


  not
  g216
  (
    n197,
    n37
  );


  not
  g217
  (
    n176,
    n51
  );


  not
  g218
  (
    n241,
    n76
  );


  buf
  g219
  (
    n219,
    n45
  );


  not
  g220
  (
    n154,
    n57
  );


  buf
  g221
  (
    n245,
    n50
  );


  buf
  g222
  (
    KeyWire_0_13,
    n59
  );


  buf
  g223
  (
    n216,
    n60
  );


  not
  g224
  (
    n161,
    n48
  );


  not
  g225
  (
    n286,
    n75
  );


  not
  g226
  (
    n280,
    n35
  );


  buf
  g227
  (
    n269,
    n69
  );


  buf
  g228
  (
    n121,
    n64
  );


  not
  g229
  (
    n168,
    n42
  );


  not
  g230
  (
    n249,
    n60
  );


  buf
  g231
  (
    n258,
    n62
  );


  buf
  g232
  (
    n194,
    n52
  );


  buf
  g233
  (
    n265,
    n73
  );


  buf
  g234
  (
    n130,
    n47
  );


  buf
  g235
  (
    n136,
    n67
  );


  buf
  g236
  (
    n173,
    n77
  );


  buf
  g237
  (
    n275,
    n68
  );


  not
  g238
  (
    n285,
    n55
  );


  not
  g239
  (
    n235,
    n33
  );


  not
  g240
  (
    n174,
    n58
  );


  not
  g241
  (
    n287,
    n58
  );


  not
  g242
  (
    n179,
    n56
  );


  not
  g243
  (
    n190,
    n39
  );


  buf
  g244
  (
    n233,
    n54
  );


  not
  g245
  (
    n231,
    n64
  );


  not
  g246
  (
    n267,
    n43
  );


  not
  g247
  (
    n240,
    n61
  );


  buf
  g248
  (
    n126,
    n73
  );


  buf
  g249
  (
    n210,
    n41
  );


  not
  g250
  (
    n295,
    n59
  );


  not
  g251
  (
    n188,
    n37
  );


  not
  g252
  (
    n272,
    n49
  );


  not
  g253
  (
    n226,
    n40
  );


  buf
  g254
  (
    n288,
    n43
  );


  buf
  g255
  (
    n239,
    n41
  );


  not
  g256
  (
    n294,
    n64
  );


  not
  g257
  (
    n257,
    n75
  );


  not
  g258
  (
    n270,
    n67
  );


  buf
  g259
  (
    n166,
    n38
  );


  buf
  g260
  (
    n140,
    n51
  );


  buf
  g261
  (
    n224,
    n44
  );


  buf
  g262
  (
    n134,
    n67
  );


  not
  g263
  (
    n198,
    n54
  );


  buf
  g264
  (
    n238,
    n68
  );


  not
  g265
  (
    n302,
    n259
  );


  not
  g266
  (
    n555,
    n160
  );


  not
  g267
  (
    n316,
    n274
  );


  not
  g268
  (
    n315,
    n166
  );


  not
  g269
  (
    n359,
    n264
  );


  not
  g270
  (
    n496,
    n194
  );


  buf
  g271
  (
    n367,
    n261
  );


  not
  g272
  (
    n509,
    n266
  );


  buf
  g273
  (
    n401,
    n267
  );


  buf
  g274
  (
    n567,
    n193
  );


  not
  g275
  (
    n545,
    n174
  );


  not
  g276
  (
    n331,
    n199
  );


  not
  g277
  (
    n422,
    n213
  );


  buf
  g278
  (
    n395,
    n263
  );


  not
  g279
  (
    n369,
    n204
  );


  not
  g280
  (
    n341,
    n276
  );


  buf
  g281
  (
    n488,
    n264
  );


  buf
  g282
  (
    n404,
    n219
  );


  not
  g283
  (
    n571,
    n291
  );


  buf
  g284
  (
    n343,
    n274
  );


  buf
  g285
  (
    n423,
    n158
  );


  buf
  g286
  (
    n410,
    n272
  );


  buf
  g287
  (
    n531,
    n287
  );


  not
  g288
  (
    n564,
    n292
  );


  not
  g289
  (
    n500,
    n257
  );


  not
  g290
  (
    n476,
    n273
  );


  not
  g291
  (
    n510,
    n275
  );


  buf
  g292
  (
    n480,
    n136
  );


  not
  g293
  (
    n419,
    n138
  );


  not
  g294
  (
    n346,
    n133
  );


  not
  g295
  (
    n335,
    n269
  );


  buf
  g296
  (
    n308,
    n134
  );


  not
  g297
  (
    n319,
    n152
  );


  buf
  g298
  (
    n578,
    n225
  );


  not
  g299
  (
    n378,
    n263
  );


  not
  g300
  (
    n455,
    n151
  );


  not
  g301
  (
    n396,
    n256
  );


  buf
  g302
  (
    n458,
    n271
  );


  not
  g303
  (
    n533,
    n241
  );


  buf
  g304
  (
    n324,
    n272
  );


  buf
  g305
  (
    n390,
    n279
  );


  buf
  g306
  (
    n358,
    n275
  );


  not
  g307
  (
    n537,
    n263
  );


  not
  g308
  (
    n575,
    n146
  );


  not
  g309
  (
    n362,
    n248
  );


  not
  g310
  (
    n321,
    n282
  );


  buf
  g311
  (
    n393,
    n282
  );


  buf
  g312
  (
    n377,
    n234
  );


  not
  g313
  (
    n303,
    n252
  );


  buf
  g314
  (
    n546,
    n232
  );


  not
  g315
  (
    n351,
    n226
  );


  not
  g316
  (
    n439,
    n171
  );


  buf
  g317
  (
    n498,
    n282
  );


  not
  g318
  (
    n322,
    n266
  );


  buf
  g319
  (
    n492,
    n127
  );


  buf
  g320
  (
    n364,
    n290
  );


  not
  g321
  (
    n443,
    n242
  );


  not
  g322
  (
    n317,
    n292
  );


  buf
  g323
  (
    n483,
    n277
  );


  buf
  g324
  (
    n549,
    n126
  );


  not
  g325
  (
    n415,
    n235
  );


  buf
  g326
  (
    n334,
    n164
  );


  not
  g327
  (
    n327,
    n256
  );


  not
  g328
  (
    n421,
    n265
  );


  buf
  g329
  (
    n428,
    n150
  );


  not
  g330
  (
    n583,
    n208
  );


  not
  g331
  (
    n576,
    n195
  );


  not
  g332
  (
    n445,
    n184
  );


  not
  g333
  (
    n389,
    n285
  );


  not
  g334
  (
    n543,
    n182
  );


  not
  g335
  (
    n298,
    n200
  );


  not
  g336
  (
    n536,
    n254
  );


  buf
  g337
  (
    n357,
    n132
  );


  not
  g338
  (
    n526,
    n217
  );


  not
  g339
  (
    n552,
    n255
  );


  not
  g340
  (
    n484,
    n287
  );


  not
  g341
  (
    n352,
    n272
  );


  buf
  g342
  (
    n407,
    n270
  );


  buf
  g343
  (
    n425,
    n190
  );


  not
  g344
  (
    n568,
    n220
  );


  not
  g345
  (
    n508,
    n269
  );


  not
  g346
  (
    n414,
    n264
  );


  not
  g347
  (
    n538,
    n212
  );


  buf
  g348
  (
    n311,
    n288
  );


  buf
  g349
  (
    n363,
    n180
  );


  not
  g350
  (
    n465,
    n163
  );


  not
  g351
  (
    n519,
    n144
  );


  not
  g352
  (
    n332,
    n291
  );


  buf
  g353
  (
    n547,
    n266
  );


  not
  g354
  (
    n548,
    n250
  );


  not
  g355
  (
    n350,
    n161
  );


  buf
  g356
  (
    n456,
    n211
  );


  not
  g357
  (
    n444,
    n222
  );


  not
  g358
  (
    n386,
    n279
  );


  not
  g359
  (
    n562,
    n268
  );


  not
  g360
  (
    n521,
    n280
  );


  buf
  g361
  (
    n482,
    n267
  );


  buf
  g362
  (
    n345,
    n215
  );


  not
  g363
  (
    n307,
    n276
  );


  buf
  g364
  (
    n540,
    n196
  );


  buf
  g365
  (
    n323,
    n145
  );


  buf
  g366
  (
    n494,
    n187
  );


  buf
  g367
  (
    n318,
    n256
  );


  not
  g368
  (
    n513,
    n272
  );


  not
  g369
  (
    KeyWire_0_9,
    n261
  );


  buf
  g370
  (
    n398,
    n262
  );


  not
  g371
  (
    n330,
    n246
  );


  buf
  g372
  (
    n372,
    n262
  );


  not
  g373
  (
    n581,
    n261
  );


  buf
  g374
  (
    n418,
    n277
  );


  buf
  g375
  (
    n512,
    n287
  );


  buf
  g376
  (
    KeyWire_0_2,
    n269
  );


  buf
  g377
  (
    n557,
    n273
  );


  buf
  g378
  (
    n577,
    n256
  );


  not
  g379
  (
    n544,
    n153
  );


  not
  g380
  (
    n355,
    n178
  );


  not
  g381
  (
    n515,
    n276
  );


  buf
  g382
  (
    n388,
    n189
  );


  not
  g383
  (
    n551,
    n277
  );


  buf
  g384
  (
    n329,
    n121
  );


  buf
  g385
  (
    n374,
    n125
  );


  not
  g386
  (
    n481,
    n279
  );


  not
  g387
  (
    n313,
    n289
  );


  buf
  g388
  (
    n520,
    n282
  );


  not
  g389
  (
    n559,
    n259
  );


  buf
  g390
  (
    n470,
    n284
  );


  not
  g391
  (
    n522,
    n147
  );


  not
  g392
  (
    n493,
    n257
  );


  buf
  g393
  (
    n347,
    n175
  );


  not
  g394
  (
    n572,
    n283
  );


  not
  g395
  (
    n495,
    n201
  );


  buf
  g396
  (
    n530,
    n293
  );


  buf
  g397
  (
    n447,
    n188
  );


  not
  g398
  (
    n527,
    n286
  );


  buf
  g399
  (
    n382,
    n271
  );


  buf
  g400
  (
    n349,
    n244
  );


  not
  g401
  (
    n460,
    n284
  );


  buf
  g402
  (
    n457,
    n142
  );


  not
  g403
  (
    n504,
    n274
  );


  not
  g404
  (
    n475,
    n286
  );


  not
  g405
  (
    n365,
    n270
  );


  buf
  g406
  (
    n429,
    n139
  );


  buf
  g407
  (
    n535,
    n224
  );


  not
  g408
  (
    n394,
    n245
  );


  not
  g409
  (
    n333,
    n261
  );


  not
  g410
  (
    n477,
    n249
  );


  buf
  g411
  (
    n400,
    n230
  );


  buf
  g412
  (
    n406,
    n185
  );


  buf
  g413
  (
    n381,
    n172
  );


  not
  g414
  (
    n342,
    n258
  );


  not
  g415
  (
    n437,
    n262
  );


  buf
  g416
  (
    n325,
    n165
  );


  not
  g417
  (
    n405,
    n198
  );


  not
  g418
  (
    n353,
    n280
  );


  buf
  g419
  (
    n474,
    n216
  );


  buf
  g420
  (
    n497,
    n238
  );


  buf
  g421
  (
    n573,
    n169
  );


  not
  g422
  (
    n397,
    n237
  );


  not
  g423
  (
    n556,
    n258
  );


  not
  g424
  (
    n517,
    n260
  );


  not
  g425
  (
    n542,
    n271
  );


  not
  g426
  (
    n469,
    n168
  );


  buf
  g427
  (
    n301,
    n278
  );


  not
  g428
  (
    n448,
    n281
  );


  buf
  g429
  (
    n574,
    n275
  );


  not
  g430
  (
    n501,
    n271
  );


  not
  g431
  (
    n487,
    n285
  );


  not
  g432
  (
    n340,
    n289
  );


  not
  g433
  (
    n507,
    n130
  );


  buf
  g434
  (
    n503,
    n197
  );


  buf
  g435
  (
    n464,
    n231
  );


  not
  g436
  (
    n408,
    n119
  );


  buf
  g437
  (
    n385,
    n257
  );


  not
  g438
  (
    n499,
    n131
  );


  buf
  g439
  (
    n360,
    n278
  );


  buf
  g440
  (
    n413,
    n183
  );


  not
  g441
  (
    n454,
    n154
  );


  not
  g442
  (
    n471,
    n203
  );


  buf
  g443
  (
    n561,
    n283
  );


  buf
  g444
  (
    n361,
    n287
  );


  not
  g445
  (
    n433,
    n290
  );


  not
  g446
  (
    KeyWire_0_10,
    n291
  );


  buf
  g447
  (
    n514,
    n124
  );


  buf
  g448
  (
    n370,
    n273
  );


  buf
  g449
  (
    n441,
    n157
  );


  buf
  g450
  (
    n305,
    n240
  );


  not
  g451
  (
    n534,
    n191
  );


  not
  g452
  (
    n384,
    n265
  );


  not
  g453
  (
    n339,
    n275
  );


  buf
  g454
  (
    n468,
    n283
  );


  not
  g455
  (
    n579,
    n202
  );


  buf
  g456
  (
    n452,
    n258
  );


  buf
  g457
  (
    n326,
    n260
  );


  buf
  g458
  (
    n449,
    n159
  );


  buf
  g459
  (
    n336,
    n292
  );


  buf
  g460
  (
    n434,
    n262
  );


  not
  g461
  (
    n344,
    n143
  );


  buf
  g462
  (
    n430,
    n268
  );


  not
  g463
  (
    n461,
    n278
  );


  not
  g464
  (
    n417,
    n288
  );


  buf
  g465
  (
    n320,
    n284
  );


  not
  g466
  (
    n442,
    n274
  );


  buf
  g467
  (
    n523,
    n167
  );


  not
  g468
  (
    n467,
    n277
  );


  buf
  g469
  (
    n354,
    n290
  );


  buf
  g470
  (
    n424,
    n279
  );


  not
  g471
  (
    n565,
    n264
  );


  buf
  g472
  (
    n314,
    n156
  );


  not
  g473
  (
    n373,
    n267
  );


  buf
  g474
  (
    n511,
    n290
  );


  not
  g475
  (
    n462,
    n206
  );


  not
  g476
  (
    n582,
    n192
  );


  buf
  g477
  (
    n516,
    n283
  );


  buf
  g478
  (
    n402,
    n268
  );


  not
  g479
  (
    n554,
    n135
  );


  not
  g480
  (
    n356,
    n181
  );


  buf
  g481
  (
    n309,
    n276
  );


  not
  g482
  (
    n485,
    n247
  );


  not
  g483
  (
    n478,
    n236
  );


  buf
  g484
  (
    n506,
    n269
  );


  not
  g485
  (
    n420,
    n259
  );


  buf
  g486
  (
    n306,
    n148
  );


  buf
  g487
  (
    n524,
    n260
  );


  buf
  g488
  (
    n532,
    n289
  );


  not
  g489
  (
    n489,
    n278
  );


  buf
  g490
  (
    n399,
    n288
  );


  buf
  g491
  (
    n529,
    n284
  );


  not
  g492
  (
    n463,
    n141
  );


  buf
  g493
  (
    n392,
    n286
  );


  not
  g494
  (
    n375,
    n285
  );


  buf
  g495
  (
    n348,
    n162
  );


  not
  g496
  (
    n432,
    n122
  );


  buf
  g497
  (
    n438,
    n265
  );


  buf
  g498
  (
    n376,
    n267
  );


  buf
  g499
  (
    n558,
    n209
  );


  not
  g500
  (
    n436,
    n258
  );


  not
  g501
  (
    n440,
    n280
  );


  not
  g502
  (
    n391,
    n289
  );


  not
  g503
  (
    n379,
    n292
  );


  not
  g504
  (
    n337,
    n229
  );


  not
  g505
  (
    n409,
    n155
  );


  buf
  g506
  (
    n371,
    n228
  );


  not
  g507
  (
    n310,
    n129
  );


  not
  g508
  (
    n490,
    n281
  );


  buf
  g509
  (
    n380,
    n173
  );


  buf
  g510
  (
    n412,
    n281
  );


  buf
  g511
  (
    n569,
    n207
  );


  not
  g512
  (
    KeyWire_0_5,
    n280
  );


  not
  g513
  (
    n560,
    n281
  );


  buf
  g514
  (
    n426,
    n218
  );


  buf
  g515
  (
    n472,
    n286
  );


  not
  g516
  (
    n505,
    n273
  );


  buf
  g517
  (
    n580,
    n239
  );


  buf
  g518
  (
    n416,
    n214
  );


  not
  g519
  (
    n466,
    n243
  );


  buf
  g520
  (
    n525,
    n137
  );


  not
  g521
  (
    n563,
    n170
  );


  not
  g522
  (
    n450,
    n266
  );


  buf
  g523
  (
    n431,
    n186
  );


  buf
  g524
  (
    KeyWire_0_0,
    n140
  );


  buf
  g525
  (
    n479,
    n223
  );


  buf
  g526
  (
    n553,
    n288
  );


  not
  g527
  (
    n486,
    n179
  );


  not
  g528
  (
    n491,
    n128
  );


  buf
  g529
  (
    n459,
    n265
  );


  buf
  g530
  (
    n453,
    n268
  );


  not
  g531
  (
    n566,
    n285
  );


  not
  g532
  (
    n338,
    n221
  );


  buf
  g533
  (
    n299,
    n176
  );


  buf
  g534
  (
    n427,
    n233
  );


  not
  g535
  (
    n502,
    n270
  );


  not
  g536
  (
    n328,
    n263
  );


  not
  g537
  (
    n518,
    n251
  );


  not
  g538
  (
    n383,
    n177
  );


  buf
  g539
  (
    n528,
    n253
  );


  not
  g540
  (
    n368,
    n259
  );


  buf
  g541
  (
    n435,
    n227
  );


  buf
  g542
  (
    n451,
    n120
  );


  buf
  g543
  (
    n403,
    n270
  );


  buf
  g544
  (
    n570,
    n205
  );


  not
  g545
  (
    n300,
    n149
  );


  buf
  g546
  (
    n550,
    n260
  );


  buf
  g547
  (
    n366,
    n210
  );


  not
  g548
  (
    n539,
    n291
  );


  buf
  g549
  (
    n411,
    n123
  );


  buf
  g550
  (
    n446,
    n257
  );


  buf
  g551
  (
    n616,
    n333
  );


  buf
  g552
  (
    n609,
    n308
  );


  buf
  g553
  (
    n624,
    n327
  );


  not
  g554
  (
    n618,
    n348
  );


  buf
  g555
  (
    n645,
    n359
  );


  not
  g556
  (
    n593,
    n331
  );


  buf
  g557
  (
    n622,
    n324
  );


  buf
  g558
  (
    n617,
    n311
  );


  not
  g559
  (
    n628,
    n319
  );


  not
  g560
  (
    n646,
    n316
  );


  not
  g561
  (
    n637,
    n332
  );


  buf
  g562
  (
    n640,
    n361
  );


  buf
  g563
  (
    n607,
    n306
  );


  not
  g564
  (
    n601,
    n350
  );


  buf
  g565
  (
    n627,
    n337
  );


  buf
  g566
  (
    n610,
    n339
  );


  not
  g567
  (
    n633,
    n307
  );


  buf
  g568
  (
    n625,
    n347
  );


  not
  g569
  (
    n634,
    n355
  );


  buf
  g570
  (
    n591,
    n360
  );


  buf
  g571
  (
    n600,
    n330
  );


  buf
  g572
  (
    n619,
    n349
  );


  not
  g573
  (
    n636,
    n321
  );


  buf
  g574
  (
    n613,
    n336
  );


  buf
  g575
  (
    KeyWire_0_4,
    n303
  );


  not
  g576
  (
    n635,
    n342
  );


  buf
  g577
  (
    n588,
    n343
  );


  not
  g578
  (
    n596,
    n313
  );


  buf
  g579
  (
    n595,
    n358
  );


  not
  g580
  (
    n602,
    n299
  );


  not
  g581
  (
    n639,
    n312
  );


  buf
  g582
  (
    n586,
    n325
  );


  buf
  g583
  (
    n604,
    n329
  );


  not
  g584
  (
    n620,
    n300
  );


  not
  g585
  (
    n585,
    n326
  );


  buf
  g586
  (
    n611,
    n310
  );


  not
  g587
  (
    n608,
    n314
  );


  not
  g588
  (
    n597,
    n335
  );


  buf
  g589
  (
    n647,
    n315
  );


  not
  g590
  (
    n642,
    n340
  );


  buf
  g591
  (
    n598,
    n352
  );


  buf
  g592
  (
    n615,
    n346
  );


  buf
  g593
  (
    n641,
    n338
  );


  buf
  g594
  (
    n612,
    n357
  );


  not
  g595
  (
    n631,
    n341
  );


  not
  g596
  (
    n594,
    n328
  );


  buf
  g597
  (
    n643,
    n317
  );


  buf
  g598
  (
    n606,
    n334
  );


  buf
  g599
  (
    n605,
    n304
  );


  buf
  g600
  (
    n590,
    n351
  );


  buf
  g601
  (
    n587,
    n322
  );


  buf
  g602
  (
    n603,
    n305
  );


  not
  g603
  (
    n638,
    n318
  );


  not
  g604
  (
    n584,
    n301
  );


  buf
  g605
  (
    n626,
    n354
  );


  buf
  g606
  (
    n592,
    n345
  );


  not
  g607
  (
    n599,
    n356
  );


  buf
  g608
  (
    n621,
    n298
  );


  buf
  g609
  (
    n614,
    n320
  );


  buf
  g610
  (
    n630,
    n323
  );


  buf
  g611
  (
    n623,
    n344
  );


  not
  g612
  (
    n644,
    n353
  );


  buf
  g613
  (
    n589,
    n309
  );


  buf
  g614
  (
    n632,
    n302
  );


  buf
  g615
  (
    n658,
    n587
  );


  not
  g616
  (
    n659,
    n599
  );


  not
  g617
  (
    n650,
    n597
  );


  not
  g618
  (
    n674,
    n599
  );


  not
  g619
  (
    n649,
    n591
  );


  buf
  g620
  (
    n666,
    n597
  );


  not
  g621
  (
    n667,
    n592
  );


  buf
  g622
  (
    n648,
    n593
  );


  buf
  g623
  (
    n668,
    n584
  );


  not
  g624
  (
    n677,
    n596
  );


  not
  g625
  (
    n665,
    n585
  );


  buf
  g626
  (
    KeyWire_0_6,
    n598
  );


  not
  g627
  (
    n673,
    n595
  );


  buf
  g628
  (
    n661,
    n596
  );


  buf
  g629
  (
    n652,
    n597
  );


  buf
  g630
  (
    n664,
    n597
  );


  not
  g631
  (
    n670,
    n589
  );


  not
  g632
  (
    n662,
    n586
  );


  buf
  g633
  (
    n653,
    n599
  );


  buf
  g634
  (
    n654,
    n600
  );


  not
  g635
  (
    n671,
    n595
  );


  not
  g636
  (
    n663,
    n588
  );


  not
  g637
  (
    n675,
    n599
  );


  not
  g638
  (
    n655,
    n598
  );


  buf
  g639
  (
    n676,
    n598
  );


  not
  g640
  (
    n651,
    n596
  );


  not
  g641
  (
    n656,
    n590
  );


  not
  g642
  (
    n672,
    n598
  );


  buf
  g643
  (
    n657,
    n594
  );


  buf
  g644
  (
    n660,
    n596
  );


  nor
  g645
  (
    n729,
    n26,
    n398,
    n458,
    n441
  );


  and
  g646
  (
    n683,
    n365,
    n380,
    n651,
    n409
  );


  nor
  g647
  (
    n687,
    n482,
    n454,
    n384,
    n455
  );


  and
  g648
  (
    n726,
    n30,
    n665,
    n25,
    n666
  );


  or
  g649
  (
    n696,
    n435,
    n28,
    n29,
    n432
  );


  nor
  g650
  (
    n711,
    n464,
    n427,
    n470,
    n367
  );


  and
  g651
  (
    n698,
    n658,
    n481,
    n668,
    n394
  );


  nor
  g652
  (
    n715,
    n667,
    n376,
    n418,
    n26
  );


  xor
  g653
  (
    n704,
    n32,
    n450,
    n392,
    n404
  );


  or
  g654
  (
    n721,
    n661,
    n662,
    n421,
    n461
  );


  or
  g655
  (
    n731,
    n28,
    n370,
    n456,
    n663
  );


  or
  g656
  (
    n682,
    n467,
    n665,
    n438,
    n22
  );


  or
  g657
  (
    n680,
    n476,
    n660,
    n24,
    n433
  );


  and
  g658
  (
    n679,
    n420,
    n668,
    n452,
    n661
  );


  xnor
  g659
  (
    n690,
    n480,
    n664,
    n24,
    n31
  );


  and
  g660
  (
    n697,
    n652,
    n32,
    n414,
    n25
  );


  nor
  g661
  (
    n691,
    n664,
    n663,
    n406,
    n373
  );


  or
  g662
  (
    n727,
    n666,
    n419,
    n29,
    n483
  );


  nor
  g663
  (
    n725,
    n366,
    n449,
    n402,
    n408
  );


  or
  g664
  (
    n681,
    n473,
    n29,
    n665,
    n417
  );


  xor
  g665
  (
    n706,
    n428,
    n23,
    n386,
    n375
  );


  nor
  g666
  (
    n700,
    n654,
    n478,
    n383,
    n405
  );


  or
  g667
  (
    n699,
    n388,
    n451,
    n660,
    n391
  );


  xor
  g668
  (
    n730,
    n400,
    n393,
    n649,
    n474
  );


  xnor
  g669
  (
    n689,
    n442,
    n443,
    n410,
    n378
  );


  nor
  g670
  (
    n684,
    n379,
    n371,
    n377,
    n466
  );


  nand
  g671
  (
    n707,
    n436,
    n31,
    n656,
    n445
  );


  and
  g672
  (
    n716,
    n662,
    n413,
    n660,
    n430
  );


  and
  g673
  (
    n724,
    n30,
    n477,
    n440,
    n23
  );


  nand
  g674
  (
    n723,
    n659,
    n664,
    n25,
    n471
  );


  xnor
  g675
  (
    n694,
    n653,
    n395,
    n23,
    n368
  );


  nand
  g676
  (
    n710,
    n479,
    n668,
    n27,
    n667
  );


  and
  g677
  (
    n693,
    n661,
    n28,
    n659,
    n24
  );


  nor
  g678
  (
    n718,
    n658,
    n22,
    n27,
    n659
  );


  xor
  g679
  (
    n695,
    n389,
    n364,
    n472,
    n484
  );


  xnor
  g680
  (
    n678,
    n469,
    n666,
    n667,
    n363
  );


  nor
  g681
  (
    n701,
    n403,
    n439,
    n385,
    n663
  );


  nand
  g682
  (
    n708,
    n669,
    n666,
    n659,
    n457
  );


  and
  g683
  (
    n709,
    n663,
    n369,
    n426,
    n30
  );


  or
  g684
  (
    n686,
    n423,
    n669,
    n650,
    n381
  );


  xor
  g685
  (
    n728,
    n668,
    n416,
    n429,
    n434
  );


  nand
  g686
  (
    n720,
    n27,
    n655,
    n397,
    n453
  );


  or
  g687
  (
    n703,
    n372,
    n660,
    n648,
    n448
  );


  xor
  g688
  (
    n722,
    n28,
    n669,
    n657,
    n437
  );


  and
  g689
  (
    n688,
    n665,
    n412,
    n465,
    n459
  );


  xor
  g690
  (
    n713,
    n444,
    n390,
    n431,
    n382
  );


  nand
  g691
  (
    n732,
    n387,
    n475,
    n26,
    n463
  );


  xnor
  g692
  (
    n705,
    n23,
    n32,
    n30
  );


  nor
  g693
  (
    n719,
    n462,
    n399,
    n31,
    n446
  );


  xor
  g694
  (
    n717,
    n407,
    n29,
    n422,
    n662
  );


  and
  g695
  (
    n714,
    n26,
    n25,
    n460,
    n425
  );


  xnor
  g696
  (
    n702,
    n415,
    n661,
    n447,
    n662
  );


  nand
  g697
  (
    n712,
    n664,
    n27,
    n411,
    n401
  );


  nor
  g698
  (
    n685,
    n424,
    n24,
    n396,
    n362
  );


  or
  g699
  (
    n692,
    n468,
    n31,
    n667,
    n374
  );


  nand
  g700
  (
    n775,
    n97,
    n95,
    n81,
    n688
  );


  nand
  g701
  (
    n748,
    n702,
    n86,
    n687,
    n689
  );


  xor
  g702
  (
    n759,
    n697,
    n90,
    n95,
    n91
  );


  and
  g703
  (
    n747,
    n708,
    n707,
    n98,
    n700
  );


  xor
  g704
  (
    n740,
    n85,
    n90,
    n698,
    n94
  );


  or
  g705
  (
    n767,
    n678,
    n698,
    n79,
    n687
  );


  nand
  g706
  (
    n769,
    n699,
    n96,
    n98,
    n707
  );


  or
  g707
  (
    n754,
    n78,
    n694,
    n686,
    n89
  );


  xnor
  g708
  (
    n749,
    n92,
    n81,
    n701,
    n686
  );


  xnor
  g709
  (
    n772,
    n697,
    n692,
    n79,
    n91
  );


  nor
  g710
  (
    n771,
    n693,
    n696,
    n79,
    n94
  );


  nor
  g711
  (
    n745,
    n693,
    n92,
    n94,
    n690
  );


  or
  g712
  (
    n739,
    n97,
    n695,
    n91,
    n77
  );


  xor
  g713
  (
    n742,
    n82,
    n691,
    n80,
    n81
  );


  and
  g714
  (
    n757,
    n699,
    n84,
    n86,
    n691
  );


  xor
  g715
  (
    n744,
    n687,
    n82,
    n696,
    n87
  );


  or
  g716
  (
    n773,
    n81,
    n704,
    n705,
    n91
  );


  or
  g717
  (
    n750,
    n97,
    n689,
    n86,
    n679
  );


  or
  g718
  (
    n763,
    n700,
    n87,
    n685,
    n705
  );


  nand
  g719
  (
    n761,
    n705,
    n80,
    n89
  );


  and
  g720
  (
    n743,
    n92,
    n97,
    n98,
    n84
  );


  xnor
  g721
  (
    n736,
    n85,
    n706,
    n80,
    n695
  );


  or
  g722
  (
    n776,
    n701,
    n90,
    n96,
    n694
  );


  xor
  g723
  (
    n779,
    n86,
    n88,
    n691,
    n702
  );


  xnor
  g724
  (
    n778,
    n696,
    n78,
    n84,
    n682
  );


  or
  g725
  (
    n735,
    n90,
    n83,
    n708,
    n87
  );


  nand
  g726
  (
    n738,
    n88,
    n702,
    n706,
    n701
  );


  xor
  g727
  (
    n777,
    n95,
    n95,
    n87,
    n93
  );


  xnor
  g728
  (
    n770,
    n697,
    n78,
    n703,
    n93
  );


  nand
  g729
  (
    n768,
    n685,
    n693,
    n692,
    n707
  );


  or
  g730
  (
    n766,
    n690,
    n79,
    n93,
    n695
  );


  nand
  g731
  (
    n774,
    n690,
    n89,
    n684,
    n85
  );


  xnor
  g732
  (
    n746,
    n88,
    n680,
    n699,
    n85
  );


  xor
  g733
  (
    n737,
    n704,
    n88,
    n688,
    n701
  );


  or
  g734
  (
    n758,
    n707,
    n94,
    n697,
    n693
  );


  or
  g735
  (
    n752,
    n99,
    n686,
    n690,
    n96
  );


  nand
  g736
  (
    n762,
    n600,
    n696,
    n703,
    n93
  );


  xor
  g737
  (
    n760,
    n83,
    n84,
    n82,
    n78
  );


  xor
  g738
  (
    n741,
    n83,
    n699,
    n689,
    n698
  );


  and
  g739
  (
    n755,
    n687,
    n691,
    n703,
    n688
  );


  or
  g740
  (
    n753,
    n99,
    n689,
    n694,
    n82
  );


  xor
  g741
  (
    n734,
    n692,
    n700,
    n704,
    n703
  );


  nor
  g742
  (
    n756,
    n694,
    n681,
    n695,
    n692
  );


  nor
  g743
  (
    n765,
    n83,
    n92,
    n706,
    n96
  );


  or
  g744
  (
    n733,
    n702,
    n686,
    n698,
    n704
  );


  and
  g745
  (
    n751,
    n705,
    n688,
    n89,
    n706
  );


  xnor
  g746
  (
    n764,
    n683,
    n700,
    n98,
    n600
  );


  xor
  g747
  (
    n787,
    n605,
    n607,
    n604,
    n601
  );


  nand
  g748
  (
    n783,
    n763,
    n293,
    n760
  );


  xor
  g749
  (
    n790,
    n297,
    n607,
    n709,
    n766
  );


  xnor
  g750
  (
    n797,
    n770,
    n602,
    n710,
    n295
  );


  xnor
  g751
  (
    n794,
    n601,
    n709,
    n710,
    n711
  );


  nand
  g752
  (
    n789,
    n755,
    n294,
    n606,
    n602
  );


  xor
  g753
  (
    n798,
    n294,
    n709,
    n711,
    n603
  );


  xor
  g754
  (
    KeyWire_0_14,
    n757,
    n294,
    n710
  );


  xor
  g755
  (
    n781,
    n762,
    n295,
    n603,
    n605
  );


  or
  g756
  (
    n786,
    n297,
    n296,
    n604,
    n772
  );


  and
  g757
  (
    n785,
    n605,
    n708,
    n754,
    n709
  );


  and
  g758
  (
    n793,
    n603,
    n293,
    n296,
    n602
  );


  or
  g759
  (
    n780,
    n765,
    n761,
    n297,
    n759
  );


  nor
  g760
  (
    n791,
    n602,
    n601,
    n603,
    n771
  );


  or
  g761
  (
    n792,
    n296,
    n604,
    n756,
    n295
  );


  and
  g762
  (
    n788,
    n606,
    n604,
    n601,
    n758
  );


  nor
  g763
  (
    n796,
    n296,
    n768,
    n764,
    n773
  );


  nand
  g764
  (
    n795,
    n769,
    n605,
    n295,
    n607
  );


  and
  g765
  (
    n784,
    n600,
    n294,
    n607,
    n708
  );


  xnor
  g766
  (
    n782,
    n606,
    n606,
    n297,
    n767
  );


  xnor
  g767
  (
    n802,
    n549,
    n555,
    n792,
    n783
  );


  and
  g768
  (
    n807,
    n560,
    n541,
    n556,
    n531
  );


  nor
  g769
  (
    n801,
    n559,
    n505,
    n519,
    n523
  );


  and
  g770
  (
    n819,
    n506,
    n542,
    n500,
    n522
  );


  or
  g771
  (
    n820,
    n503,
    n543,
    n711,
    n547
  );


  or
  g772
  (
    n806,
    n791,
    n540,
    n784,
    n495
  );


  nand
  g773
  (
    n817,
    n497,
    n535,
    n537,
    n780
  );


  nor
  g774
  (
    n800,
    n538,
    n533,
    n510,
    n790
  );


  xor
  g775
  (
    n815,
    n791,
    n554,
    n485,
    n496
  );


  nand
  g776
  (
    n824,
    n498,
    n787,
    n504,
    n552
  );


  xor
  g777
  (
    n803,
    n544,
    n507,
    n527,
    n550
  );


  nor
  g778
  (
    n805,
    n539,
    n509,
    n789,
    n516
  );


  and
  g779
  (
    n812,
    n524,
    n532,
    n515,
    n790
  );


  xor
  g780
  (
    n825,
    n488,
    n712,
    n781,
    n526
  );


  xor
  g781
  (
    n810,
    n513,
    n521,
    n551,
    n512
  );


  or
  g782
  (
    n811,
    n490,
    n782,
    n712,
    n557
  );


  or
  g783
  (
    n809,
    n502,
    n530,
    n786,
    n514
  );


  nor
  g784
  (
    n826,
    n791,
    n499,
    n493,
    n789
  );


  nand
  g785
  (
    n823,
    n791,
    n790,
    n789,
    n494
  );


  xnor
  g786
  (
    n822,
    n788,
    n487,
    n711,
    n534
  );


  xnor
  g787
  (
    n813,
    n545,
    n520,
    n792,
    n536
  );


  xnor
  g788
  (
    n816,
    n712,
    n787,
    n528,
    n788
  );


  nor
  g789
  (
    n821,
    n789,
    n501,
    n517,
    n529
  );


  xnor
  g790
  (
    n804,
    n792,
    n548,
    n492,
    n558
  );


  and
  g791
  (
    n814,
    n491,
    n790,
    n792,
    n525
  );


  and
  g792
  (
    n818,
    n553,
    n486,
    n511,
    n785
  );


  or
  g793
  (
    n808,
    n546,
    n508,
    n489,
    n518
  );


  not
  g794
  (
    n830,
    n818
  );


  buf
  g795
  (
    n836,
    n608
  );


  not
  g796
  (
    n840,
    n609
  );


  buf
  g797
  (
    n847,
    n812
  );


  not
  g798
  (
    n835,
    n806
  );


  buf
  g799
  (
    n833,
    n805
  );


  not
  g800
  (
    n828,
    n807
  );


  not
  g801
  (
    n832,
    n813
  );


  buf
  g802
  (
    n827,
    n610
  );


  buf
  g803
  (
    n846,
    n815
  );


  not
  g804
  (
    n850,
    n822
  );


  buf
  g805
  (
    n838,
    n816
  );


  buf
  g806
  (
    n843,
    n811
  );


  buf
  g807
  (
    n837,
    n810
  );


  buf
  g808
  (
    n829,
    n801
  );


  buf
  g809
  (
    n848,
    n610
  );


  not
  g810
  (
    n842,
    n809
  );


  buf
  g811
  (
    n839,
    n608
  );


  buf
  g812
  (
    n845,
    n808
  );


  buf
  g813
  (
    n841,
    n814
  );


  and
  g814
  (
    n834,
    n610,
    n802,
    n817,
    n803
  );


  or
  g815
  (
    n844,
    n610,
    n823,
    n804,
    n820
  );


  and
  g816
  (
    n849,
    n819,
    n821,
    n608,
    n609
  );


  nand
  g817
  (
    n831,
    n800,
    n608,
    n609
  );


  xor
  g818
  (
    n858,
    n566,
    n721
  );


  and
  g819
  (
    n852,
    n612,
    n564
  );


  nor
  g820
  (
    n936,
    n612,
    n836,
    n832,
    n619
  );


  or
  g821
  (
    n902,
    n639,
    n848,
    n614,
    n846
  );


  xnor
  g822
  (
    n938,
    n840,
    n634,
    n847,
    n844
  );


  or
  g823
  (
    n914,
    n794,
    n632,
    n672,
    n842
  );


  xor
  g824
  (
    n860,
    n568,
    n799,
    n716,
    n640
  );


  xnor
  g825
  (
    n886,
    n799,
    n616,
    n674,
    n719
  );


  xor
  g826
  (
    n923,
    n831,
    n828,
    n625,
    n633
  );


  and
  g827
  (
    n911,
    n622,
    n716,
    n844,
    n717
  );


  xnor
  g828
  (
    n888,
    n614,
    n673,
    n675,
    n616
  );


  xor
  g829
  (
    n865,
    n798,
    n574,
    n577,
    n718
  );


  nand
  g830
  (
    n929,
    n623,
    n619,
    n632,
    n725
  );


  nand
  g831
  (
    n855,
    n629,
    n715,
    n621,
    n620
  );


  or
  g832
  (
    n916,
    n837,
    n635,
    n638,
    n726
  );


  and
  g833
  (
    n900,
    n615,
    n846,
    n628,
    n834
  );


  xnor
  g834
  (
    n935,
    n831,
    n674,
    n620,
    n617
  );


  and
  g835
  (
    n862,
    n845,
    n836,
    n674,
    n614
  );


  nor
  g836
  (
    n878,
    n724,
    n570,
    n841,
    n670
  );


  xor
  g837
  (
    n875,
    n846,
    n794,
    n676,
    n848
  );


  xor
  g838
  (
    n895,
    n843,
    n840,
    n617,
    n572
  );


  xor
  g839
  (
    n925,
    n828,
    n845,
    n576,
    n847
  );


  nor
  g840
  (
    n941,
    n578,
    n672,
    n842,
    n675
  );


  xnor
  g841
  (
    n937,
    n641,
    n631,
    n848,
    n629
  );


  xor
  g842
  (
    n861,
    n631,
    n830,
    n718,
    n617
  );


  or
  g843
  (
    n920,
    n842,
    n611,
    n672,
    n563
  );


  xnor
  g844
  (
    n879,
    n630,
    n720,
    n799,
    n562
  );


  xnor
  g845
  (
    n898,
    n627,
    n835,
    n722,
    n828
  );


  xnor
  g846
  (
    n868,
    n712,
    n793,
    n637,
    n721
  );


  xnor
  g847
  (
    n896,
    n674,
    n832,
    n833,
    n713
  );


  or
  g848
  (
    n870,
    n101,
    n671,
    n835
  );


  xor
  g849
  (
    n921,
    n677,
    n621,
    n633,
    n640
  );


  and
  g850
  (
    n857,
    n841,
    n841,
    n613,
    n845
  );


  nor
  g851
  (
    n871,
    n722,
    n627,
    n673,
    n677
  );


  nand
  g852
  (
    n910,
    n834,
    n642,
    n717,
    n845
  );


  or
  g853
  (
    n851,
    n638,
    n796,
    n636,
    n613
  );


  nand
  g854
  (
    KeyWire_0_3,
    n617,
    n793,
    n641,
    n796
  );


  or
  g855
  (
    n872,
    n624,
    n638,
    n726,
    n794
  );


  and
  g856
  (
    n905,
    n628,
    n838,
    n626,
    n621
  );


  nor
  g857
  (
    n913,
    n673,
    n846,
    n832,
    n100
  );


  and
  g858
  (
    n931,
    n632,
    n633,
    n628,
    n840
  );


  xnor
  g859
  (
    n928,
    n839,
    n641,
    n636,
    n642
  );


  or
  g860
  (
    n891,
    n616,
    n848,
    n724,
    n676
  );


  nor
  g861
  (
    n934,
    n834,
    n722,
    n843,
    n828
  );


  nand
  g862
  (
    n932,
    n839,
    n714,
    n670,
    n720
  );


  nor
  g863
  (
    n899,
    n844,
    n626,
    n723,
    n575
  );


  xnor
  g864
  (
    n924,
    n849,
    n795,
    n671,
    n639
  );


  or
  g865
  (
    n893,
    n623,
    n796,
    n850,
    n673
  );


  nand
  g866
  (
    n880,
    n718,
    n615,
    n849,
    n619
  );


  xor
  g867
  (
    n892,
    n637,
    n795,
    n831,
    n99
  );


  and
  g868
  (
    n942,
    n677,
    n850,
    n720,
    n582
  );


  nor
  g869
  (
    n853,
    n672,
    n621,
    n849,
    n797
  );


  xnor
  g870
  (
    n890,
    n629,
    n640,
    n571,
    n624
  );


  and
  g871
  (
    n906,
    n622,
    n631,
    n794,
    n625
  );


  nor
  g872
  (
    n856,
    n716,
    n723,
    n626,
    n847
  );


  and
  g873
  (
    n922,
    n837,
    n618,
    n713,
    n714
  );


  xor
  g874
  (
    n926,
    n727,
    n642,
    n849,
    n829
  );


  nor
  g875
  (
    n907,
    n716,
    n629,
    n721,
    n623
  );


  nor
  g876
  (
    n854,
    n714,
    n634,
    n630,
    n622
  );


  xor
  g877
  (
    n915,
    n625,
    n635,
    n638,
    n723
  );


  nor
  g878
  (
    n864,
    n715,
    n834,
    n827,
    n632
  );


  xor
  g879
  (
    n877,
    n833,
    n639,
    n724,
    n827
  );


  and
  g880
  (
    n882,
    n830,
    n613,
    n796,
    n618
  );


  xor
  g881
  (
    n889,
    n713,
    n99,
    n850,
    n630
  );


  and
  g882
  (
    n919,
    n798,
    n832,
    n623,
    n634
  );


  nor
  g883
  (
    n887,
    n627,
    n569,
    n714,
    n612
  );


  or
  g884
  (
    n912,
    n831,
    n611,
    n615,
    n850
  );


  and
  g885
  (
    n930,
    n625,
    n612,
    n100,
    n627
  );


  xor
  g886
  (
    n908,
    n836,
    n719,
    n830,
    n725
  );


  nor
  g887
  (
    n944,
    n833,
    n622,
    n829,
    n100
  );


  nor
  g888
  (
    n918,
    n641,
    n726,
    n626,
    n573
  );


  and
  g889
  (
    n939,
    n636,
    n567,
    n799,
    n797
  );


  nor
  g890
  (
    n897,
    n620,
    n624,
    n671,
    n615
  );


  or
  g891
  (
    n884,
    n634,
    n793,
    n677,
    n636
  );


  xnor
  g892
  (
    n866,
    n725,
    n620,
    n727,
    n675
  );


  or
  g893
  (
    n909,
    n829,
    n842,
    n843,
    n635
  );


  and
  g894
  (
    n885,
    n639,
    n613,
    n713,
    n725
  );


  xor
  g895
  (
    n943,
    n637,
    n841,
    n721,
    n840
  );


  or
  g896
  (
    n883,
    n793,
    n628,
    n611,
    n614
  );


  nand
  g897
  (
    n933,
    n797,
    n795,
    n836,
    n838
  );


  and
  g898
  (
    n901,
    n724,
    n676,
    n795,
    n835
  );


  and
  g899
  (
    n940,
    n839,
    n833,
    n581,
    n637
  );


  and
  g900
  (
    n863,
    n838,
    n669,
    n797,
    n642
  );


  nor
  g901
  (
    n917,
    n726,
    n670,
    n830,
    n619
  );


  or
  g902
  (
    n859,
    n565,
    n618,
    n640,
    n722
  );


  and
  g903
  (
    n873,
    n670,
    n847,
    n839,
    n837
  );


  or
  g904
  (
    n903,
    n838,
    n843,
    n844,
    n580
  );


  xor
  g905
  (
    n869,
    n100,
    n676,
    n719,
    n723
  );


  and
  g906
  (
    n927,
    n616,
    n618,
    n837,
    n579
  );


  or
  g907
  (
    n876,
    n718,
    n631,
    n715,
    n624
  );


  xnor
  g908
  (
    n904,
    n798,
    n630,
    n675,
    n829
  );


  or
  g909
  (
    n874,
    n720,
    n717,
    n633,
    n719
  );


  nor
  g910
  (
    n867,
    n611,
    n635,
    n717,
    n101
  );


  and
  g911
  (
    n894,
    n798,
    n715,
    n561,
    n835
  );


  not
  g912
  (
    n945,
    n858
  );


  buf
  g913
  (
    n946,
    n854
  );


  not
  g914
  (
    n954,
    n727
  );


  buf
  g915
  (
    n947,
    n855
  );


  buf
  g916
  (
    n950,
    n859
  );


  buf
  g917
  (
    n948,
    n852
  );


  buf
  g918
  (
    n953,
    n857
  );


  not
  g919
  (
    n951,
    n727
  );


  not
  g920
  (
    n952,
    n856
  );


  xnor
  g921
  (
    n949,
    n860,
    n851,
    n853
  );


  nor
  g922
  (
    n966,
    n645,
    n947,
    n730,
    n946
  );


  xnor
  g923
  (
    n974,
    n644,
    n110,
    n105,
    n108
  );


  xnor
  g924
  (
    n973,
    n729,
    n117,
    n105,
    n948
  );


  xor
  g925
  (
    n981,
    n730,
    n103,
    n107,
    n104
  );


  nor
  g926
  (
    n979,
    n950,
    n107,
    n949,
    n948
  );


  or
  g927
  (
    n989,
    n115,
    n111,
    n950,
    n103
  );


  nand
  g928
  (
    n983,
    n728,
    n646,
    n949,
    n643
  );


  nor
  g929
  (
    n955,
    n102,
    n104,
    n113
  );


  nor
  g930
  (
    n991,
    n108,
    n106,
    n643,
    n647
  );


  or
  g931
  (
    n980,
    n118,
    n112,
    n111,
    n946
  );


  xor
  g932
  (
    n984,
    n948,
    n117,
    n107,
    n728
  );


  nor
  g933
  (
    KeyWire_0_15,
    n953,
    n102,
    n644
  );


  xnor
  g934
  (
    n978,
    n646,
    n949,
    n116
  );


  nor
  g935
  (
    n965,
    n646,
    n947,
    n729,
    n775
  );


  nand
  g936
  (
    n971,
    n105,
    n107,
    n948,
    n952
  );


  or
  g937
  (
    n987,
    n777,
    n950,
    n114,
    n104
  );


  or
  g938
  (
    n957,
    n954,
    n109,
    n108,
    n952
  );


  xor
  g939
  (
    n962,
    n645,
    n111,
    n114,
    n947
  );


  nand
  g940
  (
    n990,
    n106,
    n951,
    n731
  );


  nand
  g941
  (
    n982,
    n731,
    n113,
    n103,
    n952
  );


  nand
  g942
  (
    n967,
    n774,
    n954,
    n946,
    n729
  );


  nand
  g943
  (
    n970,
    n945,
    n111,
    n731,
    n112
  );


  xor
  g944
  (
    n988,
    n647,
    n118,
    n779,
    n953
  );


  or
  g945
  (
    KeyWire_0_7,
    n116,
    n108,
    n106,
    n101
  );


  xor
  g946
  (
    n976,
    n110,
    n728,
    n117,
    n954
  );


  or
  g947
  (
    n985,
    n115,
    n110,
    n101,
    n949
  );


  xnor
  g948
  (
    n968,
    n954,
    n730,
    n109,
    n118
  );


  nand
  g949
  (
    n986,
    n113,
    n730,
    n112,
    n109
  );


  or
  g950
  (
    n959,
    n953,
    n114,
    n946,
    n646
  );


  xor
  g951
  (
    n964,
    n114,
    n109,
    n729,
    n644
  );


  and
  g952
  (
    n977,
    n110,
    n643,
    n951,
    n947
  );


  nand
  g953
  (
    n956,
    n102,
    n103,
    n644,
    n113
  );


  xor
  g954
  (
    n961,
    n950,
    n952,
    n117,
    n778
  );


  or
  g955
  (
    n972,
    n105,
    n106,
    n115
  );


  xnor
  g956
  (
    n963,
    n116,
    n112,
    n953,
    n643
  );


  xor
  g957
  (
    n958,
    n645,
    n951,
    n776,
    n731
  );


  nor
  g958
  (
    n975,
    n645,
    n647,
    n728
  );


  xor
  g959
  (
    n996,
    n732,
    n975,
    n960,
    n963
  );


  xor
  g960
  (
    n992,
    n912,
    n900,
    n932,
    n918
  );


  or
  g961
  (
    n1013,
    n902,
    n940,
    n890,
    n982
  );


  xor
  g962
  (
    n1006,
    n898,
    n882,
    n583,
    n961
  );


  or
  g963
  (
    n1017,
    n732,
    n910,
    n985,
    n892
  );


  xnor
  g964
  (
    n1011,
    n916,
    n894,
    n964,
    n974
  );


  xnor
  g965
  (
    n1018,
    n965,
    n938,
    n939,
    n906
  );


  nand
  g966
  (
    n1010,
    n970,
    n862,
    n891,
    n986
  );


  nand
  g967
  (
    n1009,
    n929,
    n958,
    n887,
    n903
  );


  and
  g968
  (
    n1005,
    n899,
    n914,
    n959,
    n927
  );


  nor
  g969
  (
    n999,
    n880,
    n989,
    n864,
    n981
  );


  nor
  g970
  (
    n1020,
    n878,
    n926,
    n913,
    n941
  );


  or
  g971
  (
    n1012,
    n978,
    n872,
    n943,
    n922
  );


  nor
  g972
  (
    n1004,
    n583,
    n920,
    n930,
    n935
  );


  xnor
  g973
  (
    n1021,
    n869,
    n988,
    n921,
    n861
  );


  xor
  g974
  (
    n998,
    n908,
    n917,
    n972,
    n934
  );


  and
  g975
  (
    n1016,
    n968,
    n889,
    n937,
    n990
  );


  xnor
  g976
  (
    n993,
    n911,
    n886,
    n871,
    n944
  );


  nand
  g977
  (
    n1002,
    n969,
    n732,
    n919,
    n987
  );


  nor
  g978
  (
    n1003,
    n883,
    n955,
    n866,
    n976
  );


  nor
  g979
  (
    n994,
    n973,
    n896,
    n925,
    n881
  );


  nor
  g980
  (
    n1007,
    n909,
    n924,
    n991,
    n867
  );


  xnor
  g981
  (
    n1015,
    n983,
    n868,
    n984,
    n876
  );


  nor
  g982
  (
    n1001,
    n732,
    n865,
    n888,
    n933
  );


  nor
  g983
  (
    n997,
    n863,
    n956,
    n877,
    n875
  );


  or
  g984
  (
    n1000,
    n879,
    n923,
    n897,
    n971
  );


  or
  g985
  (
    n1014,
    n870,
    n967,
    n901,
    n966
  );


  and
  g986
  (
    n1008,
    n942,
    n907,
    n931,
    n118
  );


  or
  g987
  (
    n1022,
    n928,
    n905,
    n979,
    n873
  );


  xnor
  g988
  (
    n1023,
    n915,
    n895,
    n962,
    n893
  );


  nor
  g989
  (
    n995,
    n874,
    n980,
    n904,
    n936
  );


  nand
  g990
  (
    n1019,
    n884,
    n885,
    n957,
    n977
  );


  xor
  g991
  (
    n1027,
    n1012,
    n995,
    n826,
    n1020
  );


  xnor
  g992
  (
    n1032,
    n1008,
    n1010,
    n997,
    n1004
  );


  nor
  g993
  (
    n1024,
    n1009,
    n1015,
    n1000,
    n1023
  );


  nor
  g994
  (
    n1030,
    n1016,
    n993,
    n1007,
    n1021
  );


  xor
  g995
  (
    n1029,
    n1014,
    n998,
    n1017,
    n1006
  );


  and
  g996
  (
    n1028,
    n1001,
    n1018,
    n1002,
    n1005
  );


  or
  g997
  (
    n1026,
    n1003,
    n826,
    n1011,
    n994
  );


  nand
  g998
  (
    n1031,
    n996,
    n992,
    n1019,
    n1013
  );


  xnor
  g999
  (
    n1025,
    n825,
    n999,
    n1022,
    n824
  );


  xor
  KeyGate_0_0
  (
    n312,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n255,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n473,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n881,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n629,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n387,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n669,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n969,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n292,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n541,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n304,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n137,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n75,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n125,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n799,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n960,
    KeyNOTWire_0_15
  );


endmodule


